magic
tech sky130B
magscale 1 2
timestamp 1680009009
<< metal1 >>
rect 397454 700680 397460 700732
rect 397512 700720 397518 700732
rect 418798 700720 418804 700732
rect 397512 700692 418804 700720
rect 397512 700680 397518 700692
rect 418798 700680 418804 700692
rect 418856 700680 418862 700732
rect 444282 700680 444288 700732
rect 444340 700720 444346 700732
rect 478506 700720 478512 700732
rect 444340 700692 478512 700720
rect 444340 700680 444346 700692
rect 478506 700680 478512 700692
rect 478564 700680 478570 700732
rect 364978 700612 364984 700664
rect 365036 700652 365042 700664
rect 446398 700652 446404 700664
rect 365036 700624 446404 700652
rect 365036 700612 365042 700624
rect 446398 700612 446404 700624
rect 446456 700612 446462 700664
rect 332502 700544 332508 700596
rect 332560 700584 332566 700596
rect 445018 700584 445024 700596
rect 332560 700556 445024 700584
rect 332560 700544 332566 700556
rect 445018 700544 445024 700556
rect 445076 700544 445082 700596
rect 218974 700476 218980 700528
rect 219032 700516 219038 700528
rect 416038 700516 416044 700528
rect 219032 700488 416044 700516
rect 219032 700476 219038 700488
rect 416038 700476 416044 700488
rect 416096 700476 416102 700528
rect 444190 700476 444196 700528
rect 444248 700516 444254 700528
rect 494790 700516 494796 700528
rect 444248 700488 494796 700516
rect 444248 700476 444254 700488
rect 494790 700476 494796 700488
rect 494848 700476 494854 700528
rect 235166 700408 235172 700460
rect 235224 700448 235230 700460
rect 446490 700448 446496 700460
rect 235224 700420 446496 700448
rect 235224 700408 235230 700420
rect 446490 700408 446496 700420
rect 446548 700408 446554 700460
rect 170306 700340 170312 700392
rect 170364 700380 170370 700392
rect 449158 700380 449164 700392
rect 170364 700352 449164 700380
rect 170364 700340 170370 700352
rect 449158 700340 449164 700352
rect 449216 700340 449222 700392
rect 137830 700272 137836 700324
rect 137888 700312 137894 700324
rect 445110 700312 445116 700324
rect 137888 700284 445116 700312
rect 137888 700272 137894 700284
rect 445110 700272 445116 700284
rect 445168 700272 445174 700324
rect 527174 700272 527180 700324
rect 527232 700312 527238 700324
rect 543734 700312 543740 700324
rect 527232 700284 543740 700312
rect 527232 700272 527238 700284
rect 543734 700272 543740 700284
rect 543792 700272 543798 700324
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 446582 683176 446588 683188
rect 3476 683148 446588 683176
rect 3476 683136 3482 683148
rect 446582 683136 446588 683148
rect 446640 683136 446646 683188
rect 570598 683136 570604 683188
rect 570656 683176 570662 683188
rect 579614 683176 579620 683188
rect 570656 683148 579620 683176
rect 570656 683136 570662 683148
rect 579614 683136 579620 683148
rect 579672 683136 579678 683188
rect 448422 679600 448428 679652
rect 448480 679640 448486 679652
rect 462314 679640 462320 679652
rect 448480 679612 462320 679640
rect 448480 679600 448486 679612
rect 462314 679600 462320 679612
rect 462372 679600 462378 679652
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 446766 670732 446772 670744
rect 3568 670704 446772 670732
rect 3568 670692 3574 670704
rect 446766 670692 446772 670704
rect 446824 670692 446830 670744
rect 573358 670692 573364 670744
rect 573416 670732 573422 670744
rect 580166 670732 580172 670744
rect 573416 670704 580172 670732
rect 573416 670692 573422 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 348786 670216 348792 670268
rect 348844 670256 348850 670268
rect 446858 670256 446864 670268
rect 348844 670228 446864 670256
rect 348844 670216 348850 670228
rect 446858 670216 446864 670228
rect 446916 670216 446922 670268
rect 283834 670148 283840 670200
rect 283892 670188 283898 670200
rect 445202 670188 445208 670200
rect 283892 670160 445208 670188
rect 283892 670148 283898 670160
rect 445202 670148 445208 670160
rect 445260 670148 445266 670200
rect 154114 670080 154120 670132
rect 154172 670120 154178 670132
rect 446674 670120 446680 670132
rect 154172 670092 446680 670120
rect 154172 670080 154178 670092
rect 446674 670080 446680 670092
rect 446732 670080 446738 670132
rect 89162 670012 89168 670064
rect 89220 670052 89226 670064
rect 413278 670052 413284 670064
rect 89220 670024 413284 670052
rect 89220 670012 89226 670024
rect 413278 670012 413284 670024
rect 413336 670012 413342 670064
rect 72970 669944 72976 669996
rect 73028 669984 73034 669996
rect 418890 669984 418896 669996
rect 73028 669956 418896 669984
rect 73028 669944 73034 669956
rect 418890 669944 418896 669956
rect 418948 669944 418954 669996
rect 267642 668788 267648 668840
rect 267700 668828 267706 668840
rect 445294 668828 445300 668840
rect 267700 668800 445300 668828
rect 267700 668788 267706 668800
rect 445294 668788 445300 668800
rect 445352 668788 445358 668840
rect 23474 668720 23480 668772
rect 23532 668760 23538 668772
rect 380434 668760 380440 668772
rect 23532 668732 380440 668760
rect 23532 668720 23538 668732
rect 380434 668720 380440 668732
rect 380492 668720 380498 668772
rect 20714 668652 20720 668704
rect 20772 668692 20778 668704
rect 378318 668692 378324 668704
rect 20772 668664 378324 668692
rect 20772 668652 20778 668664
rect 378318 668652 378324 668664
rect 378376 668652 378382 668704
rect 20990 668584 20996 668636
rect 21048 668624 21054 668636
rect 378134 668624 378140 668636
rect 21048 668596 378140 668624
rect 21048 668584 21054 668596
rect 378134 668584 378140 668596
rect 378192 668584 378198 668636
rect 21082 668516 21088 668568
rect 21140 668556 21146 668568
rect 380342 668556 380348 668568
rect 21140 668528 380348 668556
rect 21140 668516 21146 668528
rect 380342 668516 380348 668528
rect 380400 668516 380406 668568
rect 20898 668448 20904 668500
rect 20956 668488 20962 668500
rect 380618 668488 380624 668500
rect 20956 668460 380624 668488
rect 20956 668448 20962 668460
rect 380618 668448 380624 668460
rect 380676 668448 380682 668500
rect 18874 668380 18880 668432
rect 18932 668420 18938 668432
rect 378226 668420 378232 668432
rect 18932 668392 378232 668420
rect 18932 668380 18938 668392
rect 378226 668380 378232 668392
rect 378284 668380 378290 668432
rect 20806 668312 20812 668364
rect 20864 668352 20870 668364
rect 381814 668352 381820 668364
rect 20864 668324 381820 668352
rect 20864 668312 20870 668324
rect 381814 668312 381820 668324
rect 381872 668312 381878 668364
rect 19334 668244 19340 668296
rect 19392 668284 19398 668296
rect 381538 668284 381544 668296
rect 19392 668256 381544 668284
rect 19392 668244 19398 668256
rect 381538 668244 381544 668256
rect 381596 668244 381602 668296
rect 18782 668176 18788 668228
rect 18840 668216 18846 668228
rect 380158 668216 380164 668228
rect 18840 668188 380164 668216
rect 18840 668176 18846 668188
rect 380158 668176 380164 668188
rect 380216 668176 380222 668228
rect 17862 668108 17868 668160
rect 17920 668148 17926 668160
rect 381630 668148 381636 668160
rect 17920 668120 381636 668148
rect 17920 668108 17926 668120
rect 381630 668108 381636 668120
rect 381688 668108 381694 668160
rect 7558 668040 7564 668092
rect 7616 668080 7622 668092
rect 381906 668080 381912 668092
rect 7616 668052 381912 668080
rect 7616 668040 7622 668052
rect 381906 668040 381912 668052
rect 381964 668040 381970 668092
rect 3786 667972 3792 668024
rect 3844 668012 3850 668024
rect 447042 668012 447048 668024
rect 3844 667984 447048 668012
rect 3844 667972 3850 667984
rect 447042 667972 447048 667984
rect 447100 667972 447106 668024
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 446950 667944 446956 667956
rect 3476 667916 446956 667944
rect 3476 667904 3482 667916
rect 446950 667904 446956 667916
rect 447008 667904 447014 667956
rect 378134 667836 378140 667888
rect 378192 667876 378198 667888
rect 380250 667876 380256 667888
rect 378192 667848 380256 667876
rect 378192 667836 378198 667848
rect 380250 667836 380256 667848
rect 380308 667836 380314 667888
rect 19886 667768 19892 667820
rect 19944 667808 19950 667820
rect 23474 667808 23480 667820
rect 19944 667780 23480 667808
rect 19944 667768 19950 667780
rect 23474 667768 23480 667780
rect 23532 667768 23538 667820
rect 378226 667768 378232 667820
rect 378284 667808 378290 667820
rect 381722 667808 381728 667820
rect 378284 667780 381728 667808
rect 378284 667768 378290 667780
rect 381722 667768 381728 667780
rect 381780 667768 381786 667820
rect 19794 667700 19800 667752
rect 19852 667740 19858 667752
rect 20990 667740 20996 667752
rect 19852 667712 20996 667740
rect 19852 667700 19858 667712
rect 20990 667700 20996 667712
rect 21048 667700 21054 667752
rect 378318 667700 378324 667752
rect 378376 667740 378382 667752
rect 380526 667740 380532 667752
rect 378376 667712 380532 667740
rect 378376 667700 378382 667712
rect 380526 667700 380532 667712
rect 380584 667700 380590 667752
rect 18690 667632 18696 667684
rect 18748 667672 18754 667684
rect 21082 667672 21088 667684
rect 18748 667644 21088 667672
rect 18748 667632 18754 667644
rect 21082 667632 21088 667644
rect 21140 667632 21146 667684
rect 21358 667632 21364 667684
rect 21416 667672 21422 667684
rect 420178 667672 420184 667684
rect 21416 667644 420184 667672
rect 21416 667632 21422 667644
rect 420178 667632 420184 667644
rect 420236 667632 420242 667684
rect 3694 667564 3700 667616
rect 3752 667604 3758 667616
rect 418982 667604 418988 667616
rect 3752 667576 418988 667604
rect 3752 667564 3758 667576
rect 418982 667564 418988 667576
rect 419040 667564 419046 667616
rect 18414 666680 18420 666732
rect 18472 666720 18478 666732
rect 20806 666720 20812 666732
rect 18472 666692 20812 666720
rect 18472 666680 18478 666692
rect 20806 666680 20812 666692
rect 20864 666680 20870 666732
rect 17678 666612 17684 666664
rect 17736 666652 17742 666664
rect 19334 666652 19340 666664
rect 17736 666624 19340 666652
rect 17736 666612 17742 666624
rect 19334 666612 19340 666624
rect 19392 666612 19398 666664
rect 20070 666612 20076 666664
rect 20128 666652 20134 666664
rect 20714 666652 20720 666664
rect 20128 666624 20720 666652
rect 20128 666612 20134 666624
rect 20714 666612 20720 666624
rect 20772 666612 20778 666664
rect 19978 666544 19984 666596
rect 20036 666584 20042 666596
rect 20898 666584 20904 666596
rect 20036 666556 20904 666584
rect 20036 666544 20042 666556
rect 20898 666544 20904 666556
rect 20956 666544 20962 666596
rect 16574 665456 16580 665508
rect 16632 665496 16638 665508
rect 19886 665496 19892 665508
rect 16632 665468 19892 665496
rect 16632 665456 16638 665468
rect 19886 665456 19892 665468
rect 19944 665456 19950 665508
rect 13814 665252 13820 665304
rect 13872 665292 13878 665304
rect 17862 665292 17868 665304
rect 13872 665264 17868 665292
rect 13872 665252 13878 665264
rect 17862 665252 17868 665264
rect 17920 665252 17926 665304
rect 17678 665224 17684 665236
rect 13832 665196 17684 665224
rect 10962 665116 10968 665168
rect 11020 665156 11026 665168
rect 13832 665156 13860 665196
rect 17678 665184 17684 665196
rect 17736 665184 17742 665236
rect 11020 665128 13860 665156
rect 11020 665116 11026 665128
rect 18598 664640 18604 664692
rect 18656 664680 18662 664692
rect 19794 664680 19800 664692
rect 18656 664652 19800 664680
rect 18656 664640 18662 664652
rect 19794 664640 19800 664652
rect 19852 664640 19858 664692
rect 11054 663756 11060 663808
rect 11112 663796 11118 663808
rect 16574 663796 16580 663808
rect 11112 663768 16580 663796
rect 11112 663756 11118 663768
rect 16574 663756 16580 663768
rect 16632 663756 16638 663808
rect 18414 663796 18420 663808
rect 16684 663768 18420 663796
rect 15286 663688 15292 663740
rect 15344 663728 15350 663740
rect 16684 663728 16712 663768
rect 18414 663756 18420 663768
rect 18472 663756 18478 663808
rect 15344 663700 16712 663728
rect 15344 663688 15350 663700
rect 17954 662464 17960 662516
rect 18012 662504 18018 662516
rect 20070 662504 20076 662516
rect 18012 662476 20076 662504
rect 18012 662464 18018 662476
rect 20070 662464 20076 662476
rect 20128 662464 20134 662516
rect 8662 662396 8668 662448
rect 8720 662436 8726 662448
rect 10962 662436 10968 662448
rect 8720 662408 10968 662436
rect 8720 662396 8726 662408
rect 10962 662396 10968 662408
rect 11020 662396 11026 662448
rect 13906 662396 13912 662448
rect 13964 662436 13970 662448
rect 18690 662436 18696 662448
rect 13964 662408 18696 662436
rect 13964 662396 13970 662408
rect 18690 662396 18696 662408
rect 18748 662396 18754 662448
rect 14458 661648 14464 661700
rect 14516 661688 14522 661700
rect 18782 661688 18788 661700
rect 14516 661660 18788 661688
rect 14516 661648 14522 661660
rect 18782 661648 18788 661660
rect 18840 661648 18846 661700
rect 18874 661144 18880 661156
rect 16546 661116 18880 661144
rect 15286 661076 15292 661088
rect 13832 661048 15292 661076
rect 11698 660968 11704 661020
rect 11756 661008 11762 661020
rect 13832 661008 13860 661048
rect 15286 661036 15292 661048
rect 15344 661036 15350 661088
rect 11756 660980 13860 661008
rect 11756 660968 11762 660980
rect 15194 660968 15200 661020
rect 15252 661008 15258 661020
rect 16546 661008 16574 661116
rect 18874 661104 18880 661116
rect 18932 661104 18938 661156
rect 18690 661036 18696 661088
rect 18748 661076 18754 661088
rect 19978 661076 19984 661088
rect 18748 661048 19984 661076
rect 18748 661036 18754 661048
rect 19978 661036 19984 661048
rect 20036 661036 20042 661088
rect 382274 661036 382280 661088
rect 382332 661076 382338 661088
rect 403618 661076 403624 661088
rect 382332 661048 403624 661076
rect 382332 661036 382338 661048
rect 403618 661036 403624 661048
rect 403676 661036 403682 661088
rect 15252 660980 16574 661008
rect 15252 660968 15258 660980
rect 5626 660288 5632 660340
rect 5684 660328 5690 660340
rect 7558 660328 7564 660340
rect 5684 660300 7564 660328
rect 5684 660288 5690 660300
rect 7558 660288 7564 660300
rect 7616 660288 7622 660340
rect 5534 659744 5540 659796
rect 5592 659784 5598 659796
rect 8662 659784 8668 659796
rect 5592 659756 8668 659784
rect 5592 659744 5598 659756
rect 8662 659744 8668 659756
rect 8720 659744 8726 659796
rect 9582 659676 9588 659728
rect 9640 659716 9646 659728
rect 13814 659716 13820 659728
rect 9640 659688 13820 659716
rect 9640 659676 9646 659688
rect 13814 659676 13820 659688
rect 13872 659676 13878 659728
rect 11054 658288 11060 658300
rect 9692 658260 11060 658288
rect 8938 658180 8944 658232
rect 8996 658220 9002 658232
rect 9692 658220 9720 658260
rect 11054 658248 11060 658260
rect 11112 658248 11118 658300
rect 8996 658192 9720 658220
rect 8996 658180 9002 658192
rect 14642 657296 14648 657348
rect 14700 657336 14706 657348
rect 15194 657336 15200 657348
rect 14700 657308 15200 657336
rect 14700 657296 14706 657308
rect 15194 657296 15200 657308
rect 15252 657296 15258 657348
rect 10042 656344 10048 656396
rect 10100 656384 10106 656396
rect 13906 656384 13912 656396
rect 10100 656356 13912 656384
rect 10100 656344 10106 656356
rect 13906 656344 13912 656356
rect 13964 656344 13970 656396
rect 7098 656276 7104 656328
rect 7156 656316 7162 656328
rect 9582 656316 9588 656328
rect 7156 656288 9588 656316
rect 7156 656276 7162 656288
rect 9582 656276 9588 656288
rect 9640 656276 9646 656328
rect 460474 655800 460480 655852
rect 460532 655840 460538 655852
rect 460658 655840 460664 655852
rect 460532 655812 460664 655840
rect 460532 655800 460538 655812
rect 460658 655800 460664 655812
rect 460716 655800 460722 655852
rect 5626 655568 5632 655580
rect 4172 655540 5632 655568
rect 3418 655460 3424 655512
rect 3476 655500 3482 655512
rect 4172 655500 4200 655540
rect 5626 655528 5632 655540
rect 5684 655528 5690 655580
rect 15930 655528 15936 655580
rect 15988 655568 15994 655580
rect 17862 655568 17868 655580
rect 15988 655540 17868 655568
rect 15988 655528 15994 655540
rect 17862 655528 17868 655540
rect 17920 655528 17926 655580
rect 3476 655472 4200 655500
rect 3476 655460 3482 655472
rect 4798 654440 4804 654492
rect 4856 654480 4862 654492
rect 5534 654480 5540 654492
rect 4856 654452 5540 654480
rect 4856 654440 4862 654452
rect 5534 654440 5540 654452
rect 5592 654440 5598 654492
rect 8294 652876 8300 652928
rect 8352 652916 8358 652928
rect 14458 652916 14464 652928
rect 8352 652888 14464 652916
rect 8352 652876 8358 652888
rect 14458 652876 14464 652888
rect 14516 652876 14522 652928
rect 5626 652808 5632 652860
rect 5684 652848 5690 652860
rect 8938 652848 8944 652860
rect 5684 652820 8944 652848
rect 5684 652808 5690 652820
rect 8938 652808 8944 652820
rect 8996 652808 9002 652860
rect 7098 652780 7104 652792
rect 6886 652752 7104 652780
rect 5074 652672 5080 652724
rect 5132 652712 5138 652724
rect 6886 652712 6914 652752
rect 7098 652740 7104 652752
rect 7156 652740 7162 652792
rect 9214 652740 9220 652792
rect 9272 652780 9278 652792
rect 11698 652780 11704 652792
rect 9272 652752 11704 652780
rect 9272 652740 9278 652752
rect 11698 652740 11704 652752
rect 11756 652740 11762 652792
rect 17034 652740 17040 652792
rect 17092 652780 17098 652792
rect 18690 652780 18696 652792
rect 17092 652752 18696 652780
rect 17092 652740 17098 652752
rect 18690 652740 18696 652752
rect 18748 652740 18754 652792
rect 5132 652684 6914 652712
rect 5132 652672 5138 652684
rect 3510 651992 3516 652044
rect 3568 652032 3574 652044
rect 10042 652032 10048 652044
rect 3568 652004 10048 652032
rect 3568 651992 3574 652004
rect 10042 651992 10048 652004
rect 10100 651992 10106 652044
rect 12434 651448 12440 651500
rect 12492 651488 12498 651500
rect 14642 651488 14648 651500
rect 12492 651460 14648 651488
rect 12492 651448 12498 651460
rect 14642 651448 14648 651460
rect 14700 651448 14706 651500
rect 13814 651380 13820 651432
rect 13872 651420 13878 651432
rect 15930 651420 15936 651432
rect 13872 651392 15936 651420
rect 13872 651380 13878 651392
rect 15930 651380 15936 651392
rect 15988 651380 15994 651432
rect 382274 651380 382280 651432
rect 382332 651420 382338 651432
rect 396718 651420 396724 651432
rect 382332 651392 396724 651420
rect 382332 651380 382338 651392
rect 396718 651380 396724 651392
rect 396776 651380 396782 651432
rect 5534 650224 5540 650276
rect 5592 650264 5598 650276
rect 9214 650264 9220 650276
rect 5592 650236 9220 650264
rect 5592 650224 5598 650236
rect 9214 650224 9220 650236
rect 9272 650224 9278 650276
rect 5626 650060 5632 650072
rect 4172 650032 5632 650060
rect 3602 649952 3608 650004
rect 3660 649992 3666 650004
rect 4172 649992 4200 650032
rect 5626 650020 5632 650032
rect 5684 650020 5690 650072
rect 3660 649964 4200 649992
rect 3660 649952 3666 649964
rect 4890 649680 4896 649732
rect 4948 649720 4954 649732
rect 8202 649720 8208 649732
rect 4948 649692 8208 649720
rect 4948 649680 4954 649692
rect 8202 649680 8208 649692
rect 8260 649680 8266 649732
rect 12434 648632 12440 648644
rect 11072 648604 12440 648632
rect 8938 648524 8944 648576
rect 8996 648564 9002 648576
rect 11072 648564 11100 648604
rect 12434 648592 12440 648604
rect 12492 648592 12498 648644
rect 18598 648632 18604 648644
rect 16546 648604 18604 648632
rect 8996 648536 11100 648564
rect 8996 648524 9002 648536
rect 15194 648524 15200 648576
rect 15252 648564 15258 648576
rect 16546 648564 16574 648604
rect 18598 648592 18604 648604
rect 18656 648592 18662 648644
rect 15252 648536 16574 648564
rect 15252 648524 15258 648536
rect 11054 646552 11060 646604
rect 11112 646592 11118 646604
rect 13814 646592 13820 646604
rect 11112 646564 13820 646592
rect 11112 646552 11118 646564
rect 13814 646552 13820 646564
rect 13872 646552 13878 646604
rect 13078 645940 13084 645992
rect 13136 645980 13142 645992
rect 17034 645980 17040 645992
rect 13136 645952 17040 645980
rect 13136 645940 13142 645952
rect 17034 645940 17040 645952
rect 17092 645940 17098 645992
rect 12434 645464 12440 645516
rect 12492 645504 12498 645516
rect 15194 645504 15200 645516
rect 12492 645476 15200 645504
rect 12492 645464 12498 645476
rect 15194 645464 15200 645476
rect 15252 645464 15258 645516
rect 460290 643696 460296 643748
rect 460348 643736 460354 643748
rect 460750 643736 460756 643748
rect 460348 643708 460756 643736
rect 460348 643696 460354 643708
rect 460750 643696 460756 643708
rect 460808 643696 460814 643748
rect 8938 643124 8944 643136
rect 6886 643096 8944 643124
rect 4982 643016 4988 643068
rect 5040 643056 5046 643068
rect 6886 643056 6914 643096
rect 8938 643084 8944 643096
rect 8996 643084 9002 643136
rect 5040 643028 6914 643056
rect 5040 643016 5046 643028
rect 11054 640336 11060 640348
rect 9692 640308 11060 640336
rect 8938 640228 8944 640280
rect 8996 640268 9002 640280
rect 9692 640268 9720 640308
rect 11054 640296 11060 640308
rect 11112 640296 11118 640348
rect 8996 640240 9720 640268
rect 8996 640228 9002 640240
rect 9674 637712 9680 637764
rect 9732 637752 9738 637764
rect 12342 637752 12348 637764
rect 9732 637724 12348 637752
rect 9732 637712 9738 637724
rect 12342 637712 12348 637724
rect 12400 637712 12406 637764
rect 6914 636148 6920 636200
rect 6972 636188 6978 636200
rect 9674 636188 9680 636200
rect 6972 636160 9680 636188
rect 6972 636148 6978 636160
rect 9674 636148 9680 636160
rect 9732 636148 9738 636200
rect 13078 632108 13084 632120
rect 11072 632080 13084 632108
rect 10686 632000 10692 632052
rect 10744 632040 10750 632052
rect 11072 632040 11100 632080
rect 13078 632068 13084 632080
rect 13136 632068 13142 632120
rect 10744 632012 11100 632040
rect 10744 632000 10750 632012
rect 7926 631660 7932 631712
rect 7984 631700 7990 631712
rect 8938 631700 8944 631712
rect 7984 631672 8944 631700
rect 7984 631660 7990 631672
rect 8938 631660 8944 631672
rect 8996 631660 9002 631712
rect 3694 630640 3700 630692
rect 3752 630680 3758 630692
rect 6822 630680 6828 630692
rect 3752 630652 6828 630680
rect 3752 630640 3758 630652
rect 6822 630640 6828 630652
rect 6880 630640 6886 630692
rect 577498 630640 577504 630692
rect 577556 630680 577562 630692
rect 580442 630680 580448 630692
rect 577556 630652 580448 630680
rect 577556 630640 577562 630652
rect 580442 630640 580448 630652
rect 580500 630640 580506 630692
rect 382274 629280 382280 629332
rect 382332 629320 382338 629332
rect 395338 629320 395344 629332
rect 382332 629292 395344 629320
rect 382332 629280 382338 629292
rect 395338 629280 395344 629292
rect 395396 629280 395402 629332
rect 5534 628736 5540 628788
rect 5592 628776 5598 628788
rect 7926 628776 7932 628788
rect 5592 628748 7932 628776
rect 5592 628736 5598 628748
rect 7926 628736 7932 628748
rect 7984 628736 7990 628788
rect 4154 626900 4160 626952
rect 4212 626940 4218 626952
rect 5534 626940 5540 626952
rect 4212 626912 5540 626940
rect 4212 626900 4218 626912
rect 5534 626900 5540 626912
rect 5592 626900 5598 626952
rect 8938 625880 8944 625932
rect 8996 625920 9002 625932
rect 10686 625920 10692 625932
rect 8996 625892 10692 625920
rect 8996 625880 9002 625892
rect 10686 625880 10692 625892
rect 10744 625880 10750 625932
rect 382274 619624 382280 619676
rect 382332 619664 382338 619676
rect 399478 619664 399484 619676
rect 382332 619636 399484 619664
rect 382332 619624 382338 619636
rect 399478 619624 399484 619636
rect 399536 619624 399542 619676
rect 3142 619556 3148 619608
rect 3200 619596 3206 619608
rect 20898 619596 20904 619608
rect 3200 619568 20904 619596
rect 3200 619556 3206 619568
rect 20898 619556 20904 619568
rect 20956 619556 20962 619608
rect 7558 617924 7564 617976
rect 7616 617964 7622 617976
rect 8938 617964 8944 617976
rect 7616 617936 8944 617964
rect 7616 617924 7622 617936
rect 8938 617924 8944 617936
rect 8996 617924 9002 617976
rect 571978 616836 571984 616888
rect 572036 616876 572042 616888
rect 580166 616876 580172 616888
rect 572036 616848 580172 616876
rect 572036 616836 572042 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 457530 610648 457536 610700
rect 457588 610688 457594 610700
rect 457898 610688 457904 610700
rect 457588 610660 457904 610688
rect 457588 610648 457594 610660
rect 457898 610648 457904 610660
rect 457956 610648 457962 610700
rect 382274 608608 382280 608660
rect 382332 608648 382338 608660
rect 393958 608648 393964 608660
rect 382332 608620 393964 608648
rect 382332 608608 382338 608620
rect 393958 608608 393964 608620
rect 394016 608608 394022 608660
rect 460474 602896 460480 602948
rect 460532 602896 460538 602948
rect 460492 602676 460520 602896
rect 460474 602624 460480 602676
rect 460532 602624 460538 602676
rect 6178 601604 6184 601656
rect 6236 601644 6242 601656
rect 7558 601644 7564 601656
rect 6236 601616 7564 601644
rect 6236 601604 6242 601616
rect 7558 601604 7564 601616
rect 7616 601604 7622 601656
rect 460566 600652 460572 600704
rect 460624 600692 460630 600704
rect 461578 600692 461584 600704
rect 460624 600664 461584 600692
rect 460624 600652 460630 600664
rect 461578 600652 461584 600664
rect 461636 600652 461642 600704
rect 457898 600244 457904 600296
rect 457956 600284 457962 600296
rect 462958 600284 462964 600296
rect 457956 600256 462964 600284
rect 457956 600244 457962 600256
rect 462958 600244 462964 600256
rect 463016 600244 463022 600296
rect 457254 600176 457260 600228
rect 457312 600216 457318 600228
rect 463050 600216 463056 600228
rect 457312 600188 463056 600216
rect 457312 600176 457318 600188
rect 463050 600176 463056 600188
rect 463108 600176 463114 600228
rect 457530 599700 457536 599752
rect 457588 599740 457594 599752
rect 464338 599740 464344 599752
rect 457588 599712 464344 599740
rect 457588 599700 457594 599712
rect 464338 599700 464344 599712
rect 464396 599700 464402 599752
rect 457438 599632 457444 599684
rect 457496 599672 457502 599684
rect 467098 599672 467104 599684
rect 457496 599644 467104 599672
rect 457496 599632 457502 599644
rect 467098 599632 467104 599644
rect 467156 599632 467162 599684
rect 518158 599632 518164 599684
rect 518216 599672 518222 599684
rect 543734 599672 543740 599684
rect 518216 599644 543740 599672
rect 518216 599632 518222 599644
rect 543734 599632 543740 599644
rect 543792 599632 543798 599684
rect 460382 599564 460388 599616
rect 460440 599604 460446 599616
rect 503714 599604 503720 599616
rect 460440 599576 503720 599604
rect 460440 599564 460446 599576
rect 503714 599564 503720 599576
rect 503772 599564 503778 599616
rect 515398 599564 515404 599616
rect 515456 599604 515462 599616
rect 580350 599604 580356 599616
rect 515456 599576 580356 599604
rect 515456 599564 515462 599576
rect 580350 599564 580356 599576
rect 580408 599564 580414 599616
rect 457346 598408 457352 598460
rect 457404 598448 457410 598460
rect 468478 598448 468484 598460
rect 457404 598420 468484 598448
rect 457404 598408 457410 598420
rect 468478 598408 468484 598420
rect 468536 598408 468542 598460
rect 457806 598340 457812 598392
rect 457864 598380 457870 598392
rect 471238 598380 471244 598392
rect 457864 598352 471244 598380
rect 457864 598340 457870 598352
rect 471238 598340 471244 598352
rect 471296 598340 471302 598392
rect 459094 598272 459100 598324
rect 459152 598312 459158 598324
rect 502334 598312 502340 598324
rect 459152 598284 502340 598312
rect 459152 598272 459158 598284
rect 502334 598272 502340 598284
rect 502392 598272 502398 598324
rect 460290 598204 460296 598256
rect 460348 598244 460354 598256
rect 495434 598244 495440 598256
rect 460348 598216 495440 598244
rect 460348 598204 460354 598216
rect 495434 598204 495440 598216
rect 495492 598204 495498 598256
rect 496078 598204 496084 598256
rect 496136 598244 496142 598256
rect 540514 598244 540520 598256
rect 496136 598216 540520 598244
rect 496136 598204 496142 598216
rect 540514 598204 540520 598216
rect 540572 598204 540578 598256
rect 382274 597524 382280 597576
rect 382332 597564 382338 597576
rect 406378 597564 406384 597576
rect 382332 597536 406384 597564
rect 382332 597524 382338 597536
rect 406378 597524 406384 597536
rect 406436 597524 406442 597576
rect 457622 596844 457628 596896
rect 457680 596884 457686 596896
rect 467190 596884 467196 596896
rect 457680 596856 467196 596884
rect 457680 596844 457686 596856
rect 467190 596844 467196 596856
rect 467248 596844 467254 596896
rect 459002 596776 459008 596828
rect 459060 596816 459066 596828
rect 496814 596816 496820 596828
rect 459060 596788 496820 596816
rect 459060 596776 459066 596788
rect 496814 596776 496820 596788
rect 496872 596776 496878 596828
rect 457714 595484 457720 595536
rect 457772 595524 457778 595536
rect 468570 595524 468576 595536
rect 457772 595496 468576 595524
rect 457772 595484 457778 595496
rect 468570 595484 468576 595496
rect 468628 595484 468634 595536
rect 460474 595416 460480 595468
rect 460532 595456 460538 595468
rect 500954 595456 500960 595468
rect 460532 595428 500960 595456
rect 460532 595416 460538 595428
rect 500954 595416 500960 595428
rect 501012 595416 501018 595468
rect 458910 592628 458916 592680
rect 458968 592668 458974 592680
rect 494054 592668 494060 592680
rect 458968 592640 494060 592668
rect 458968 592628 458974 592640
rect 494054 592628 494060 592640
rect 494112 592628 494118 592680
rect 459278 591268 459284 591320
rect 459336 591308 459342 591320
rect 503806 591308 503812 591320
rect 459336 591280 503812 591308
rect 459336 591268 459342 591280
rect 503806 591268 503812 591280
rect 503864 591268 503870 591320
rect 459186 589908 459192 589960
rect 459244 589948 459250 589960
rect 499574 589948 499580 589960
rect 459244 589920 499580 589948
rect 459244 589908 459250 589920
rect 499574 589908 499580 589920
rect 499632 589908 499638 589960
rect 6178 587908 6184 587920
rect 4172 587880 6184 587908
rect 3786 587800 3792 587852
rect 3844 587840 3850 587852
rect 4172 587840 4200 587880
rect 6178 587868 6184 587880
rect 6236 587868 6242 587920
rect 382274 587868 382280 587920
rect 382332 587908 382338 587920
rect 392578 587908 392584 587920
rect 382332 587880 392584 587908
rect 382332 587868 382338 587880
rect 392578 587868 392584 587880
rect 392636 587868 392642 587920
rect 3844 587812 4200 587840
rect 3844 587800 3850 587812
rect 3602 578416 3608 578468
rect 3660 578456 3666 578468
rect 5166 578456 5172 578468
rect 3660 578428 5172 578456
rect 3660 578416 3666 578428
rect 5166 578416 5172 578428
rect 5224 578416 5230 578468
rect 382274 576852 382280 576904
rect 382332 576892 382338 576904
rect 419074 576892 419080 576904
rect 382332 576864 419080 576892
rect 382332 576852 382338 576864
rect 419074 576852 419080 576864
rect 419132 576852 419138 576904
rect 518250 576852 518256 576904
rect 518308 576892 518314 576904
rect 579614 576892 579620 576904
rect 518308 576864 579620 576892
rect 518308 576852 518314 576864
rect 579614 576852 579620 576864
rect 579672 576852 579678 576904
rect 381906 573996 381912 574048
rect 381964 574036 381970 574048
rect 384298 574036 384304 574048
rect 381964 574008 384304 574036
rect 381964 573996 381970 574008
rect 384298 573996 384304 574008
rect 384356 573996 384362 574048
rect 381814 572160 381820 572212
rect 381872 572200 381878 572212
rect 383010 572200 383016 572212
rect 381872 572172 383016 572200
rect 381872 572160 381878 572172
rect 383010 572160 383016 572172
rect 383068 572160 383074 572212
rect 3878 565836 3884 565888
rect 3936 565876 3942 565888
rect 5074 565876 5080 565888
rect 3936 565848 5080 565876
rect 3936 565836 3942 565848
rect 5074 565836 5080 565848
rect 5132 565836 5138 565888
rect 382274 565088 382280 565140
rect 382332 565128 382338 565140
rect 407758 565128 407764 565140
rect 382332 565100 407764 565128
rect 382332 565088 382338 565100
rect 407758 565088 407764 565100
rect 407816 565088 407822 565140
rect 515490 563048 515496 563100
rect 515548 563088 515554 563100
rect 580166 563088 580172 563100
rect 515548 563060 580172 563088
rect 515548 563048 515554 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 383010 559512 383016 559564
rect 383068 559552 383074 559564
rect 387610 559552 387616 559564
rect 383068 559524 387616 559552
rect 383068 559512 383074 559524
rect 387610 559512 387616 559524
rect 387668 559512 387674 559564
rect 384298 556588 384304 556640
rect 384356 556628 384362 556640
rect 385034 556628 385040 556640
rect 384356 556600 385040 556628
rect 384356 556588 384362 556600
rect 385034 556588 385040 556600
rect 385092 556588 385098 556640
rect 382274 556180 382280 556232
rect 382332 556220 382338 556232
rect 391198 556220 391204 556232
rect 382332 556192 391204 556220
rect 382332 556180 382338 556192
rect 391198 556180 391204 556192
rect 391256 556180 391262 556232
rect 385034 554344 385040 554396
rect 385092 554384 385098 554396
rect 387150 554384 387156 554396
rect 385092 554356 387156 554384
rect 385092 554344 385098 554356
rect 387150 554344 387156 554356
rect 387208 554344 387214 554396
rect 3786 553392 3792 553444
rect 3844 553432 3850 553444
rect 4982 553432 4988 553444
rect 3844 553404 4988 553432
rect 3844 553392 3850 553404
rect 4982 553392 4988 553404
rect 5040 553392 5046 553444
rect 380618 553392 380624 553444
rect 380676 553432 380682 553444
rect 380676 553404 380940 553432
rect 380676 553392 380682 553404
rect 380912 553364 380940 553404
rect 383010 553364 383016 553376
rect 380912 553336 383016 553364
rect 383010 553324 383016 553336
rect 383068 553324 383074 553376
rect 387610 552644 387616 552696
rect 387668 552684 387674 552696
rect 389910 552684 389916 552696
rect 387668 552656 389916 552684
rect 387668 552644 387674 552656
rect 389910 552644 389916 552656
rect 389968 552644 389974 552696
rect 382274 545096 382280 545148
rect 382332 545136 382338 545148
rect 389818 545136 389824 545148
rect 382332 545108 389824 545136
rect 382332 545096 382338 545108
rect 389818 545096 389824 545108
rect 389876 545096 389882 545148
rect 389910 543668 389916 543720
rect 389968 543708 389974 543720
rect 394050 543708 394056 543720
rect 389968 543680 394056 543708
rect 389968 543668 389974 543680
rect 394050 543668 394056 543680
rect 394108 543668 394114 543720
rect 380526 543192 380532 543244
rect 380584 543232 380590 543244
rect 381814 543232 381820 543244
rect 380584 543204 381820 543232
rect 380584 543192 380590 543204
rect 381814 543192 381820 543204
rect 381872 543192 381878 543244
rect 381722 537480 381728 537532
rect 381780 537520 381786 537532
rect 389174 537520 389180 537532
rect 381780 537492 389180 537520
rect 381780 537480 381786 537492
rect 389174 537480 389180 537492
rect 389232 537480 389238 537532
rect 460658 537480 460664 537532
rect 460716 537520 460722 537532
rect 498194 537520 498200 537532
rect 460716 537492 498200 537520
rect 460716 537480 460722 537492
rect 498194 537480 498200 537492
rect 498252 537480 498258 537532
rect 518342 536800 518348 536852
rect 518400 536840 518406 536852
rect 580166 536840 580172 536852
rect 518400 536812 580172 536840
rect 518400 536800 518406 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 383010 536596 383016 536648
rect 383068 536636 383074 536648
rect 384114 536636 384120 536648
rect 383068 536608 384120 536636
rect 383068 536596 383074 536608
rect 384114 536596 384120 536608
rect 384172 536596 384178 536648
rect 389174 535780 389180 535832
rect 389232 535820 389238 535832
rect 391934 535820 391940 535832
rect 389232 535792 391940 535820
rect 389232 535780 389238 535792
rect 391934 535780 391940 535792
rect 391992 535780 391998 535832
rect 382274 534080 382280 534132
rect 382332 534120 382338 534132
rect 387058 534120 387064 534132
rect 382332 534092 387064 534120
rect 382332 534080 382338 534092
rect 387058 534080 387064 534092
rect 387116 534080 387122 534132
rect 391934 534012 391940 534064
rect 391992 534052 391998 534064
rect 394878 534052 394884 534064
rect 391992 534024 394884 534052
rect 391992 534012 391998 534024
rect 394878 534012 394884 534024
rect 394936 534012 394942 534064
rect 381814 533536 381820 533588
rect 381872 533576 381878 533588
rect 383010 533576 383016 533588
rect 381872 533548 383016 533576
rect 381872 533536 381878 533548
rect 383010 533536 383016 533548
rect 383068 533536 383074 533588
rect 384114 532720 384120 532772
rect 384172 532760 384178 532772
rect 384172 532732 385080 532760
rect 384172 532720 384178 532732
rect 385052 532692 385080 532732
rect 389174 532692 389180 532704
rect 385052 532664 389180 532692
rect 389174 532652 389180 532664
rect 389232 532652 389238 532704
rect 394050 531224 394056 531276
rect 394108 531264 394114 531276
rect 396810 531264 396816 531276
rect 394108 531236 396816 531264
rect 394108 531224 394114 531236
rect 396810 531224 396816 531236
rect 396868 531224 396874 531276
rect 389174 529932 389180 529984
rect 389232 529972 389238 529984
rect 389232 529944 390600 529972
rect 389232 529932 389238 529944
rect 390572 529904 390600 529944
rect 394050 529904 394056 529916
rect 390572 529876 394056 529904
rect 394050 529864 394056 529876
rect 394108 529864 394114 529916
rect 394878 529864 394884 529916
rect 394936 529904 394942 529916
rect 397086 529904 397092 529916
rect 394936 529876 397092 529904
rect 394936 529864 394942 529876
rect 397086 529864 397092 529876
rect 397144 529864 397150 529916
rect 381630 529524 381636 529576
rect 381688 529564 381694 529576
rect 385770 529564 385776 529576
rect 381688 529536 385776 529564
rect 381688 529524 381694 529536
rect 385770 529524 385776 529536
rect 385828 529524 385834 529576
rect 3510 525784 3516 525836
rect 3568 525824 3574 525836
rect 4890 525824 4896 525836
rect 3568 525796 4896 525824
rect 3568 525784 3574 525796
rect 4890 525784 4896 525796
rect 4948 525784 4954 525836
rect 382274 524424 382280 524476
rect 382332 524464 382338 524476
rect 385678 524464 385684 524476
rect 382332 524436 385684 524464
rect 382332 524424 382338 524436
rect 385678 524424 385684 524436
rect 385736 524424 385742 524476
rect 458082 522248 458088 522300
rect 458140 522288 458146 522300
rect 467282 522288 467288 522300
rect 458140 522260 467288 522288
rect 458140 522248 458146 522260
rect 467282 522248 467288 522260
rect 467340 522248 467346 522300
rect 397454 521568 397460 521620
rect 397512 521608 397518 521620
rect 402238 521608 402244 521620
rect 397512 521580 402244 521608
rect 397512 521568 397518 521580
rect 402238 521568 402244 521580
rect 402296 521568 402302 521620
rect 482922 520888 482928 520940
rect 482980 520928 482986 520940
rect 531314 520928 531320 520940
rect 482980 520900 531320 520928
rect 482980 520888 482986 520900
rect 531314 520888 531320 520900
rect 531372 520888 531378 520940
rect 461670 520276 461676 520328
rect 461728 520316 461734 520328
rect 488626 520316 488632 520328
rect 461728 520288 488632 520316
rect 461728 520276 461734 520288
rect 488626 520276 488632 520288
rect 488684 520276 488690 520328
rect 460750 519528 460756 519580
rect 460808 519568 460814 519580
rect 493042 519568 493048 519580
rect 460808 519540 493048 519568
rect 460808 519528 460814 519540
rect 493042 519528 493048 519540
rect 493100 519528 493106 519580
rect 457990 518168 457996 518220
rect 458048 518208 458054 518220
rect 469858 518208 469864 518220
rect 458048 518180 469864 518208
rect 458048 518168 458054 518180
rect 469858 518168 469864 518180
rect 469916 518168 469922 518220
rect 387150 518032 387156 518084
rect 387208 518072 387214 518084
rect 391934 518072 391940 518084
rect 387208 518044 391940 518072
rect 387208 518032 387214 518044
rect 391934 518032 391940 518044
rect 391992 518032 391998 518084
rect 394050 517964 394056 518016
rect 394108 518004 394114 518016
rect 394694 518004 394700 518016
rect 394108 517976 394700 518004
rect 394108 517964 394114 517976
rect 394694 517964 394700 517976
rect 394752 517964 394758 518016
rect 450354 517556 450360 517608
rect 450412 517596 450418 517608
rect 491846 517596 491852 517608
rect 450412 517568 491852 517596
rect 450412 517556 450418 517568
rect 491846 517556 491852 517568
rect 491904 517556 491910 517608
rect 450538 517488 450544 517540
rect 450596 517528 450602 517540
rect 514754 517528 514760 517540
rect 450596 517500 514760 517528
rect 450596 517488 450602 517500
rect 514754 517488 514760 517500
rect 514812 517488 514818 517540
rect 489178 517420 489184 517472
rect 489236 517420 489242 517472
rect 450170 516808 450176 516860
rect 450228 516848 450234 516860
rect 480438 516848 480444 516860
rect 450228 516820 480444 516848
rect 450228 516808 450234 516820
rect 480438 516808 480444 516820
rect 480496 516808 480502 516860
rect 450630 516740 450636 516792
rect 450688 516780 450694 516792
rect 489196 516780 489224 517420
rect 494146 516780 494152 516792
rect 450688 516752 494152 516780
rect 450688 516740 450694 516752
rect 494146 516740 494152 516752
rect 494204 516740 494210 516792
rect 383010 516060 383016 516112
rect 383068 516100 383074 516112
rect 384942 516100 384948 516112
rect 383068 516072 384948 516100
rect 383068 516060 383074 516072
rect 384942 516060 384948 516072
rect 385000 516060 385006 516112
rect 391934 516060 391940 516112
rect 391992 516100 391998 516112
rect 395062 516100 395068 516112
rect 391992 516072 395068 516100
rect 391992 516060 391998 516072
rect 395062 516060 395068 516072
rect 395120 516060 395126 516112
rect 494790 515924 494796 515976
rect 494848 515964 494854 515976
rect 498286 515964 498292 515976
rect 494848 515936 498292 515964
rect 494848 515924 494854 515936
rect 498286 515924 498292 515936
rect 498344 515924 498350 515976
rect 396810 514768 396816 514820
rect 396868 514808 396874 514820
rect 396868 514780 398880 514808
rect 396868 514768 396874 514780
rect 398852 514740 398880 514780
rect 400214 514740 400220 514752
rect 398852 514712 400220 514740
rect 400214 514700 400220 514712
rect 400272 514700 400278 514752
rect 514754 514020 514760 514072
rect 514812 514060 514818 514072
rect 547874 514060 547880 514072
rect 514812 514032 547880 514060
rect 514812 514020 514818 514032
rect 547874 514020 547880 514032
rect 547932 514020 547938 514072
rect 382274 513544 382280 513596
rect 382332 513584 382338 513596
rect 384298 513584 384304 513596
rect 382332 513556 384304 513584
rect 382332 513544 382338 513556
rect 384298 513544 384304 513556
rect 384356 513544 384362 513596
rect 395062 513340 395068 513392
rect 395120 513380 395126 513392
rect 399570 513380 399576 513392
rect 395120 513352 399576 513380
rect 395120 513340 395126 513352
rect 399570 513340 399576 513352
rect 399628 513340 399634 513392
rect 506566 512660 506572 512712
rect 506624 512700 506630 512712
rect 543734 512700 543740 512712
rect 506624 512672 543740 512700
rect 506624 512660 506630 512672
rect 543734 512660 543740 512672
rect 543792 512660 543798 512712
rect 494146 512592 494152 512644
rect 494204 512632 494210 512644
rect 538214 512632 538220 512644
rect 494204 512604 538220 512632
rect 494204 512592 494210 512604
rect 538214 512592 538220 512604
rect 538272 512592 538278 512644
rect 519538 510620 519544 510672
rect 519596 510660 519602 510672
rect 580166 510660 580172 510672
rect 519596 510632 580172 510660
rect 519596 510620 519602 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 385770 510552 385776 510604
rect 385828 510592 385834 510604
rect 387150 510592 387156 510604
rect 385828 510564 387156 510592
rect 385828 510552 385834 510564
rect 387150 510552 387156 510564
rect 387208 510552 387214 510604
rect 394694 510552 394700 510604
rect 394752 510592 394758 510604
rect 397178 510592 397184 510604
rect 394752 510564 397184 510592
rect 394752 510552 394758 510564
rect 397178 510552 397184 510564
rect 397236 510552 397242 510604
rect 400214 510552 400220 510604
rect 400272 510592 400278 510604
rect 402146 510592 402152 510604
rect 400272 510564 402152 510592
rect 400272 510552 400278 510564
rect 402146 510552 402152 510564
rect 402204 510552 402210 510604
rect 385034 510484 385040 510536
rect 385092 510524 385098 510536
rect 388070 510524 388076 510536
rect 385092 510496 388076 510524
rect 385092 510484 385098 510496
rect 388070 510484 388076 510496
rect 388128 510484 388134 510536
rect 498286 509872 498292 509924
rect 498344 509912 498350 509924
rect 540974 509912 540980 509924
rect 498344 509884 540980 509912
rect 498344 509872 498350 509884
rect 540974 509872 540980 509884
rect 541032 509872 541038 509924
rect 397178 509192 397184 509244
rect 397236 509232 397242 509244
rect 403986 509232 403992 509244
rect 397236 509204 403992 509232
rect 397236 509192 397242 509204
rect 403986 509192 403992 509204
rect 404044 509192 404050 509244
rect 492122 508512 492128 508564
rect 492180 508552 492186 508564
rect 534074 508552 534080 508564
rect 492180 508524 534080 508552
rect 492180 508512 492186 508524
rect 534074 508512 534080 508524
rect 534132 508512 534138 508564
rect 3694 507832 3700 507884
rect 3752 507872 3758 507884
rect 4798 507872 4804 507884
rect 3752 507844 4804 507872
rect 3752 507832 3758 507844
rect 4798 507832 4804 507844
rect 4856 507832 4862 507884
rect 494146 505112 494152 505164
rect 494204 505152 494210 505164
rect 531314 505152 531320 505164
rect 494204 505124 531320 505152
rect 494204 505112 494210 505124
rect 531314 505112 531320 505124
rect 531372 505112 531378 505164
rect 388070 504636 388076 504688
rect 388128 504676 388134 504688
rect 389174 504676 389180 504688
rect 388128 504648 389180 504676
rect 388128 504636 388134 504648
rect 389174 504636 389180 504648
rect 389232 504636 389238 504688
rect 402146 503684 402152 503736
rect 402204 503724 402210 503736
rect 402204 503696 402974 503724
rect 402204 503684 402210 503696
rect 402946 503656 402974 503696
rect 404722 503656 404728 503668
rect 402946 503628 404728 503656
rect 404722 503616 404728 503628
rect 404780 503616 404786 503668
rect 382274 502324 382280 502376
rect 382332 502364 382338 502376
rect 410518 502364 410524 502376
rect 382332 502336 410524 502364
rect 382332 502324 382338 502336
rect 410518 502324 410524 502336
rect 410576 502324 410582 502376
rect 389174 502256 389180 502308
rect 389232 502296 389238 502308
rect 392670 502296 392676 502308
rect 389232 502268 392676 502296
rect 389232 502256 389238 502268
rect 392670 502256 392676 502268
rect 392728 502256 392734 502308
rect 403986 502256 403992 502308
rect 404044 502296 404050 502308
rect 404998 502296 405004 502308
rect 404044 502268 405004 502296
rect 404044 502256 404050 502268
rect 404998 502256 405004 502268
rect 405056 502256 405062 502308
rect 387150 500896 387156 500948
rect 387208 500936 387214 500948
rect 389910 500936 389916 500948
rect 387208 500908 389916 500936
rect 387208 500896 387214 500908
rect 389910 500896 389916 500908
rect 389968 500896 389974 500948
rect 404722 500896 404728 500948
rect 404780 500936 404786 500948
rect 406562 500936 406568 500948
rect 404780 500908 406568 500936
rect 404780 500896 404786 500908
rect 406562 500896 406568 500908
rect 406620 500896 406626 500948
rect 450538 500896 450544 500948
rect 450596 500936 450602 500948
rect 472618 500936 472624 500948
rect 450596 500908 472624 500936
rect 450596 500896 450602 500908
rect 472618 500896 472624 500908
rect 472676 500936 472682 500948
rect 494146 500936 494152 500948
rect 472676 500908 494152 500936
rect 472676 500896 472682 500908
rect 494146 500896 494152 500908
rect 494204 500896 494210 500948
rect 464430 497564 464436 497616
rect 464488 497604 464494 497616
rect 485038 497604 485044 497616
rect 464488 497576 485044 497604
rect 464488 497564 464494 497576
rect 485038 497564 485044 497576
rect 485096 497564 485102 497616
rect 454678 497496 454684 497548
rect 454736 497536 454742 497548
rect 486234 497536 486240 497548
rect 454736 497508 486240 497536
rect 454736 497496 454742 497508
rect 486234 497496 486240 497508
rect 486292 497496 486298 497548
rect 453298 497428 453304 497480
rect 453356 497468 453362 497480
rect 489914 497468 489920 497480
rect 453356 497440 489920 497468
rect 453356 497428 453362 497440
rect 489914 497428 489920 497440
rect 489972 497428 489978 497480
rect 399570 497156 399576 497208
rect 399628 497196 399634 497208
rect 400858 497196 400864 497208
rect 399628 497168 400864 497196
rect 399628 497156 399634 497168
rect 400858 497156 400864 497168
rect 400916 497156 400922 497208
rect 461394 494708 461400 494760
rect 461452 494748 461458 494760
rect 461762 494748 461768 494760
rect 461452 494720 461768 494748
rect 461452 494708 461458 494720
rect 461762 494708 461768 494720
rect 461820 494708 461826 494760
rect 382274 492668 382280 492720
rect 382332 492708 382338 492720
rect 411898 492708 411904 492720
rect 382332 492680 411904 492708
rect 382332 492668 382338 492680
rect 411898 492668 411904 492680
rect 411956 492668 411962 492720
rect 404998 492600 405004 492652
rect 405056 492640 405062 492652
rect 406746 492640 406752 492652
rect 405056 492612 406752 492640
rect 405056 492600 405062 492612
rect 406746 492600 406752 492612
rect 406804 492600 406810 492652
rect 481634 490424 481640 490476
rect 481692 490464 481698 490476
rect 482646 490464 482652 490476
rect 481692 490436 482652 490464
rect 481692 490424 481698 490436
rect 482646 490424 482652 490436
rect 482704 490424 482710 490476
rect 380434 489880 380440 489932
rect 380492 489920 380498 489932
rect 380492 489892 380940 489920
rect 380492 489880 380498 489892
rect 380912 489852 380940 489892
rect 383010 489852 383016 489864
rect 380912 489824 383016 489852
rect 383010 489812 383016 489824
rect 383068 489812 383074 489864
rect 392670 488860 392676 488912
rect 392728 488900 392734 488912
rect 395614 488900 395620 488912
rect 392728 488872 395620 488900
rect 392728 488860 392734 488872
rect 395614 488860 395620 488872
rect 395672 488860 395678 488912
rect 395614 485596 395620 485648
rect 395672 485636 395678 485648
rect 400214 485636 400220 485648
rect 395672 485608 400220 485636
rect 395672 485596 395678 485608
rect 400214 485596 400220 485608
rect 400272 485596 400278 485648
rect 400858 485052 400864 485104
rect 400916 485092 400922 485104
rect 406654 485092 406660 485104
rect 400916 485064 406660 485092
rect 400916 485052 400922 485064
rect 406654 485052 406660 485064
rect 406712 485052 406718 485104
rect 402238 484304 402244 484356
rect 402296 484344 402302 484356
rect 403710 484344 403716 484356
rect 402296 484316 403716 484344
rect 402296 484304 402302 484316
rect 403710 484304 403716 484316
rect 403768 484304 403774 484356
rect 406746 484304 406752 484356
rect 406804 484344 406810 484356
rect 407850 484344 407856 484356
rect 406804 484316 407856 484344
rect 406804 484304 406810 484316
rect 407850 484304 407856 484316
rect 407908 484304 407914 484356
rect 382274 481652 382280 481704
rect 382332 481692 382338 481704
rect 414658 481692 414664 481704
rect 382332 481664 414664 481692
rect 382332 481652 382338 481664
rect 414658 481652 414664 481664
rect 414716 481652 414722 481704
rect 400214 480224 400220 480276
rect 400272 480264 400278 480276
rect 400272 480236 401640 480264
rect 400272 480224 400278 480236
rect 401612 480196 401640 480236
rect 403894 480196 403900 480208
rect 401612 480168 403900 480196
rect 403894 480156 403900 480168
rect 403952 480156 403958 480208
rect 380342 478796 380348 478848
rect 380400 478836 380406 478848
rect 381354 478836 381360 478848
rect 380400 478808 381360 478836
rect 380400 478796 380406 478808
rect 381354 478796 381360 478808
rect 381412 478796 381418 478848
rect 389910 477504 389916 477556
rect 389968 477544 389974 477556
rect 389968 477516 393314 477544
rect 389968 477504 389974 477516
rect 393286 477476 393314 477516
rect 394602 477476 394608 477488
rect 393286 477448 394608 477476
rect 394602 477436 394608 477448
rect 394660 477436 394666 477488
rect 403894 476076 403900 476128
rect 403952 476116 403958 476128
rect 403952 476088 404400 476116
rect 403952 476076 403958 476088
rect 404372 476048 404400 476088
rect 406470 476048 406476 476060
rect 404372 476020 406476 476048
rect 406470 476008 406476 476020
rect 406528 476008 406534 476060
rect 380250 473356 380256 473408
rect 380308 473396 380314 473408
rect 380308 473368 380940 473396
rect 380308 473356 380314 473368
rect 380912 473328 380940 473368
rect 394694 473356 394700 473408
rect 394752 473396 394758 473408
rect 394752 473368 398880 473396
rect 394752 473356 394758 473368
rect 382274 473328 382280 473340
rect 380912 473300 382280 473328
rect 382274 473288 382280 473300
rect 382332 473288 382338 473340
rect 398852 473328 398880 473368
rect 401502 473328 401508 473340
rect 398852 473300 401508 473328
rect 401502 473288 401508 473300
rect 401560 473288 401566 473340
rect 381354 470568 381360 470620
rect 381412 470608 381418 470620
rect 381412 470580 382320 470608
rect 381412 470568 381418 470580
rect 382292 470540 382320 470580
rect 382366 470568 382372 470620
rect 382424 470608 382430 470620
rect 419166 470608 419172 470620
rect 382424 470580 419172 470608
rect 382424 470568 382430 470580
rect 419166 470568 419172 470580
rect 419224 470568 419230 470620
rect 514018 470568 514024 470620
rect 514076 470608 514082 470620
rect 579982 470608 579988 470620
rect 514076 470580 579988 470608
rect 514076 470568 514082 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 384758 470540 384764 470552
rect 382292 470512 384764 470540
rect 384758 470500 384764 470512
rect 384816 470500 384822 470552
rect 382274 469208 382280 469260
rect 382332 469248 382338 469260
rect 382332 469220 383654 469248
rect 382332 469208 382338 469220
rect 383626 469180 383654 469220
rect 385034 469180 385040 469192
rect 383626 469152 385040 469180
rect 385034 469140 385040 469152
rect 385092 469140 385098 469192
rect 384758 468120 384764 468172
rect 384816 468160 384822 468172
rect 387150 468160 387156 468172
rect 384816 468132 387156 468160
rect 384816 468120 384822 468132
rect 387150 468120 387156 468132
rect 387208 468120 387214 468172
rect 401594 467780 401600 467832
rect 401652 467820 401658 467832
rect 403802 467820 403808 467832
rect 401652 467792 403808 467820
rect 401652 467780 401658 467792
rect 403802 467780 403808 467792
rect 403860 467780 403866 467832
rect 494790 466488 494796 466540
rect 494848 466528 494854 466540
rect 528370 466528 528376 466540
rect 494848 466500 528376 466528
rect 494848 466488 494854 466500
rect 528370 466488 528376 466500
rect 528428 466488 528434 466540
rect 385034 466420 385040 466472
rect 385092 466460 385098 466472
rect 385092 466432 386460 466460
rect 385092 466420 385098 466432
rect 386432 466392 386460 466432
rect 406562 466420 406568 466472
rect 406620 466460 406626 466472
rect 406620 466432 407160 466460
rect 406620 466420 406626 466432
rect 388162 466392 388168 466404
rect 386432 466364 388168 466392
rect 388162 466352 388168 466364
rect 388220 466352 388226 466404
rect 407132 466392 407160 466432
rect 454770 466420 454776 466472
rect 454828 466460 454834 466472
rect 525058 466460 525064 466472
rect 454828 466432 525064 466460
rect 454828 466420 454834 466432
rect 525058 466420 525064 466432
rect 525116 466420 525122 466472
rect 408494 466392 408500 466404
rect 407132 466364 408500 466392
rect 408494 466352 408500 466364
rect 408552 466352 408558 466404
rect 511258 465672 511264 465724
rect 511316 465712 511322 465724
rect 580258 465712 580264 465724
rect 511316 465684 580264 465712
rect 511316 465672 511322 465684
rect 580258 465672 580264 465684
rect 580316 465672 580322 465724
rect 464522 465128 464528 465180
rect 464580 465168 464586 465180
rect 554866 465168 554872 465180
rect 464580 465140 554872 465168
rect 464580 465128 464586 465140
rect 554866 465128 554872 465140
rect 554924 465128 554930 465180
rect 458818 465060 458824 465112
rect 458876 465100 458882 465112
rect 558178 465100 558184 465112
rect 458876 465072 558184 465100
rect 458876 465060 458882 465072
rect 558178 465060 558184 465072
rect 558236 465060 558242 465112
rect 406654 464992 406660 465044
rect 406712 465032 406718 465044
rect 407942 465032 407948 465044
rect 406712 465004 407948 465032
rect 406712 464992 406718 465004
rect 407942 464992 407948 465004
rect 408000 464992 408006 465044
rect 388162 463700 388168 463752
rect 388220 463740 388226 463752
rect 388220 463712 389220 463740
rect 388220 463700 388226 463712
rect 389192 463672 389220 463712
rect 408494 463700 408500 463752
rect 408552 463740 408558 463752
rect 408552 463712 409920 463740
rect 408552 463700 408558 463712
rect 391934 463672 391940 463684
rect 389192 463644 391940 463672
rect 391934 463632 391940 463644
rect 391992 463632 391998 463684
rect 407850 463632 407856 463684
rect 407908 463672 407914 463684
rect 409322 463672 409328 463684
rect 407908 463644 409328 463672
rect 407908 463632 407914 463644
rect 409322 463632 409328 463644
rect 409380 463632 409386 463684
rect 409892 463672 409920 463712
rect 412082 463672 412088 463684
rect 409892 463644 412088 463672
rect 412082 463632 412088 463644
rect 412140 463632 412146 463684
rect 391934 461592 391940 461644
rect 391992 461632 391998 461644
rect 400766 461632 400772 461644
rect 391992 461604 400772 461632
rect 391992 461592 391998 461604
rect 400766 461592 400772 461604
rect 400824 461592 400830 461644
rect 449066 461592 449072 461644
rect 449124 461632 449130 461644
rect 487154 461632 487160 461644
rect 449124 461604 487160 461632
rect 449124 461592 449130 461604
rect 487154 461592 487160 461604
rect 487212 461592 487218 461644
rect 383010 460844 383016 460896
rect 383068 460884 383074 460896
rect 384574 460884 384580 460896
rect 383068 460856 384580 460884
rect 383068 460844 383074 460856
rect 384574 460844 384580 460856
rect 384632 460844 384638 460896
rect 400766 460232 400772 460284
rect 400824 460272 400830 460284
rect 404262 460272 404268 460284
rect 400824 460244 404268 460272
rect 400824 460232 400830 460244
rect 404262 460232 404268 460244
rect 404320 460232 404326 460284
rect 449618 460164 449624 460216
rect 449676 460204 449682 460216
rect 488534 460204 488540 460216
rect 449676 460176 488540 460204
rect 449676 460164 449682 460176
rect 488534 460164 488540 460176
rect 488592 460164 488598 460216
rect 382274 459552 382280 459604
rect 382332 459592 382338 459604
rect 400858 459592 400864 459604
rect 382332 459564 400864 459592
rect 382332 459552 382338 459564
rect 400858 459552 400864 459564
rect 400916 459552 400922 459604
rect 404262 458464 404268 458516
rect 404320 458504 404326 458516
rect 405918 458504 405924 458516
rect 404320 458476 405924 458504
rect 404320 458464 404326 458476
rect 405918 458464 405924 458476
rect 405976 458464 405982 458516
rect 468662 458328 468668 458380
rect 468720 458368 468726 458380
rect 473998 458368 474004 458380
rect 468720 458340 474004 458368
rect 468720 458328 468726 458340
rect 473998 458328 474004 458340
rect 474056 458368 474062 458380
rect 478138 458368 478144 458380
rect 474056 458340 478144 458368
rect 474056 458328 474062 458340
rect 478138 458328 478144 458340
rect 478196 458328 478202 458380
rect 456058 458260 456064 458312
rect 456116 458300 456122 458312
rect 482002 458300 482008 458312
rect 456116 458272 482008 458300
rect 456116 458260 456122 458272
rect 482002 458260 482008 458272
rect 482060 458260 482066 458312
rect 384574 458192 384580 458244
rect 384632 458232 384638 458244
rect 384632 458204 385080 458232
rect 384632 458192 384638 458204
rect 385052 458164 385080 458204
rect 403710 458192 403716 458244
rect 403768 458232 403774 458244
rect 403768 458204 404400 458232
rect 403768 458192 403774 458204
rect 387702 458164 387708 458176
rect 385052 458136 387708 458164
rect 387702 458124 387708 458136
rect 387760 458124 387766 458176
rect 404372 458164 404400 458204
rect 409322 458192 409328 458244
rect 409380 458232 409386 458244
rect 410610 458232 410616 458244
rect 409380 458204 410616 458232
rect 409380 458192 409386 458204
rect 410610 458192 410616 458204
rect 410668 458192 410674 458244
rect 457438 458192 457444 458244
rect 457496 458232 457502 458244
rect 490006 458232 490012 458244
rect 457496 458204 490012 458232
rect 457496 458192 457502 458204
rect 490006 458192 490012 458204
rect 490064 458232 490070 458244
rect 494790 458232 494796 458244
rect 490064 458204 494796 458232
rect 490064 458192 490070 458204
rect 494790 458192 494796 458204
rect 494848 458192 494854 458244
rect 407850 458164 407856 458176
rect 404372 458136 407856 458164
rect 407850 458124 407856 458136
rect 407908 458124 407914 458176
rect 449710 457512 449716 457564
rect 449768 457552 449774 457564
rect 481726 457552 481732 457564
rect 449768 457524 481732 457552
rect 449768 457512 449774 457524
rect 481726 457512 481732 457524
rect 481784 457512 481790 457564
rect 449526 457444 449532 457496
rect 449584 457484 449590 457496
rect 481634 457484 481640 457496
rect 449584 457456 481640 457484
rect 449584 457444 449590 457456
rect 481634 457444 481640 457456
rect 481692 457444 481698 457496
rect 405918 456764 405924 456816
rect 405976 456804 405982 456816
rect 405976 456776 407160 456804
rect 405976 456764 405982 456776
rect 407132 456736 407160 456776
rect 570690 456764 570696 456816
rect 570748 456804 570754 456816
rect 580166 456804 580172 456816
rect 570748 456776 580172 456804
rect 570748 456764 570754 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 410794 456736 410800 456748
rect 407132 456708 410800 456736
rect 410794 456696 410800 456708
rect 410852 456696 410858 456748
rect 449434 456152 449440 456204
rect 449492 456192 449498 456204
rect 480254 456192 480260 456204
rect 449492 456164 480260 456192
rect 449492 456152 449498 456164
rect 480254 456152 480260 456164
rect 480312 456152 480318 456204
rect 407850 456084 407856 456136
rect 407908 456124 407914 456136
rect 411990 456124 411996 456136
rect 407908 456096 411996 456124
rect 407908 456084 407914 456096
rect 411990 456084 411996 456096
rect 412048 456084 412054 456136
rect 449342 456084 449348 456136
rect 449400 456124 449406 456136
rect 483106 456124 483112 456136
rect 449400 456096 483112 456124
rect 449400 456084 449406 456096
rect 483106 456084 483112 456096
rect 483164 456084 483170 456136
rect 449250 456016 449256 456068
rect 449308 456056 449314 456068
rect 491294 456056 491300 456068
rect 449308 456028 491300 456056
rect 449308 456016 449314 456028
rect 491294 456016 491300 456028
rect 491352 456016 491358 456068
rect 403802 453976 403808 454028
rect 403860 454016 403866 454028
rect 406562 454016 406568 454028
rect 403860 453988 406568 454016
rect 403860 453976 403866 453988
rect 406562 453976 406568 453988
rect 406620 453976 406626 454028
rect 387794 452548 387800 452600
rect 387852 452588 387858 452600
rect 389910 452588 389916 452600
rect 387852 452560 389916 452588
rect 387852 452548 387858 452560
rect 389910 452548 389916 452560
rect 389968 452548 389974 452600
rect 382274 449896 382280 449948
rect 382332 449936 382338 449948
rect 399570 449936 399576 449948
rect 382332 449908 399576 449936
rect 382332 449896 382338 449908
rect 399570 449896 399576 449908
rect 399628 449896 399634 449948
rect 387150 449556 387156 449608
rect 387208 449596 387214 449608
rect 390278 449596 390284 449608
rect 387208 449568 390284 449596
rect 387208 449556 387214 449568
rect 390278 449556 390284 449568
rect 390336 449556 390342 449608
rect 389910 448536 389916 448588
rect 389968 448576 389974 448588
rect 391290 448576 391296 448588
rect 389968 448548 391296 448576
rect 389968 448536 389974 448548
rect 391290 448536 391296 448548
rect 391348 448536 391354 448588
rect 407942 448536 407948 448588
rect 408000 448576 408006 448588
rect 408000 448548 408540 448576
rect 408000 448536 408006 448548
rect 408512 448508 408540 448548
rect 410702 448508 410708 448520
rect 408512 448480 410708 448508
rect 410702 448468 410708 448480
rect 410760 448468 410766 448520
rect 410794 448468 410800 448520
rect 410852 448508 410858 448520
rect 413462 448508 413468 448520
rect 410852 448480 413468 448508
rect 410852 448468 410858 448480
rect 413462 448468 413468 448480
rect 413520 448468 413526 448520
rect 447870 447924 447876 447976
rect 447928 447964 447934 447976
rect 458818 447964 458824 447976
rect 447928 447936 458824 447964
rect 447928 447924 447934 447936
rect 458818 447924 458824 447936
rect 458876 447924 458882 447976
rect 447134 447856 447140 447908
rect 447192 447896 447198 447908
rect 447778 447896 447784 447908
rect 447192 447868 447784 447896
rect 447192 447856 447198 447868
rect 447778 447856 447784 447868
rect 447836 447896 447842 447908
rect 464522 447896 464528 447908
rect 447836 447868 464528 447896
rect 447836 447856 447842 447868
rect 464522 447856 464528 447868
rect 464580 447856 464586 447908
rect 449894 447788 449900 447840
rect 449952 447828 449958 447840
rect 450630 447828 450636 447840
rect 449952 447800 450636 447828
rect 449952 447788 449958 447800
rect 450630 447788 450636 447800
rect 450688 447828 450694 447840
rect 468662 447828 468668 447840
rect 450688 447800 468668 447828
rect 450688 447788 450694 447800
rect 468662 447788 468668 447800
rect 468720 447788 468726 447840
rect 437382 447312 437388 447364
rect 437440 447352 437446 447364
rect 447870 447352 447876 447364
rect 437440 447324 447876 447352
rect 437440 447312 437446 447324
rect 447870 447312 447876 447324
rect 447928 447352 447934 447364
rect 448238 447352 448244 447364
rect 447928 447324 448244 447352
rect 447928 447312 447934 447324
rect 448238 447312 448244 447324
rect 448296 447312 448302 447364
rect 432414 447244 432420 447296
rect 432472 447284 432478 447296
rect 447134 447284 447140 447296
rect 432472 447256 447140 447284
rect 432472 447244 432478 447256
rect 447134 447244 447140 447256
rect 447192 447244 447198 447296
rect 427446 447176 427452 447228
rect 427504 447216 427510 447228
rect 446214 447216 446220 447228
rect 427504 447188 446220 447216
rect 427504 447176 427510 447188
rect 446214 447176 446220 447188
rect 446272 447176 446278 447228
rect 390278 447108 390284 447160
rect 390336 447148 390342 447160
rect 390336 447120 393314 447148
rect 390336 447108 390342 447120
rect 393286 447080 393314 447120
rect 422478 447108 422484 447160
rect 422536 447148 422542 447160
rect 449894 447148 449900 447160
rect 422536 447120 449900 447148
rect 422536 447108 422542 447120
rect 449894 447108 449900 447120
rect 449952 447108 449958 447160
rect 395154 447080 395160 447092
rect 393286 447052 395160 447080
rect 395154 447040 395160 447052
rect 395212 447040 395218 447092
rect 410610 445680 410616 445732
rect 410668 445720 410674 445732
rect 411254 445720 411260 445732
rect 410668 445692 411260 445720
rect 410668 445680 410674 445692
rect 411254 445680 411260 445692
rect 411312 445680 411318 445732
rect 429838 445000 429844 445052
rect 429896 445040 429902 445052
rect 445478 445040 445484 445052
rect 429896 445012 445484 445040
rect 429896 445000 429902 445012
rect 445478 445000 445484 445012
rect 445536 445000 445542 445052
rect 442626 444388 442632 444440
rect 442684 444428 442690 444440
rect 446306 444428 446312 444440
rect 442684 444400 446312 444428
rect 442684 444388 442690 444400
rect 446306 444388 446312 444400
rect 446364 444388 446370 444440
rect 395154 444320 395160 444372
rect 395212 444360 395218 444372
rect 402238 444360 402244 444372
rect 395212 444332 402244 444360
rect 395212 444320 395218 444332
rect 402238 444320 402244 444332
rect 402296 444320 402302 444372
rect 411990 442960 411996 443012
rect 412048 443000 412054 443012
rect 413370 443000 413376 443012
rect 412048 442972 413376 443000
rect 412048 442960 412054 442972
rect 413370 442960 413376 442972
rect 413428 442960 413434 443012
rect 411254 441804 411260 441856
rect 411312 441844 411318 441856
rect 413554 441844 413560 441856
rect 411312 441816 413560 441844
rect 411312 441804 411318 441816
rect 413554 441804 413560 441816
rect 413612 441804 413618 441856
rect 391290 440240 391296 440292
rect 391348 440280 391354 440292
rect 392670 440280 392676 440292
rect 391348 440252 392676 440280
rect 391348 440240 391354 440252
rect 392670 440240 392676 440252
rect 392728 440240 392734 440292
rect 406470 440240 406476 440292
rect 406528 440280 406534 440292
rect 406528 440252 407160 440280
rect 406528 440240 406534 440252
rect 407132 440212 407160 440252
rect 409138 440212 409144 440224
rect 407132 440184 409144 440212
rect 409138 440172 409144 440184
rect 409196 440172 409202 440224
rect 413462 439356 413468 439408
rect 413520 439396 413526 439408
rect 415854 439396 415860 439408
rect 413520 439368 415860 439396
rect 413520 439356 413526 439368
rect 415854 439356 415860 439368
rect 415912 439356 415918 439408
rect 406562 439084 406568 439136
rect 406620 439124 406626 439136
rect 408678 439124 408684 439136
rect 406620 439096 408684 439124
rect 406620 439084 406626 439096
rect 408678 439084 408684 439096
rect 408736 439084 408742 439136
rect 413554 437724 413560 437776
rect 413612 437764 413618 437776
rect 414750 437764 414756 437776
rect 413612 437736 414756 437764
rect 413612 437724 413618 437736
rect 414750 437724 414756 437736
rect 414808 437724 414814 437776
rect 410702 436908 410708 436960
rect 410760 436948 410766 436960
rect 411990 436948 411996 436960
rect 410760 436920 411996 436948
rect 410760 436908 410766 436920
rect 411990 436908 411996 436920
rect 412048 436908 412054 436960
rect 408678 436772 408684 436824
rect 408736 436812 408742 436824
rect 410610 436812 410616 436824
rect 408736 436784 410616 436812
rect 408736 436772 408742 436784
rect 410610 436772 410616 436784
rect 410668 436772 410674 436824
rect 415854 436704 415860 436756
rect 415912 436744 415918 436756
rect 418154 436744 418160 436756
rect 415912 436716 418160 436744
rect 415912 436704 415918 436716
rect 418154 436704 418160 436716
rect 418212 436704 418218 436756
rect 418154 434664 418160 434716
rect 418212 434704 418218 434716
rect 420270 434704 420276 434716
rect 418212 434676 420276 434704
rect 418212 434664 418218 434676
rect 420270 434664 420276 434676
rect 420328 434664 420334 434716
rect 414750 431060 414756 431112
rect 414808 431100 414814 431112
rect 416682 431100 416688 431112
rect 414808 431072 416688 431100
rect 414808 431060 414814 431072
rect 416682 431060 416688 431072
rect 416740 431060 416746 431112
rect 411990 430584 411996 430636
rect 412048 430624 412054 430636
rect 412048 430596 412634 430624
rect 412048 430584 412054 430596
rect 412606 430556 412634 430596
rect 414750 430556 414756 430568
rect 412606 430528 414756 430556
rect 414750 430516 414756 430528
rect 414808 430516 414814 430568
rect 464982 429972 464988 430024
rect 465040 430012 465046 430024
rect 474642 430012 474648 430024
rect 465040 429984 474648 430012
rect 465040 429972 465046 429984
rect 474642 429972 474648 429984
rect 474700 429972 474706 430024
rect 466270 429904 466276 429956
rect 466328 429944 466334 429956
rect 477586 429944 477592 429956
rect 466328 429916 477592 429944
rect 466328 429904 466334 429916
rect 477586 429904 477592 429916
rect 477644 429904 477650 429956
rect 479518 429904 479524 429956
rect 479576 429944 479582 429956
rect 489362 429944 489368 429956
rect 479576 429916 489368 429944
rect 479576 429904 479582 429916
rect 489362 429904 489368 429916
rect 489420 429904 489426 429956
rect 466362 429836 466368 429888
rect 466420 429876 466426 429888
rect 480530 429876 480536 429888
rect 466420 429848 480536 429876
rect 466420 429836 466426 429848
rect 480530 429836 480536 429848
rect 480588 429836 480594 429888
rect 485038 429156 485044 429208
rect 485096 429196 485102 429208
rect 486418 429196 486424 429208
rect 485096 429168 486424 429196
rect 485096 429156 485102 429168
rect 486418 429156 486424 429168
rect 486476 429156 486482 429208
rect 490558 429156 490564 429208
rect 490616 429196 490622 429208
rect 492306 429196 492312 429208
rect 490616 429168 492312 429196
rect 490616 429156 490622 429168
rect 492306 429156 492312 429168
rect 492364 429156 492370 429208
rect 402238 429088 402244 429140
rect 402296 429128 402302 429140
rect 404906 429128 404912 429140
rect 402296 429100 404912 429128
rect 402296 429088 402302 429100
rect 404906 429088 404912 429100
rect 404964 429088 404970 429140
rect 409138 428476 409144 428528
rect 409196 428516 409202 428528
rect 411990 428516 411996 428528
rect 409196 428488 411996 428516
rect 409196 428476 409202 428488
rect 411990 428476 411996 428488
rect 412048 428476 412054 428528
rect 416774 427524 416780 427576
rect 416832 427564 416838 427576
rect 419350 427564 419356 427576
rect 416832 427536 419356 427564
rect 416832 427524 416838 427536
rect 419350 427524 419356 427536
rect 419408 427524 419414 427576
rect 463602 427048 463608 427100
rect 463660 427088 463666 427100
rect 471698 427088 471704 427100
rect 463660 427060 471704 427088
rect 463660 427048 463666 427060
rect 471698 427048 471704 427060
rect 471756 427048 471762 427100
rect 412082 426368 412088 426420
rect 412140 426408 412146 426420
rect 413922 426408 413928 426420
rect 412140 426380 413928 426408
rect 412140 426368 412146 426380
rect 413922 426368 413928 426380
rect 413980 426368 413986 426420
rect 410610 424328 410616 424380
rect 410668 424368 410674 424380
rect 416682 424368 416688 424380
rect 410668 424340 416688 424368
rect 410668 424328 410674 424340
rect 416682 424328 416688 424340
rect 416740 424328 416746 424380
rect 413922 423648 413928 423700
rect 413980 423688 413986 423700
rect 413980 423660 414060 423688
rect 413980 423648 413986 423660
rect 404906 423580 404912 423632
rect 404964 423620 404970 423632
rect 407022 423620 407028 423632
rect 404964 423592 407028 423620
rect 404964 423580 404970 423592
rect 407022 423580 407028 423592
rect 407080 423580 407086 423632
rect 414032 423620 414060 423660
rect 415946 423620 415952 423632
rect 414032 423592 415952 423620
rect 415946 423580 415952 423592
rect 416004 423580 416010 423632
rect 536098 423376 536104 423428
rect 536156 423416 536162 423428
rect 545850 423416 545856 423428
rect 536156 423388 545856 423416
rect 536156 423376 536162 423388
rect 545850 423376 545856 423388
rect 545908 423376 545914 423428
rect 537478 423308 537484 423360
rect 537536 423348 537542 423360
rect 547322 423348 547328 423360
rect 537536 423320 547328 423348
rect 537536 423308 537542 423320
rect 547322 423308 547328 423320
rect 547380 423308 547386 423360
rect 533338 423240 533344 423292
rect 533396 423280 533402 423292
rect 544378 423280 544384 423292
rect 533396 423252 544384 423280
rect 533396 423240 533402 423252
rect 544378 423240 544384 423252
rect 544436 423240 544442 423292
rect 544470 423240 544476 423292
rect 544528 423280 544534 423292
rect 553210 423280 553216 423292
rect 544528 423252 553216 423280
rect 544528 423240 544534 423252
rect 553210 423240 553216 423252
rect 553268 423240 553274 423292
rect 523678 423172 523684 423224
rect 523736 423212 523742 423224
rect 532602 423212 532608 423224
rect 523736 423184 532608 423212
rect 523736 423172 523742 423184
rect 532602 423172 532608 423184
rect 532660 423172 532666 423224
rect 540238 423172 540244 423224
rect 540296 423212 540302 423224
rect 551738 423212 551744 423224
rect 540296 423184 551744 423212
rect 540296 423172 540302 423184
rect 551738 423172 551744 423184
rect 551796 423172 551802 423224
rect 518434 423104 518440 423156
rect 518492 423144 518498 423156
rect 528186 423144 528192 423156
rect 518492 423116 528192 423144
rect 518492 423104 518498 423116
rect 528186 423104 528192 423116
rect 528244 423104 528250 423156
rect 538858 423104 538864 423156
rect 538916 423144 538922 423156
rect 550266 423144 550272 423156
rect 538916 423116 550272 423144
rect 538916 423104 538922 423116
rect 550266 423104 550272 423116
rect 550324 423104 550330 423156
rect 512638 423036 512644 423088
rect 512696 423076 512702 423088
rect 556154 423076 556160 423088
rect 512696 423048 556160 423076
rect 512696 423036 512702 423048
rect 556154 423036 556160 423048
rect 556212 423036 556218 423088
rect 512822 422968 512828 423020
rect 512880 423008 512886 423020
rect 557626 423008 557632 423020
rect 512880 422980 557632 423008
rect 512880 422968 512886 422980
rect 557626 422968 557632 422980
rect 557684 422968 557690 423020
rect 512730 422900 512736 422952
rect 512788 422940 512794 422952
rect 559098 422940 559104 422952
rect 512788 422912 559104 422940
rect 512788 422900 512794 422912
rect 559098 422900 559104 422912
rect 559156 422900 559162 422952
rect 522390 422764 522396 422816
rect 522448 422804 522454 422816
rect 529658 422804 529664 422816
rect 522448 422776 529664 422804
rect 522448 422764 522454 422776
rect 529658 422764 529664 422776
rect 529716 422764 529722 422816
rect 519630 422356 519636 422408
rect 519688 422396 519694 422408
rect 525242 422396 525248 422408
rect 519688 422368 525248 422396
rect 519688 422356 519694 422368
rect 525242 422356 525248 422368
rect 525300 422356 525306 422408
rect 515582 421880 515588 421932
rect 515640 421920 515646 421932
rect 520826 421920 520832 421932
rect 515640 421892 520832 421920
rect 515640 421880 515646 421892
rect 520826 421880 520832 421892
rect 520884 421880 520890 421932
rect 547138 421540 547144 421592
rect 547196 421580 547202 421592
rect 554682 421580 554688 421592
rect 547196 421552 554688 421580
rect 547196 421540 547202 421552
rect 554682 421540 554688 421552
rect 554740 421540 554746 421592
rect 416774 420316 416780 420368
rect 416832 420356 416838 420368
rect 419442 420356 419448 420368
rect 416832 420328 419448 420356
rect 416832 420316 416838 420328
rect 419442 420316 419448 420328
rect 419500 420316 419506 420368
rect 518526 420180 518532 420232
rect 518584 420220 518590 420232
rect 541434 420220 541440 420232
rect 518584 420192 541440 420220
rect 518584 420180 518590 420192
rect 541434 420180 541440 420192
rect 541492 420180 541498 420232
rect 419350 419704 419356 419756
rect 419408 419744 419414 419756
rect 421650 419744 421656 419756
rect 419408 419716 421656 419744
rect 419408 419704 419414 419716
rect 421650 419704 421656 419716
rect 421708 419704 421714 419756
rect 415946 419500 415952 419552
rect 416004 419540 416010 419552
rect 420914 419540 420920 419552
rect 416004 419512 420920 419540
rect 416004 419500 416010 419512
rect 420914 419500 420920 419512
rect 420972 419500 420978 419552
rect 382918 418752 382924 418804
rect 382976 418792 382982 418804
rect 439498 418792 439504 418804
rect 382976 418764 439504 418792
rect 382976 418752 382982 418764
rect 439498 418752 439504 418764
rect 439556 418752 439562 418804
rect 407114 418616 407120 418668
rect 407172 418656 407178 418668
rect 408862 418656 408868 418668
rect 407172 418628 408868 418656
rect 407172 418616 407178 418628
rect 408862 418616 408868 418628
rect 408920 418616 408926 418668
rect 413370 418140 413376 418192
rect 413428 418180 413434 418192
rect 413428 418152 415440 418180
rect 413428 418140 413434 418152
rect 415412 418112 415440 418152
rect 417418 418112 417424 418124
rect 415412 418084 417424 418112
rect 417418 418072 417424 418084
rect 417476 418072 417482 418124
rect 420270 418072 420276 418124
rect 420328 418112 420334 418124
rect 424318 418112 424324 418124
rect 420328 418084 424324 418112
rect 420328 418072 420334 418084
rect 424318 418072 424324 418084
rect 424376 418072 424382 418124
rect 424042 417392 424048 417444
rect 424100 417432 424106 417444
rect 443638 417432 443644 417444
rect 424100 417404 443644 417432
rect 424100 417392 424106 417404
rect 443638 417392 443644 417404
rect 443696 417392 443702 417444
rect 408862 416712 408868 416764
rect 408920 416752 408926 416764
rect 410610 416752 410616 416764
rect 408920 416724 410616 416752
rect 408920 416712 408926 416724
rect 410610 416712 410616 416724
rect 410668 416712 410674 416764
rect 414750 416712 414756 416764
rect 414808 416752 414814 416764
rect 421558 416752 421564 416764
rect 414808 416724 421564 416752
rect 414808 416712 414814 416724
rect 421558 416712 421564 416724
rect 421616 416712 421622 416764
rect 421834 416304 421840 416356
rect 421892 416344 421898 416356
rect 422202 416344 422208 416356
rect 421892 416316 422208 416344
rect 421892 416304 421898 416316
rect 422202 416304 422208 416316
rect 422260 416304 422266 416356
rect 423122 416304 423128 416356
rect 423180 416344 423186 416356
rect 423582 416344 423588 416356
rect 423180 416316 423588 416344
rect 423180 416304 423186 416316
rect 423582 416304 423588 416316
rect 423640 416304 423646 416356
rect 392670 416032 392676 416084
rect 392728 416072 392734 416084
rect 398098 416072 398104 416084
rect 392728 416044 398104 416072
rect 392728 416032 392734 416044
rect 398098 416032 398104 416044
rect 398156 416032 398162 416084
rect 381538 414672 381544 414724
rect 381596 414712 381602 414724
rect 386598 414712 386604 414724
rect 381596 414684 386604 414712
rect 381596 414672 381602 414684
rect 386598 414672 386604 414684
rect 386656 414672 386662 414724
rect 419442 413244 419448 413296
rect 419500 413284 419506 413296
rect 428458 413284 428464 413296
rect 419500 413256 428464 413284
rect 419500 413244 419506 413256
rect 428458 413244 428464 413256
rect 428516 413244 428522 413296
rect 420914 412972 420920 413024
rect 420972 413012 420978 413024
rect 423674 413012 423680 413024
rect 420972 412984 423680 413012
rect 420972 412972 420978 412984
rect 423674 412972 423680 412984
rect 423732 412972 423738 413024
rect 522298 411884 522304 411936
rect 522356 411924 522362 411936
rect 580442 411924 580448 411936
rect 522356 411896 580448 411924
rect 522356 411884 522362 411896
rect 580442 411884 580448 411896
rect 580500 411884 580506 411936
rect 398098 411748 398104 411800
rect 398156 411788 398162 411800
rect 398834 411788 398840 411800
rect 398156 411760 398840 411788
rect 398156 411748 398162 411760
rect 398834 411748 398840 411760
rect 398892 411748 398898 411800
rect 424318 411748 424324 411800
rect 424376 411788 424382 411800
rect 425790 411788 425796 411800
rect 424376 411760 425796 411788
rect 424376 411748 424382 411760
rect 425790 411748 425796 411760
rect 425848 411748 425854 411800
rect 421650 411544 421656 411596
rect 421708 411584 421714 411596
rect 424410 411584 424416 411596
rect 421708 411556 424416 411584
rect 421708 411544 421714 411556
rect 424410 411544 424416 411556
rect 424468 411544 424474 411596
rect 386598 410524 386604 410576
rect 386656 410564 386662 410576
rect 403710 410564 403716 410576
rect 386656 410536 403716 410564
rect 386656 410524 386662 410536
rect 403710 410524 403716 410536
rect 403768 410524 403774 410576
rect 410610 409300 410616 409352
rect 410668 409340 410674 409352
rect 412082 409340 412088 409352
rect 410668 409312 412088 409340
rect 410668 409300 410674 409312
rect 412082 409300 412088 409312
rect 412140 409300 412146 409352
rect 423674 408484 423680 408536
rect 423732 408524 423738 408536
rect 423732 408496 426480 408524
rect 423732 408484 423738 408496
rect 426452 408456 426480 408496
rect 428550 408456 428556 408468
rect 426452 408428 428556 408456
rect 428550 408416 428556 408428
rect 428608 408416 428614 408468
rect 425790 408348 425796 408400
rect 425848 408388 425854 408400
rect 427078 408388 427084 408400
rect 425848 408360 427084 408388
rect 425848 408348 425854 408360
rect 427078 408348 427084 408360
rect 427136 408348 427142 408400
rect 382274 407124 382280 407176
rect 382332 407164 382338 407176
rect 435358 407164 435364 407176
rect 382332 407136 435364 407164
rect 382332 407124 382338 407136
rect 435358 407124 435364 407136
rect 435416 407124 435422 407176
rect 461578 406376 461584 406428
rect 461636 406416 461642 406428
rect 473354 406416 473360 406428
rect 461636 406388 473360 406416
rect 461636 406376 461642 406388
rect 473354 406376 473360 406388
rect 473412 406376 473418 406428
rect 398834 405628 398840 405680
rect 398892 405668 398898 405680
rect 401502 405668 401508 405680
rect 398892 405640 401508 405668
rect 398892 405628 398898 405640
rect 401502 405628 401508 405640
rect 401560 405628 401566 405680
rect 380158 404948 380164 405000
rect 380216 404988 380222 405000
rect 389910 404988 389916 405000
rect 380216 404960 389916 404988
rect 380216 404948 380222 404960
rect 389910 404948 389916 404960
rect 389968 404948 389974 405000
rect 421558 404540 421564 404592
rect 421616 404580 421622 404592
rect 424318 404580 424324 404592
rect 421616 404552 424324 404580
rect 421616 404540 421622 404552
rect 424318 404540 424324 404552
rect 424376 404540 424382 404592
rect 401502 401616 401508 401668
rect 401560 401656 401566 401668
rect 401560 401628 402974 401656
rect 401560 401616 401566 401628
rect 402946 401588 402974 401628
rect 404998 401588 405004 401600
rect 402946 401560 405004 401588
rect 404998 401548 405004 401560
rect 405056 401548 405062 401600
rect 412082 400120 412088 400172
rect 412140 400160 412146 400172
rect 415302 400160 415308 400172
rect 412140 400132 415308 400160
rect 412140 400120 412146 400132
rect 415302 400120 415308 400132
rect 415360 400120 415366 400172
rect 382274 396040 382280 396092
rect 382332 396080 382338 396092
rect 436738 396080 436744 396092
rect 382332 396052 436744 396080
rect 382332 396040 382338 396052
rect 436738 396040 436744 396052
rect 436796 396040 436802 396092
rect 417418 394748 417424 394800
rect 417476 394788 417482 394800
rect 417476 394760 419580 394788
rect 417476 394748 417482 394760
rect 415394 394612 415400 394664
rect 415452 394652 415458 394664
rect 417418 394652 417424 394664
rect 415452 394624 417424 394652
rect 415452 394612 415458 394624
rect 417418 394612 417424 394624
rect 417476 394612 417482 394664
rect 419552 394652 419580 394760
rect 421558 394652 421564 394664
rect 419552 394624 421564 394652
rect 421558 394612 421564 394624
rect 421616 394612 421622 394664
rect 411990 391892 411996 391944
rect 412048 391932 412054 391944
rect 414566 391932 414572 391944
rect 412048 391904 414572 391932
rect 412048 391892 412054 391904
rect 414566 391892 414572 391904
rect 414624 391892 414630 391944
rect 424410 390804 424416 390856
rect 424468 390844 424474 390856
rect 425790 390844 425796 390856
rect 424468 390816 425796 390844
rect 424468 390804 424474 390816
rect 425790 390804 425796 390816
rect 425848 390804 425854 390856
rect 414566 389172 414572 389224
rect 414624 389212 414630 389224
rect 417510 389212 417516 389224
rect 414624 389184 417516 389212
rect 414624 389172 414630 389184
rect 417510 389172 417516 389184
rect 417568 389172 417574 389224
rect 403710 388900 403716 388952
rect 403768 388940 403774 388952
rect 406470 388940 406476 388952
rect 403768 388912 406476 388940
rect 403768 388900 403774 388912
rect 406470 388900 406476 388912
rect 406528 388900 406534 388952
rect 427078 387812 427084 387864
rect 427136 387852 427142 387864
rect 427136 387824 427860 387852
rect 427136 387812 427142 387824
rect 427832 387784 427860 387824
rect 429838 387784 429844 387796
rect 427832 387756 429844 387784
rect 429838 387744 429844 387756
rect 429896 387744 429902 387796
rect 471882 387064 471888 387116
rect 471940 387104 471946 387116
rect 490558 387104 490564 387116
rect 471940 387076 490564 387104
rect 471940 387064 471946 387076
rect 490558 387064 490564 387076
rect 490616 387064 490622 387116
rect 382274 386384 382280 386436
rect 382332 386424 382338 386436
rect 443730 386424 443736 386436
rect 382332 386396 443736 386424
rect 382332 386384 382338 386396
rect 443730 386384 443736 386396
rect 443788 386384 443794 386436
rect 389910 385636 389916 385688
rect 389968 385676 389974 385688
rect 398098 385676 398104 385688
rect 389968 385648 398104 385676
rect 389968 385636 389974 385648
rect 398098 385636 398104 385648
rect 398156 385636 398162 385688
rect 468938 385636 468944 385688
rect 468996 385676 469002 385688
rect 485038 385676 485044 385688
rect 468996 385648 485044 385676
rect 468996 385636 469002 385648
rect 485038 385636 485044 385648
rect 485096 385636 485102 385688
rect 515674 385636 515680 385688
rect 515732 385676 515738 385688
rect 547874 385676 547880 385688
rect 515732 385648 547880 385676
rect 515732 385636 515738 385648
rect 547874 385636 547880 385648
rect 547932 385636 547938 385688
rect 470226 384344 470232 384396
rect 470284 384384 470290 384396
rect 479518 384384 479524 384396
rect 470284 384356 479524 384384
rect 470284 384344 470290 384356
rect 479518 384344 479524 384356
rect 479576 384344 479582 384396
rect 447594 384276 447600 384328
rect 447652 384316 447658 384328
rect 454770 384316 454776 384328
rect 447652 384288 454776 384316
rect 447652 384276 447658 384288
rect 454770 384276 454776 384288
rect 454828 384276 454834 384328
rect 467650 384276 467656 384328
rect 467708 384316 467714 384328
rect 483014 384316 483020 384328
rect 467708 384288 483020 384316
rect 467708 384276 467714 384288
rect 483014 384276 483020 384288
rect 483072 384276 483078 384328
rect 519722 384276 519728 384328
rect 519780 384316 519786 384328
rect 542354 384316 542360 384328
rect 519780 384288 542360 384316
rect 519780 384276 519786 384288
rect 542354 384276 542360 384288
rect 542412 384276 542418 384328
rect 468478 383596 468484 383648
rect 468536 383636 468542 383648
rect 477954 383636 477960 383648
rect 468536 383608 477960 383636
rect 468536 383596 468542 383608
rect 477954 383596 477960 383608
rect 478012 383596 478018 383648
rect 467098 383528 467104 383580
rect 467156 383568 467162 383580
rect 479242 383568 479248 383580
rect 467156 383540 479248 383568
rect 467156 383528 467162 383540
rect 479242 383528 479248 383540
rect 479300 383528 479306 383580
rect 469858 383460 469864 383512
rect 469916 383500 469922 383512
rect 481818 383500 481824 383512
rect 469916 383472 481824 383500
rect 469916 383460 469922 383472
rect 481818 383460 481824 383472
rect 481876 383460 481882 383512
rect 462958 383392 462964 383444
rect 463016 383432 463022 383444
rect 476666 383432 476672 383444
rect 463016 383404 476672 383432
rect 463016 383392 463022 383404
rect 476666 383392 476672 383404
rect 476724 383392 476730 383444
rect 471238 383324 471244 383376
rect 471296 383364 471302 383376
rect 486970 383364 486976 383376
rect 471296 383336 486976 383364
rect 471296 383324 471302 383336
rect 486970 383324 486976 383336
rect 487028 383324 487034 383376
rect 468570 383256 468576 383308
rect 468628 383296 468634 383308
rect 485682 383296 485688 383308
rect 468628 383268 485688 383296
rect 468628 383256 468634 383268
rect 485682 383256 485688 383268
rect 485740 383256 485746 383308
rect 467190 383188 467196 383240
rect 467248 383228 467254 383240
rect 483106 383228 483112 383240
rect 467248 383200 483112 383228
rect 467248 383188 467254 383200
rect 483106 383188 483112 383200
rect 483164 383188 483170 383240
rect 463050 383120 463056 383172
rect 463108 383160 463114 383172
rect 480530 383160 480536 383172
rect 463108 383132 480536 383160
rect 463108 383120 463114 383132
rect 480530 383120 480536 383132
rect 480588 383120 480594 383172
rect 424318 383052 424324 383104
rect 424376 383092 424382 383104
rect 425698 383092 425704 383104
rect 424376 383064 425704 383092
rect 424376 383052 424382 383064
rect 425698 383052 425704 383064
rect 425756 383052 425762 383104
rect 467282 383052 467288 383104
rect 467340 383092 467346 383104
rect 484394 383092 484400 383104
rect 467340 383064 484400 383092
rect 467340 383052 467346 383064
rect 484394 383052 484400 383064
rect 484452 383052 484458 383104
rect 448054 382984 448060 383036
rect 448112 383024 448118 383036
rect 456058 383024 456064 383036
rect 448112 382996 456064 383024
rect 448112 382984 448118 382996
rect 456058 382984 456064 382996
rect 456116 382984 456122 383036
rect 464338 382984 464344 383036
rect 464396 383024 464402 383036
rect 488258 383024 488264 383036
rect 464396 382996 488264 383024
rect 464396 382984 464402 382996
rect 488258 382984 488264 382996
rect 488316 382984 488322 383036
rect 494698 382984 494704 383036
rect 494756 383024 494762 383036
rect 506290 383024 506296 383036
rect 494756 382996 506296 383024
rect 494756 382984 494762 382996
rect 506290 382984 506296 382996
rect 506348 382984 506354 383036
rect 450630 382916 450636 382968
rect 450688 382956 450694 382968
rect 554958 382956 554964 382968
rect 450688 382928 554964 382956
rect 450688 382916 450694 382928
rect 554958 382916 554964 382928
rect 555016 382916 555022 382968
rect 404998 382372 405004 382424
rect 405056 382412 405062 382424
rect 408402 382412 408408 382424
rect 405056 382384 408408 382412
rect 405056 382372 405062 382384
rect 408402 382372 408408 382384
rect 408460 382372 408466 382424
rect 442902 382236 442908 382288
rect 442960 382276 442966 382288
rect 450630 382276 450636 382288
rect 442960 382248 450636 382276
rect 442960 382236 442966 382248
rect 450630 382236 450636 382248
rect 450688 382236 450694 382288
rect 452562 382236 452568 382288
rect 452620 382276 452626 382288
rect 453482 382276 453488 382288
rect 452620 382248 453488 382276
rect 452620 382236 452626 382248
rect 453482 382236 453488 382248
rect 453540 382236 453546 382288
rect 455322 382236 455328 382288
rect 455380 382276 455386 382288
rect 456058 382276 456064 382288
rect 455380 382248 456064 382276
rect 455380 382236 455386 382248
rect 456058 382236 456064 382248
rect 456116 382236 456122 382288
rect 450630 381624 450636 381676
rect 450688 381664 450694 381676
rect 457438 381664 457444 381676
rect 450688 381636 457444 381664
rect 450688 381624 450694 381636
rect 457438 381624 457444 381636
rect 457496 381624 457502 381676
rect 447962 381556 447968 381608
rect 448020 381596 448026 381608
rect 461670 381596 461676 381608
rect 448020 381568 461676 381596
rect 448020 381556 448026 381568
rect 461670 381556 461676 381568
rect 461728 381556 461734 381608
rect 448146 381488 448152 381540
rect 448204 381528 448210 381540
rect 496078 381528 496084 381540
rect 448204 381500 496084 381528
rect 448204 381488 448210 381500
rect 496078 381488 496084 381500
rect 496136 381488 496142 381540
rect 514110 381488 514116 381540
rect 514168 381528 514174 381540
rect 539594 381528 539600 381540
rect 514168 381500 539600 381528
rect 514168 381488 514174 381500
rect 539594 381488 539600 381500
rect 539652 381488 539658 381540
rect 428458 381012 428464 381064
rect 428516 381052 428522 381064
rect 431218 381052 431224 381064
rect 428516 381024 431224 381052
rect 428516 381012 428522 381024
rect 431218 381012 431224 381024
rect 431276 381012 431282 381064
rect 428550 380944 428556 380996
rect 428608 380984 428614 380996
rect 429930 380984 429936 380996
rect 428608 380956 429936 380984
rect 428608 380944 428614 380956
rect 429930 380944 429936 380956
rect 429988 380944 429994 380996
rect 464430 380440 464436 380452
rect 460906 380412 464436 380440
rect 447410 380196 447416 380248
rect 447468 380236 447474 380248
rect 454678 380236 454684 380248
rect 447468 380208 454684 380236
rect 447468 380196 447474 380208
rect 454678 380196 454684 380208
rect 454736 380196 454742 380248
rect 447870 380128 447876 380180
rect 447928 380168 447934 380180
rect 460906 380168 460934 380412
rect 464430 380400 464436 380412
rect 464488 380400 464494 380452
rect 447928 380140 460934 380168
rect 447928 380128 447934 380140
rect 515766 380128 515772 380180
rect 515824 380168 515830 380180
rect 535454 380168 535460 380180
rect 515824 380140 535460 380168
rect 515824 380128 515830 380140
rect 535454 380128 535460 380140
rect 535512 380128 535518 380180
rect 542998 380128 543004 380180
rect 543056 380168 543062 380180
rect 561674 380168 561680 380180
rect 543056 380140 561680 380168
rect 543056 380128 543062 380140
rect 561674 380128 561680 380140
rect 561732 380128 561738 380180
rect 448330 379788 448336 379840
rect 448388 379828 448394 379840
rect 453298 379828 453304 379840
rect 448388 379800 453304 379828
rect 448388 379788 448394 379800
rect 453298 379788 453304 379800
rect 453356 379788 453362 379840
rect 449802 379516 449808 379568
rect 449860 379556 449866 379568
rect 564526 379556 564532 379568
rect 449860 379528 564532 379556
rect 449860 379516 449866 379528
rect 564526 379516 564532 379528
rect 564584 379516 564590 379568
rect 398098 379448 398104 379500
rect 398156 379488 398162 379500
rect 403710 379488 403716 379500
rect 398156 379460 403716 379488
rect 398156 379448 398162 379460
rect 403710 379448 403716 379460
rect 403768 379448 403774 379500
rect 512822 379448 512828 379500
rect 512880 379488 512886 379500
rect 542998 379488 543004 379500
rect 512880 379460 543004 379488
rect 512880 379448 512886 379460
rect 542998 379448 543004 379460
rect 543056 379448 543062 379500
rect 570782 378156 570788 378208
rect 570840 378196 570846 378208
rect 579614 378196 579620 378208
rect 570840 378168 579620 378196
rect 570840 378156 570846 378168
rect 579614 378156 579620 378168
rect 579672 378156 579678 378208
rect 512270 378088 512276 378140
rect 512328 378128 512334 378140
rect 547138 378128 547144 378140
rect 512328 378100 547144 378128
rect 512328 378088 512334 378100
rect 547138 378088 547144 378100
rect 547196 378088 547202 378140
rect 512730 377408 512736 377460
rect 512788 377448 512794 377460
rect 536834 377448 536840 377460
rect 512788 377420 536840 377448
rect 512788 377408 512794 377420
rect 536834 377408 536840 377420
rect 536892 377408 536898 377460
rect 406470 376660 406476 376712
rect 406528 376700 406534 376712
rect 411990 376700 411996 376712
rect 406528 376672 411996 376700
rect 406528 376660 406534 376672
rect 411990 376660 411996 376672
rect 412048 376660 412054 376712
rect 447134 376700 447140 376712
rect 412606 376672 447140 376700
rect 403618 376592 403624 376644
rect 403676 376632 403682 376644
rect 412606 376632 412634 376672
rect 447134 376660 447140 376672
rect 447192 376660 447198 376712
rect 403676 376604 412634 376632
rect 403676 376592 403682 376604
rect 417510 376592 417516 376644
rect 417568 376632 417574 376644
rect 420730 376632 420736 376644
rect 417568 376604 420736 376632
rect 417568 376592 417574 376604
rect 420730 376592 420736 376604
rect 420788 376592 420794 376644
rect 513190 376592 513196 376644
rect 513248 376632 513254 376644
rect 540238 376632 540244 376644
rect 513248 376604 540244 376632
rect 513248 376592 513254 376604
rect 540238 376592 540244 376604
rect 540296 376592 540302 376644
rect 408494 376524 408500 376576
rect 408552 376564 408558 376576
rect 412266 376564 412272 376576
rect 408552 376536 412272 376564
rect 408552 376524 408558 376536
rect 412266 376524 412272 376536
rect 412324 376524 412330 376576
rect 513098 376524 513104 376576
rect 513156 376564 513162 376576
rect 538858 376564 538864 376576
rect 513156 376536 538864 376564
rect 513156 376524 513162 376536
rect 538858 376524 538864 376536
rect 538916 376524 538922 376576
rect 513282 376456 513288 376508
rect 513340 376496 513346 376508
rect 544378 376496 544384 376508
rect 513340 376468 544384 376496
rect 513340 376456 513346 376468
rect 544378 376456 544384 376468
rect 544436 376456 544442 376508
rect 512270 375912 512276 375964
rect 512328 375952 512334 375964
rect 515674 375952 515680 375964
rect 512328 375924 515680 375952
rect 512328 375912 512334 375924
rect 515674 375912 515680 375924
rect 515732 375912 515738 375964
rect 382274 375368 382280 375420
rect 382332 375408 382338 375420
rect 439590 375408 439596 375420
rect 382332 375380 439596 375408
rect 382332 375368 382338 375380
rect 439590 375368 439596 375380
rect 439648 375368 439654 375420
rect 395338 375300 395344 375352
rect 395396 375340 395402 375352
rect 447318 375340 447324 375352
rect 395396 375312 447324 375340
rect 395396 375300 395402 375312
rect 447318 375300 447324 375312
rect 447376 375300 447382 375352
rect 512086 375300 512092 375352
rect 512144 375340 512150 375352
rect 537478 375340 537484 375352
rect 512144 375312 537484 375340
rect 512144 375300 512150 375312
rect 537478 375300 537484 375312
rect 537536 375300 537542 375352
rect 396718 375232 396724 375284
rect 396776 375272 396782 375284
rect 447134 375272 447140 375284
rect 396776 375244 447140 375272
rect 396776 375232 396782 375244
rect 447134 375232 447140 375244
rect 447192 375232 447198 375284
rect 513282 375232 513288 375284
rect 513340 375272 513346 375284
rect 536098 375272 536104 375284
rect 513340 375244 536104 375272
rect 513340 375232 513346 375244
rect 536098 375232 536104 375244
rect 536156 375232 536162 375284
rect 439498 375164 439504 375216
rect 439556 375204 439562 375216
rect 447226 375204 447232 375216
rect 439556 375176 447232 375204
rect 439556 375164 439562 375176
rect 447226 375164 447232 375176
rect 447284 375164 447290 375216
rect 512822 375164 512828 375216
rect 512880 375204 512886 375216
rect 533338 375204 533344 375216
rect 512880 375176 533344 375204
rect 512880 375164 512886 375176
rect 533338 375164 533344 375176
rect 533396 375164 533402 375216
rect 393958 373940 393964 373992
rect 394016 373980 394022 373992
rect 447226 373980 447232 373992
rect 394016 373952 447232 373980
rect 394016 373940 394022 373952
rect 447226 373940 447232 373952
rect 447284 373940 447290 373992
rect 513282 373940 513288 373992
rect 513340 373980 513346 373992
rect 519722 373980 519728 373992
rect 513340 373952 519728 373980
rect 513340 373940 513346 373952
rect 519722 373940 519728 373952
rect 519780 373940 519786 373992
rect 399478 373872 399484 373924
rect 399536 373912 399542 373924
rect 447134 373912 447140 373924
rect 399536 373884 447140 373912
rect 399536 373872 399542 373884
rect 447134 373872 447140 373884
rect 447192 373872 447198 373924
rect 513282 373464 513288 373516
rect 513340 373504 513346 373516
rect 518526 373504 518532 373516
rect 513340 373476 518532 373504
rect 513340 373464 513346 373476
rect 518526 373464 518532 373476
rect 518584 373464 518590 373516
rect 511994 373328 512000 373380
rect 512052 373368 512058 373380
rect 514110 373368 514116 373380
rect 512052 373340 514116 373368
rect 512052 373328 512058 373340
rect 514110 373328 514116 373340
rect 514168 373328 514174 373380
rect 517514 373260 517520 373312
rect 517572 373300 517578 373312
rect 538214 373300 538220 373312
rect 517572 373272 538220 373300
rect 517572 373260 517578 373272
rect 538214 373260 538220 373272
rect 538272 373260 538278 373312
rect 429930 373124 429936 373176
rect 429988 373164 429994 373176
rect 430942 373164 430948 373176
rect 429988 373136 430948 373164
rect 429988 373124 429994 373136
rect 430942 373124 430948 373136
rect 431000 373124 431006 373176
rect 412266 372580 412272 372632
rect 412324 372620 412330 372632
rect 415118 372620 415124 372632
rect 412324 372592 415124 372620
rect 412324 372580 412330 372592
rect 415118 372580 415124 372592
rect 415176 372580 415182 372632
rect 392578 372512 392584 372564
rect 392636 372552 392642 372564
rect 447318 372552 447324 372564
rect 392636 372524 447324 372552
rect 392636 372512 392642 372524
rect 447318 372512 447324 372524
rect 447376 372512 447382 372564
rect 513282 372512 513288 372564
rect 513340 372552 513346 372564
rect 517514 372552 517520 372564
rect 513340 372524 517520 372552
rect 513340 372512 513346 372524
rect 517514 372512 517520 372524
rect 517572 372512 517578 372564
rect 534074 372552 534080 372564
rect 518866 372524 534080 372552
rect 406378 372444 406384 372496
rect 406436 372484 406442 372496
rect 447134 372484 447140 372496
rect 406436 372456 447140 372484
rect 406436 372444 406442 372456
rect 447134 372444 447140 372456
rect 447192 372444 447198 372496
rect 513190 372444 513196 372496
rect 513248 372484 513254 372496
rect 518866 372484 518894 372524
rect 534074 372512 534080 372524
rect 534132 372512 534138 372564
rect 513248 372456 518894 372484
rect 513248 372444 513254 372456
rect 419074 372376 419080 372428
rect 419132 372416 419138 372428
rect 447226 372416 447232 372428
rect 419132 372388 447232 372416
rect 419132 372376 419138 372388
rect 447226 372376 447232 372388
rect 447284 372376 447290 372428
rect 421558 371900 421564 371952
rect 421616 371940 421622 371952
rect 422938 371940 422944 371952
rect 421616 371912 422944 371940
rect 421616 371900 421622 371912
rect 422938 371900 422944 371912
rect 422996 371900 423002 371952
rect 512454 371764 512460 371816
rect 512512 371804 512518 371816
rect 515766 371804 515772 371816
rect 512512 371776 515772 371804
rect 512512 371764 512518 371776
rect 515766 371764 515772 371776
rect 515824 371764 515830 371816
rect 417418 371492 417424 371544
rect 417476 371532 417482 371544
rect 418706 371532 418712 371544
rect 417476 371504 418712 371532
rect 417476 371492 417482 371504
rect 418706 371492 418712 371504
rect 418764 371492 418770 371544
rect 425790 371492 425796 371544
rect 425848 371532 425854 371544
rect 427078 371532 427084 371544
rect 425848 371504 427084 371532
rect 425848 371492 425854 371504
rect 427078 371492 427084 371504
rect 427136 371492 427142 371544
rect 389818 371152 389824 371204
rect 389876 371192 389882 371204
rect 447318 371192 447324 371204
rect 389876 371164 447324 371192
rect 389876 371152 389882 371164
rect 447318 371152 447324 371164
rect 447376 371152 447382 371204
rect 513190 371152 513196 371204
rect 513248 371192 513254 371204
rect 529934 371192 529940 371204
rect 513248 371164 529940 371192
rect 513248 371152 513254 371164
rect 529934 371152 529940 371164
rect 529992 371152 529998 371204
rect 391198 371084 391204 371136
rect 391256 371124 391262 371136
rect 447226 371124 447232 371136
rect 391256 371096 447232 371124
rect 391256 371084 391262 371096
rect 447226 371084 447232 371096
rect 447284 371084 447290 371136
rect 513282 371084 513288 371136
rect 513340 371124 513346 371136
rect 523678 371124 523684 371136
rect 513340 371096 523684 371124
rect 513340 371084 513346 371096
rect 523678 371084 523684 371096
rect 523736 371084 523742 371136
rect 407758 371016 407764 371068
rect 407816 371056 407822 371068
rect 447134 371056 447140 371068
rect 407816 371028 447140 371056
rect 407816 371016 407822 371028
rect 447134 371016 447140 371028
rect 447192 371016 447198 371068
rect 513098 371016 513104 371068
rect 513156 371056 513162 371068
rect 522390 371056 522396 371068
rect 513156 371028 522396 371056
rect 513156 371016 513162 371028
rect 522390 371016 522396 371028
rect 522448 371016 522454 371068
rect 418706 370948 418712 371000
rect 418764 370988 418770 371000
rect 420270 370988 420276 371000
rect 418764 370960 420276 370988
rect 418764 370948 418770 370960
rect 420270 370948 420276 370960
rect 420328 370948 420334 371000
rect 420730 370948 420736 371000
rect 420788 370988 420794 371000
rect 423306 370988 423312 371000
rect 420788 370960 423312 370988
rect 420788 370948 420794 370960
rect 423306 370948 423312 370960
rect 423364 370948 423370 371000
rect 385678 369792 385684 369844
rect 385736 369832 385742 369844
rect 447226 369832 447232 369844
rect 385736 369804 447232 369832
rect 385736 369792 385742 369804
rect 447226 369792 447232 369804
rect 447284 369792 447290 369844
rect 513282 369792 513288 369844
rect 513340 369832 513346 369844
rect 525794 369832 525800 369844
rect 513340 369804 525800 369832
rect 513340 369792 513346 369804
rect 525794 369792 525800 369804
rect 525852 369792 525858 369844
rect 387058 369724 387064 369776
rect 387116 369764 387122 369776
rect 447134 369764 447140 369776
rect 387116 369736 447140 369764
rect 387116 369724 387122 369736
rect 447134 369724 447140 369736
rect 447192 369724 447198 369776
rect 513190 369724 513196 369776
rect 513248 369764 513254 369776
rect 523034 369764 523040 369776
rect 513248 369736 523040 369764
rect 513248 369724 513254 369736
rect 523034 369724 523040 369736
rect 523092 369724 523098 369776
rect 430942 369656 430948 369708
rect 431000 369696 431006 369708
rect 432690 369696 432696 369708
rect 431000 369668 432696 369696
rect 431000 369656 431006 369668
rect 432690 369656 432696 369668
rect 432748 369656 432754 369708
rect 513098 369656 513104 369708
rect 513156 369696 513162 369708
rect 518434 369696 518440 369708
rect 513156 369668 518440 369696
rect 513156 369656 513162 369668
rect 518434 369656 518440 369668
rect 518492 369656 518498 369708
rect 403710 369520 403716 369572
rect 403768 369560 403774 369572
rect 409138 369560 409144 369572
rect 403768 369532 409144 369560
rect 403768 369520 403774 369532
rect 409138 369520 409144 369532
rect 409196 369520 409202 369572
rect 513282 369044 513288 369096
rect 513340 369084 513346 369096
rect 519630 369084 519636 369096
rect 513340 369056 519636 369084
rect 513340 369044 513346 369056
rect 519630 369044 519636 369056
rect 519688 369044 519694 369096
rect 423306 368568 423312 368620
rect 423364 368608 423370 368620
rect 424318 368608 424324 368620
rect 423364 368580 424324 368608
rect 423364 368568 423370 368580
rect 424318 368568 424324 368580
rect 424376 368568 424382 368620
rect 384298 368432 384304 368484
rect 384356 368472 384362 368484
rect 447134 368472 447140 368484
rect 384356 368444 447140 368472
rect 384356 368432 384362 368444
rect 447134 368432 447140 368444
rect 447192 368432 447198 368484
rect 512178 368432 512184 368484
rect 512236 368472 512242 368484
rect 521654 368472 521660 368484
rect 512236 368444 521660 368472
rect 512236 368432 512242 368444
rect 521654 368432 521660 368444
rect 521712 368432 521718 368484
rect 410518 368364 410524 368416
rect 410576 368404 410582 368416
rect 447226 368404 447232 368416
rect 410576 368376 447232 368404
rect 410576 368364 410582 368376
rect 447226 368364 447232 368376
rect 447284 368364 447290 368416
rect 411898 368296 411904 368348
rect 411956 368336 411962 368348
rect 447318 368336 447324 368348
rect 411956 368308 447324 368336
rect 411956 368296 411962 368308
rect 447318 368296 447324 368308
rect 447376 368296 447382 368348
rect 415118 368228 415124 368280
rect 415176 368268 415182 368280
rect 420914 368268 420920 368280
rect 415176 368240 420920 368268
rect 415176 368228 415182 368240
rect 420914 368228 420920 368240
rect 420972 368228 420978 368280
rect 512270 367752 512276 367804
rect 512328 367792 512334 367804
rect 515582 367792 515588 367804
rect 512328 367764 515588 367792
rect 512328 367752 512334 367764
rect 515582 367752 515588 367764
rect 515640 367752 515646 367804
rect 513282 367072 513288 367124
rect 513340 367112 513346 367124
rect 547138 367112 547144 367124
rect 513340 367084 547144 367112
rect 513340 367072 513346 367084
rect 547138 367072 547144 367084
rect 547196 367072 547202 367124
rect 414658 367004 414664 367056
rect 414716 367044 414722 367056
rect 447134 367044 447140 367056
rect 414716 367016 447140 367044
rect 414716 367004 414722 367016
rect 447134 367004 447140 367016
rect 447192 367004 447198 367056
rect 419166 366936 419172 366988
rect 419224 366976 419230 366988
rect 447226 366976 447232 366988
rect 419224 366948 447232 366976
rect 419224 366936 419230 366948
rect 447226 366936 447232 366948
rect 447284 366936 447290 366988
rect 513190 366256 513196 366308
rect 513248 366296 513254 366308
rect 518894 366296 518900 366308
rect 513248 366268 518900 366296
rect 513248 366256 513254 366268
rect 518894 366256 518900 366268
rect 518952 366256 518958 366308
rect 513006 365712 513012 365764
rect 513064 365752 513070 365764
rect 547966 365752 547972 365764
rect 513064 365724 547972 365752
rect 513064 365712 513070 365724
rect 547966 365712 547972 365724
rect 548024 365712 548030 365764
rect 383010 365644 383016 365696
rect 383068 365684 383074 365696
rect 447318 365684 447324 365696
rect 383068 365656 447324 365684
rect 383068 365644 383074 365656
rect 447318 365644 447324 365656
rect 447376 365644 447382 365696
rect 399570 365576 399576 365628
rect 399628 365616 399634 365628
rect 447226 365616 447232 365628
rect 399628 365588 447232 365616
rect 399628 365576 399634 365588
rect 447226 365576 447232 365588
rect 447284 365576 447290 365628
rect 400858 365508 400864 365560
rect 400916 365548 400922 365560
rect 447134 365548 447140 365560
rect 400916 365520 447140 365548
rect 400916 365508 400922 365520
rect 447134 365508 447140 365520
rect 447192 365508 447198 365560
rect 420914 364964 420920 365016
rect 420972 365004 420978 365016
rect 425790 365004 425796 365016
rect 420972 364976 425796 365004
rect 420972 364964 420978 364976
rect 425790 364964 425796 364976
rect 425848 364964 425854 365016
rect 512914 364420 512920 364472
rect 512972 364460 512978 364472
rect 548058 364460 548064 364472
rect 512972 364432 548064 364460
rect 512972 364420 512978 364432
rect 548058 364420 548064 364432
rect 548116 364420 548122 364472
rect 431218 364352 431224 364404
rect 431276 364392 431282 364404
rect 432598 364392 432604 364404
rect 431276 364364 432604 364392
rect 431276 364352 431282 364364
rect 432598 364352 432604 364364
rect 432656 364352 432662 364404
rect 513282 364352 513288 364404
rect 513340 364392 513346 364404
rect 549346 364392 549352 364404
rect 513340 364364 549352 364392
rect 513340 364352 513346 364364
rect 549346 364352 549352 364364
rect 549404 364352 549410 364404
rect 572070 364352 572076 364404
rect 572128 364392 572134 364404
rect 580166 364392 580172 364404
rect 572128 364364 580172 364392
rect 572128 364352 572134 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 383194 364284 383200 364336
rect 383252 364324 383258 364336
rect 447226 364324 447232 364336
rect 383252 364296 447232 364324
rect 383252 364284 383258 364296
rect 447226 364284 447232 364296
rect 447284 364284 447290 364336
rect 383102 364216 383108 364268
rect 383160 364256 383166 364268
rect 447134 364256 447140 364268
rect 383160 364228 447140 364256
rect 383160 364216 383166 364228
rect 447134 364216 447140 364228
rect 447192 364216 447198 364268
rect 512086 363808 512092 363860
rect 512144 363848 512150 363860
rect 514754 363848 514760 363860
rect 512144 363820 514760 363848
rect 512144 363808 512150 363820
rect 514754 363808 514760 363820
rect 514812 363808 514818 363860
rect 382642 363604 382648 363656
rect 382700 363644 382706 363656
rect 443914 363644 443920 363656
rect 382700 363616 443920 363644
rect 382700 363604 382706 363616
rect 443914 363604 443920 363616
rect 443972 363604 443978 363656
rect 513006 363128 513012 363180
rect 513064 363168 513070 363180
rect 514846 363168 514852 363180
rect 513064 363140 514852 363168
rect 513064 363128 513070 363140
rect 514846 363128 514852 363140
rect 514904 363128 514910 363180
rect 420270 362924 420276 362976
rect 420328 362964 420334 362976
rect 421558 362964 421564 362976
rect 420328 362936 421564 362964
rect 420328 362924 420334 362936
rect 421558 362924 421564 362936
rect 421616 362924 421622 362976
rect 513282 362924 513288 362976
rect 513340 362964 513346 362976
rect 550542 362964 550548 362976
rect 513340 362936 550548 362964
rect 513340 362924 513346 362936
rect 550542 362924 550548 362936
rect 550600 362924 550606 362976
rect 435358 362856 435364 362908
rect 435416 362896 435422 362908
rect 447134 362896 447140 362908
rect 435416 362868 447140 362896
rect 435416 362856 435422 362868
rect 447134 362856 447140 362868
rect 447192 362856 447198 362908
rect 436738 362788 436744 362840
rect 436796 362828 436802 362840
rect 447226 362828 447232 362840
rect 436796 362800 447232 362828
rect 436796 362788 436802 362800
rect 447226 362788 447232 362800
rect 447284 362788 447290 362840
rect 443730 362720 443736 362772
rect 443788 362760 443794 362772
rect 447318 362760 447324 362772
rect 443788 362732 447324 362760
rect 443788 362720 443794 362732
rect 447318 362720 447324 362732
rect 447376 362720 447382 362772
rect 513190 362176 513196 362228
rect 513248 362216 513254 362228
rect 549162 362216 549168 362228
rect 513248 362188 549168 362216
rect 513248 362176 513254 362188
rect 549162 362176 549168 362188
rect 549220 362176 549226 362228
rect 512086 361904 512092 361956
rect 512144 361944 512150 361956
rect 514938 361944 514944 361956
rect 512144 361916 514944 361944
rect 512144 361904 512150 361916
rect 514938 361904 514944 361916
rect 514996 361904 515002 361956
rect 513282 361700 513288 361752
rect 513340 361740 513346 361752
rect 523034 361740 523040 361752
rect 513340 361712 523040 361740
rect 513340 361700 513346 361712
rect 523034 361700 523040 361712
rect 523092 361700 523098 361752
rect 512638 361632 512644 361684
rect 512696 361672 512702 361684
rect 517514 361672 517520 361684
rect 512696 361644 517520 361672
rect 512696 361632 512702 361644
rect 517514 361632 517520 361644
rect 517572 361632 517578 361684
rect 439590 361496 439596 361548
rect 439648 361536 439654 361548
rect 447134 361536 447140 361548
rect 439648 361508 447140 361536
rect 439648 361496 439654 361508
rect 447134 361496 447140 361508
rect 447192 361496 447198 361548
rect 443914 361428 443920 361480
rect 443972 361468 443978 361480
rect 447226 361468 447232 361480
rect 443972 361440 447232 361468
rect 443972 361428 443978 361440
rect 447226 361428 447232 361440
rect 447284 361428 447290 361480
rect 512822 360884 512828 360936
rect 512880 360924 512886 360936
rect 550726 360924 550732 360936
rect 512880 360896 550732 360924
rect 512880 360884 512886 360896
rect 550726 360884 550732 360896
rect 550784 360884 550790 360936
rect 513098 360816 513104 360868
rect 513156 360856 513162 360868
rect 513156 360828 547874 360856
rect 513156 360816 513162 360828
rect 409138 360748 409144 360800
rect 409196 360788 409202 360800
rect 411898 360788 411904 360800
rect 409196 360760 411904 360788
rect 409196 360748 409202 360760
rect 411898 360748 411904 360760
rect 411956 360748 411962 360800
rect 429838 360748 429844 360800
rect 429896 360788 429902 360800
rect 431310 360788 431316 360800
rect 429896 360760 431316 360788
rect 429896 360748 429902 360760
rect 431310 360748 431316 360760
rect 431368 360748 431374 360800
rect 547846 360720 547874 360828
rect 551922 360720 551928 360732
rect 547846 360692 551928 360720
rect 551922 360680 551928 360692
rect 551980 360680 551986 360732
rect 550726 360612 550732 360664
rect 550784 360652 550790 360664
rect 551462 360652 551468 360664
rect 550784 360624 551468 360652
rect 550784 360612 550790 360624
rect 551462 360612 551468 360624
rect 551520 360612 551526 360664
rect 513098 360204 513104 360256
rect 513156 360244 513162 360256
rect 520274 360244 520280 360256
rect 513156 360216 520280 360244
rect 513156 360204 513162 360216
rect 520274 360204 520280 360216
rect 520332 360204 520338 360256
rect 549346 360136 549352 360188
rect 549404 360176 549410 360188
rect 557166 360176 557172 360188
rect 549404 360148 557172 360176
rect 549404 360136 549410 360148
rect 557166 360136 557172 360148
rect 557224 360136 557230 360188
rect 517514 360068 517520 360120
rect 517572 360108 517578 360120
rect 550634 360108 550640 360120
rect 517572 360080 550640 360108
rect 517572 360068 517578 360080
rect 550634 360068 550640 360080
rect 550692 360068 550698 360120
rect 547138 360000 547144 360052
rect 547196 360040 547202 360052
rect 568758 360040 568764 360052
rect 547196 360012 568764 360040
rect 547196 360000 547202 360012
rect 568758 360000 568764 360012
rect 568816 360000 568822 360052
rect 550542 359932 550548 359984
rect 550600 359972 550606 359984
rect 553854 359972 553860 359984
rect 550600 359944 553860 359972
rect 550600 359932 550606 359944
rect 553854 359932 553860 359944
rect 553912 359932 553918 359984
rect 514754 359864 514760 359916
rect 514812 359904 514818 359916
rect 555786 359904 555792 359916
rect 514812 359876 555792 359904
rect 514812 359864 514818 359876
rect 555786 359864 555792 359876
rect 555844 359864 555850 359916
rect 547966 359796 547972 359848
rect 548024 359836 548030 359848
rect 567378 359836 567384 359848
rect 548024 359808 567384 359836
rect 548024 359796 548030 359808
rect 567378 359796 567384 359808
rect 567436 359796 567442 359848
rect 425790 359456 425796 359508
rect 425848 359496 425854 359508
rect 427262 359496 427268 359508
rect 425848 359468 427268 359496
rect 425848 359456 425854 359468
rect 427262 359456 427268 359468
rect 427320 359456 427326 359508
rect 444006 358912 444012 358964
rect 444064 358952 444070 358964
rect 447318 358952 447324 358964
rect 444064 358924 447324 358952
rect 444064 358912 444070 358924
rect 447318 358912 447324 358924
rect 447376 358912 447382 358964
rect 439774 358844 439780 358896
rect 439832 358884 439838 358896
rect 447134 358884 447140 358896
rect 439832 358856 447140 358884
rect 439832 358844 439838 358856
rect 447134 358844 447140 358856
rect 447192 358844 447198 358896
rect 433978 358776 433984 358828
rect 434036 358816 434042 358828
rect 447226 358816 447232 358828
rect 434036 358788 447232 358816
rect 434036 358776 434042 358788
rect 447226 358776 447232 358788
rect 447284 358776 447290 358828
rect 513006 358776 513012 358828
rect 513064 358816 513070 358828
rect 523126 358816 523132 358828
rect 513064 358788 523132 358816
rect 513064 358776 513070 358788
rect 523126 358776 523132 358788
rect 523184 358776 523190 358828
rect 425698 358708 425704 358760
rect 425756 358748 425762 358760
rect 427170 358748 427176 358760
rect 425756 358720 427176 358748
rect 425756 358708 425762 358720
rect 427170 358708 427176 358720
rect 427228 358708 427234 358760
rect 551922 358708 551928 358760
rect 551980 358748 551986 358760
rect 559098 358748 559104 358760
rect 551980 358720 559104 358748
rect 551980 358708 551986 358720
rect 559098 358708 559104 358720
rect 559156 358708 559162 358760
rect 424318 358640 424324 358692
rect 424376 358680 424382 358692
rect 426434 358680 426440 358692
rect 424376 358652 426440 358680
rect 424376 358640 424382 358652
rect 426434 358640 426440 358652
rect 426492 358640 426498 358692
rect 514846 358640 514852 358692
rect 514904 358680 514910 358692
rect 552474 358680 552480 358692
rect 514904 358652 552480 358680
rect 514904 358640 514910 358652
rect 552474 358640 552480 358652
rect 552532 358640 552538 358692
rect 548058 358572 548064 358624
rect 548116 358612 548122 358624
rect 562410 358612 562416 358624
rect 548116 358584 562416 358612
rect 548116 358572 548122 358584
rect 562410 358572 562416 358584
rect 562468 358572 562474 358624
rect 549162 358504 549168 358556
rect 549220 358544 549226 358556
rect 560754 358544 560760 358556
rect 549220 358516 560760 358544
rect 549220 358504 549226 358516
rect 560754 358504 560760 358516
rect 560812 358504 560818 358556
rect 518894 358436 518900 358488
rect 518952 358476 518958 358488
rect 565722 358476 565728 358488
rect 518952 358448 565728 358476
rect 518952 358436 518958 358448
rect 565722 358436 565728 358448
rect 565780 358436 565786 358488
rect 551462 358368 551468 358420
rect 551520 358408 551526 358420
rect 564066 358408 564072 358420
rect 551520 358380 564072 358408
rect 551520 358368 551526 358380
rect 564066 358368 564072 358380
rect 564124 358368 564130 358420
rect 513006 357960 513012 358012
rect 513064 358000 513070 358012
rect 520366 358000 520372 358012
rect 513064 357972 520372 358000
rect 513064 357960 513070 357972
rect 520366 357960 520372 357972
rect 520424 357960 520430 358012
rect 512086 357688 512092 357740
rect 512144 357728 512150 357740
rect 514938 357728 514944 357740
rect 512144 357700 514944 357728
rect 512144 357688 512150 357700
rect 514938 357688 514944 357700
rect 514996 357688 515002 357740
rect 440970 357484 440976 357536
rect 441028 357524 441034 357536
rect 447226 357524 447232 357536
rect 441028 357496 447232 357524
rect 441028 357484 441034 357496
rect 447226 357484 447232 357496
rect 447284 357484 447290 357536
rect 435450 357416 435456 357468
rect 435508 357456 435514 357468
rect 447134 357456 447140 357468
rect 435508 357428 447140 357456
rect 435508 357416 435514 357428
rect 447134 357416 447140 357428
rect 447192 357416 447198 357468
rect 513282 357416 513288 357468
rect 513340 357456 513346 357468
rect 523218 357456 523224 357468
rect 513340 357428 523224 357456
rect 513340 357416 513346 357428
rect 523218 357416 523224 357428
rect 523276 357416 523282 357468
rect 443730 356192 443736 356244
rect 443788 356232 443794 356244
rect 447318 356232 447324 356244
rect 443788 356204 447324 356232
rect 443788 356192 443794 356204
rect 447318 356192 447324 356204
rect 447376 356192 447382 356244
rect 512178 356192 512184 356244
rect 512236 356232 512242 356244
rect 514846 356232 514852 356244
rect 512236 356204 514852 356232
rect 512236 356192 512242 356204
rect 514846 356192 514852 356204
rect 514904 356192 514910 356244
rect 439682 356124 439688 356176
rect 439740 356164 439746 356176
rect 447134 356164 447140 356176
rect 439740 356136 447140 356164
rect 439740 356124 439746 356136
rect 447134 356124 447140 356136
rect 447192 356124 447198 356176
rect 436922 356056 436928 356108
rect 436980 356096 436986 356108
rect 447226 356096 447232 356108
rect 436980 356068 447232 356096
rect 436980 356056 436986 356068
rect 447226 356056 447232 356068
rect 447284 356056 447290 356108
rect 512638 356056 512644 356108
rect 512696 356096 512702 356108
rect 516226 356096 516232 356108
rect 512696 356068 516232 356096
rect 512696 356056 512702 356068
rect 516226 356056 516232 356068
rect 516284 356056 516290 356108
rect 512730 354968 512736 355020
rect 512788 355008 512794 355020
rect 517514 355008 517520 355020
rect 512788 354980 517520 355008
rect 512788 354968 512794 354980
rect 517514 354968 517520 354980
rect 517572 354968 517578 355020
rect 426434 354696 426440 354748
rect 426492 354736 426498 354748
rect 426492 354708 427860 354736
rect 426492 354696 426498 354708
rect 427832 354668 427860 354708
rect 513282 354696 513288 354748
rect 513340 354736 513346 354748
rect 523310 354736 523316 354748
rect 513340 354708 523316 354736
rect 513340 354696 513346 354708
rect 523310 354696 523316 354708
rect 523368 354696 523374 354748
rect 430574 354668 430580 354680
rect 427832 354640 430580 354668
rect 430574 354628 430580 354640
rect 430632 354628 430638 354680
rect 432598 354220 432604 354272
rect 432656 354260 432662 354272
rect 434070 354260 434076 354272
rect 432656 354232 434076 354260
rect 432656 354220 432662 354232
rect 434070 354220 434076 354232
rect 434128 354220 434134 354272
rect 512546 354084 512552 354136
rect 512604 354124 512610 354136
rect 517606 354124 517612 354136
rect 512604 354096 517612 354124
rect 512604 354084 512610 354096
rect 517606 354084 517612 354096
rect 517664 354084 517670 354136
rect 411898 353948 411904 354000
rect 411956 353988 411962 354000
rect 423582 353988 423588 354000
rect 411956 353960 423588 353988
rect 411956 353948 411962 353960
rect 423582 353948 423588 353960
rect 423640 353948 423646 354000
rect 513098 353268 513104 353320
rect 513156 353308 513162 353320
rect 518894 353308 518900 353320
rect 513156 353280 518900 353308
rect 513156 353268 513162 353280
rect 518894 353268 518900 353280
rect 518952 353268 518958 353320
rect 512270 352248 512276 352300
rect 512328 352288 512334 352300
rect 520642 352288 520648 352300
rect 512328 352260 520648 352288
rect 512328 352248 512334 352260
rect 520642 352248 520648 352260
rect 520700 352248 520706 352300
rect 513282 351908 513288 351960
rect 513340 351948 513346 351960
rect 523402 351948 523408 351960
rect 513340 351920 523408 351948
rect 513340 351908 513346 351920
rect 523402 351908 523408 351920
rect 523460 351908 523466 351960
rect 430574 351840 430580 351892
rect 430632 351880 430638 351892
rect 434162 351880 434168 351892
rect 430632 351852 434168 351880
rect 430632 351840 430638 351852
rect 434162 351840 434168 351852
rect 434220 351840 434226 351892
rect 512638 351704 512644 351756
rect 512696 351744 512702 351756
rect 516318 351744 516324 351756
rect 512696 351716 516324 351744
rect 512696 351704 512702 351716
rect 516318 351704 516324 351716
rect 516376 351704 516382 351756
rect 513282 351024 513288 351076
rect 513340 351064 513346 351076
rect 520458 351064 520464 351076
rect 513340 351036 520464 351064
rect 513340 351024 513346 351036
rect 520458 351024 520464 351036
rect 520516 351024 520522 351076
rect 423582 350888 423588 350940
rect 423640 350928 423646 350940
rect 431218 350928 431224 350940
rect 423640 350900 431224 350928
rect 423640 350888 423646 350900
rect 431218 350888 431224 350900
rect 431276 350888 431282 350940
rect 512638 350888 512644 350940
rect 512696 350928 512702 350940
rect 516962 350928 516968 350940
rect 512696 350900 516968 350928
rect 512696 350888 512702 350900
rect 516962 350888 516968 350900
rect 517020 350888 517026 350940
rect 422938 350820 422944 350872
rect 422996 350860 423002 350872
rect 425698 350860 425704 350872
rect 422996 350832 425704 350860
rect 422996 350820 423002 350832
rect 425698 350820 425704 350832
rect 425756 350820 425762 350872
rect 513282 350548 513288 350600
rect 513340 350588 513346 350600
rect 517698 350588 517704 350600
rect 513340 350560 517704 350588
rect 513340 350548 513346 350560
rect 517698 350548 517704 350560
rect 517756 350548 517762 350600
rect 421558 350480 421564 350532
rect 421616 350520 421622 350532
rect 423582 350520 423588 350532
rect 421616 350492 423588 350520
rect 421616 350480 421622 350492
rect 423582 350480 423588 350492
rect 423640 350480 423646 350532
rect 424962 350480 424968 350532
rect 425020 350520 425026 350532
rect 447318 350520 447324 350532
rect 425020 350492 447324 350520
rect 425020 350480 425026 350492
rect 447318 350480 447324 350492
rect 447376 350480 447382 350532
rect 431310 350412 431316 350464
rect 431368 350452 431374 350464
rect 433702 350452 433708 350464
rect 431368 350424 433708 350452
rect 431368 350412 431374 350424
rect 433702 350412 433708 350424
rect 433760 350412 433766 350464
rect 447134 350452 447140 350464
rect 436756 350424 447140 350452
rect 426342 350344 426348 350396
rect 426400 350384 426406 350396
rect 436756 350384 436784 350424
rect 447134 350412 447140 350424
rect 447192 350412 447198 350464
rect 447226 350384 447232 350396
rect 426400 350356 436784 350384
rect 441586 350356 447232 350384
rect 426400 350344 426406 350356
rect 427262 350276 427268 350328
rect 427320 350316 427326 350328
rect 428550 350316 428556 350328
rect 427320 350288 428556 350316
rect 427320 350276 427326 350288
rect 428550 350276 428556 350288
rect 428608 350276 428614 350328
rect 426250 350208 426256 350260
rect 426308 350248 426314 350260
rect 441586 350248 441614 350356
rect 447226 350344 447232 350356
rect 447284 350344 447290 350396
rect 426308 350220 441614 350248
rect 426308 350208 426314 350220
rect 513282 349528 513288 349580
rect 513340 349568 513346 349580
rect 518986 349568 518992 349580
rect 513340 349540 518992 349568
rect 513340 349528 513346 349540
rect 518986 349528 518992 349540
rect 519044 349528 519050 349580
rect 512822 349256 512828 349308
rect 512880 349296 512886 349308
rect 520550 349296 520556 349308
rect 512880 349268 520556 349296
rect 512880 349256 512886 349268
rect 520550 349256 520556 349268
rect 520608 349256 520614 349308
rect 512178 349188 512184 349240
rect 512236 349228 512242 349240
rect 515030 349228 515036 349240
rect 512236 349200 515036 349228
rect 512236 349188 512242 349200
rect 515030 349188 515036 349200
rect 515088 349188 515094 349240
rect 427170 349052 427176 349104
rect 427228 349092 427234 349104
rect 428458 349092 428464 349104
rect 427228 349064 428464 349092
rect 427228 349052 427234 349064
rect 428458 349052 428464 349064
rect 428516 349052 428522 349104
rect 447134 349092 447140 349104
rect 431926 349064 447140 349092
rect 423306 348984 423312 349036
rect 423364 349024 423370 349036
rect 431926 349024 431954 349064
rect 447134 349052 447140 349064
rect 447192 349052 447198 349104
rect 423364 348996 431954 349024
rect 423364 348984 423370 348996
rect 443638 348984 443644 349036
rect 443696 349024 443702 349036
rect 447226 349024 447232 349036
rect 443696 348996 447232 349024
rect 443696 348984 443702 348996
rect 447226 348984 447232 348996
rect 447284 348984 447290 349036
rect 513282 348168 513288 348220
rect 513340 348208 513346 348220
rect 520734 348208 520740 348220
rect 513340 348180 520740 348208
rect 513340 348168 513346 348180
rect 520734 348168 520740 348180
rect 520792 348168 520798 348220
rect 513190 347760 513196 347812
rect 513248 347800 513254 347812
rect 521654 347800 521660 347812
rect 513248 347772 521660 347800
rect 513248 347760 513254 347772
rect 521654 347760 521660 347772
rect 521712 347760 521718 347812
rect 422110 347692 422116 347744
rect 422168 347732 422174 347744
rect 447226 347732 447232 347744
rect 422168 347704 447232 347732
rect 422168 347692 422174 347704
rect 447226 347692 447232 347704
rect 447284 347692 447290 347744
rect 422202 347624 422208 347676
rect 422260 347664 422266 347676
rect 447318 347664 447324 347676
rect 422260 347636 447324 347664
rect 422260 347624 422266 347636
rect 447318 347624 447324 347636
rect 447376 347624 447382 347676
rect 428550 347556 428556 347608
rect 428608 347596 428614 347608
rect 429562 347596 429568 347608
rect 428608 347568 429568 347596
rect 428608 347556 428614 347568
rect 429562 347556 429568 347568
rect 429620 347556 429626 347608
rect 447134 347596 447140 347608
rect 431926 347568 447140 347596
rect 423490 347488 423496 347540
rect 423548 347528 423554 347540
rect 431926 347528 431954 347568
rect 447134 347556 447140 347568
rect 447192 347556 447198 347608
rect 423548 347500 431954 347528
rect 423548 347488 423554 347500
rect 512822 346672 512828 346724
rect 512880 346712 512886 346724
rect 519078 346712 519084 346724
rect 512880 346684 519084 346712
rect 512880 346672 512886 346684
rect 519078 346672 519084 346684
rect 519136 346672 519142 346724
rect 513006 346536 513012 346588
rect 513064 346576 513070 346588
rect 521746 346576 521752 346588
rect 513064 346548 521752 346576
rect 513064 346536 513070 346548
rect 521746 346536 521752 346548
rect 521804 346536 521810 346588
rect 427078 346400 427084 346452
rect 427136 346440 427142 346452
rect 427136 346412 429240 346440
rect 427136 346400 427142 346412
rect 429212 346372 429240 346412
rect 512178 346400 512184 346452
rect 512236 346440 512242 346452
rect 513742 346440 513748 346452
rect 512236 346412 513748 346440
rect 512236 346400 512242 346412
rect 513742 346400 513748 346412
rect 513800 346400 513806 346452
rect 430574 346372 430580 346384
rect 429212 346344 430580 346372
rect 430574 346332 430580 346344
rect 430632 346332 430638 346384
rect 433702 346332 433708 346384
rect 433760 346372 433766 346384
rect 435634 346372 435640 346384
rect 433760 346344 435640 346372
rect 433760 346332 433766 346344
rect 435634 346332 435640 346344
rect 435692 346332 435698 346384
rect 513190 345176 513196 345228
rect 513248 345216 513254 345228
rect 519170 345216 519176 345228
rect 513248 345188 519176 345216
rect 513248 345176 513254 345188
rect 519170 345176 519176 345188
rect 519228 345176 519234 345228
rect 407022 345040 407028 345092
rect 407080 345080 407086 345092
rect 447134 345080 447140 345092
rect 407080 345052 447140 345080
rect 407080 345040 407086 345052
rect 447134 345040 447140 345052
rect 447192 345040 447198 345092
rect 513282 345040 513288 345092
rect 513340 345080 513346 345092
rect 521838 345080 521844 345092
rect 513340 345052 521844 345080
rect 513340 345040 513346 345052
rect 521838 345040 521844 345052
rect 521896 345040 521902 345092
rect 446214 344428 446220 344480
rect 446272 344468 446278 344480
rect 447870 344468 447876 344480
rect 446272 344440 447876 344468
rect 446272 344428 446278 344440
rect 447870 344428 447876 344440
rect 447928 344428 447934 344480
rect 513282 344360 513288 344412
rect 513340 344400 513346 344412
rect 520826 344400 520832 344412
rect 513340 344372 520832 344400
rect 513340 344360 513346 344372
rect 520826 344360 520832 344372
rect 520884 344360 520890 344412
rect 423674 344156 423680 344208
rect 423732 344196 423738 344208
rect 426342 344196 426348 344208
rect 423732 344168 426348 344196
rect 423732 344156 423738 344168
rect 426342 344156 426348 344168
rect 426400 344156 426406 344208
rect 512270 343952 512276 344004
rect 512328 343992 512334 344004
rect 515122 343992 515128 344004
rect 512328 343964 515128 343992
rect 512328 343952 512334 343964
rect 515122 343952 515128 343964
rect 515180 343952 515186 344004
rect 425698 343884 425704 343936
rect 425756 343924 425762 343936
rect 427722 343924 427728 343936
rect 425756 343896 427728 343924
rect 425756 343884 425762 343896
rect 427722 343884 427728 343896
rect 427780 343884 427786 343936
rect 512822 343748 512828 343800
rect 512880 343788 512886 343800
rect 521930 343788 521936 343800
rect 512880 343760 521936 343788
rect 512880 343748 512886 343760
rect 521930 343748 521936 343760
rect 521988 343748 521994 343800
rect 382274 343680 382280 343732
rect 382332 343720 382338 343732
rect 386322 343720 386328 343732
rect 382332 343692 386328 343720
rect 382332 343680 382338 343692
rect 386322 343680 386328 343692
rect 386380 343680 386386 343732
rect 382918 343544 382924 343596
rect 382976 343584 382982 343596
rect 447134 343584 447140 343596
rect 382976 343556 447140 343584
rect 382976 343544 382982 343556
rect 447134 343544 447140 343556
rect 447192 343544 447198 343596
rect 426342 343476 426348 343528
rect 426400 343516 426406 343528
rect 429102 343516 429108 343528
rect 426400 343488 429108 343516
rect 426400 343476 426406 343488
rect 429102 343476 429108 343488
rect 429160 343476 429166 343528
rect 411990 342864 411996 342916
rect 412048 342904 412054 342916
rect 418154 342904 418160 342916
rect 412048 342876 418160 342904
rect 412048 342864 412054 342876
rect 418154 342864 418160 342876
rect 418212 342864 418218 342916
rect 512362 342864 512368 342916
rect 512420 342904 512426 342916
rect 515214 342904 515220 342916
rect 512420 342876 515220 342904
rect 512420 342864 512426 342876
rect 515214 342864 515220 342876
rect 515272 342864 515278 342916
rect 513282 342320 513288 342372
rect 513340 342360 513346 342372
rect 519262 342360 519268 342372
rect 513340 342332 519268 342360
rect 513340 342320 513346 342332
rect 519262 342320 519268 342332
rect 519320 342320 519326 342372
rect 428458 342252 428464 342304
rect 428516 342292 428522 342304
rect 428516 342264 431954 342292
rect 428516 342252 428522 342264
rect 431926 342224 431954 342264
rect 434254 342224 434260 342236
rect 431926 342196 434260 342224
rect 434254 342184 434260 342196
rect 434312 342184 434318 342236
rect 386322 341504 386328 341556
rect 386380 341544 386386 341556
rect 402146 341544 402152 341556
rect 386380 341516 402152 341544
rect 386380 341504 386386 341516
rect 402146 341504 402152 341516
rect 402204 341504 402210 341556
rect 512270 341368 512276 341420
rect 512328 341408 512334 341420
rect 513834 341408 513840 341420
rect 512328 341380 513840 341408
rect 512328 341368 512334 341380
rect 513834 341368 513840 341380
rect 513892 341368 513898 341420
rect 512270 341232 512276 341284
rect 512328 341272 512334 341284
rect 519446 341272 519452 341284
rect 512328 341244 519452 341272
rect 512328 341232 512334 341244
rect 519446 341232 519452 341244
rect 519504 341232 519510 341284
rect 435634 341164 435640 341216
rect 435692 341204 435698 341216
rect 438118 341204 438124 341216
rect 435692 341176 438124 341204
rect 435692 341164 435698 341176
rect 438118 341164 438124 341176
rect 438176 341164 438182 341216
rect 513282 340892 513288 340944
rect 513340 340932 513346 340944
rect 522022 340932 522028 340944
rect 513340 340904 522028 340932
rect 513340 340892 513346 340904
rect 522022 340892 522028 340904
rect 522080 340892 522086 340944
rect 427722 340824 427728 340876
rect 427780 340864 427786 340876
rect 430666 340864 430672 340876
rect 427780 340836 430672 340864
rect 427780 340824 427786 340836
rect 430666 340824 430672 340836
rect 430724 340824 430730 340876
rect 430574 340756 430580 340808
rect 430632 340796 430638 340808
rect 432966 340796 432972 340808
rect 430632 340768 432972 340796
rect 430632 340756 430638 340768
rect 432966 340756 432972 340768
rect 433024 340756 433030 340808
rect 418154 340212 418160 340264
rect 418212 340252 418218 340264
rect 432782 340252 432788 340264
rect 418212 340224 432788 340252
rect 418212 340212 418218 340224
rect 432782 340212 432788 340224
rect 432840 340212 432846 340264
rect 413646 340144 413652 340196
rect 413704 340184 413710 340196
rect 449342 340184 449348 340196
rect 413704 340156 449348 340184
rect 413704 340144 413710 340156
rect 449342 340144 449348 340156
rect 449400 340144 449406 340196
rect 513282 339872 513288 339924
rect 513340 339912 513346 339924
rect 517790 339912 517796 339924
rect 513340 339884 517796 339912
rect 513340 339872 513346 339884
rect 517790 339872 517796 339884
rect 517848 339872 517854 339924
rect 513006 339736 513012 339788
rect 513064 339776 513070 339788
rect 518066 339776 518072 339788
rect 513064 339748 518072 339776
rect 513064 339736 513070 339748
rect 518066 339736 518072 339748
rect 518124 339736 518130 339788
rect 512362 339668 512368 339720
rect 512420 339708 512426 339720
rect 515306 339708 515312 339720
rect 512420 339680 515312 339708
rect 512420 339668 512426 339680
rect 515306 339668 515312 339680
rect 515364 339668 515370 339720
rect 512362 339464 512368 339516
rect 512420 339504 512426 339516
rect 514110 339504 514116 339516
rect 512420 339476 514116 339504
rect 512420 339464 512426 339476
rect 514110 339464 514116 339476
rect 514168 339464 514174 339516
rect 429562 339396 429568 339448
rect 429620 339436 429626 339448
rect 433242 339436 433248 339448
rect 429620 339408 433248 339436
rect 429620 339396 429626 339408
rect 433242 339396 433248 339408
rect 433300 339396 433306 339448
rect 449986 339396 449992 339448
rect 450044 339436 450050 339448
rect 450354 339436 450360 339448
rect 450044 339408 450360 339436
rect 450044 339396 450050 339408
rect 450354 339396 450360 339408
rect 450412 339396 450418 339448
rect 450078 339328 450084 339380
rect 450136 339368 450142 339380
rect 450446 339368 450452 339380
rect 450136 339340 450452 339368
rect 450136 339328 450142 339340
rect 450446 339328 450452 339340
rect 450504 339328 450510 339380
rect 449618 339260 449624 339312
rect 449676 339300 449682 339312
rect 450630 339300 450636 339312
rect 449676 339272 450636 339300
rect 449676 339260 449682 339272
rect 450630 339260 450636 339272
rect 450688 339260 450694 339312
rect 447870 339056 447876 339108
rect 447928 339096 447934 339108
rect 450078 339096 450084 339108
rect 447928 339068 450084 339096
rect 447928 339056 447934 339068
rect 450078 339056 450084 339068
rect 450136 339056 450142 339108
rect 450078 338920 450084 338972
rect 450136 338960 450142 338972
rect 450538 338960 450544 338972
rect 450136 338932 450544 338960
rect 450136 338920 450142 338932
rect 450538 338920 450544 338932
rect 450596 338920 450602 338972
rect 383102 338512 383108 338564
rect 383160 338552 383166 338564
rect 447134 338552 447140 338564
rect 383160 338524 447140 338552
rect 383160 338512 383166 338524
rect 447134 338512 447140 338524
rect 447192 338512 447198 338564
rect 429838 338444 429844 338496
rect 429896 338484 429902 338496
rect 450354 338484 450360 338496
rect 429896 338456 450360 338484
rect 429896 338444 429902 338456
rect 450354 338444 450360 338456
rect 450412 338444 450418 338496
rect 425882 338376 425888 338428
rect 425940 338416 425946 338428
rect 450446 338416 450452 338428
rect 425940 338388 450452 338416
rect 425940 338376 425946 338388
rect 450446 338376 450452 338388
rect 450504 338376 450510 338428
rect 513190 338376 513196 338428
rect 513248 338416 513254 338428
rect 517882 338416 517888 338428
rect 513248 338388 517888 338416
rect 513248 338376 513254 338388
rect 517882 338376 517888 338388
rect 517940 338376 517946 338428
rect 417970 338308 417976 338360
rect 418028 338348 418034 338360
rect 450170 338348 450176 338360
rect 418028 338320 450176 338348
rect 418028 338308 418034 338320
rect 450170 338308 450176 338320
rect 450228 338308 450234 338360
rect 414014 338240 414020 338292
rect 414072 338280 414078 338292
rect 450078 338280 450084 338292
rect 414072 338252 450084 338280
rect 414072 338240 414078 338252
rect 450078 338240 450084 338252
rect 450136 338240 450142 338292
rect 512546 338240 512552 338292
rect 512604 338280 512610 338292
rect 515582 338280 515588 338292
rect 512604 338252 515588 338280
rect 512604 338240 512610 338252
rect 515582 338240 515588 338252
rect 515640 338240 515646 338292
rect 410058 338172 410064 338224
rect 410116 338212 410122 338224
rect 449618 338212 449624 338224
rect 410116 338184 449624 338212
rect 410116 338172 410122 338184
rect 449618 338172 449624 338184
rect 449676 338172 449682 338224
rect 513282 338104 513288 338156
rect 513340 338144 513346 338156
rect 522114 338144 522120 338156
rect 513340 338116 522120 338144
rect 513340 338104 513346 338116
rect 522114 338104 522120 338116
rect 522172 338104 522178 338156
rect 434162 338036 434168 338088
rect 434220 338076 434226 338088
rect 437014 338076 437020 338088
rect 434220 338048 437020 338076
rect 434220 338036 434226 338048
rect 437014 338036 437020 338048
rect 437072 338036 437078 338088
rect 420178 337696 420184 337748
rect 420236 337736 420242 337748
rect 439958 337736 439964 337748
rect 420236 337708 439964 337736
rect 420236 337696 420242 337708
rect 439958 337696 439964 337708
rect 440016 337696 440022 337748
rect 418890 337628 418896 337680
rect 418948 337668 418954 337680
rect 442350 337668 442356 337680
rect 418948 337640 442356 337668
rect 418948 337628 418954 337640
rect 442350 337628 442356 337640
rect 442408 337628 442414 337680
rect 416038 337560 416044 337612
rect 416096 337600 416102 337612
rect 440050 337600 440056 337612
rect 416096 337572 440056 337600
rect 416096 337560 416102 337572
rect 440050 337560 440056 337572
rect 440108 337560 440114 337612
rect 418982 337492 418988 337544
rect 419040 337532 419046 337544
rect 445570 337532 445576 337544
rect 419040 337504 445576 337532
rect 419040 337492 419046 337504
rect 445570 337492 445576 337504
rect 445628 337492 445634 337544
rect 413278 337424 413284 337476
rect 413336 337464 413342 337476
rect 439866 337464 439872 337476
rect 413336 337436 439872 337464
rect 413336 337424 413342 337436
rect 439866 337424 439872 337436
rect 439924 337424 439930 337476
rect 418798 337356 418804 337408
rect 418856 337396 418862 337408
rect 449250 337396 449256 337408
rect 418856 337368 449256 337396
rect 418856 337356 418862 337368
rect 449250 337356 449256 337368
rect 449308 337356 449314 337408
rect 512914 337016 512920 337068
rect 512972 337056 512978 337068
rect 516594 337056 516600 337068
rect 512972 337028 516600 337056
rect 512972 337016 512978 337028
rect 516594 337016 516600 337028
rect 516652 337016 516658 337068
rect 430666 336880 430672 336932
rect 430724 336920 430730 336932
rect 432874 336920 432880 336932
rect 430724 336892 432880 336920
rect 430724 336880 430730 336892
rect 432874 336880 432880 336892
rect 432932 336880 432938 336932
rect 382918 336812 382924 336864
rect 382976 336852 382982 336864
rect 447134 336852 447140 336864
rect 382976 336824 447140 336852
rect 382976 336812 382982 336824
rect 447134 336812 447140 336824
rect 447192 336812 447198 336864
rect 383010 336744 383016 336796
rect 383068 336784 383074 336796
rect 447226 336784 447232 336796
rect 383068 336756 447232 336784
rect 383068 336744 383074 336756
rect 447226 336744 447232 336756
rect 447284 336744 447290 336796
rect 513006 336744 513012 336796
rect 513064 336784 513070 336796
rect 522206 336784 522212 336796
rect 513064 336756 522212 336784
rect 513064 336744 513070 336756
rect 522206 336744 522212 336756
rect 522264 336744 522270 336796
rect 402238 336676 402244 336728
rect 402296 336716 402302 336728
rect 442902 336716 442908 336728
rect 402296 336688 442908 336716
rect 402296 336676 402302 336688
rect 442902 336676 442908 336688
rect 442960 336716 442966 336728
rect 447870 336716 447876 336728
rect 442960 336688 447876 336716
rect 442960 336676 442966 336688
rect 447870 336676 447876 336688
rect 447928 336676 447934 336728
rect 429194 336608 429200 336660
rect 429252 336648 429258 336660
rect 431862 336648 431868 336660
rect 429252 336620 431868 336648
rect 429252 336608 429258 336620
rect 431862 336608 431868 336620
rect 431920 336608 431926 336660
rect 513190 335928 513196 335980
rect 513248 335968 513254 335980
rect 517974 335968 517980 335980
rect 513248 335940 517980 335968
rect 513248 335928 513254 335940
rect 517974 335928 517980 335940
rect 518032 335928 518038 335980
rect 442258 335792 442264 335844
rect 442316 335832 442322 335844
rect 447226 335832 447232 335844
rect 442316 335804 447232 335832
rect 442316 335792 442322 335804
rect 447226 335792 447232 335804
rect 447284 335792 447290 335844
rect 443914 335724 443920 335776
rect 443972 335764 443978 335776
rect 447134 335764 447140 335776
rect 443972 335736 447140 335764
rect 443972 335724 443978 335736
rect 447134 335724 447140 335736
rect 447192 335724 447198 335776
rect 513282 335656 513288 335708
rect 513340 335696 513346 335708
rect 519354 335696 519360 335708
rect 513340 335668 519360 335696
rect 513340 335656 513346 335668
rect 519354 335656 519360 335668
rect 519412 335656 519418 335708
rect 512730 335384 512736 335436
rect 512788 335424 512794 335436
rect 516134 335424 516140 335436
rect 512788 335396 516140 335424
rect 512788 335384 512794 335396
rect 516134 335384 516140 335396
rect 516192 335384 516198 335436
rect 431862 335044 431868 335096
rect 431920 335084 431926 335096
rect 434622 335084 434628 335096
rect 431920 335056 434628 335084
rect 431920 335044 431926 335056
rect 434622 335044 434628 335056
rect 434680 335044 434686 335096
rect 439590 334568 439596 334620
rect 439648 334608 439654 334620
rect 447318 334608 447324 334620
rect 439648 334580 447324 334608
rect 439648 334568 439654 334580
rect 447318 334568 447324 334580
rect 447376 334568 447382 334620
rect 434070 334500 434076 334552
rect 434128 334540 434134 334552
rect 435726 334540 435732 334552
rect 434128 334512 435732 334540
rect 434128 334500 434134 334512
rect 435726 334500 435732 334512
rect 435784 334500 435790 334552
rect 513006 334160 513012 334212
rect 513064 334200 513070 334212
rect 516686 334200 516692 334212
rect 513064 334172 516692 334200
rect 513064 334160 513070 334172
rect 516686 334160 516692 334172
rect 516744 334160 516750 334212
rect 433426 334024 433432 334076
rect 433484 334064 433490 334076
rect 433484 334036 434852 334064
rect 433484 334024 433490 334036
rect 434254 333956 434260 334008
rect 434312 333996 434318 334008
rect 434824 333996 434852 334036
rect 435358 334024 435364 334076
rect 435416 334064 435422 334076
rect 435416 334036 436600 334064
rect 435416 334024 435422 334036
rect 436572 333996 436600 334036
rect 436830 334024 436836 334076
rect 436888 334064 436894 334076
rect 447226 334064 447232 334076
rect 436888 334036 447232 334064
rect 436888 334024 436894 334036
rect 447226 334024 447232 334036
rect 447284 334024 447290 334076
rect 512822 334024 512828 334076
rect 512880 334064 512886 334076
rect 516410 334064 516416 334076
rect 512880 334036 516416 334064
rect 512880 334024 512886 334036
rect 516410 334024 516416 334036
rect 516468 334024 516474 334076
rect 447134 333996 447140 334008
rect 434312 333968 434760 333996
rect 434824 333968 436508 333996
rect 436572 333968 447140 333996
rect 434312 333956 434318 333968
rect 434732 333928 434760 333968
rect 436370 333928 436376 333940
rect 434732 333900 436376 333928
rect 436370 333888 436376 333900
rect 436428 333888 436434 333940
rect 436480 333928 436508 333968
rect 447134 333956 447140 333968
rect 447192 333956 447198 334008
rect 437382 333928 437388 333940
rect 436480 333900 437388 333928
rect 437382 333888 437388 333900
rect 437440 333888 437446 333940
rect 512914 332800 512920 332852
rect 512972 332840 512978 332852
rect 516502 332840 516508 332852
rect 512972 332812 516508 332840
rect 512972 332800 512978 332812
rect 516502 332800 516508 332812
rect 516560 332800 516566 332852
rect 513282 332732 513288 332784
rect 513340 332772 513346 332784
rect 519630 332772 519636 332784
rect 513340 332744 519636 332772
rect 513340 332732 513346 332744
rect 519630 332732 519636 332744
rect 519688 332732 519694 332784
rect 440878 332664 440884 332716
rect 440936 332704 440942 332716
rect 447134 332704 447140 332716
rect 440936 332676 447140 332704
rect 440936 332664 440942 332676
rect 447134 332664 447140 332676
rect 447192 332664 447198 332716
rect 432598 332596 432604 332648
rect 432656 332636 432662 332648
rect 447226 332636 447232 332648
rect 432656 332608 447232 332636
rect 432656 332596 432662 332608
rect 447226 332596 447232 332608
rect 447284 332596 447290 332648
rect 512822 332596 512828 332648
rect 512880 332636 512886 332648
rect 523494 332636 523500 332648
rect 512880 332608 523500 332636
rect 512880 332596 512886 332608
rect 523494 332596 523500 332608
rect 523552 332596 523558 332648
rect 433426 331984 433432 332036
rect 433484 332024 433490 332036
rect 439774 332024 439780 332036
rect 433484 331996 439780 332024
rect 433484 331984 433490 331996
rect 439774 331984 439780 331996
rect 439832 331984 439838 332036
rect 434438 331848 434444 331900
rect 434496 331888 434502 331900
rect 444006 331888 444012 331900
rect 434496 331860 444012 331888
rect 434496 331848 434502 331860
rect 444006 331848 444012 331860
rect 444064 331848 444070 331900
rect 513282 331440 513288 331492
rect 513340 331480 513346 331492
rect 519722 331480 519728 331492
rect 513340 331452 519728 331480
rect 513340 331440 513346 331452
rect 519722 331440 519728 331452
rect 519780 331440 519786 331492
rect 443822 331372 443828 331424
rect 443880 331412 443886 331424
rect 447410 331412 447416 331424
rect 443880 331384 447416 331412
rect 443880 331372 443886 331384
rect 447410 331372 447416 331384
rect 447468 331372 447474 331424
rect 443638 331304 443644 331356
rect 443696 331344 443702 331356
rect 447226 331344 447232 331356
rect 443696 331316 447232 331344
rect 443696 331304 443702 331316
rect 447226 331304 447232 331316
rect 447284 331304 447290 331356
rect 432690 331236 432696 331288
rect 432748 331276 432754 331288
rect 432748 331248 433380 331276
rect 432748 331236 432754 331248
rect 433352 331208 433380 331248
rect 439498 331236 439504 331288
rect 439556 331276 439562 331288
rect 447134 331276 447140 331288
rect 439556 331248 447140 331276
rect 439556 331236 439562 331248
rect 447134 331236 447140 331248
rect 447192 331236 447198 331288
rect 512822 331236 512828 331288
rect 512880 331276 512886 331288
rect 516870 331276 516876 331288
rect 512880 331248 516876 331276
rect 512880 331236 512886 331248
rect 516870 331236 516876 331248
rect 516928 331236 516934 331288
rect 435082 331208 435088 331220
rect 433352 331180 435088 331208
rect 435082 331168 435088 331180
rect 435140 331168 435146 331220
rect 436370 331100 436376 331152
rect 436428 331140 436434 331152
rect 438302 331140 438308 331152
rect 436428 331112 438308 331140
rect 436428 331100 436434 331112
rect 438302 331100 438308 331112
rect 438360 331100 438366 331152
rect 432966 330556 432972 330608
rect 433024 330596 433030 330608
rect 436002 330596 436008 330608
rect 433024 330568 436008 330596
rect 433024 330556 433030 330568
rect 436002 330556 436008 330568
rect 436060 330556 436066 330608
rect 436738 330488 436744 330540
rect 436796 330528 436802 330540
rect 447318 330528 447324 330540
rect 436796 330500 447324 330528
rect 436796 330488 436802 330500
rect 447318 330488 447324 330500
rect 447376 330488 447382 330540
rect 434714 329740 434720 329792
rect 434772 329780 434778 329792
rect 438210 329780 438216 329792
rect 434772 329752 438216 329780
rect 434772 329740 434778 329752
rect 438210 329740 438216 329752
rect 438268 329740 438274 329792
rect 446306 329604 446312 329656
rect 446364 329644 446370 329656
rect 448238 329644 448244 329656
rect 446364 329616 448244 329644
rect 446364 329604 446370 329616
rect 448238 329604 448244 329616
rect 448296 329604 448302 329656
rect 431218 329060 431224 329112
rect 431276 329100 431282 329112
rect 435634 329100 435640 329112
rect 431276 329072 435640 329100
rect 431276 329060 431282 329072
rect 435634 329060 435640 329072
rect 435692 329060 435698 329112
rect 512546 328992 512552 329044
rect 512604 329032 512610 329044
rect 514202 329032 514208 329044
rect 512604 329004 514208 329032
rect 512604 328992 512610 329004
rect 514202 328992 514208 329004
rect 514260 328992 514266 329044
rect 512546 328720 512552 328772
rect 512604 328760 512610 328772
rect 513926 328760 513932 328772
rect 512604 328732 513932 328760
rect 512604 328720 512610 328732
rect 513926 328720 513932 328732
rect 513984 328720 513990 328772
rect 442902 328448 442908 328500
rect 442960 328488 442966 328500
rect 447778 328488 447784 328500
rect 442960 328460 447784 328488
rect 442960 328448 442966 328460
rect 447778 328448 447784 328460
rect 447836 328488 447842 328500
rect 448238 328488 448244 328500
rect 447836 328460 448244 328488
rect 447836 328448 447842 328460
rect 448238 328448 448244 328460
rect 448296 328448 448302 328500
rect 513282 328448 513288 328500
rect 513340 328488 513346 328500
rect 523586 328488 523592 328500
rect 513340 328460 523592 328488
rect 513340 328448 513346 328460
rect 523586 328448 523592 328460
rect 523644 328448 523650 328500
rect 432874 328380 432880 328432
rect 432932 328420 432938 328432
rect 433794 328420 433800 328432
rect 432932 328392 433800 328420
rect 432932 328380 432938 328392
rect 433794 328380 433800 328392
rect 433852 328380 433858 328432
rect 435082 328380 435088 328432
rect 435140 328420 435146 328432
rect 437382 328420 437388 328432
rect 435140 328392 437388 328420
rect 435140 328380 435146 328392
rect 437382 328380 437388 328392
rect 437440 328380 437446 328432
rect 513282 327360 513288 327412
rect 513340 327400 513346 327412
rect 520918 327400 520924 327412
rect 513340 327372 520924 327400
rect 513340 327360 513346 327372
rect 520918 327360 520924 327372
rect 520976 327360 520982 327412
rect 438762 327088 438768 327140
rect 438820 327128 438826 327140
rect 448514 327128 448520 327140
rect 438820 327100 448520 327128
rect 438820 327088 438826 327100
rect 448514 327088 448520 327100
rect 448572 327088 448578 327140
rect 435726 327020 435732 327072
rect 435784 327060 435790 327072
rect 437290 327060 437296 327072
rect 435784 327032 437296 327060
rect 435784 327020 435790 327032
rect 437290 327020 437296 327032
rect 437348 327020 437354 327072
rect 437474 327020 437480 327072
rect 437532 327060 437538 327072
rect 439774 327060 439780 327072
rect 437532 327032 439780 327060
rect 437532 327020 437538 327032
rect 439774 327020 439780 327032
rect 439832 327020 439838 327072
rect 447686 327020 447692 327072
rect 447744 327060 447750 327072
rect 450262 327060 450268 327072
rect 447744 327032 450268 327060
rect 447744 327020 447750 327032
rect 450262 327020 450268 327032
rect 450320 327020 450326 327072
rect 438118 325116 438124 325168
rect 438176 325156 438182 325168
rect 440234 325156 440240 325168
rect 438176 325128 440240 325156
rect 438176 325116 438182 325128
rect 440234 325116 440240 325128
rect 440292 325116 440298 325168
rect 434070 324300 434076 324352
rect 434128 324340 434134 324352
rect 440970 324340 440976 324352
rect 434128 324312 440976 324340
rect 434128 324300 434134 324312
rect 440970 324300 440976 324312
rect 441028 324300 441034 324352
rect 437014 323620 437020 323672
rect 437072 323660 437078 323672
rect 440326 323660 440332 323672
rect 437072 323632 440332 323660
rect 437072 323620 437078 323632
rect 440326 323620 440332 323632
rect 440384 323620 440390 323672
rect 433794 323484 433800 323536
rect 433852 323524 433858 323536
rect 436186 323524 436192 323536
rect 433852 323496 436192 323524
rect 433852 323484 433858 323496
rect 436186 323484 436192 323496
rect 436244 323484 436250 323536
rect 436094 322872 436100 322924
rect 436152 322912 436158 322924
rect 442718 322912 442724 322924
rect 436152 322884 442724 322912
rect 436152 322872 436158 322884
rect 442718 322872 442724 322884
rect 442776 322872 442782 322924
rect 435634 322328 435640 322380
rect 435692 322368 435698 322380
rect 440418 322368 440424 322380
rect 435692 322340 440424 322368
rect 435692 322328 435698 322340
rect 440418 322328 440424 322340
rect 440476 322328 440482 322380
rect 433978 322192 433984 322244
rect 434036 322232 434042 322244
rect 443730 322232 443736 322244
rect 434036 322204 443736 322232
rect 434036 322192 434042 322204
rect 443730 322192 443736 322204
rect 443788 322192 443794 322244
rect 511902 322192 511908 322244
rect 511960 322232 511966 322244
rect 580350 322232 580356 322244
rect 511960 322204 580356 322232
rect 511960 322192 511966 322204
rect 580350 322192 580356 322204
rect 580408 322192 580414 322244
rect 438302 321512 438308 321564
rect 438360 321552 438366 321564
rect 438854 321552 438860 321564
rect 438360 321524 438860 321552
rect 438360 321512 438366 321524
rect 438854 321512 438860 321524
rect 438912 321512 438918 321564
rect 439774 321512 439780 321564
rect 439832 321552 439838 321564
rect 440694 321552 440700 321564
rect 439832 321524 440700 321552
rect 439832 321512 439838 321524
rect 440694 321512 440700 321524
rect 440752 321512 440758 321564
rect 511350 320900 511356 320952
rect 511408 320940 511414 320952
rect 580534 320940 580540 320952
rect 511408 320912 580540 320940
rect 511408 320900 511414 320912
rect 580534 320900 580540 320912
rect 580592 320900 580598 320952
rect 509970 320832 509976 320884
rect 510028 320872 510034 320884
rect 580626 320872 580632 320884
rect 510028 320844 580632 320872
rect 510028 320832 510034 320844
rect 580626 320832 580632 320844
rect 580684 320832 580690 320884
rect 437290 320152 437296 320204
rect 437348 320192 437354 320204
rect 442534 320192 442540 320204
rect 437348 320164 442540 320192
rect 437348 320152 437354 320164
rect 442534 320152 442540 320164
rect 442592 320152 442598 320204
rect 440234 320084 440240 320136
rect 440292 320124 440298 320136
rect 441982 320124 441988 320136
rect 440292 320096 441988 320124
rect 440292 320084 440298 320096
rect 441982 320084 441988 320096
rect 442040 320084 442046 320136
rect 442718 320084 442724 320136
rect 442776 320124 442782 320136
rect 445754 320124 445760 320136
rect 442776 320096 445760 320124
rect 442776 320084 442782 320096
rect 445754 320084 445760 320096
rect 445812 320084 445818 320136
rect 449158 319948 449164 320000
rect 449216 319988 449222 320000
rect 461578 319988 461584 320000
rect 449216 319960 461584 319988
rect 449216 319948 449222 319960
rect 461578 319948 461584 319960
rect 461636 319948 461642 320000
rect 572070 319988 572076 320000
rect 468588 319960 572076 319988
rect 468588 319932 468616 319960
rect 572070 319948 572076 319960
rect 572128 319948 572134 320000
rect 446582 319880 446588 319932
rect 446640 319920 446646 319932
rect 462498 319920 462504 319932
rect 446640 319892 462504 319920
rect 446640 319880 446646 319892
rect 462498 319880 462504 319892
rect 462556 319880 462562 319932
rect 468570 319880 468576 319932
rect 468628 319880 468634 319932
rect 470226 319880 470232 319932
rect 470284 319920 470290 319932
rect 570598 319920 570604 319932
rect 470284 319892 570604 319920
rect 470284 319880 470290 319892
rect 570598 319880 570604 319892
rect 570656 319880 570662 319932
rect 432782 319812 432788 319864
rect 432840 319852 432846 319864
rect 451734 319852 451740 319864
rect 432840 319824 451740 319852
rect 432840 319812 432846 319824
rect 451734 319812 451740 319824
rect 451792 319812 451798 319864
rect 451918 319812 451924 319864
rect 451976 319852 451982 319864
rect 474366 319852 474372 319864
rect 451976 319824 474372 319852
rect 451976 319812 451982 319824
rect 474366 319812 474372 319824
rect 474424 319812 474430 319864
rect 485038 319812 485044 319864
rect 485096 319852 485102 319864
rect 570782 319852 570788 319864
rect 485096 319824 570788 319852
rect 485096 319812 485102 319824
rect 570782 319812 570788 319824
rect 570840 319812 570846 319864
rect 451826 319744 451832 319796
rect 451884 319784 451890 319796
rect 461394 319784 461400 319796
rect 451884 319756 461400 319784
rect 451884 319744 451890 319756
rect 461394 319744 461400 319756
rect 461452 319744 461458 319796
rect 469674 319744 469680 319796
rect 469732 319784 469738 319796
rect 518250 319784 518256 319796
rect 469732 319756 518256 319784
rect 469732 319744 469738 319756
rect 518250 319744 518256 319756
rect 518308 319744 518314 319796
rect 436186 319676 436192 319728
rect 436244 319716 436250 319728
rect 451734 319716 451740 319728
rect 436244 319688 451740 319716
rect 436244 319676 436250 319688
rect 451734 319676 451740 319688
rect 451792 319676 451798 319728
rect 451918 319676 451924 319728
rect 451976 319716 451982 319728
rect 484578 319716 484584 319728
rect 451976 319688 484584 319716
rect 451976 319676 451982 319688
rect 484578 319676 484584 319688
rect 484636 319676 484642 319728
rect 437474 319608 437480 319660
rect 437532 319648 437538 319660
rect 446306 319648 446312 319660
rect 437532 319620 446312 319648
rect 437532 319608 437538 319620
rect 446306 319608 446312 319620
rect 446364 319608 446370 319660
rect 446490 319608 446496 319660
rect 446548 319648 446554 319660
rect 451826 319648 451832 319660
rect 446548 319620 451832 319648
rect 446548 319608 446554 319620
rect 451826 319608 451832 319620
rect 451884 319608 451890 319660
rect 469122 319608 469128 319660
rect 469180 319648 469186 319660
rect 514018 319648 514024 319660
rect 469180 319620 514024 319648
rect 469180 319608 469186 319620
rect 514018 319608 514024 319620
rect 514076 319608 514082 319660
rect 440326 319540 440332 319592
rect 440384 319580 440390 319592
rect 484026 319580 484032 319592
rect 440384 319552 484032 319580
rect 440384 319540 440390 319552
rect 484026 319540 484032 319552
rect 484084 319540 484090 319592
rect 445110 319472 445116 319524
rect 445168 319512 445174 319524
rect 471238 319512 471244 319524
rect 445168 319484 471244 319512
rect 445168 319472 445174 319484
rect 471238 319472 471244 319484
rect 471296 319472 471302 319524
rect 500218 319472 500224 319524
rect 500276 319512 500282 319524
rect 580258 319512 580264 319524
rect 500276 319484 580264 319512
rect 500276 319472 500282 319484
rect 580258 319472 580264 319484
rect 580316 319472 580322 319524
rect 438210 319404 438216 319456
rect 438268 319444 438274 319456
rect 446398 319444 446404 319456
rect 438268 319416 446404 319444
rect 438268 319404 438274 319416
rect 446398 319404 446404 319416
rect 446456 319404 446462 319456
rect 481450 319404 481456 319456
rect 481508 319444 481514 319456
rect 579982 319444 579988 319456
rect 481508 319416 579988 319444
rect 481508 319404 481514 319416
rect 579982 319404 579988 319416
rect 580040 319404 580046 319456
rect 447042 319336 447048 319388
rect 447100 319376 447106 319388
rect 483750 319376 483756 319388
rect 447100 319348 483756 319376
rect 447100 319336 447106 319348
rect 483750 319336 483756 319348
rect 483808 319336 483814 319388
rect 446490 319268 446496 319320
rect 446548 319308 446554 319320
rect 460842 319308 460848 319320
rect 446548 319280 460848 319308
rect 446548 319268 446554 319280
rect 460842 319268 460848 319280
rect 460900 319268 460906 319320
rect 433518 319200 433524 319252
rect 433576 319240 433582 319252
rect 435450 319240 435456 319252
rect 433576 319212 435456 319240
rect 433576 319200 433582 319212
rect 435450 319200 435456 319212
rect 435508 319200 435514 319252
rect 446766 319200 446772 319252
rect 446824 319240 446830 319252
rect 446824 319212 458864 319240
rect 446824 319200 446830 319212
rect 438854 319132 438860 319184
rect 438912 319172 438918 319184
rect 438912 319144 447134 319172
rect 438912 319132 438918 319144
rect 447106 319104 447134 319144
rect 458836 319104 458864 319212
rect 479058 319200 479064 319252
rect 479116 319240 479122 319252
rect 485038 319240 485044 319252
rect 479116 319212 485044 319240
rect 479116 319200 479122 319212
rect 485038 319200 485044 319212
rect 485096 319200 485102 319252
rect 461026 319132 461032 319184
rect 461084 319172 461090 319184
rect 484302 319172 484308 319184
rect 461084 319144 484308 319172
rect 461084 319132 461090 319144
rect 484302 319132 484308 319144
rect 484360 319132 484366 319184
rect 472986 319104 472992 319116
rect 447106 319076 454034 319104
rect 458836 319076 472992 319104
rect 454006 319036 454034 319076
rect 472986 319064 472992 319076
rect 473044 319064 473050 319116
rect 461026 319036 461032 319048
rect 454006 319008 461032 319036
rect 461026 318996 461032 319008
rect 461084 318996 461090 319048
rect 471238 318996 471244 319048
rect 471296 319036 471302 319048
rect 482646 319036 482652 319048
rect 471296 319008 482652 319036
rect 471296 318996 471302 319008
rect 482646 318996 482652 319008
rect 482704 318996 482710 319048
rect 442534 318792 442540 318844
rect 442592 318832 442598 318844
rect 481450 318832 481456 318844
rect 442592 318804 443040 318832
rect 442592 318792 442598 318804
rect 443012 318764 443040 318804
rect 480226 318804 481456 318832
rect 445846 318764 445852 318776
rect 443012 318736 445852 318764
rect 445846 318724 445852 318736
rect 445904 318724 445910 318776
rect 446398 318724 446404 318776
rect 446456 318764 446462 318776
rect 463326 318764 463332 318776
rect 446456 318736 463332 318764
rect 446456 318724 446462 318736
rect 463326 318724 463332 318736
rect 463384 318724 463390 318776
rect 478782 318724 478788 318776
rect 478840 318764 478846 318776
rect 480226 318764 480254 318804
rect 481450 318792 481456 318804
rect 481508 318792 481514 318844
rect 478840 318736 480254 318764
rect 478840 318724 478846 318736
rect 480438 318724 480444 318776
rect 480496 318764 480502 318776
rect 489638 318764 489644 318776
rect 480496 318736 489644 318764
rect 480496 318724 480502 318736
rect 489638 318724 489644 318736
rect 489696 318724 489702 318776
rect 458358 318656 458364 318708
rect 458416 318696 458422 318708
rect 580442 318696 580448 318708
rect 458416 318668 580448 318696
rect 458416 318656 458422 318668
rect 580442 318656 580448 318668
rect 580500 318656 580506 318708
rect 445478 318588 445484 318640
rect 445536 318628 445542 318640
rect 460566 318628 460572 318640
rect 445536 318600 460572 318628
rect 445536 318588 445542 318600
rect 460566 318588 460572 318600
rect 460624 318588 460630 318640
rect 469950 318588 469956 318640
rect 470008 318628 470014 318640
rect 577498 318628 577504 318640
rect 470008 318600 577504 318628
rect 470008 318588 470014 318600
rect 577498 318588 577504 318600
rect 577556 318588 577562 318640
rect 444190 318520 444196 318572
rect 444248 318560 444254 318572
rect 460290 318560 460296 318572
rect 444248 318532 460296 318560
rect 444248 318520 444254 318532
rect 460290 318520 460296 318532
rect 460348 318520 460354 318572
rect 470502 318520 470508 318572
rect 470560 318560 470566 318572
rect 516778 318560 516784 318572
rect 470560 318532 516784 318560
rect 470560 318520 470566 318532
rect 516778 318520 516784 318532
rect 516836 318520 516842 318572
rect 441982 318452 441988 318504
rect 442040 318492 442046 318504
rect 444650 318492 444656 318504
rect 442040 318464 444656 318492
rect 442040 318452 442046 318464
rect 444650 318452 444656 318464
rect 444708 318452 444714 318504
rect 449342 318452 449348 318504
rect 449400 318492 449406 318504
rect 471054 318492 471060 318504
rect 449400 318464 471060 318492
rect 449400 318452 449406 318464
rect 471054 318452 471060 318464
rect 471112 318452 471118 318504
rect 480162 318452 480168 318504
rect 480220 318492 480226 318504
rect 522298 318492 522304 318504
rect 480220 318464 522304 318492
rect 480220 318452 480226 318464
rect 522298 318452 522304 318464
rect 522356 318452 522362 318504
rect 468846 318384 468852 318436
rect 468904 318424 468910 318436
rect 509970 318424 509976 318436
rect 468904 318396 509976 318424
rect 468904 318384 468910 318396
rect 509970 318384 509976 318396
rect 510028 318384 510034 318436
rect 469398 318316 469404 318368
rect 469456 318356 469462 318368
rect 511902 318356 511908 318368
rect 469456 318328 511908 318356
rect 469456 318316 469462 318328
rect 511902 318316 511908 318328
rect 511960 318316 511966 318368
rect 445570 318248 445576 318300
rect 445628 318288 445634 318300
rect 462774 318288 462780 318300
rect 445628 318260 462780 318288
rect 445628 318248 445634 318260
rect 462774 318248 462780 318260
rect 462832 318248 462838 318300
rect 479886 318248 479892 318300
rect 479944 318288 479950 318300
rect 518342 318288 518348 318300
rect 479944 318260 518348 318288
rect 479944 318248 479950 318260
rect 518342 318248 518348 318260
rect 518400 318248 518406 318300
rect 446674 318180 446680 318232
rect 446732 318220 446738 318232
rect 472158 318220 472164 318232
rect 446732 318192 472164 318220
rect 446732 318180 446738 318192
rect 472158 318180 472164 318192
rect 472216 318180 472222 318232
rect 479334 318180 479340 318232
rect 479392 318220 479398 318232
rect 479392 318192 480254 318220
rect 479392 318180 479398 318192
rect 458082 318112 458088 318164
rect 458140 318152 458146 318164
rect 462222 318152 462228 318164
rect 458140 318124 462228 318152
rect 458140 318112 458146 318124
rect 462222 318112 462228 318124
rect 462280 318112 462286 318164
rect 478506 318112 478512 318164
rect 478564 318152 478570 318164
rect 479518 318152 479524 318164
rect 478564 318124 479524 318152
rect 478564 318112 478570 318124
rect 479518 318112 479524 318124
rect 479576 318112 479582 318164
rect 480226 318152 480254 318192
rect 480990 318180 480996 318232
rect 481048 318220 481054 318232
rect 481450 318220 481456 318232
rect 481048 318192 481456 318220
rect 481048 318180 481054 318192
rect 481450 318180 481456 318192
rect 481508 318180 481514 318232
rect 487154 318180 487160 318232
rect 487212 318220 487218 318232
rect 488442 318220 488448 318232
rect 487212 318192 488448 318220
rect 487212 318180 487218 318192
rect 488442 318180 488448 318192
rect 488500 318180 488506 318232
rect 489914 318180 489920 318232
rect 489972 318220 489978 318232
rect 491202 318220 491208 318232
rect 489972 318192 491208 318220
rect 489972 318180 489978 318192
rect 491202 318180 491208 318192
rect 491260 318180 491266 318232
rect 494146 318180 494152 318232
rect 494204 318220 494210 318232
rect 494790 318220 494796 318232
rect 494204 318192 494796 318220
rect 494204 318180 494210 318192
rect 494790 318180 494796 318192
rect 494848 318180 494854 318232
rect 498378 318180 498384 318232
rect 498436 318220 498442 318232
rect 542998 318220 543004 318232
rect 498436 318192 543004 318220
rect 498436 318180 498442 318192
rect 542998 318180 543004 318192
rect 543056 318180 543062 318232
rect 500218 318152 500224 318164
rect 480226 318124 500224 318152
rect 500218 318112 500224 318124
rect 500276 318112 500282 318164
rect 503070 318112 503076 318164
rect 503128 318152 503134 318164
rect 548518 318152 548524 318164
rect 503128 318124 548524 318152
rect 503128 318112 503134 318124
rect 548518 318112 548524 318124
rect 548576 318112 548582 318164
rect 440694 318044 440700 318096
rect 440752 318084 440758 318096
rect 444466 318084 444472 318096
rect 440752 318056 444472 318084
rect 440752 318044 440758 318056
rect 444466 318044 444472 318056
rect 444524 318044 444530 318096
rect 461578 318044 461584 318096
rect 461636 318084 461642 318096
rect 461636 318056 476114 318084
rect 461636 318044 461642 318056
rect 445754 317976 445760 318028
rect 445812 318016 445818 318028
rect 473538 318016 473544 318028
rect 445812 317988 473544 318016
rect 445812 317976 445818 317988
rect 473538 317976 473544 317988
rect 473596 317976 473602 318028
rect 445202 317908 445208 317960
rect 445260 317948 445266 317960
rect 471606 317948 471612 317960
rect 445260 317920 471612 317948
rect 445260 317908 445266 317920
rect 471606 317908 471612 317920
rect 471664 317908 471670 317960
rect 476086 317948 476114 318056
rect 477954 318044 477960 318096
rect 478012 318084 478018 318096
rect 478598 318084 478604 318096
rect 478012 318056 478604 318084
rect 478012 318044 478018 318056
rect 478598 318044 478604 318056
rect 478656 318044 478662 318096
rect 484486 318044 484492 318096
rect 484544 318084 484550 318096
rect 485406 318084 485412 318096
rect 484544 318056 485412 318084
rect 484544 318044 484550 318056
rect 485406 318044 485412 318056
rect 485464 318044 485470 318096
rect 485866 318044 485872 318096
rect 485924 318084 485930 318096
rect 486786 318084 486792 318096
rect 485924 318056 486792 318084
rect 485924 318044 485930 318056
rect 486786 318044 486792 318056
rect 486844 318044 486850 318096
rect 487614 318044 487620 318096
rect 487672 318084 487678 318096
rect 488350 318084 488356 318096
rect 487672 318056 488356 318084
rect 487672 318044 487678 318056
rect 488350 318044 488356 318056
rect 488408 318044 488414 318096
rect 490006 318044 490012 318096
rect 490064 318084 490070 318096
rect 490374 318084 490380 318096
rect 490064 318056 490380 318084
rect 490064 318044 490070 318056
rect 490374 318044 490380 318056
rect 490432 318044 490438 318096
rect 494054 318044 494060 318096
rect 494112 318084 494118 318096
rect 494514 318084 494520 318096
rect 494112 318056 494520 318084
rect 494112 318044 494118 318056
rect 494514 318044 494520 318056
rect 494572 318044 494578 318096
rect 497274 318044 497280 318096
rect 497332 318084 497338 318096
rect 548610 318084 548616 318096
rect 497332 318056 548616 318084
rect 497332 318044 497338 318056
rect 548610 318044 548616 318056
rect 548668 318044 548674 318096
rect 477678 317976 477684 318028
rect 477736 318016 477742 318028
rect 478690 318016 478696 318028
rect 477736 317988 478696 318016
rect 477736 317976 477742 317988
rect 478690 317976 478696 317988
rect 478748 317976 478754 318028
rect 481450 317976 481456 318028
rect 481508 318016 481514 318028
rect 481508 317988 487752 318016
rect 481508 317976 481514 317988
rect 476298 317948 476304 317960
rect 476086 317920 476304 317948
rect 476298 317908 476304 317920
rect 476356 317908 476362 317960
rect 477126 317908 477132 317960
rect 477184 317948 477190 317960
rect 477494 317948 477500 317960
rect 477184 317920 477500 317948
rect 477184 317908 477190 317920
rect 477494 317908 477500 317920
rect 477552 317908 477558 317960
rect 480346 317908 480352 317960
rect 480404 317948 480410 317960
rect 481542 317948 481548 317960
rect 480404 317920 481548 317948
rect 480404 317908 480410 317920
rect 481542 317908 481548 317920
rect 481600 317908 481606 317960
rect 484670 317908 484676 317960
rect 484728 317948 484734 317960
rect 485682 317948 485688 317960
rect 484728 317920 485688 317948
rect 484728 317908 484734 317920
rect 485682 317908 485688 317920
rect 485740 317908 485746 317960
rect 485958 317908 485964 317960
rect 486016 317948 486022 317960
rect 486510 317948 486516 317960
rect 486016 317920 486516 317948
rect 486016 317908 486022 317920
rect 486510 317908 486516 317920
rect 486568 317908 486574 317960
rect 487724 317948 487752 317988
rect 487890 317976 487896 318028
rect 487948 318016 487954 318028
rect 488442 318016 488448 318028
rect 487948 317988 488448 318016
rect 487948 317976 487954 317988
rect 488442 317976 488448 317988
rect 488500 317976 488506 318028
rect 518158 318016 518164 318028
rect 488552 317988 518164 318016
rect 488552 317948 488580 317988
rect 518158 317976 518164 317988
rect 518216 317976 518222 318028
rect 487724 317920 488580 317948
rect 488626 317908 488632 317960
rect 488684 317948 488690 317960
rect 489546 317948 489552 317960
rect 488684 317920 489552 317948
rect 488684 317908 488690 317920
rect 489546 317908 489552 317920
rect 489604 317908 489610 317960
rect 489638 317908 489644 317960
rect 489696 317948 489702 317960
rect 515398 317948 515404 317960
rect 489696 317920 515404 317948
rect 489696 317908 489702 317920
rect 515398 317908 515404 317920
rect 515456 317908 515462 317960
rect 456334 317840 456340 317892
rect 456392 317880 456398 317892
rect 461578 317880 461584 317892
rect 456392 317852 461584 317880
rect 456392 317840 456398 317852
rect 461578 317840 461584 317852
rect 461636 317840 461642 317892
rect 462222 317840 462228 317892
rect 462280 317880 462286 317892
rect 580718 317880 580724 317892
rect 462280 317852 580724 317880
rect 462280 317840 462286 317852
rect 580718 317840 580724 317852
rect 580776 317840 580782 317892
rect 446858 317772 446864 317824
rect 446916 317812 446922 317824
rect 471330 317812 471336 317824
rect 446916 317784 471336 317812
rect 446916 317772 446922 317784
rect 471330 317772 471336 317784
rect 471388 317772 471394 317824
rect 479610 317772 479616 317824
rect 479668 317812 479674 317824
rect 511350 317812 511356 317824
rect 479668 317784 511356 317812
rect 479668 317772 479674 317784
rect 511350 317772 511356 317784
rect 511408 317772 511414 317824
rect 445294 317704 445300 317756
rect 445352 317744 445358 317756
rect 482094 317744 482100 317756
rect 445352 317716 482100 317744
rect 445352 317704 445358 317716
rect 482094 317704 482100 317716
rect 482152 317704 482158 317756
rect 486050 317704 486056 317756
rect 486108 317744 486114 317756
rect 487062 317744 487068 317756
rect 486108 317716 487068 317744
rect 486108 317704 486114 317716
rect 487062 317704 487068 317716
rect 487120 317704 487126 317756
rect 490190 317704 490196 317756
rect 490248 317744 490254 317756
rect 490650 317744 490656 317756
rect 490248 317716 490656 317744
rect 490248 317704 490254 317716
rect 490650 317704 490656 317716
rect 490708 317704 490714 317756
rect 491386 317704 491392 317756
rect 491444 317744 491450 317756
rect 492030 317744 492036 317756
rect 491444 317716 492036 317744
rect 491444 317704 491450 317716
rect 492030 317704 492036 317716
rect 492088 317704 492094 317756
rect 492766 317704 492772 317756
rect 492824 317744 492830 317756
rect 493962 317744 493968 317756
rect 492824 317716 493968 317744
rect 492824 317704 492830 317716
rect 493962 317704 493968 317716
rect 494020 317704 494026 317756
rect 444282 317636 444288 317688
rect 444340 317676 444346 317688
rect 470778 317676 470784 317688
rect 444340 317648 470784 317676
rect 444340 317636 444346 317648
rect 470778 317636 470784 317648
rect 470836 317636 470842 317688
rect 485038 317636 485044 317688
rect 485096 317676 485102 317688
rect 486234 317676 486240 317688
rect 485096 317648 486240 317676
rect 485096 317636 485102 317648
rect 486234 317636 486240 317648
rect 486292 317636 486298 317688
rect 490098 317636 490104 317688
rect 490156 317676 490162 317688
rect 490926 317676 490932 317688
rect 490156 317648 490932 317676
rect 490156 317636 490162 317648
rect 490926 317636 490932 317648
rect 490984 317636 490990 317688
rect 491478 317636 491484 317688
rect 491536 317676 491542 317688
rect 492306 317676 492312 317688
rect 491536 317648 492312 317676
rect 491536 317636 491542 317648
rect 492306 317636 492312 317648
rect 492364 317636 492370 317688
rect 471974 317500 471980 317552
rect 472032 317540 472038 317552
rect 474918 317540 474924 317552
rect 472032 317512 474924 317540
rect 472032 317500 472038 317512
rect 474918 317500 474924 317512
rect 474976 317500 474982 317552
rect 460198 317432 460204 317484
rect 460256 317472 460262 317484
rect 465810 317472 465816 317484
rect 460256 317444 465816 317472
rect 460256 317432 460262 317444
rect 465810 317432 465816 317444
rect 465868 317432 465874 317484
rect 472710 317432 472716 317484
rect 472768 317472 472774 317484
rect 475194 317472 475200 317484
rect 472768 317444 475200 317472
rect 472768 317432 472774 317444
rect 475194 317432 475200 317444
rect 475252 317432 475258 317484
rect 446398 317364 446404 317416
rect 446456 317404 446462 317416
rect 447962 317404 447968 317416
rect 446456 317376 447968 317404
rect 446456 317364 446462 317376
rect 447962 317364 447968 317376
rect 448020 317364 448026 317416
rect 459462 317364 459468 317416
rect 459520 317404 459526 317416
rect 571978 317404 571984 317416
rect 459520 317376 571984 317404
rect 459520 317364 459526 317376
rect 571978 317364 571984 317376
rect 572036 317364 572042 317416
rect 459738 317296 459744 317348
rect 459796 317336 459802 317348
rect 573358 317336 573364 317348
rect 459796 317308 573364 317336
rect 459796 317296 459802 317308
rect 573358 317296 573364 317308
rect 573416 317296 573422 317348
rect 458634 317228 458640 317280
rect 458692 317268 458698 317280
rect 570690 317268 570696 317280
rect 458692 317240 570696 317268
rect 458692 317228 458698 317240
rect 570690 317228 570696 317240
rect 570748 317228 570754 317280
rect 458910 317160 458916 317212
rect 458968 317200 458974 317212
rect 519538 317200 519544 317212
rect 458968 317172 519544 317200
rect 458968 317160 458974 317172
rect 519538 317160 519544 317172
rect 519596 317160 519602 317212
rect 459186 317092 459192 317144
rect 459244 317132 459250 317144
rect 515490 317132 515496 317144
rect 459244 317104 515496 317132
rect 459244 317092 459250 317104
rect 515490 317092 515496 317104
rect 515548 317092 515554 317144
rect 445018 317024 445024 317076
rect 445076 317064 445082 317076
rect 481818 317064 481824 317076
rect 445076 317036 481824 317064
rect 445076 317024 445082 317036
rect 481818 317024 481824 317036
rect 481876 317024 481882 317076
rect 440050 316956 440056 317008
rect 440108 316996 440114 317008
rect 471882 316996 471888 317008
rect 440108 316968 471888 316996
rect 440108 316956 440114 316968
rect 471882 316956 471888 316968
rect 471940 316956 471946 317008
rect 444650 316888 444656 316940
rect 444708 316928 444714 316940
rect 473814 316928 473820 316940
rect 444708 316900 473820 316928
rect 444708 316888 444714 316900
rect 473814 316888 473820 316900
rect 473872 316888 473878 316940
rect 439958 316820 439964 316872
rect 440016 316860 440022 316872
rect 473262 316860 473268 316872
rect 440016 316832 473268 316860
rect 440016 316820 440022 316832
rect 473262 316820 473268 316832
rect 473320 316820 473326 316872
rect 481634 316820 481640 316872
rect 481692 316860 481698 316872
rect 485130 316860 485136 316872
rect 481692 316832 485136 316860
rect 481692 316820 481698 316832
rect 485130 316820 485136 316832
rect 485188 316820 485194 316872
rect 446306 316752 446312 316804
rect 446364 316792 446370 316804
rect 474090 316792 474096 316804
rect 446364 316764 474096 316792
rect 446364 316752 446370 316764
rect 474090 316752 474096 316764
rect 474148 316752 474154 316804
rect 494238 316752 494244 316804
rect 494296 316792 494302 316804
rect 495342 316792 495348 316804
rect 494296 316764 495348 316792
rect 494296 316752 494302 316764
rect 495342 316752 495348 316764
rect 495400 316752 495406 316804
rect 450446 316684 450452 316736
rect 450504 316724 450510 316736
rect 451918 316724 451924 316736
rect 450504 316696 451924 316724
rect 450504 316684 450510 316696
rect 451918 316684 451924 316696
rect 451976 316684 451982 316736
rect 439866 316616 439872 316668
rect 439924 316656 439930 316668
rect 472434 316656 472440 316668
rect 439924 316628 472440 316656
rect 439924 316616 439930 316628
rect 472434 316616 472440 316628
rect 472492 316616 472498 316668
rect 440418 316548 440424 316600
rect 440476 316588 440482 316600
rect 463878 316588 463884 316600
rect 440476 316560 463884 316588
rect 440476 316548 440482 316560
rect 463878 316548 463884 316560
rect 463936 316548 463942 316600
rect 445846 316480 445852 316532
rect 445904 316520 445910 316532
rect 463602 316520 463608 316532
rect 445904 316492 463608 316520
rect 445904 316480 445910 316492
rect 463602 316480 463608 316492
rect 463660 316480 463666 316532
rect 444466 316412 444472 316464
rect 444524 316452 444530 316464
rect 463050 316452 463056 316464
rect 444524 316424 463056 316452
rect 444524 316412 444530 316424
rect 463050 316412 463056 316424
rect 463108 316412 463114 316464
rect 456978 316072 456984 316124
rect 457036 316112 457042 316124
rect 457898 316112 457904 316124
rect 457036 316084 457904 316112
rect 457036 316072 457042 316084
rect 457898 316072 457904 316084
rect 457956 316072 457962 316124
rect 457254 316004 457260 316056
rect 457312 316044 457318 316056
rect 457990 316044 457996 316056
rect 457312 316016 457996 316044
rect 457312 316004 457318 316016
rect 457990 316004 457996 316016
rect 458048 316004 458054 316056
rect 442350 315936 442356 315988
rect 442408 315976 442414 315988
rect 481818 315976 481824 315988
rect 442408 315948 481824 315976
rect 442408 315936 442414 315948
rect 481818 315936 481824 315948
rect 481876 315936 481882 315988
rect 498654 315936 498660 315988
rect 498712 315976 498718 315988
rect 499390 315976 499396 315988
rect 498712 315948 499396 315976
rect 498712 315936 498718 315948
rect 499390 315936 499396 315948
rect 499448 315936 499454 315988
rect 501414 315936 501420 315988
rect 501472 315976 501478 315988
rect 502058 315976 502064 315988
rect 501472 315948 502064 315976
rect 501472 315936 501478 315948
rect 502058 315936 502064 315948
rect 502116 315936 502122 315988
rect 450630 315868 450636 315920
rect 450688 315908 450694 315920
rect 452010 315908 452016 315920
rect 450688 315880 452016 315908
rect 450688 315868 450694 315880
rect 452010 315868 452016 315880
rect 452068 315868 452074 315920
rect 480254 315908 480260 315920
rect 453500 315880 480260 315908
rect 450814 315800 450820 315852
rect 450872 315840 450878 315852
rect 453298 315840 453304 315852
rect 450872 315812 453304 315840
rect 450872 315800 450878 315812
rect 453298 315800 453304 315812
rect 453356 315800 453362 315852
rect 448422 315664 448428 315716
rect 448480 315704 448486 315716
rect 453500 315704 453528 315880
rect 480254 315868 480260 315880
rect 480312 315868 480318 315920
rect 497550 315868 497556 315920
rect 497608 315908 497614 315920
rect 498010 315908 498016 315920
rect 497608 315880 498016 315908
rect 497608 315868 497614 315880
rect 498010 315868 498016 315880
rect 498068 315868 498074 315920
rect 500586 315868 500592 315920
rect 500644 315908 500650 315920
rect 500770 315908 500776 315920
rect 500644 315880 500776 315908
rect 500644 315868 500650 315880
rect 500770 315868 500776 315880
rect 500828 315868 500834 315920
rect 501690 315868 501696 315920
rect 501748 315908 501754 315920
rect 502242 315908 502248 315920
rect 501748 315880 502248 315908
rect 501748 315868 501754 315880
rect 502242 315868 502248 315880
rect 502300 315868 502306 315920
rect 480346 315840 480352 315852
rect 448480 315676 453528 315704
rect 453592 315812 480352 315840
rect 448480 315664 448486 315676
rect 449250 315596 449256 315648
rect 449308 315636 449314 315648
rect 453592 315636 453620 315812
rect 480346 315800 480352 315812
rect 480404 315800 480410 315852
rect 455138 315732 455144 315784
rect 455196 315772 455202 315784
rect 476022 315772 476028 315784
rect 455196 315744 476028 315772
rect 455196 315732 455202 315744
rect 476022 315732 476028 315744
rect 476080 315732 476086 315784
rect 500034 315732 500040 315784
rect 500092 315772 500098 315784
rect 500586 315772 500592 315784
rect 500092 315744 500592 315772
rect 500092 315732 500098 315744
rect 500586 315732 500592 315744
rect 500644 315732 500650 315784
rect 454862 315664 454868 315716
rect 454920 315704 454926 315716
rect 510798 315704 510804 315716
rect 454920 315676 510804 315704
rect 454920 315664 454926 315676
rect 510798 315664 510804 315676
rect 510856 315664 510862 315716
rect 449308 315608 453620 315636
rect 449308 315596 449314 315608
rect 456058 315596 456064 315648
rect 456116 315636 456122 315648
rect 512730 315636 512736 315648
rect 456116 315608 512736 315636
rect 456116 315596 456122 315608
rect 512730 315596 512736 315608
rect 512788 315596 512794 315648
rect 456242 315528 456248 315580
rect 456300 315568 456306 315580
rect 512546 315568 512552 315580
rect 456300 315540 512552 315568
rect 456300 315528 456306 315540
rect 512546 315528 512552 315540
rect 512604 315528 512610 315580
rect 454678 315460 454684 315512
rect 454736 315500 454742 315512
rect 512178 315500 512184 315512
rect 454736 315472 512184 315500
rect 454736 315460 454742 315472
rect 512178 315460 512184 315472
rect 512236 315460 512242 315512
rect 454954 315392 454960 315444
rect 455012 315432 455018 315444
rect 513650 315432 513656 315444
rect 455012 315404 513656 315432
rect 455012 315392 455018 315404
rect 513650 315392 513656 315404
rect 513708 315392 513714 315444
rect 448514 315324 448520 315376
rect 448572 315364 448578 315376
rect 471974 315364 471980 315376
rect 448572 315336 471980 315364
rect 448572 315324 448578 315336
rect 471974 315324 471980 315336
rect 472032 315324 472038 315376
rect 478598 315324 478604 315376
rect 478656 315364 478662 315376
rect 538858 315364 538864 315376
rect 478656 315336 538864 315364
rect 478656 315324 478662 315336
rect 538858 315324 538864 315336
rect 538916 315324 538922 315376
rect 455046 315256 455052 315308
rect 455104 315296 455110 315308
rect 516134 315296 516140 315308
rect 455104 315268 516140 315296
rect 455104 315256 455110 315268
rect 516134 315256 516140 315268
rect 516192 315256 516198 315308
rect 456426 315188 456432 315240
rect 456484 315228 456490 315240
rect 456702 315228 456708 315240
rect 456484 315200 456708 315228
rect 456484 315188 456490 315200
rect 456702 315188 456708 315200
rect 456760 315188 456766 315240
rect 457806 315188 457812 315240
rect 457864 315228 457870 315240
rect 461578 315228 461584 315240
rect 457864 315200 461584 315228
rect 457864 315188 457870 315200
rect 461578 315188 461584 315200
rect 461636 315188 461642 315240
rect 463602 315188 463608 315240
rect 463660 315228 463666 315240
rect 464154 315228 464160 315240
rect 463660 315200 464160 315228
rect 463660 315188 463666 315200
rect 464154 315188 464160 315200
rect 464212 315188 464218 315240
rect 473354 315188 473360 315240
rect 473412 315228 473418 315240
rect 486142 315228 486148 315240
rect 473412 315200 486148 315228
rect 473412 315188 473418 315200
rect 486142 315188 486148 315200
rect 486200 315188 486206 315240
rect 455230 315120 455236 315172
rect 455288 315160 455294 315172
rect 465534 315160 465540 315172
rect 455288 315132 465540 315160
rect 455288 315120 455294 315132
rect 465534 315120 465540 315132
rect 465592 315120 465598 315172
rect 434254 315052 434260 315104
rect 434312 315092 434318 315104
rect 436922 315092 436928 315104
rect 434312 315064 436928 315092
rect 434312 315052 434318 315064
rect 436922 315052 436928 315064
rect 436980 315052 436986 315104
rect 456150 314848 456156 314900
rect 456208 314888 456214 314900
rect 456610 314888 456616 314900
rect 456208 314860 456616 314888
rect 456208 314848 456214 314860
rect 456610 314848 456616 314860
rect 456668 314848 456674 314900
rect 481634 314684 481640 314696
rect 480226 314656 481640 314684
rect 462222 314576 462228 314628
rect 462280 314616 462286 314628
rect 464982 314616 464988 314628
rect 462280 314588 464988 314616
rect 462280 314576 462286 314588
rect 464982 314576 464988 314588
rect 465040 314576 465046 314628
rect 479610 314576 479616 314628
rect 479668 314616 479674 314628
rect 480226 314616 480254 314656
rect 481634 314644 481640 314656
rect 481692 314644 481698 314696
rect 484578 314684 484584 314696
rect 481744 314656 484584 314684
rect 479668 314588 480254 314616
rect 479668 314576 479674 314588
rect 481542 314576 481548 314628
rect 481600 314616 481606 314628
rect 481744 314616 481772 314656
rect 484578 314644 484584 314656
rect 484636 314644 484642 314696
rect 481600 314588 481772 314616
rect 481600 314576 481606 314588
rect 467558 314168 467564 314220
rect 467616 314208 467622 314220
rect 467742 314208 467748 314220
rect 467616 314180 467748 314208
rect 467616 314168 467622 314180
rect 467742 314168 467748 314180
rect 467800 314168 467806 314220
rect 460474 314100 460480 314152
rect 460532 314140 460538 314152
rect 491294 314140 491300 314152
rect 460532 314112 491300 314140
rect 460532 314100 460538 314112
rect 491294 314100 491300 314112
rect 491352 314100 491358 314152
rect 440970 314032 440976 314084
rect 441028 314072 441034 314084
rect 475746 314072 475752 314084
rect 441028 314044 475752 314072
rect 441028 314032 441034 314044
rect 475746 314032 475752 314044
rect 475804 314032 475810 314084
rect 499758 314032 499764 314084
rect 499816 314072 499822 314084
rect 550910 314072 550916 314084
rect 499816 314044 550916 314072
rect 499816 314032 499822 314044
rect 550910 314032 550916 314044
rect 550968 314032 550974 314084
rect 459002 313964 459008 314016
rect 459060 314004 459066 314016
rect 495894 314004 495900 314016
rect 459060 313976 495900 314004
rect 459060 313964 459066 313976
rect 495894 313964 495900 313976
rect 495952 313964 495958 314016
rect 496170 313964 496176 314016
rect 496228 314004 496234 314016
rect 550634 314004 550640 314016
rect 496228 313976 550640 314004
rect 496228 313964 496234 313976
rect 550634 313964 550640 313976
rect 550692 313964 550698 314016
rect 455966 313896 455972 313948
rect 456024 313936 456030 313948
rect 566458 313936 566464 313948
rect 456024 313908 566464 313936
rect 456024 313896 456030 313908
rect 566458 313896 566464 313908
rect 566516 313896 566522 313948
rect 466914 313828 466920 313880
rect 466972 313868 466978 313880
rect 467558 313868 467564 313880
rect 466972 313840 467564 313868
rect 466972 313828 466978 313840
rect 467558 313828 467564 313840
rect 467616 313828 467622 313880
rect 468294 313216 468300 313268
rect 468352 313256 468358 313268
rect 580166 313256 580172 313268
rect 468352 313228 580172 313256
rect 468352 313216 468358 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 472618 313012 472624 313064
rect 472676 313052 472682 313064
rect 474642 313052 474648 313064
rect 472676 313024 474648 313052
rect 472676 313012 472682 313024
rect 474642 313012 474648 313024
rect 474700 313012 474706 313064
rect 465810 312808 465816 312860
rect 465868 312848 465874 312860
rect 473354 312848 473360 312860
rect 465868 312820 473360 312848
rect 465868 312808 465874 312820
rect 473354 312808 473360 312820
rect 473412 312808 473418 312860
rect 460290 312740 460296 312792
rect 460348 312780 460354 312792
rect 488534 312780 488540 312792
rect 460348 312752 488540 312780
rect 460348 312740 460354 312752
rect 488534 312740 488540 312752
rect 488592 312740 488598 312792
rect 499482 312740 499488 312792
rect 499540 312780 499546 312792
rect 499540 312752 502288 312780
rect 499540 312740 499546 312752
rect 460382 312672 460388 312724
rect 460440 312712 460446 312724
rect 488810 312712 488816 312724
rect 460440 312684 488816 312712
rect 460440 312672 460446 312684
rect 488810 312672 488816 312684
rect 488868 312672 488874 312724
rect 501138 312672 501144 312724
rect 501196 312712 501202 312724
rect 501966 312712 501972 312724
rect 501196 312684 501972 312712
rect 501196 312672 501202 312684
rect 501966 312672 501972 312684
rect 502024 312672 502030 312724
rect 502260 312712 502288 312752
rect 502518 312740 502524 312792
rect 502576 312780 502582 312792
rect 549530 312780 549536 312792
rect 502576 312752 549536 312780
rect 502576 312740 502582 312752
rect 549530 312740 549536 312752
rect 549588 312740 549594 312792
rect 550818 312712 550824 312724
rect 502260 312684 550824 312712
rect 550818 312672 550824 312684
rect 550876 312672 550882 312724
rect 458818 312604 458824 312656
rect 458876 312644 458882 312656
rect 492674 312644 492680 312656
rect 458876 312616 492680 312644
rect 458876 312604 458882 312616
rect 492674 312604 492680 312616
rect 492732 312604 492738 312656
rect 498930 312604 498936 312656
rect 498988 312644 498994 312656
rect 550726 312644 550732 312656
rect 498988 312616 550732 312644
rect 498988 312604 498994 312616
rect 550726 312604 550732 312616
rect 550784 312604 550790 312656
rect 456242 312536 456248 312588
rect 456300 312576 456306 312588
rect 518066 312576 518072 312588
rect 456300 312548 518072 312576
rect 456300 312536 456306 312548
rect 518066 312536 518072 312548
rect 518124 312536 518130 312588
rect 460566 311312 460572 311364
rect 460624 311352 460630 311364
rect 465166 311352 465172 311364
rect 460624 311324 465172 311352
rect 460624 311312 460630 311324
rect 465166 311312 465172 311324
rect 465224 311312 465230 311364
rect 461762 311244 461768 311296
rect 461820 311284 461826 311296
rect 463602 311284 463608 311296
rect 461820 311256 463608 311284
rect 461820 311244 461826 311256
rect 463602 311244 463608 311256
rect 463660 311244 463666 311296
rect 500586 311244 500592 311296
rect 500644 311284 500650 311296
rect 551002 311284 551008 311296
rect 500644 311256 551008 311284
rect 500644 311244 500650 311256
rect 551002 311244 551008 311256
rect 551060 311244 551066 311296
rect 458910 311176 458916 311228
rect 458968 311216 458974 311228
rect 494422 311216 494428 311228
rect 458968 311188 494428 311216
rect 458968 311176 458974 311188
rect 494422 311176 494428 311188
rect 494480 311176 494486 311228
rect 501874 311176 501880 311228
rect 501932 311216 501938 311228
rect 552474 311216 552480 311228
rect 501932 311188 552480 311216
rect 501932 311176 501938 311188
rect 552474 311176 552480 311188
rect 552532 311176 552538 311228
rect 456518 311108 456524 311160
rect 456576 311148 456582 311160
rect 558178 311148 558184 311160
rect 456576 311120 558184 311148
rect 456576 311108 456582 311120
rect 558178 311108 558184 311120
rect 558236 311108 558242 311160
rect 481542 310536 481548 310548
rect 480226 310508 481548 310536
rect 477218 310428 477224 310480
rect 477276 310468 477282 310480
rect 480226 310468 480254 310508
rect 481542 310496 481548 310508
rect 481600 310496 481606 310548
rect 477276 310440 480254 310468
rect 477276 310428 477282 310440
rect 443730 310088 443736 310140
rect 443788 310128 443794 310140
rect 448514 310128 448520 310140
rect 443788 310100 448520 310128
rect 443788 310088 443794 310100
rect 448514 310088 448520 310100
rect 448572 310088 448578 310140
rect 459094 309816 459100 309868
rect 459152 309856 459158 309868
rect 495434 309856 495440 309868
rect 459152 309828 495440 309856
rect 459152 309816 459158 309828
rect 495434 309816 495440 309828
rect 495492 309816 495498 309868
rect 501966 309816 501972 309868
rect 502024 309856 502030 309868
rect 552750 309856 552756 309868
rect 502024 309828 552756 309856
rect 502024 309816 502030 309828
rect 552750 309816 552756 309828
rect 552808 309816 552814 309868
rect 452194 309748 452200 309800
rect 452252 309788 452258 309800
rect 463970 309788 463976 309800
rect 452252 309760 463976 309788
rect 452252 309748 452258 309760
rect 463970 309748 463976 309760
rect 464028 309748 464034 309800
rect 477126 309748 477132 309800
rect 477184 309788 477190 309800
rect 562318 309788 562324 309800
rect 477184 309760 562324 309788
rect 477184 309748 477190 309760
rect 562318 309748 562324 309760
rect 562376 309748 562382 309800
rect 502058 308524 502064 308576
rect 502116 308564 502122 308576
rect 552290 308564 552296 308576
rect 502116 308536 552296 308564
rect 502116 308524 502122 308536
rect 552290 308524 552296 308536
rect 552348 308524 552354 308576
rect 497826 308456 497832 308508
rect 497884 308496 497890 308508
rect 549346 308496 549352 308508
rect 497884 308468 549352 308496
rect 497884 308456 497890 308468
rect 549346 308456 549352 308468
rect 549404 308456 549410 308508
rect 456610 308388 456616 308440
rect 456668 308428 456674 308440
rect 569218 308428 569224 308440
rect 456668 308400 569224 308428
rect 456668 308388 456674 308400
rect 569218 308388 569224 308400
rect 569276 308388 569282 308440
rect 457438 307776 457444 307828
rect 457496 307816 457502 307828
rect 462222 307816 462228 307828
rect 457496 307788 462228 307816
rect 457496 307776 457502 307788
rect 462222 307776 462228 307788
rect 462280 307776 462286 307828
rect 465718 307776 465724 307828
rect 465776 307816 465782 307828
rect 472710 307816 472716 307828
rect 465776 307788 472716 307816
rect 465776 307776 465782 307788
rect 472710 307776 472716 307788
rect 472768 307776 472774 307828
rect 433886 307708 433892 307760
rect 433944 307748 433950 307760
rect 439682 307748 439688 307760
rect 433944 307720 439688 307748
rect 433944 307708 433950 307720
rect 439682 307708 439688 307720
rect 439740 307708 439746 307760
rect 483750 307708 483756 307760
rect 483808 307748 483814 307760
rect 485038 307748 485044 307760
rect 483808 307720 485044 307748
rect 483808 307708 483814 307720
rect 485038 307708 485044 307720
rect 485096 307708 485102 307760
rect 488166 307164 488172 307216
rect 488224 307204 488230 307216
rect 529934 307204 529940 307216
rect 488224 307176 529940 307204
rect 488224 307164 488230 307176
rect 529934 307164 529940 307176
rect 529992 307164 529998 307216
rect 496630 307096 496636 307148
rect 496688 307136 496694 307148
rect 549254 307136 549260 307148
rect 496688 307108 549260 307136
rect 496688 307096 496694 307108
rect 549254 307096 549260 307108
rect 549312 307096 549318 307148
rect 478690 307028 478696 307080
rect 478748 307068 478754 307080
rect 544378 307068 544384 307080
rect 478748 307040 544384 307068
rect 478748 307028 478754 307040
rect 544378 307028 544384 307040
rect 544436 307028 544442 307080
rect 477218 306388 477224 306400
rect 474752 306360 477224 306388
rect 473354 306280 473360 306332
rect 473412 306320 473418 306332
rect 474752 306320 474780 306360
rect 477218 306348 477224 306360
rect 477276 306348 477282 306400
rect 473412 306292 474780 306320
rect 473412 306280 473418 306292
rect 458174 306076 458180 306128
rect 458232 306116 458238 306128
rect 461762 306116 461768 306128
rect 458232 306088 461768 306116
rect 458232 306076 458238 306088
rect 461762 306076 461768 306088
rect 461820 306076 461826 306128
rect 438118 306008 438124 306060
rect 438176 306048 438182 306060
rect 460566 306048 460572 306060
rect 438176 306020 460572 306048
rect 438176 306008 438182 306020
rect 460566 306008 460572 306020
rect 460624 306008 460630 306060
rect 473998 306008 474004 306060
rect 474056 306048 474062 306060
rect 484486 306048 484492 306060
rect 474056 306020 484492 306048
rect 474056 306008 474062 306020
rect 484486 306008 484492 306020
rect 484544 306008 484550 306060
rect 406470 305940 406476 305992
rect 406528 305980 406534 305992
rect 485958 305980 485964 305992
rect 406528 305952 485964 305980
rect 406528 305940 406534 305952
rect 485958 305940 485964 305952
rect 486016 305940 486022 305992
rect 383286 305872 383292 305924
rect 383344 305912 383350 305924
rect 443914 305912 443920 305924
rect 383344 305884 443920 305912
rect 383344 305872 383350 305884
rect 443914 305872 443920 305884
rect 443972 305872 443978 305924
rect 477310 305872 477316 305924
rect 477368 305912 477374 305924
rect 570598 305912 570604 305924
rect 477368 305884 570604 305912
rect 477368 305872 477374 305884
rect 570598 305872 570604 305884
rect 570656 305872 570662 305924
rect 403894 305804 403900 305856
rect 403952 305844 403958 305856
rect 511534 305844 511540 305856
rect 403952 305816 511540 305844
rect 403952 305804 403958 305816
rect 511534 305804 511540 305816
rect 511592 305804 511598 305856
rect 403710 305736 403716 305788
rect 403768 305776 403774 305788
rect 511166 305776 511172 305788
rect 403768 305748 511172 305776
rect 403768 305736 403774 305748
rect 511166 305736 511172 305748
rect 511224 305736 511230 305788
rect 380158 305668 380164 305720
rect 380216 305708 380222 305720
rect 512638 305708 512644 305720
rect 380216 305680 512644 305708
rect 380216 305668 380222 305680
rect 512638 305668 512644 305680
rect 512696 305668 512702 305720
rect 380250 305600 380256 305652
rect 380308 305640 380314 305652
rect 512362 305640 512368 305652
rect 380308 305612 512368 305640
rect 380308 305600 380314 305612
rect 512362 305600 512368 305612
rect 512420 305600 512426 305652
rect 438210 304988 438216 305040
rect 438268 305028 438274 305040
rect 440970 305028 440976 305040
rect 438268 305000 440976 305028
rect 438268 304988 438274 305000
rect 440970 304988 440976 305000
rect 441028 304988 441034 305040
rect 488258 304512 488264 304564
rect 488316 304552 488322 304564
rect 531406 304552 531412 304564
rect 488316 304524 531412 304552
rect 488316 304512 488322 304524
rect 531406 304512 531412 304524
rect 531464 304512 531470 304564
rect 410518 304444 410524 304496
rect 410576 304484 410582 304496
rect 514938 304484 514944 304496
rect 410576 304456 514944 304484
rect 410576 304444 410582 304456
rect 514938 304444 514944 304456
rect 514996 304444 515002 304496
rect 382274 304376 382280 304428
rect 382332 304416 382338 304428
rect 442258 304416 442264 304428
rect 382332 304388 442264 304416
rect 382332 304376 382338 304388
rect 442258 304376 442264 304388
rect 442316 304376 442322 304428
rect 448422 304376 448428 304428
rect 448480 304416 448486 304428
rect 458174 304416 458180 304428
rect 448480 304388 458180 304416
rect 448480 304376 448486 304388
rect 458174 304376 458180 304388
rect 458232 304376 458238 304428
rect 467374 304376 467380 304428
rect 467432 304416 467438 304428
rect 573358 304416 573364 304428
rect 467432 304388 573364 304416
rect 467432 304376 467438 304388
rect 573358 304376 573364 304388
rect 573416 304376 573422 304428
rect 407942 304308 407948 304360
rect 408000 304348 408006 304360
rect 516226 304348 516232 304360
rect 408000 304320 516232 304348
rect 408000 304308 408006 304320
rect 516226 304308 516232 304320
rect 516284 304308 516290 304360
rect 381538 304240 381544 304292
rect 381596 304280 381602 304292
rect 512454 304280 512460 304292
rect 381596 304252 512460 304280
rect 381596 304240 381602 304252
rect 512454 304240 512460 304252
rect 512512 304240 512518 304292
rect 481266 303764 481272 303816
rect 481324 303804 481330 303816
rect 483750 303804 483756 303816
rect 481324 303776 483756 303804
rect 481324 303764 481330 303776
rect 483750 303764 483756 303776
rect 483808 303764 483814 303816
rect 472710 303628 472716 303680
rect 472768 303668 472774 303680
rect 475010 303668 475016 303680
rect 472768 303640 475016 303668
rect 472768 303628 472774 303640
rect 475010 303628 475016 303640
rect 475068 303628 475074 303680
rect 401134 303560 401140 303612
rect 401192 303600 401198 303612
rect 510890 303600 510896 303612
rect 401192 303572 510896 303600
rect 401192 303560 401198 303572
rect 510890 303560 510896 303572
rect 510948 303560 510954 303612
rect 404078 303492 404084 303544
rect 404136 303532 404142 303544
rect 514110 303532 514116 303544
rect 404136 303504 514116 303532
rect 404136 303492 404142 303504
rect 514110 303492 514116 303504
rect 514168 303492 514174 303544
rect 403986 303424 403992 303476
rect 404044 303464 404050 303476
rect 515306 303464 515312 303476
rect 404044 303436 515312 303464
rect 404044 303424 404050 303436
rect 515306 303424 515312 303436
rect 515364 303424 515370 303476
rect 403802 303356 403808 303408
rect 403860 303396 403866 303408
rect 515582 303396 515588 303408
rect 403860 303368 515588 303396
rect 403860 303356 403866 303368
rect 515582 303356 515588 303368
rect 515640 303356 515646 303408
rect 401318 303288 401324 303340
rect 401376 303328 401382 303340
rect 513834 303328 513840 303340
rect 401376 303300 513840 303328
rect 401376 303288 401382 303300
rect 513834 303288 513840 303300
rect 513892 303288 513898 303340
rect 401226 303220 401232 303272
rect 401284 303260 401290 303272
rect 513742 303260 513748 303272
rect 401284 303232 513748 303260
rect 401284 303220 401290 303232
rect 513742 303220 513748 303232
rect 513800 303220 513806 303272
rect 398098 303152 398104 303204
rect 398156 303192 398162 303204
rect 510706 303192 510712 303204
rect 398156 303164 510712 303192
rect 398156 303152 398162 303164
rect 510706 303152 510712 303164
rect 510764 303152 510770 303204
rect 401042 303084 401048 303136
rect 401100 303124 401106 303136
rect 515122 303124 515128 303136
rect 401100 303096 515128 303124
rect 401100 303084 401106 303096
rect 515122 303084 515128 303096
rect 515180 303084 515186 303136
rect 400950 303016 400956 303068
rect 401008 303056 401014 303068
rect 515214 303056 515220 303068
rect 401008 303028 515220 303056
rect 401008 303016 401014 303028
rect 515214 303016 515220 303028
rect 515272 303016 515278 303068
rect 381722 302948 381728 303000
rect 381780 302988 381786 303000
rect 512086 302988 512092 303000
rect 381780 302960 512092 302988
rect 381780 302948 381786 302960
rect 512086 302948 512092 302960
rect 512144 302948 512150 303000
rect 381630 302880 381636 302932
rect 381688 302920 381694 302932
rect 511994 302920 512000 302932
rect 381688 302892 512000 302920
rect 381688 302880 381694 302892
rect 511994 302880 512000 302892
rect 512052 302880 512058 302932
rect 456702 302812 456708 302864
rect 456760 302852 456766 302864
rect 555418 302852 555424 302864
rect 456760 302824 555424 302852
rect 456760 302812 456766 302824
rect 555418 302812 555424 302824
rect 555476 302812 555482 302864
rect 400858 302744 400864 302796
rect 400916 302784 400922 302796
rect 465350 302784 465356 302796
rect 400916 302756 465356 302784
rect 400916 302744 400922 302756
rect 465350 302744 465356 302756
rect 465408 302744 465414 302796
rect 440970 302404 440976 302456
rect 441028 302444 441034 302456
rect 443730 302444 443736 302456
rect 441028 302416 443736 302444
rect 441028 302404 441034 302416
rect 443730 302404 443736 302416
rect 443788 302404 443794 302456
rect 446490 302200 446496 302252
rect 446548 302240 446554 302252
rect 448422 302240 448428 302252
rect 446548 302212 448428 302240
rect 446548 302200 446554 302212
rect 448422 302200 448428 302212
rect 448480 302200 448486 302252
rect 478138 302200 478144 302252
rect 478196 302240 478202 302252
rect 479610 302240 479616 302252
rect 478196 302212 479616 302240
rect 478196 302200 478202 302212
rect 479610 302200 479616 302212
rect 479668 302200 479674 302252
rect 3602 302064 3608 302116
rect 3660 302104 3666 302116
rect 4890 302104 4896 302116
rect 3660 302076 4896 302104
rect 3660 302064 3666 302076
rect 4890 302064 4896 302076
rect 4948 302064 4954 302116
rect 477494 301928 477500 301980
rect 477552 301968 477558 301980
rect 481266 301968 481272 301980
rect 477552 301940 481272 301968
rect 477552 301928 477558 301940
rect 481266 301928 481272 301940
rect 481324 301928 481330 301980
rect 457898 301452 457904 301504
rect 457956 301492 457962 301504
rect 536098 301492 536104 301504
rect 457956 301464 536104 301492
rect 457956 301452 457962 301464
rect 536098 301452 536104 301464
rect 536156 301452 536162 301504
rect 395338 300772 395344 300824
rect 395396 300812 395402 300824
rect 510246 300812 510252 300824
rect 395396 300784 510252 300812
rect 395396 300772 395402 300784
rect 510246 300772 510252 300784
rect 510304 300772 510310 300824
rect 395706 300704 395712 300756
rect 395764 300744 395770 300756
rect 509878 300744 509884 300756
rect 395764 300716 509884 300744
rect 395764 300704 395770 300716
rect 509878 300704 509884 300716
rect 509936 300704 509942 300756
rect 398374 300636 398380 300688
rect 398432 300676 398438 300688
rect 515030 300676 515036 300688
rect 398432 300648 515036 300676
rect 398432 300636 398438 300648
rect 515030 300636 515036 300648
rect 515088 300636 515094 300688
rect 392670 300568 392676 300620
rect 392728 300608 392734 300620
rect 510338 300608 510344 300620
rect 392728 300580 510344 300608
rect 392728 300568 392734 300580
rect 510338 300568 510344 300580
rect 510396 300568 510402 300620
rect 395522 300500 395528 300552
rect 395580 300540 395586 300552
rect 513558 300540 513564 300552
rect 395580 300512 513564 300540
rect 395580 300500 395586 300512
rect 513558 300500 513564 300512
rect 513616 300500 513622 300552
rect 398282 300432 398288 300484
rect 398340 300472 398346 300484
rect 517698 300472 517704 300484
rect 398340 300444 517704 300472
rect 398340 300432 398346 300444
rect 517698 300432 517704 300444
rect 517756 300432 517762 300484
rect 395798 300364 395804 300416
rect 395856 300404 395862 300416
rect 516318 300404 516324 300416
rect 395856 300376 516324 300404
rect 395856 300364 395862 300376
rect 516318 300364 516324 300376
rect 516376 300364 516382 300416
rect 392578 300296 392584 300348
rect 392636 300336 392642 300348
rect 514202 300336 514208 300348
rect 392636 300308 514208 300336
rect 392636 300296 392642 300308
rect 514202 300296 514208 300308
rect 514260 300296 514266 300348
rect 395614 300228 395620 300280
rect 395672 300268 395678 300280
rect 517606 300268 517612 300280
rect 395672 300240 517612 300268
rect 395672 300228 395678 300240
rect 517606 300228 517612 300240
rect 517664 300228 517670 300280
rect 395430 300160 395436 300212
rect 395488 300200 395494 300212
rect 517514 300200 517520 300212
rect 395488 300172 517520 300200
rect 395488 300160 395494 300172
rect 517514 300160 517520 300172
rect 517572 300160 517578 300212
rect 392762 300092 392768 300144
rect 392820 300132 392826 300144
rect 516870 300132 516876 300144
rect 392820 300104 516876 300132
rect 392820 300092 392826 300104
rect 516870 300092 516876 300104
rect 516928 300092 516934 300144
rect 448054 300024 448060 300076
rect 448112 300064 448118 300076
rect 546494 300064 546500 300076
rect 448112 300036 546500 300064
rect 448112 300024 448118 300036
rect 546494 300024 546500 300036
rect 546552 300024 546558 300076
rect 477402 299956 477408 300008
rect 477460 299996 477466 300008
rect 559558 299996 559564 300008
rect 477460 299968 559564 299996
rect 477460 299956 477466 299968
rect 559558 299956 559564 299968
rect 559616 299956 559622 300008
rect 461578 299412 461584 299464
rect 461636 299452 461642 299464
rect 580166 299452 580172 299464
rect 461636 299424 580172 299452
rect 461636 299412 461642 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 435450 299344 435456 299396
rect 435508 299384 435514 299396
rect 438210 299384 438216 299396
rect 435508 299356 438216 299384
rect 435508 299344 435514 299356
rect 438210 299344 438216 299356
rect 438268 299344 438274 299396
rect 470594 298936 470600 298988
rect 470652 298976 470658 298988
rect 473354 298976 473360 298988
rect 470652 298948 473360 298976
rect 470652 298936 470658 298948
rect 473354 298936 473360 298948
rect 473412 298936 473418 298988
rect 475102 298936 475108 298988
rect 475160 298976 475166 298988
rect 477494 298976 477500 298988
rect 475160 298948 477500 298976
rect 475160 298936 475166 298948
rect 477494 298936 477500 298948
rect 477552 298936 477558 298988
rect 387426 298052 387432 298104
rect 387484 298092 387490 298104
rect 510614 298092 510620 298104
rect 387484 298064 510620 298092
rect 387484 298052 387490 298064
rect 510614 298052 510620 298064
rect 510672 298052 510678 298104
rect 390094 297984 390100 298036
rect 390152 298024 390158 298036
rect 516594 298024 516600 298036
rect 390152 297996 516600 298024
rect 390152 297984 390158 297996
rect 516594 297984 516600 297996
rect 516652 297984 516658 298036
rect 390186 297916 390192 297968
rect 390244 297956 390250 297968
rect 516686 297956 516692 297968
rect 390244 297928 516692 297956
rect 390244 297916 390250 297928
rect 516686 297916 516692 297928
rect 516744 297916 516750 297968
rect 390278 297848 390284 297900
rect 390336 297888 390342 297900
rect 517974 297888 517980 297900
rect 390336 297860 517980 297888
rect 390336 297848 390342 297860
rect 517974 297848 517980 297860
rect 518032 297848 518038 297900
rect 390002 297780 390008 297832
rect 390060 297820 390066 297832
rect 517882 297820 517888 297832
rect 390060 297792 517888 297820
rect 390060 297780 390066 297792
rect 517882 297780 517888 297792
rect 517940 297780 517946 297832
rect 389910 297712 389916 297764
rect 389968 297752 389974 297764
rect 517790 297752 517796 297764
rect 389968 297724 517796 297752
rect 389968 297712 389974 297724
rect 517790 297712 517796 297724
rect 517848 297712 517854 297764
rect 387518 297644 387524 297696
rect 387576 297684 387582 297696
rect 519262 297684 519268 297696
rect 387576 297656 519268 297684
rect 387576 297644 387582 297656
rect 519262 297644 519268 297656
rect 519320 297644 519326 297696
rect 387242 297576 387248 297628
rect 387300 297616 387306 297628
rect 519078 297616 519084 297628
rect 387300 297588 519084 297616
rect 387300 297576 387306 297588
rect 519078 297576 519084 297588
rect 519136 297576 519142 297628
rect 387150 297508 387156 297560
rect 387208 297548 387214 297560
rect 519170 297548 519176 297560
rect 387208 297520 519176 297548
rect 387208 297508 387214 297520
rect 519170 297508 519176 297520
rect 519228 297508 519234 297560
rect 387334 297440 387340 297492
rect 387392 297480 387398 297492
rect 519446 297480 519452 297492
rect 387392 297452 519452 297480
rect 387392 297440 387398 297452
rect 519446 297440 519452 297452
rect 519504 297440 519510 297492
rect 387058 297372 387064 297424
rect 387116 297412 387122 297424
rect 520826 297412 520832 297424
rect 387116 297384 520832 297412
rect 387116 297372 387122 297384
rect 520826 297372 520832 297384
rect 520884 297372 520890 297424
rect 452102 297304 452108 297356
rect 452160 297344 452166 297356
rect 457438 297344 457444 297356
rect 452160 297316 457444 297344
rect 452160 297304 452166 297316
rect 457438 297304 457444 297316
rect 457496 297304 457502 297356
rect 457990 297304 457996 297356
rect 458048 297344 458054 297356
rect 533338 297344 533344 297356
rect 458048 297316 533344 297344
rect 458048 297304 458054 297316
rect 533338 297304 533344 297316
rect 533396 297304 533402 297356
rect 457806 296012 457812 296064
rect 457864 296052 457870 296064
rect 537478 296052 537484 296064
rect 457864 296024 537484 296052
rect 457864 296012 457870 296024
rect 537478 296012 537484 296024
rect 537536 296012 537542 296064
rect 380342 295944 380348 295996
rect 380400 295984 380406 295996
rect 512270 295984 512276 295996
rect 380400 295956 512276 295984
rect 380400 295944 380406 295956
rect 512270 295944 512276 295956
rect 512328 295944 512334 295996
rect 394326 295264 394332 295316
rect 394384 295304 394390 295316
rect 513466 295304 513472 295316
rect 394384 295276 513472 295304
rect 394384 295264 394390 295276
rect 513466 295264 513472 295276
rect 513524 295264 513530 295316
rect 393958 295196 393964 295248
rect 394016 295236 394022 295248
rect 513374 295236 513380 295248
rect 394016 295208 513380 295236
rect 394016 295196 394022 295208
rect 513374 295196 513380 295208
rect 513432 295196 513438 295248
rect 399478 295128 399484 295180
rect 399536 295168 399542 295180
rect 520274 295168 520280 295180
rect 399536 295140 520280 295168
rect 399536 295128 399542 295140
rect 520274 295128 520280 295140
rect 520332 295128 520338 295180
rect 382918 295060 382924 295112
rect 382976 295100 382982 295112
rect 508498 295100 508504 295112
rect 382976 295072 508504 295100
rect 382976 295060 382982 295072
rect 508498 295060 508504 295072
rect 508556 295060 508562 295112
rect 384390 294992 384396 295044
rect 384448 295032 384454 295044
rect 516962 295032 516968 295044
rect 384448 295004 516968 295032
rect 384448 294992 384454 295004
rect 516962 294992 516968 295004
rect 517020 294992 517026 295044
rect 381814 294924 381820 294976
rect 381872 294964 381878 294976
rect 514846 294964 514852 294976
rect 381872 294936 514852 294964
rect 381872 294924 381878 294936
rect 514846 294924 514852 294936
rect 514904 294924 514910 294976
rect 384574 294856 384580 294908
rect 384632 294896 384638 294908
rect 518986 294896 518992 294908
rect 384632 294868 518992 294896
rect 384632 294856 384638 294868
rect 518986 294856 518992 294868
rect 519044 294856 519050 294908
rect 384482 294788 384488 294840
rect 384540 294828 384546 294840
rect 520734 294828 520740 294840
rect 384540 294800 520740 294828
rect 384540 294788 384546 294800
rect 520734 294788 520740 294800
rect 520792 294788 520798 294840
rect 381906 294720 381912 294772
rect 381964 294760 381970 294772
rect 518894 294760 518900 294772
rect 381964 294732 518900 294760
rect 381964 294720 381970 294732
rect 518894 294720 518900 294732
rect 518952 294720 518958 294772
rect 383010 294652 383016 294704
rect 383068 294692 383074 294704
rect 520366 294692 520372 294704
rect 383068 294664 520372 294692
rect 383068 294652 383074 294664
rect 520366 294652 520372 294664
rect 520424 294652 520430 294704
rect 381998 294584 382004 294636
rect 382056 294624 382062 294636
rect 520642 294624 520648 294636
rect 382056 294596 520648 294624
rect 382056 294584 382062 294596
rect 520642 294584 520648 294596
rect 520700 294584 520706 294636
rect 478506 294516 478512 294568
rect 478564 294556 478570 294568
rect 540238 294556 540244 294568
rect 478564 294528 540244 294556
rect 478564 294516 478570 294528
rect 540238 294516 540244 294528
rect 540296 294516 540302 294568
rect 457438 294448 457444 294500
rect 457496 294488 457502 294500
rect 492950 294488 492956 294500
rect 457496 294460 492956 294488
rect 457496 294448 457502 294460
rect 492950 294448 492956 294460
rect 493008 294448 493014 294500
rect 444374 294244 444380 294296
rect 444432 294284 444438 294296
rect 446490 294284 446496 294296
rect 444432 294256 446496 294284
rect 444432 294244 444438 294256
rect 446490 294244 446496 294256
rect 446548 294244 446554 294296
rect 399754 293292 399760 293344
rect 399812 293332 399818 293344
rect 485866 293332 485872 293344
rect 399812 293304 485872 293332
rect 399812 293292 399818 293304
rect 485866 293292 485872 293304
rect 485924 293292 485930 293344
rect 488350 293292 488356 293344
rect 488408 293332 488414 293344
rect 531314 293332 531320 293344
rect 488408 293304 531320 293332
rect 488408 293292 488414 293304
rect 531314 293292 531320 293304
rect 531372 293292 531378 293344
rect 440234 293224 440240 293276
rect 440292 293264 440298 293276
rect 444374 293264 444380 293276
rect 440292 293236 444380 293264
rect 440292 293224 440298 293236
rect 444374 293224 444380 293236
rect 444432 293224 444438 293276
rect 467466 293224 467472 293276
rect 467524 293264 467530 293276
rect 576118 293264 576124 293276
rect 467524 293236 576124 293264
rect 467524 293224 467530 293236
rect 576118 293224 576124 293236
rect 576176 293224 576182 293276
rect 471974 292544 471980 292596
rect 472032 292584 472038 292596
rect 475102 292584 475108 292596
rect 472032 292556 475108 292584
rect 472032 292544 472038 292556
rect 475102 292544 475108 292556
rect 475160 292544 475166 292596
rect 476758 292544 476764 292596
rect 476816 292584 476822 292596
rect 478138 292584 478144 292596
rect 476816 292556 478144 292584
rect 476816 292544 476822 292556
rect 478138 292544 478144 292556
rect 478196 292544 478202 292596
rect 397086 292476 397092 292528
rect 397144 292516 397150 292528
rect 514754 292516 514760 292528
rect 397144 292488 514760 292516
rect 397144 292476 397150 292488
rect 514754 292476 514760 292488
rect 514812 292476 514818 292528
rect 383194 292408 383200 292460
rect 383252 292448 383258 292460
rect 510154 292448 510160 292460
rect 383252 292420 510160 292448
rect 383252 292408 383258 292420
rect 510154 292408 510160 292420
rect 510212 292408 510218 292460
rect 388530 292340 388536 292392
rect 388588 292380 388594 292392
rect 516410 292380 516416 292392
rect 388588 292352 516416 292380
rect 388588 292340 388594 292352
rect 516410 292340 516416 292352
rect 516468 292340 516474 292392
rect 385954 292272 385960 292324
rect 386012 292312 386018 292324
rect 516502 292312 516508 292324
rect 386012 292284 516508 292312
rect 386012 292272 386018 292284
rect 516502 292272 516508 292284
rect 516560 292272 516566 292324
rect 391382 292204 391388 292256
rect 391440 292244 391446 292256
rect 522022 292244 522028 292256
rect 391440 292216 522028 292244
rect 391440 292204 391446 292216
rect 522022 292204 522028 292216
rect 522080 292204 522086 292256
rect 388622 292136 388628 292188
rect 388680 292176 388686 292188
rect 519354 292176 519360 292188
rect 388680 292148 519360 292176
rect 388680 292136 388686 292148
rect 519354 292136 519360 292148
rect 519412 292136 519418 292188
rect 383102 292068 383108 292120
rect 383160 292108 383166 292120
rect 513926 292108 513932 292120
rect 383160 292080 513932 292108
rect 383160 292068 383166 292080
rect 513926 292068 513932 292080
rect 513984 292068 513990 292120
rect 391290 292000 391296 292052
rect 391348 292040 391354 292052
rect 522206 292040 522212 292052
rect 391348 292012 522212 292040
rect 391348 292000 391354 292012
rect 522206 292000 522212 292012
rect 522264 292000 522270 292052
rect 391198 291932 391204 291984
rect 391256 291972 391262 291984
rect 522114 291972 522120 291984
rect 391256 291944 522120 291972
rect 391256 291932 391262 291944
rect 522114 291932 522120 291944
rect 522172 291932 522178 291984
rect 385770 291864 385776 291916
rect 385828 291904 385834 291916
rect 519630 291904 519636 291916
rect 385828 291876 519636 291904
rect 385828 291864 385834 291876
rect 519630 291864 519636 291876
rect 519688 291864 519694 291916
rect 385678 291796 385684 291848
rect 385736 291836 385742 291848
rect 519722 291836 519728 291848
rect 385736 291808 519728 291836
rect 385736 291796 385742 291808
rect 519722 291796 519728 291808
rect 519780 291796 519786 291848
rect 467558 291728 467564 291780
rect 467616 291768 467622 291780
rect 574738 291768 574744 291780
rect 467616 291740 574744 291768
rect 467616 291728 467622 291740
rect 574738 291728 574744 291740
rect 574796 291728 574802 291780
rect 396718 291660 396724 291712
rect 396776 291700 396782 291712
rect 486050 291700 486056 291712
rect 396776 291672 486056 291700
rect 396776 291660 396782 291672
rect 486050 291660 486056 291672
rect 486108 291660 486114 291712
rect 466362 290436 466368 290488
rect 466420 290476 466426 290488
rect 571978 290476 571984 290488
rect 466420 290448 571984 290476
rect 466420 290436 466426 290448
rect 571978 290436 571984 290448
rect 572036 290436 572042 290488
rect 468478 290368 468484 290420
rect 468536 290408 468542 290420
rect 470502 290408 470508 290420
rect 468536 290380 470508 290408
rect 468536 290368 468542 290380
rect 470502 290368 470508 290380
rect 470560 290368 470566 290420
rect 405090 289756 405096 289808
rect 405148 289796 405154 289808
rect 523034 289796 523040 289808
rect 405148 289768 523040 289796
rect 405148 289756 405154 289768
rect 523034 289756 523040 289768
rect 523092 289756 523098 289808
rect 402238 289688 402244 289740
rect 402296 289728 402302 289740
rect 523126 289728 523132 289740
rect 402296 289700 523132 289728
rect 402296 289688 402302 289700
rect 523126 289688 523132 289700
rect 523184 289688 523190 289740
rect 399846 289620 399852 289672
rect 399904 289660 399910 289672
rect 523218 289660 523224 289672
rect 399904 289632 523224 289660
rect 399904 289620 399910 289632
rect 523218 289620 523224 289632
rect 523276 289620 523282 289672
rect 396902 289552 396908 289604
rect 396960 289592 396966 289604
rect 520458 289592 520464 289604
rect 396960 289564 520464 289592
rect 396960 289552 396966 289564
rect 520458 289552 520464 289564
rect 520516 289552 520522 289604
rect 396994 289484 397000 289536
rect 397052 289524 397058 289536
rect 520550 289524 520556 289536
rect 397052 289496 520556 289524
rect 397052 289484 397058 289496
rect 520550 289484 520556 289496
rect 520608 289484 520614 289536
rect 399662 289416 399668 289468
rect 399720 289456 399726 289468
rect 523402 289456 523408 289468
rect 399720 289428 523408 289456
rect 399720 289416 399726 289428
rect 523402 289416 523408 289428
rect 523460 289416 523466 289468
rect 399570 289348 399576 289400
rect 399628 289388 399634 289400
rect 523310 289388 523316 289400
rect 399628 289360 523316 289388
rect 399628 289348 399634 289360
rect 523310 289348 523316 289360
rect 523368 289348 523374 289400
rect 396810 289280 396816 289332
rect 396868 289320 396874 289332
rect 521654 289320 521660 289332
rect 396868 289292 521660 289320
rect 396868 289280 396874 289292
rect 521654 289280 521660 289292
rect 521712 289280 521718 289332
rect 394234 289212 394240 289264
rect 394292 289252 394298 289264
rect 521838 289252 521844 289264
rect 394292 289224 521844 289252
rect 394292 289212 394298 289224
rect 521838 289212 521844 289224
rect 521896 289212 521902 289264
rect 394142 289144 394148 289196
rect 394200 289184 394206 289196
rect 521746 289184 521752 289196
rect 394200 289156 521752 289184
rect 394200 289144 394206 289156
rect 521746 289144 521752 289156
rect 521804 289144 521810 289196
rect 394050 289076 394056 289128
rect 394108 289116 394114 289128
rect 521930 289116 521936 289128
rect 394108 289088 521936 289116
rect 394108 289076 394114 289088
rect 521930 289076 521936 289088
rect 521988 289076 521994 289128
rect 404998 289008 405004 289060
rect 405056 289048 405062 289060
rect 520918 289048 520924 289060
rect 405056 289020 520924 289048
rect 405056 289008 405062 289020
rect 520918 289008 520924 289020
rect 520976 289008 520982 289060
rect 432690 288940 432696 288992
rect 432748 288980 432754 288992
rect 435450 288980 435456 288992
rect 432748 288952 435456 288980
rect 432748 288940 432754 288952
rect 435450 288940 435456 288952
rect 435508 288940 435514 288992
rect 479518 288940 479524 288992
rect 479576 288980 479582 288992
rect 580350 288980 580356 288992
rect 479576 288952 580356 288980
rect 479576 288940 479582 288952
rect 580350 288940 580356 288952
rect 580408 288940 580414 288992
rect 471882 288436 471888 288448
rect 470566 288408 471888 288436
rect 467834 288328 467840 288380
rect 467892 288368 467898 288380
rect 470566 288368 470594 288408
rect 471882 288396 471888 288408
rect 471940 288396 471946 288448
rect 467892 288340 470594 288368
rect 467892 288328 467898 288340
rect 467650 287648 467656 287700
rect 467708 287688 467714 287700
rect 580258 287688 580264 287700
rect 467708 287660 580264 287688
rect 467708 287648 467714 287660
rect 580258 287648 580264 287660
rect 580316 287648 580322 287700
rect 440234 287076 440240 287088
rect 437584 287048 440240 287076
rect 436922 286968 436928 287020
rect 436980 287008 436986 287020
rect 437584 287008 437612 287048
rect 440234 287036 440240 287048
rect 440292 287036 440298 287088
rect 436980 286980 437612 287008
rect 436980 286968 436986 286980
rect 403618 286424 403624 286476
rect 403676 286464 403682 286476
rect 476206 286464 476212 286476
rect 403676 286436 476212 286464
rect 403676 286424 403682 286436
rect 476206 286424 476212 286436
rect 476264 286424 476270 286476
rect 407850 286356 407856 286408
rect 407908 286396 407914 286408
rect 523586 286396 523592 286408
rect 407908 286368 523592 286396
rect 407908 286356 407914 286368
rect 523586 286356 523592 286368
rect 523644 286356 523650 286408
rect 405182 286288 405188 286340
rect 405240 286328 405246 286340
rect 523494 286328 523500 286340
rect 405240 286300 523500 286328
rect 405240 286288 405246 286300
rect 523494 286288 523500 286300
rect 523552 286288 523558 286340
rect 449158 285676 449164 285728
rect 449216 285716 449222 285728
rect 452194 285716 452200 285728
rect 449216 285688 452200 285716
rect 449216 285676 449222 285688
rect 452194 285676 452200 285688
rect 452252 285676 452258 285728
rect 461670 285676 461676 285728
rect 461728 285716 461734 285728
rect 465810 285716 465816 285728
rect 461728 285688 465816 285716
rect 461728 285676 461734 285688
rect 465810 285676 465816 285688
rect 465868 285676 465874 285728
rect 467834 285716 467840 285728
rect 466472 285688 467840 285716
rect 466178 285608 466184 285660
rect 466236 285648 466242 285660
rect 466472 285648 466500 285688
rect 467834 285676 467840 285688
rect 467892 285676 467898 285728
rect 471514 285676 471520 285728
rect 471572 285716 471578 285728
rect 473998 285716 474004 285728
rect 471572 285688 474004 285716
rect 471572 285676 471578 285688
rect 473998 285676 474004 285688
rect 474056 285676 474062 285728
rect 466236 285620 466500 285648
rect 466236 285608 466242 285620
rect 469858 284724 469864 284776
rect 469916 284764 469922 284776
rect 472618 284764 472624 284776
rect 469916 284736 472624 284764
rect 469916 284724 469922 284736
rect 472618 284724 472624 284736
rect 472676 284724 472682 284776
rect 466454 284316 466460 284368
rect 466512 284356 466518 284368
rect 468478 284356 468484 284368
rect 466512 284328 468484 284356
rect 466512 284316 466518 284328
rect 468478 284316 468484 284328
rect 468536 284316 468542 284368
rect 436646 283636 436652 283688
rect 436704 283676 436710 283688
rect 461670 283676 461676 283688
rect 436704 283648 461676 283676
rect 436704 283636 436710 283648
rect 461670 283636 461676 283648
rect 461728 283636 461734 283688
rect 457714 283568 457720 283620
rect 457772 283608 457778 283620
rect 494330 283608 494336 283620
rect 457772 283580 494336 283608
rect 457772 283568 457778 283580
rect 494330 283568 494336 283580
rect 494388 283568 494394 283620
rect 439682 282140 439688 282192
rect 439740 282180 439746 282192
rect 472710 282180 472716 282192
rect 439740 282152 472716 282180
rect 439740 282140 439746 282152
rect 472710 282140 472716 282152
rect 472768 282140 472774 282192
rect 464338 282072 464344 282124
rect 464396 282112 464402 282124
rect 466178 282112 466184 282124
rect 464396 282084 466184 282112
rect 464396 282072 464402 282084
rect 466178 282072 466184 282084
rect 466236 282072 466242 282124
rect 382274 281460 382280 281512
rect 382332 281500 382338 281512
rect 439590 281500 439596 281512
rect 382332 281472 439596 281500
rect 382332 281460 382338 281472
rect 439590 281460 439596 281472
rect 439648 281460 439654 281512
rect 406654 280780 406660 280832
rect 406712 280820 406718 280832
rect 436646 280820 436652 280832
rect 406712 280792 436652 280820
rect 406712 280780 406718 280792
rect 436646 280780 436652 280792
rect 436704 280780 436710 280832
rect 467742 280780 467748 280832
rect 467800 280820 467806 280832
rect 543090 280820 543096 280832
rect 467800 280792 543096 280820
rect 467800 280780 467806 280792
rect 543090 280780 543096 280792
rect 543148 280780 543154 280832
rect 457806 279420 457812 279472
rect 457864 279460 457870 279472
rect 494238 279460 494244 279472
rect 457864 279432 494244 279460
rect 457864 279420 457870 279432
rect 494238 279420 494244 279432
rect 494296 279420 494302 279472
rect 458082 278060 458088 278112
rect 458140 278100 458146 278112
rect 466362 278100 466368 278112
rect 458140 278072 466368 278100
rect 458140 278060 458146 278072
rect 466362 278060 466368 278072
rect 466420 278060 466426 278112
rect 488442 278060 488448 278112
rect 488500 278100 488506 278112
rect 530026 278100 530032 278112
rect 488500 278072 530032 278100
rect 488500 278060 488506 278072
rect 530026 278060 530032 278072
rect 530084 278060 530090 278112
rect 459554 277992 459560 278044
rect 459612 278032 459618 278044
rect 471514 278032 471520 278044
rect 459612 278004 471520 278032
rect 459612 277992 459618 278004
rect 471514 277992 471520 278004
rect 471572 277992 471578 278044
rect 500678 277992 500684 278044
rect 500736 278032 500742 278044
rect 551186 278032 551192 278044
rect 500736 278004 551192 278032
rect 500736 277992 500742 278004
rect 551186 277992 551192 278004
rect 551244 277992 551250 278044
rect 400214 276632 400220 276684
rect 400272 276672 400278 276684
rect 406654 276672 406660 276684
rect 400272 276644 406660 276672
rect 400272 276632 400278 276644
rect 406654 276632 406660 276644
rect 406712 276632 406718 276684
rect 457622 276632 457628 276684
rect 457680 276672 457686 276684
rect 492858 276672 492864 276684
rect 457680 276644 492864 276672
rect 457680 276632 457686 276644
rect 492858 276632 492864 276644
rect 492916 276632 492922 276684
rect 445754 276020 445760 276072
rect 445812 276060 445818 276072
rect 449158 276060 449164 276072
rect 445812 276032 449164 276060
rect 445812 276020 445818 276032
rect 449158 276020 449164 276032
rect 449216 276020 449222 276072
rect 458174 275408 458180 275460
rect 458232 275448 458238 275460
rect 464338 275448 464344 275460
rect 458232 275420 464344 275448
rect 458232 275408 458238 275420
rect 464338 275408 464344 275420
rect 464396 275408 464402 275460
rect 460658 275340 460664 275392
rect 460716 275380 460722 275392
rect 490190 275380 490196 275392
rect 460716 275352 490196 275380
rect 460716 275340 460722 275352
rect 490190 275340 490196 275352
rect 490248 275340 490254 275392
rect 380434 275272 380440 275324
rect 380492 275312 380498 275324
rect 512822 275312 512828 275324
rect 380492 275284 512828 275312
rect 380492 275272 380498 275284
rect 512822 275272 512828 275284
rect 512880 275272 512886 275324
rect 435542 275000 435548 275052
rect 435600 275040 435606 275052
rect 440970 275040 440976 275052
rect 435600 275012 440976 275040
rect 435600 275000 435606 275012
rect 440970 275000 440976 275012
rect 441028 275000 441034 275052
rect 482462 274660 482468 274712
rect 482520 274700 482526 274712
rect 484670 274700 484676 274712
rect 482520 274672 484676 274700
rect 482520 274660 482526 274672
rect 484670 274660 484676 274672
rect 484728 274660 484734 274712
rect 452562 274116 452568 274168
rect 452620 274156 452626 274168
rect 458082 274156 458088 274168
rect 452620 274128 458088 274156
rect 452620 274116 452626 274128
rect 458082 274116 458088 274128
rect 458140 274116 458146 274168
rect 460566 273980 460572 274032
rect 460624 274020 460630 274032
rect 488902 274020 488908 274032
rect 460624 273992 488908 274020
rect 460624 273980 460630 273992
rect 488902 273980 488908 273992
rect 488960 273980 488966 274032
rect 431218 273912 431224 273964
rect 431276 273952 431282 273964
rect 438118 273952 438124 273964
rect 431276 273924 438124 273952
rect 431276 273912 431282 273924
rect 438118 273912 438124 273924
rect 438176 273912 438182 273964
rect 457530 273912 457536 273964
rect 457588 273952 457594 273964
rect 490098 273952 490104 273964
rect 457588 273924 490104 273952
rect 457588 273912 457594 273924
rect 490098 273912 490104 273924
rect 490156 273912 490162 273964
rect 497918 273912 497924 273964
rect 497976 273952 497982 273964
rect 549438 273952 549444 273964
rect 497976 273924 549444 273952
rect 497976 273912 497982 273924
rect 549438 273912 549444 273924
rect 549496 273912 549502 273964
rect 452286 273232 452292 273284
rect 452344 273272 452350 273284
rect 459554 273272 459560 273284
rect 452344 273244 459560 273272
rect 452344 273232 452350 273244
rect 459554 273232 459560 273244
rect 459612 273232 459618 273284
rect 499390 272552 499396 272604
rect 499448 272592 499454 272604
rect 549622 272592 549628 272604
rect 499448 272564 549628 272592
rect 499448 272552 499454 272564
rect 549622 272552 549628 272564
rect 549680 272552 549686 272604
rect 420178 272484 420184 272536
rect 420236 272524 420242 272536
rect 435542 272524 435548 272536
rect 420236 272496 435548 272524
rect 420236 272484 420242 272496
rect 435542 272484 435548 272496
rect 435600 272484 435606 272536
rect 458726 272484 458732 272536
rect 458784 272524 458790 272536
rect 494146 272524 494152 272536
rect 458784 272496 494152 272524
rect 458784 272484 458790 272496
rect 494146 272484 494152 272496
rect 494204 272484 494210 272536
rect 498010 272484 498016 272536
rect 498068 272524 498074 272536
rect 552382 272524 552388 272536
rect 498068 272496 552388 272524
rect 498068 272484 498074 272496
rect 552382 272484 552388 272496
rect 552440 272484 552446 272536
rect 469858 271912 469864 271924
rect 466472 271884 469864 271912
rect 463326 271804 463332 271856
rect 463384 271844 463390 271856
rect 466472 271844 466500 271884
rect 469858 271872 469864 271884
rect 469916 271872 469922 271924
rect 476758 271912 476764 271924
rect 473740 271884 476764 271912
rect 463384 271816 466500 271844
rect 463384 271804 463390 271816
rect 472710 271804 472716 271856
rect 472768 271844 472774 271856
rect 473740 271844 473768 271884
rect 476758 271872 476764 271884
rect 476816 271872 476822 271924
rect 472768 271816 473768 271844
rect 472768 271804 472774 271816
rect 449250 271396 449256 271448
rect 449308 271436 449314 271448
rect 452562 271436 452568 271448
rect 449308 271408 452568 271436
rect 449308 271396 449314 271408
rect 452562 271396 452568 271408
rect 452620 271396 452626 271448
rect 433978 271260 433984 271312
rect 434036 271300 434042 271312
rect 436922 271300 436928 271312
rect 434036 271272 436928 271300
rect 434036 271260 434042 271272
rect 436922 271260 436928 271272
rect 436980 271260 436986 271312
rect 502150 271260 502156 271312
rect 502208 271300 502214 271312
rect 549806 271300 549812 271312
rect 502208 271272 549812 271300
rect 502208 271260 502214 271272
rect 549806 271260 549812 271272
rect 549864 271260 549870 271312
rect 453022 271192 453028 271244
rect 453080 271232 453086 271244
rect 458174 271232 458180 271244
rect 453080 271204 458180 271232
rect 453080 271192 453086 271204
rect 458174 271192 458180 271204
rect 458232 271192 458238 271244
rect 459370 271192 459376 271244
rect 459428 271232 459434 271244
rect 492766 271232 492772 271244
rect 459428 271204 492772 271232
rect 459428 271192 459434 271204
rect 492766 271192 492772 271204
rect 492824 271192 492830 271244
rect 497734 271192 497740 271244
rect 497792 271232 497798 271244
rect 552198 271232 552204 271244
rect 497792 271204 552204 271232
rect 497792 271192 497798 271204
rect 552198 271192 552204 271204
rect 552256 271192 552262 271244
rect 458634 271124 458640 271176
rect 458692 271164 458698 271176
rect 494054 271164 494060 271176
rect 458692 271136 494060 271164
rect 458692 271124 458698 271136
rect 494054 271124 494060 271136
rect 494112 271124 494118 271176
rect 496722 271124 496728 271176
rect 496780 271164 496786 271176
rect 552014 271164 552020 271176
rect 496780 271136 552020 271164
rect 496780 271124 496786 271136
rect 552014 271124 552020 271136
rect 552072 271124 552078 271176
rect 443914 271056 443920 271108
rect 443972 271096 443978 271108
rect 446490 271096 446496 271108
rect 443972 271068 446496 271096
rect 443972 271056 443978 271068
rect 446490 271056 446496 271068
rect 446548 271056 446554 271108
rect 382274 270444 382280 270496
rect 382332 270484 382338 270496
rect 436830 270484 436836 270496
rect 382332 270456 436836 270484
rect 382332 270444 382338 270456
rect 436830 270444 436836 270456
rect 436888 270444 436894 270496
rect 397178 270104 397184 270156
rect 397236 270144 397242 270156
rect 400214 270144 400220 270156
rect 397236 270116 400220 270144
rect 397236 270104 397242 270116
rect 400214 270104 400220 270116
rect 400272 270104 400278 270156
rect 473262 270036 473268 270088
rect 473320 270076 473326 270088
rect 482462 270076 482468 270088
rect 473320 270048 482468 270076
rect 473320 270036 473326 270048
rect 482462 270036 482468 270048
rect 482520 270036 482526 270088
rect 460750 269968 460756 270020
rect 460808 270008 460814 270020
rect 491570 270008 491576 270020
rect 460808 269980 491576 270008
rect 460808 269968 460814 269980
rect 491570 269968 491576 269980
rect 491628 269968 491634 270020
rect 502242 269968 502248 270020
rect 502300 270008 502306 270020
rect 549714 270008 549720 270020
rect 502300 269980 549720 270008
rect 502300 269968 502306 269980
rect 549714 269968 549720 269980
rect 549772 269968 549778 270020
rect 460106 269900 460112 269952
rect 460164 269940 460170 269952
rect 491478 269940 491484 269952
rect 460164 269912 491484 269940
rect 460164 269900 460170 269912
rect 491478 269900 491484 269912
rect 491536 269900 491542 269952
rect 505002 269900 505008 269952
rect 505060 269940 505066 269952
rect 554774 269940 554780 269952
rect 505060 269912 554780 269940
rect 505060 269900 505066 269912
rect 554774 269900 554780 269912
rect 554832 269900 554838 269952
rect 459462 269832 459468 269884
rect 459520 269872 459526 269884
rect 493042 269872 493048 269884
rect 459520 269844 493048 269872
rect 459520 269832 459526 269844
rect 493042 269832 493048 269844
rect 493100 269832 493106 269884
rect 500770 269832 500776 269884
rect 500828 269872 500834 269884
rect 551370 269872 551376 269884
rect 500828 269844 551376 269872
rect 500828 269832 500834 269844
rect 551370 269832 551376 269844
rect 551428 269832 551434 269884
rect 452194 269764 452200 269816
rect 452252 269804 452258 269816
rect 463326 269804 463332 269816
rect 452252 269776 463332 269804
rect 452252 269764 452258 269776
rect 463326 269764 463332 269776
rect 463384 269764 463390 269816
rect 468938 269764 468944 269816
rect 468996 269804 469002 269816
rect 580350 269804 580356 269816
rect 468996 269776 580356 269804
rect 468996 269764 469002 269776
rect 580350 269764 580356 269776
rect 580408 269764 580414 269816
rect 451274 268744 451280 268796
rect 451332 268784 451338 268796
rect 453022 268784 453028 268796
rect 451332 268756 453028 268784
rect 451332 268744 451338 268756
rect 453022 268744 453028 268756
rect 453080 268744 453086 268796
rect 456702 268676 456708 268728
rect 456760 268716 456766 268728
rect 472710 268716 472716 268728
rect 456760 268688 472716 268716
rect 456760 268676 456766 268688
rect 472710 268676 472716 268688
rect 472768 268676 472774 268728
rect 449342 268608 449348 268660
rect 449400 268648 449406 268660
rect 465718 268648 465724 268660
rect 449400 268620 465724 268648
rect 449400 268608 449406 268620
rect 465718 268608 465724 268620
rect 465776 268608 465782 268660
rect 443730 268540 443736 268592
rect 443788 268580 443794 268592
rect 473262 268580 473268 268592
rect 443788 268552 473268 268580
rect 443788 268540 443794 268552
rect 473262 268540 473268 268552
rect 473320 268540 473326 268592
rect 457898 268472 457904 268524
rect 457956 268512 457962 268524
rect 487154 268512 487160 268524
rect 457956 268484 487160 268512
rect 457956 268472 457962 268484
rect 487154 268472 487160 268484
rect 487212 268472 487218 268524
rect 503254 268472 503260 268524
rect 503312 268512 503318 268524
rect 552566 268512 552572 268524
rect 503312 268484 552572 268512
rect 503312 268472 503318 268484
rect 552566 268472 552572 268484
rect 552624 268472 552630 268524
rect 459278 268404 459284 268456
rect 459336 268444 459342 268456
rect 491662 268444 491668 268456
rect 459336 268416 491668 268444
rect 459336 268404 459342 268416
rect 491662 268404 491668 268416
rect 491720 268404 491726 268456
rect 500494 268404 500500 268456
rect 500552 268444 500558 268456
rect 551278 268444 551284 268456
rect 500552 268416 551284 268444
rect 500552 268404 500558 268416
rect 551278 268404 551284 268416
rect 551336 268404 551342 268456
rect 440970 268336 440976 268388
rect 441028 268376 441034 268388
rect 445754 268376 445760 268388
rect 441028 268348 445760 268376
rect 441028 268336 441034 268348
rect 445754 268336 445760 268348
rect 445812 268336 445818 268388
rect 459186 268336 459192 268388
rect 459244 268376 459250 268388
rect 491386 268376 491392 268388
rect 459244 268348 491392 268376
rect 459244 268336 459250 268348
rect 491386 268336 491392 268348
rect 491444 268336 491450 268388
rect 499114 268336 499120 268388
rect 499172 268376 499178 268388
rect 551094 268376 551100 268388
rect 499172 268348 551100 268376
rect 499172 268336 499178 268348
rect 551094 268336 551100 268348
rect 551152 268336 551158 268388
rect 3694 266636 3700 266688
rect 3752 266676 3758 266688
rect 5258 266676 5264 266688
rect 3752 266648 5264 266676
rect 3752 266636 3758 266648
rect 5258 266636 5264 266648
rect 5316 266636 5322 266688
rect 413278 266364 413284 266416
rect 413336 266404 413342 266416
rect 420178 266404 420184 266416
rect 413336 266376 420184 266404
rect 413336 266364 413342 266376
rect 420178 266364 420184 266376
rect 420236 266364 420242 266416
rect 427814 266364 427820 266416
rect 427872 266404 427878 266416
rect 431218 266404 431224 266416
rect 427872 266376 431224 266404
rect 427872 266364 427878 266376
rect 431218 266364 431224 266376
rect 431276 266364 431282 266416
rect 453022 266364 453028 266416
rect 453080 266404 453086 266416
rect 456702 266404 456708 266416
rect 453080 266376 456708 266404
rect 453080 266364 453086 266376
rect 456702 266364 456708 266376
rect 456760 266364 456766 266416
rect 453022 264976 453028 264988
rect 451246 264948 453028 264976
rect 448514 264868 448520 264920
rect 448572 264908 448578 264920
rect 451246 264908 451274 264948
rect 453022 264936 453028 264948
rect 453080 264936 453086 264988
rect 448572 264880 451274 264908
rect 448572 264868 448578 264880
rect 383378 264188 383384 264240
rect 383436 264228 383442 264240
rect 443822 264228 443828 264240
rect 383436 264200 443828 264228
rect 383436 264188 383442 264200
rect 443822 264188 443828 264200
rect 443880 264188 443886 264240
rect 449710 263508 449716 263560
rect 449768 263548 449774 263560
rect 456794 263548 456800 263560
rect 449768 263520 456800 263548
rect 449768 263508 449774 263520
rect 456794 263508 456800 263520
rect 456852 263508 456858 263560
rect 447778 263440 447784 263492
rect 447836 263480 447842 263492
rect 451274 263480 451280 263492
rect 447836 263452 451280 263480
rect 447836 263440 447842 263452
rect 451274 263440 451280 263452
rect 451332 263440 451338 263492
rect 438118 262692 438124 262744
rect 438176 262732 438182 262744
rect 443914 262732 443920 262744
rect 438176 262704 443920 262732
rect 438176 262692 438182 262704
rect 443914 262692 443920 262704
rect 443972 262692 443978 262744
rect 445754 260380 445760 260432
rect 445812 260420 445818 260432
rect 448422 260420 448428 260432
rect 445812 260392 448428 260420
rect 445812 260380 445818 260392
rect 448422 260380 448428 260392
rect 448480 260380 448486 260432
rect 382274 259360 382280 259412
rect 382332 259400 382338 259412
rect 435358 259400 435364 259412
rect 382332 259372 435364 259400
rect 382332 259360 382338 259372
rect 435358 259360 435364 259372
rect 435416 259360 435422 259412
rect 425698 258952 425704 259004
rect 425756 258992 425762 259004
rect 427814 258992 427820 259004
rect 425756 258964 427820 258992
rect 425756 258952 425762 258964
rect 427814 258952 427820 258964
rect 427872 258952 427878 259004
rect 429562 258340 429568 258392
rect 429620 258380 429626 258392
rect 433978 258380 433984 258392
rect 429620 258352 433984 258380
rect 429620 258340 429626 258352
rect 433978 258340 433984 258352
rect 434036 258340 434042 258392
rect 449158 258068 449164 258120
rect 449216 258108 449222 258120
rect 452286 258108 452292 258120
rect 449216 258080 452292 258108
rect 449216 258068 449222 258080
rect 452286 258068 452292 258080
rect 452344 258068 452350 258120
rect 424134 257320 424140 257372
rect 424192 257360 424198 257372
rect 432690 257360 432696 257372
rect 424192 257332 432696 257360
rect 424192 257320 424198 257332
rect 432690 257320 432696 257332
rect 432748 257320 432754 257372
rect 437474 257320 437480 257372
rect 437532 257360 437538 257372
rect 449342 257360 449348 257372
rect 437532 257332 449348 257360
rect 437532 257320 437538 257332
rect 449342 257320 449348 257332
rect 449400 257320 449406 257372
rect 424318 255280 424324 255332
rect 424376 255320 424382 255332
rect 429562 255320 429568 255332
rect 424376 255292 429568 255320
rect 424376 255280 424382 255292
rect 429562 255280 429568 255292
rect 429620 255280 429626 255332
rect 449250 255320 449256 255332
rect 447152 255292 449256 255320
rect 446122 255212 446128 255264
rect 446180 255252 446186 255264
rect 447152 255252 447180 255292
rect 449250 255280 449256 255292
rect 449308 255280 449314 255332
rect 446180 255224 447180 255252
rect 446180 255212 446186 255224
rect 409138 254532 409144 254584
rect 409196 254572 409202 254584
rect 424134 254572 424140 254584
rect 409196 254544 424140 254572
rect 409196 254532 409202 254544
rect 424134 254532 424140 254544
rect 424192 254532 424198 254584
rect 441062 254532 441068 254584
rect 441120 254572 441126 254584
rect 445662 254572 445668 254584
rect 441120 254544 445668 254572
rect 441120 254532 441126 254544
rect 445662 254532 445668 254544
rect 445720 254532 445726 254584
rect 3510 253920 3516 253972
rect 3568 253960 3574 253972
rect 5166 253960 5172 253972
rect 3568 253932 5172 253960
rect 3568 253920 3574 253932
rect 5166 253920 5172 253932
rect 5224 253920 5230 253972
rect 394418 253920 394424 253972
rect 394476 253960 394482 253972
rect 397178 253960 397184 253972
rect 394476 253932 397184 253960
rect 394476 253920 394482 253932
rect 397178 253920 397184 253932
rect 397236 253920 397242 253972
rect 435358 252900 435364 252952
rect 435416 252940 435422 252952
rect 437474 252940 437480 252952
rect 435416 252912 437480 252940
rect 435416 252900 435422 252912
rect 437474 252900 437480 252912
rect 437532 252900 437538 252952
rect 426342 251812 426348 251864
rect 426400 251852 426406 251864
rect 438118 251852 438124 251864
rect 426400 251824 438124 251852
rect 426400 251812 426406 251824
rect 438118 251812 438124 251824
rect 438176 251812 438182 251864
rect 418798 250452 418804 250504
rect 418856 250492 418862 250504
rect 425698 250492 425704 250504
rect 418856 250464 425704 250492
rect 418856 250452 418862 250464
rect 425698 250452 425704 250464
rect 425756 250452 425762 250504
rect 443822 250384 443828 250436
rect 443880 250424 443886 250436
rect 446122 250424 446128 250436
rect 443880 250396 446128 250424
rect 443880 250384 443886 250396
rect 446122 250384 446128 250396
rect 446180 250384 446186 250436
rect 382274 249704 382280 249756
rect 382332 249744 382338 249756
rect 432598 249744 432604 249756
rect 382332 249716 432604 249744
rect 382332 249704 382338 249716
rect 432598 249704 432604 249716
rect 432656 249704 432662 249756
rect 411254 249024 411260 249076
rect 411312 249064 411318 249076
rect 426342 249064 426348 249076
rect 411312 249036 426348 249064
rect 411312 249024 411318 249036
rect 426342 249024 426348 249036
rect 426400 249024 426406 249076
rect 447870 249024 447876 249076
rect 447928 249064 447934 249076
rect 457990 249064 457996 249076
rect 447928 249036 457996 249064
rect 447928 249024 447934 249036
rect 457990 249024 457996 249036
rect 458048 249024 458054 249076
rect 436002 248480 436008 248532
rect 436060 248520 436066 248532
rect 439682 248520 439688 248532
rect 436060 248492 439688 248520
rect 436060 248480 436066 248492
rect 439682 248480 439688 248492
rect 439740 248480 439746 248532
rect 422938 246304 422944 246356
rect 422996 246344 423002 246356
rect 435358 246344 435364 246356
rect 422996 246316 435364 246344
rect 422996 246304 423002 246316
rect 435358 246304 435364 246316
rect 435416 246304 435422 246356
rect 3970 245964 3976 246016
rect 4028 246004 4034 246016
rect 5074 246004 5080 246016
rect 4028 245976 5080 246004
rect 4028 245964 4034 245976
rect 5074 245964 5080 245976
rect 5132 245964 5138 246016
rect 405274 245624 405280 245676
rect 405332 245664 405338 245676
rect 411254 245664 411260 245676
rect 405332 245636 411260 245664
rect 405332 245624 405338 245636
rect 411254 245624 411260 245636
rect 411312 245624 411318 245676
rect 446490 245624 446496 245676
rect 446548 245664 446554 245676
rect 447778 245664 447784 245676
rect 446548 245636 447784 245664
rect 446548 245624 446554 245636
rect 447778 245624 447784 245636
rect 447836 245624 447842 245676
rect 537478 245556 537484 245608
rect 537536 245596 537542 245608
rect 580166 245596 580172 245608
rect 537536 245568 580172 245596
rect 537536 245556 537542 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 390370 245148 390376 245200
rect 390428 245188 390434 245200
rect 394418 245188 394424 245200
rect 390428 245160 394424 245188
rect 390428 245148 390434 245160
rect 394418 245148 394424 245160
rect 394476 245148 394482 245200
rect 429838 244876 429844 244928
rect 429896 244916 429902 244928
rect 436002 244916 436008 244928
rect 429896 244888 436008 244916
rect 429896 244876 429902 244888
rect 436002 244876 436008 244888
rect 436060 244876 436066 244928
rect 424318 244304 424324 244316
rect 422266 244276 424324 244304
rect 420914 244196 420920 244248
rect 420972 244236 420978 244248
rect 422266 244236 422294 244276
rect 424318 244264 424324 244276
rect 424376 244264 424382 244316
rect 420972 244208 422294 244236
rect 420972 244196 420978 244208
rect 445018 243176 445024 243228
rect 445076 243216 445082 243228
rect 446490 243216 446496 243228
rect 445076 243188 446496 243216
rect 445076 243176 445082 243188
rect 446490 243176 446496 243188
rect 446548 243176 446554 243228
rect 442994 240864 443000 240916
rect 443052 240904 443058 240916
rect 449158 240904 449164 240916
rect 443052 240876 449164 240904
rect 443052 240864 443058 240876
rect 449158 240864 449164 240876
rect 449216 240864 449222 240916
rect 419534 239844 419540 239896
rect 419592 239884 419598 239896
rect 420914 239884 420920 239896
rect 419592 239856 420920 239884
rect 419592 239844 419598 239856
rect 420914 239844 420920 239856
rect 420972 239844 420978 239896
rect 395890 239368 395896 239420
rect 395948 239408 395954 239420
rect 413278 239408 413284 239420
rect 395948 239380 413284 239408
rect 395948 239368 395954 239380
rect 413278 239368 413284 239380
rect 413336 239368 413342 239420
rect 382274 238688 382280 238740
rect 382332 238728 382338 238740
rect 440878 238728 440884 238740
rect 382332 238700 440884 238728
rect 382332 238688 382338 238700
rect 440878 238688 440884 238700
rect 440936 238688 440942 238740
rect 417418 237396 417424 237448
rect 417476 237436 417482 237448
rect 419534 237436 419540 237448
rect 417476 237408 419540 237436
rect 417476 237396 417482 237408
rect 419534 237396 419540 237408
rect 419592 237396 419598 237448
rect 420178 235628 420184 235680
rect 420236 235668 420242 235680
rect 422938 235668 422944 235680
rect 420236 235640 422944 235668
rect 420236 235628 420242 235640
rect 422938 235628 422944 235640
rect 422996 235628 423002 235680
rect 434898 235424 434904 235476
rect 434956 235464 434962 235476
rect 442994 235464 443000 235476
rect 434956 235436 443000 235464
rect 434956 235424 434962 235436
rect 442994 235424 443000 235436
rect 443052 235424 443058 235476
rect 383286 235220 383292 235272
rect 383344 235260 383350 235272
rect 390370 235260 390376 235272
rect 383344 235232 390376 235260
rect 383344 235220 383350 235232
rect 390370 235220 390376 235232
rect 390428 235220 390434 235272
rect 453298 234948 453304 235000
rect 453356 234988 453362 235000
rect 457162 234988 457168 235000
rect 453356 234960 457168 234988
rect 453356 234948 453362 234960
rect 457162 234948 457168 234960
rect 457220 234948 457226 235000
rect 450078 234608 450084 234660
rect 450136 234648 450142 234660
rect 452194 234648 452200 234660
rect 450136 234620 452200 234648
rect 450136 234608 450142 234620
rect 452194 234608 452200 234620
rect 452252 234608 452258 234660
rect 416038 233860 416044 233912
rect 416096 233900 416102 233912
rect 418798 233900 418804 233912
rect 416096 233872 418804 233900
rect 416096 233860 416102 233872
rect 418798 233860 418804 233872
rect 418856 233860 418862 233912
rect 540238 233180 540244 233232
rect 540296 233220 540302 233232
rect 580166 233220 580172 233232
rect 540296 233192 580172 233220
rect 540296 233180 540302 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 449158 232704 449164 232756
rect 449216 232744 449222 232756
rect 452102 232744 452108 232756
rect 449216 232716 452108 232744
rect 449216 232704 449222 232716
rect 452102 232704 452108 232716
rect 452160 232704 452166 232756
rect 427078 232500 427084 232552
rect 427136 232540 427142 232552
rect 434898 232540 434904 232552
rect 427136 232512 434904 232540
rect 427136 232500 427142 232512
rect 434898 232500 434904 232512
rect 434956 232500 434962 232552
rect 447778 231820 447784 231872
rect 447836 231860 447842 231872
rect 450078 231860 450084 231872
rect 447836 231832 450084 231860
rect 447836 231820 447842 231832
rect 450078 231820 450084 231832
rect 450136 231820 450142 231872
rect 443822 230500 443828 230512
rect 438872 230472 443828 230500
rect 435450 230392 435456 230444
rect 435508 230432 435514 230444
rect 438872 230432 438900 230472
rect 443822 230460 443828 230472
rect 443880 230460 443886 230512
rect 435508 230404 438900 230432
rect 435508 230392 435514 230404
rect 422938 229984 422944 230036
rect 422996 230024 423002 230036
rect 429838 230024 429844 230036
rect 422996 229996 429844 230024
rect 422996 229984 423002 229996
rect 429838 229984 429844 229996
rect 429896 229984 429902 230036
rect 397178 229100 397184 229152
rect 397236 229140 397242 229152
rect 405274 229140 405280 229152
rect 397236 229112 405280 229140
rect 397236 229100 397242 229112
rect 405274 229100 405280 229112
rect 405332 229100 405338 229152
rect 387610 227740 387616 227792
rect 387668 227780 387674 227792
rect 395890 227780 395896 227792
rect 387668 227752 395896 227780
rect 387668 227740 387674 227752
rect 395890 227740 395896 227752
rect 395948 227740 395954 227792
rect 382274 227672 382280 227724
rect 382332 227712 382338 227724
rect 436738 227712 436744 227724
rect 382332 227684 436744 227712
rect 382332 227672 382338 227684
rect 436738 227672 436744 227684
rect 436796 227672 436802 227724
rect 411254 226992 411260 227044
rect 411312 227032 411318 227044
rect 416038 227032 416044 227044
rect 411312 227004 416044 227032
rect 411312 226992 411318 227004
rect 416038 226992 416044 227004
rect 416096 226992 416102 227044
rect 421558 224204 421564 224256
rect 421616 224244 421622 224256
rect 427078 224244 427084 224256
rect 421616 224216 427084 224244
rect 421616 224204 421622 224216
rect 427078 224204 427084 224216
rect 427136 224204 427142 224256
rect 438118 224204 438124 224256
rect 438176 224244 438182 224256
rect 441062 224244 441068 224256
rect 438176 224216 441068 224244
rect 438176 224204 438182 224216
rect 441062 224204 441068 224216
rect 441120 224204 441126 224256
rect 416774 223728 416780 223780
rect 416832 223768 416838 223780
rect 420178 223768 420184 223780
rect 416832 223740 420184 223768
rect 416832 223728 416838 223740
rect 420178 223728 420184 223740
rect 420236 223728 420242 223780
rect 444190 223252 444196 223304
rect 444248 223292 444254 223304
rect 449158 223292 449164 223304
rect 444248 223264 449164 223292
rect 444248 223252 444254 223264
rect 449158 223252 449164 223264
rect 449216 223252 449222 223304
rect 452010 222096 452016 222148
rect 452068 222136 452074 222148
rect 457346 222136 457352 222148
rect 452068 222108 457352 222136
rect 452068 222096 452074 222108
rect 457346 222096 457352 222108
rect 457404 222096 457410 222148
rect 433978 220736 433984 220788
rect 434036 220776 434042 220788
rect 435450 220776 435456 220788
rect 434036 220748 435456 220776
rect 434036 220736 434042 220748
rect 435450 220736 435456 220748
rect 435508 220736 435514 220788
rect 408770 220328 408776 220380
rect 408828 220368 408834 220380
rect 411254 220368 411260 220380
rect 408828 220340 411260 220368
rect 408828 220328 408834 220340
rect 411254 220328 411260 220340
rect 411312 220328 411318 220380
rect 411254 220056 411260 220108
rect 411312 220096 411318 220108
rect 416774 220096 416780 220108
rect 411312 220068 416780 220096
rect 411312 220056 411318 220068
rect 416774 220056 416780 220068
rect 416832 220056 416838 220108
rect 435358 219444 435364 219496
rect 435416 219484 435422 219496
rect 444190 219484 444196 219496
rect 435416 219456 444196 219484
rect 435416 219444 435422 219456
rect 444190 219444 444196 219456
rect 444248 219444 444254 219496
rect 442718 218084 442724 218136
rect 442776 218124 442782 218136
rect 445018 218124 445024 218136
rect 442776 218096 445024 218124
rect 442776 218084 442782 218096
rect 445018 218084 445024 218096
rect 445076 218084 445082 218136
rect 417510 216928 417516 216980
rect 417568 216968 417574 216980
rect 422938 216968 422944 216980
rect 417568 216940 422944 216968
rect 417568 216928 417574 216940
rect 422938 216928 422944 216940
rect 422996 216928 423002 216980
rect 440878 216656 440884 216708
rect 440936 216696 440942 216708
rect 442718 216696 442724 216708
rect 440936 216668 442724 216696
rect 440936 216656 440942 216668
rect 442718 216656 442724 216668
rect 442776 216656 442782 216708
rect 3418 215500 3424 215552
rect 3476 215540 3482 215552
rect 5350 215540 5356 215552
rect 3476 215512 5356 215540
rect 3476 215500 3482 215512
rect 5350 215500 5356 215512
rect 5408 215500 5414 215552
rect 406930 215296 406936 215348
rect 406988 215336 406994 215348
rect 411254 215336 411260 215348
rect 406988 215308 411260 215336
rect 406988 215296 406994 215308
rect 411254 215296 411260 215308
rect 411312 215296 411318 215348
rect 413278 215296 413284 215348
rect 413336 215336 413342 215348
rect 417418 215336 417424 215348
rect 413336 215308 417424 215336
rect 413336 215296 413342 215308
rect 417418 215296 417424 215308
rect 417476 215296 417482 215348
rect 384666 214548 384672 214600
rect 384724 214588 384730 214600
rect 397178 214588 397184 214600
rect 384724 214560 397184 214588
rect 384724 214548 384730 214560
rect 397178 214548 397184 214560
rect 397236 214548 397242 214600
rect 399938 213188 399944 213240
rect 399996 213228 400002 213240
rect 408770 213228 408776 213240
rect 399996 213200 408776 213228
rect 399996 213188 400002 213200
rect 408770 213188 408776 213200
rect 408828 213188 408834 213240
rect 3878 212440 3884 212492
rect 3936 212480 3942 212492
rect 4982 212480 4988 212492
rect 3936 212452 4988 212480
rect 3936 212440 3942 212452
rect 4982 212440 4988 212452
rect 5040 212440 5046 212492
rect 402974 212440 402980 212492
rect 403032 212480 403038 212492
rect 406930 212480 406936 212492
rect 403032 212452 406936 212480
rect 403032 212440 403038 212452
rect 406930 212440 406936 212452
rect 406988 212440 406994 212492
rect 436738 212440 436744 212492
rect 436796 212480 436802 212492
rect 438118 212480 438124 212492
rect 436796 212452 438124 212480
rect 436796 212440 436802 212452
rect 438118 212440 438124 212452
rect 438176 212440 438182 212492
rect 425698 211760 425704 211812
rect 425756 211800 425762 211812
rect 440970 211800 440976 211812
rect 425756 211772 440976 211800
rect 425756 211760 425762 211772
rect 440970 211760 440976 211772
rect 441028 211760 441034 211812
rect 443822 211284 443828 211336
rect 443880 211324 443886 211336
rect 447778 211324 447784 211336
rect 443880 211296 447784 211324
rect 443880 211284 443886 211296
rect 447778 211284 447784 211296
rect 447836 211284 447842 211336
rect 383378 207612 383384 207664
rect 383436 207652 383442 207664
rect 399938 207652 399944 207664
rect 383436 207624 399944 207652
rect 383436 207612 383442 207624
rect 399938 207612 399944 207624
rect 399996 207612 400002 207664
rect 451918 207204 451924 207256
rect 451976 207244 451982 207256
rect 456794 207244 456800 207256
rect 451976 207216 456800 207244
rect 451976 207204 451982 207216
rect 456794 207204 456800 207216
rect 456852 207204 456858 207256
rect 382274 206932 382280 206984
rect 382332 206972 382338 206984
rect 439498 206972 439504 206984
rect 382332 206944 439504 206972
rect 382332 206932 382338 206944
rect 439498 206932 439504 206944
rect 439556 206932 439562 206984
rect 533338 206932 533344 206984
rect 533396 206972 533402 206984
rect 579798 206972 579804 206984
rect 533396 206944 579804 206972
rect 533396 206932 533402 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 393130 206320 393136 206372
rect 393188 206360 393194 206372
rect 402974 206360 402980 206372
rect 393188 206332 402980 206360
rect 393188 206320 393194 206332
rect 402974 206320 402980 206332
rect 403032 206320 403038 206372
rect 395890 206252 395896 206304
rect 395948 206292 395954 206304
rect 409138 206292 409144 206304
rect 395948 206264 409144 206292
rect 395948 206252 395954 206264
rect 409138 206252 409144 206264
rect 409196 206252 409202 206304
rect 411898 205572 411904 205624
rect 411956 205612 411962 205624
rect 413278 205612 413284 205624
rect 411956 205584 413284 205612
rect 411956 205572 411962 205584
rect 413278 205572 413284 205584
rect 413336 205572 413342 205624
rect 432322 202784 432328 202836
rect 432380 202824 432386 202836
rect 435358 202824 435364 202836
rect 432380 202796 435364 202824
rect 432380 202784 432386 202796
rect 435358 202784 435364 202796
rect 435416 202784 435422 202836
rect 422938 201424 422944 201476
rect 422996 201464 423002 201476
rect 425698 201464 425704 201476
rect 422996 201436 425704 201464
rect 422996 201424 423002 201436
rect 425698 201424 425704 201436
rect 425756 201424 425762 201476
rect 438854 201424 438860 201476
rect 438912 201464 438918 201476
rect 440878 201464 440884 201476
rect 438912 201436 440884 201464
rect 438912 201424 438918 201436
rect 440878 201424 440884 201436
rect 440936 201424 440942 201476
rect 408494 199452 408500 199504
rect 408552 199492 408558 199504
rect 421558 199492 421564 199504
rect 408552 199464 421564 199492
rect 408552 199452 408558 199464
rect 421558 199452 421564 199464
rect 421616 199452 421622 199504
rect 384758 199384 384764 199436
rect 384816 199424 384822 199436
rect 395890 199424 395896 199436
rect 384816 199396 395896 199424
rect 384816 199384 384822 199396
rect 395890 199384 395896 199396
rect 395948 199384 395954 199436
rect 402422 199384 402428 199436
rect 402480 199424 402486 199436
rect 417510 199424 417516 199436
rect 402480 199396 417516 199424
rect 402480 199384 402486 199396
rect 417510 199384 417516 199396
rect 417568 199384 417574 199436
rect 432966 198704 432972 198756
rect 433024 198744 433030 198756
rect 433978 198744 433984 198756
rect 433024 198716 433984 198744
rect 433024 198704 433030 198716
rect 433978 198704 433984 198716
rect 434036 198704 434042 198756
rect 433978 197344 433984 197396
rect 434036 197384 434042 197396
rect 436738 197384 436744 197396
rect 434036 197356 436744 197384
rect 434036 197344 434042 197356
rect 436738 197344 436744 197356
rect 436796 197344 436802 197396
rect 429930 196936 429936 196988
rect 429988 196976 429994 196988
rect 432966 196976 432972 196988
rect 429988 196948 432972 196976
rect 429988 196936 429994 196948
rect 432966 196936 432972 196948
rect 433024 196936 433030 196988
rect 400766 196596 400772 196648
rect 400824 196636 400830 196648
rect 408494 196636 408500 196648
rect 400824 196608 408500 196636
rect 400824 196596 400830 196608
rect 408494 196596 408500 196608
rect 408552 196596 408558 196648
rect 436738 195984 436744 196036
rect 436796 196024 436802 196036
rect 438854 196024 438860 196036
rect 436796 195996 438860 196024
rect 436796 195984 436802 195996
rect 438854 195984 438860 195996
rect 438912 195984 438918 196036
rect 382274 195916 382280 195968
rect 382332 195956 382338 195968
rect 443638 195956 443644 195968
rect 382332 195928 443644 195956
rect 382332 195916 382338 195928
rect 443638 195916 443644 195928
rect 443696 195916 443702 195968
rect 429838 193944 429844 193996
rect 429896 193984 429902 193996
rect 432322 193984 432328 193996
rect 429896 193956 432328 193984
rect 429896 193944 429902 193956
rect 432322 193944 432328 193956
rect 432380 193944 432386 193996
rect 410610 193740 410616 193792
rect 410668 193780 410674 193792
rect 411898 193780 411904 193792
rect 410668 193752 411904 193780
rect 410668 193740 410674 193752
rect 411898 193740 411904 193752
rect 411956 193740 411962 193792
rect 538858 193128 538864 193180
rect 538916 193168 538922 193180
rect 580166 193168 580172 193180
rect 538916 193140 580172 193168
rect 538916 193128 538922 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 398466 192856 398472 192908
rect 398524 192896 398530 192908
rect 400766 192896 400772 192908
rect 398524 192868 400772 192896
rect 398524 192856 398530 192868
rect 400766 192856 400772 192868
rect 400824 192856 400830 192908
rect 440234 189048 440240 189100
rect 440292 189088 440298 189100
rect 443822 189088 443828 189100
rect 440292 189060 443828 189088
rect 440292 189048 440298 189060
rect 443822 189048 443828 189060
rect 443880 189048 443886 189100
rect 4890 188028 4896 188080
rect 4948 188068 4954 188080
rect 6178 188068 6184 188080
rect 4948 188040 6184 188068
rect 4948 188028 4954 188040
rect 6178 188028 6184 188040
rect 6236 188028 6242 188080
rect 3602 187688 3608 187740
rect 3660 187728 3666 187740
rect 4798 187728 4804 187740
rect 3660 187700 4804 187728
rect 3660 187688 3666 187700
rect 4798 187688 4804 187700
rect 4856 187688 4862 187740
rect 407114 187688 407120 187740
rect 407172 187728 407178 187740
rect 410610 187728 410616 187740
rect 407172 187700 410616 187728
rect 407172 187688 407178 187700
rect 410610 187688 410616 187700
rect 410668 187688 410674 187740
rect 416038 187076 416044 187128
rect 416096 187116 416102 187128
rect 422938 187116 422944 187128
rect 416096 187088 422944 187116
rect 416096 187076 416102 187088
rect 422938 187076 422944 187088
rect 422996 187076 423002 187128
rect 439498 186532 439504 186584
rect 439556 186572 439562 186584
rect 443730 186572 443736 186584
rect 439556 186544 443736 186572
rect 439556 186532 439562 186544
rect 443730 186532 443736 186544
rect 443788 186532 443794 186584
rect 390370 186328 390376 186380
rect 390428 186368 390434 186380
rect 393130 186368 393136 186380
rect 390428 186340 393136 186368
rect 390428 186328 390434 186340
rect 393130 186328 393136 186340
rect 393188 186328 393194 186380
rect 382274 186260 382280 186312
rect 382332 186300 382338 186312
rect 447134 186300 447140 186312
rect 382332 186272 447140 186300
rect 382332 186260 382338 186272
rect 447134 186260 447140 186272
rect 447192 186260 447198 186312
rect 382090 186192 382096 186244
rect 382148 186232 382154 186244
rect 384758 186232 384764 186244
rect 382148 186204 384764 186232
rect 382148 186192 382154 186204
rect 384758 186192 384764 186204
rect 384816 186192 384822 186244
rect 447134 185580 447140 185632
rect 447192 185620 447198 185632
rect 448146 185620 448152 185632
rect 447192 185592 448152 185620
rect 447192 185580 447198 185592
rect 448146 185580 448152 185592
rect 448204 185620 448210 185632
rect 536834 185620 536840 185632
rect 448204 185592 536840 185620
rect 448204 185580 448210 185592
rect 536834 185580 536840 185592
rect 536892 185580 536898 185632
rect 428458 185444 428464 185496
rect 428516 185484 428522 185496
rect 429930 185484 429936 185496
rect 428516 185456 429936 185484
rect 428516 185444 428522 185456
rect 429930 185444 429936 185456
rect 429988 185444 429994 185496
rect 405550 183880 405556 183932
rect 405608 183920 405614 183932
rect 407114 183920 407120 183932
rect 405608 183892 407120 183920
rect 405608 183880 405614 183892
rect 407114 183880 407120 183892
rect 407172 183880 407178 183932
rect 432782 183540 432788 183592
rect 432840 183580 432846 183592
rect 433978 183580 433984 183592
rect 432840 183552 433984 183580
rect 432840 183540 432846 183552
rect 433978 183540 433984 183552
rect 434036 183540 434042 183592
rect 438854 183064 438860 183116
rect 438912 183104 438918 183116
rect 440234 183104 440240 183116
rect 438912 183076 440240 183104
rect 438912 183064 438918 183076
rect 440234 183064 440240 183076
rect 440292 183064 440298 183116
rect 397270 182384 397276 182436
rect 397328 182424 397334 182436
rect 402422 182424 402428 182436
rect 397328 182396 402428 182424
rect 397328 182384 397334 182396
rect 402422 182384 402428 182396
rect 402480 182384 402486 182436
rect 405550 182220 405556 182232
rect 402946 182192 405556 182220
rect 397362 182112 397368 182164
rect 397420 182152 397426 182164
rect 402946 182152 402974 182192
rect 405550 182180 405556 182192
rect 405608 182180 405614 182232
rect 431218 182180 431224 182232
rect 431276 182220 431282 182232
rect 432782 182220 432788 182232
rect 431276 182192 432788 182220
rect 431276 182180 431282 182192
rect 432782 182180 432788 182192
rect 432840 182180 432846 182232
rect 397420 182124 402974 182152
rect 397420 182112 397426 182124
rect 435358 182112 435364 182164
rect 435416 182152 435422 182164
rect 436738 182152 436744 182164
rect 435416 182124 436744 182152
rect 435416 182112 435422 182124
rect 436738 182112 436744 182124
rect 436796 182112 436802 182164
rect 436094 179392 436100 179444
rect 436152 179432 436158 179444
rect 438854 179432 438860 179444
rect 436152 179404 438860 179432
rect 436152 179392 436158 179404
rect 438854 179392 438860 179404
rect 438912 179392 438918 179444
rect 543090 179324 543096 179376
rect 543148 179364 543154 179376
rect 580166 179364 580172 179376
rect 543148 179336 580172 179364
rect 543148 179324 543154 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 401410 178644 401416 178696
rect 401468 178684 401474 178696
rect 416038 178684 416044 178696
rect 401468 178656 416044 178684
rect 401468 178644 401474 178656
rect 416038 178644 416044 178656
rect 416096 178644 416102 178696
rect 393130 175924 393136 175976
rect 393188 175964 393194 175976
rect 397270 175964 397276 175976
rect 393188 175936 397276 175964
rect 393188 175924 393194 175936
rect 397270 175924 397276 175936
rect 397328 175924 397334 175976
rect 426434 175924 426440 175976
rect 426492 175964 426498 175976
rect 428458 175964 428464 175976
rect 426492 175936 428464 175964
rect 426492 175924 426498 175936
rect 428458 175924 428464 175936
rect 428516 175924 428522 175976
rect 430574 175924 430580 175976
rect 430632 175964 430638 175976
rect 436094 175964 436100 175976
rect 430632 175936 436100 175964
rect 430632 175924 430638 175936
rect 436094 175924 436100 175936
rect 436152 175924 436158 175976
rect 422938 175856 422944 175908
rect 422996 175896 423002 175908
rect 429838 175896 429844 175908
rect 422996 175868 429844 175896
rect 422996 175856 423002 175868
rect 429838 175856 429844 175868
rect 429896 175856 429902 175908
rect 382274 175176 382280 175228
rect 382332 175216 382338 175228
rect 447134 175216 447140 175228
rect 382332 175188 447140 175216
rect 382332 175176 382338 175188
rect 447134 175176 447140 175188
rect 447192 175216 447198 175228
rect 447502 175216 447508 175228
rect 447192 175188 447508 175216
rect 447192 175176 447198 175188
rect 447502 175176 447508 175188
rect 447560 175176 447566 175228
rect 447134 174496 447140 174548
rect 447192 174536 447198 174548
rect 532694 174536 532700 174548
rect 447192 174508 532700 174536
rect 447192 174496 447198 174508
rect 532694 174496 532700 174508
rect 532752 174496 532758 174548
rect 395246 173952 395252 174004
rect 395304 173992 395310 174004
rect 397362 173992 397368 174004
rect 395304 173964 397368 173992
rect 395304 173952 395310 173964
rect 397362 173952 397368 173964
rect 397420 173952 397426 174004
rect 426434 173924 426440 173936
rect 425072 173896 426440 173924
rect 423674 173816 423680 173868
rect 423732 173856 423738 173868
rect 425072 173856 425100 173896
rect 426434 173884 426440 173896
rect 426492 173884 426498 173936
rect 423732 173828 425100 173856
rect 423732 173816 423738 173828
rect 380526 173136 380532 173188
rect 380584 173176 380590 173188
rect 390370 173176 390376 173188
rect 380584 173148 390376 173176
rect 380584 173136 380590 173148
rect 390370 173136 390376 173148
rect 390428 173136 390434 173188
rect 429286 172456 429292 172508
rect 429344 172496 429350 172508
rect 431218 172496 431224 172508
rect 429344 172468 431224 172496
rect 429344 172456 429350 172468
rect 431218 172456 431224 172468
rect 431276 172456 431282 172508
rect 393314 172048 393320 172100
rect 393372 172088 393378 172100
rect 395246 172088 395252 172100
rect 393372 172060 395252 172088
rect 393372 172048 393378 172060
rect 395246 172048 395252 172060
rect 395304 172048 395310 172100
rect 429194 171776 429200 171828
rect 429252 171816 429258 171828
rect 430574 171816 430580 171828
rect 429252 171788 430580 171816
rect 429252 171776 429258 171788
rect 430574 171776 430580 171788
rect 430632 171776 430638 171828
rect 422294 169736 422300 169788
rect 422352 169776 422358 169788
rect 423674 169776 423680 169788
rect 422352 169748 423680 169776
rect 422352 169736 422358 169748
rect 423674 169736 423680 169748
rect 423732 169736 423738 169788
rect 388714 169056 388720 169108
rect 388772 169096 388778 169108
rect 393314 169096 393320 169108
rect 388772 169068 393320 169096
rect 388772 169056 388778 169068
rect 393314 169056 393320 169068
rect 393372 169056 393378 169108
rect 449802 169056 449808 169108
rect 449860 169096 449866 169108
rect 452838 169096 452844 169108
rect 449860 169068 452844 169096
rect 449860 169056 449866 169068
rect 452838 169056 452844 169068
rect 452896 169056 452902 169108
rect 386138 168988 386144 169040
rect 386196 169028 386202 169040
rect 401410 169028 401416 169040
rect 386196 169000 401416 169028
rect 386196 168988 386202 169000
rect 401410 168988 401416 169000
rect 401468 168988 401474 169040
rect 429194 168416 429200 168428
rect 423692 168388 429200 168416
rect 423122 168308 423128 168360
rect 423180 168348 423186 168360
rect 423692 168348 423720 168388
rect 429194 168376 429200 168388
rect 429252 168376 429258 168428
rect 423180 168320 423720 168348
rect 423180 168308 423186 168320
rect 449342 168036 449348 168088
rect 449400 168076 449406 168088
rect 456794 168076 456800 168088
rect 449400 168048 456800 168076
rect 449400 168036 449406 168048
rect 456794 168036 456800 168048
rect 456852 168036 456858 168088
rect 457254 167968 457260 168020
rect 457312 168008 457318 168020
rect 482370 168008 482376 168020
rect 457312 167980 482376 168008
rect 457312 167968 457318 167980
rect 482370 167968 482376 167980
rect 482428 167968 482434 168020
rect 430758 167900 430764 167952
rect 430816 167940 430822 167952
rect 439498 167940 439504 167952
rect 430816 167912 439504 167940
rect 430816 167900 430822 167912
rect 439498 167900 439504 167912
rect 439556 167900 439562 167952
rect 456886 167900 456892 167952
rect 456944 167940 456950 167952
rect 457346 167940 457352 167952
rect 456944 167912 457352 167940
rect 456944 167900 456950 167912
rect 457346 167900 457352 167912
rect 457404 167940 457410 167952
rect 487154 167940 487160 167952
rect 457404 167912 487160 167940
rect 457404 167900 457410 167912
rect 487154 167900 487160 167912
rect 487212 167900 487218 167952
rect 419718 167832 419724 167884
rect 419776 167872 419782 167884
rect 458082 167872 458088 167884
rect 419776 167844 458088 167872
rect 419776 167832 419782 167844
rect 458082 167832 458088 167844
rect 458140 167872 458146 167884
rect 458140 167844 460934 167872
rect 458140 167832 458146 167844
rect 416222 167764 416228 167816
rect 416280 167804 416286 167816
rect 456886 167804 456892 167816
rect 416280 167776 456892 167804
rect 416280 167764 416286 167776
rect 456886 167764 456892 167776
rect 456944 167764 456950 167816
rect 460906 167804 460934 167844
rect 491570 167804 491576 167816
rect 460906 167776 491576 167804
rect 491570 167764 491576 167776
rect 491628 167764 491634 167816
rect 404446 167696 404452 167748
rect 404504 167736 404510 167748
rect 422938 167736 422944 167748
rect 404504 167708 422944 167736
rect 404504 167696 404510 167708
rect 422938 167696 422944 167708
rect 422996 167696 423002 167748
rect 427078 167696 427084 167748
rect 427136 167736 427142 167748
rect 450538 167736 450544 167748
rect 427136 167708 450544 167736
rect 427136 167696 427142 167708
rect 450538 167696 450544 167708
rect 450596 167736 450602 167748
rect 500954 167736 500960 167748
rect 450596 167708 500960 167736
rect 450596 167696 450602 167708
rect 500954 167696 500960 167708
rect 501012 167696 501018 167748
rect 411898 167628 411904 167680
rect 411956 167668 411962 167680
rect 411956 167640 451274 167668
rect 411956 167628 411962 167640
rect 451246 167600 451274 167640
rect 456794 167628 456800 167680
rect 456852 167668 456858 167680
rect 457990 167668 457996 167680
rect 456852 167640 457996 167668
rect 456852 167628 456858 167640
rect 457990 167628 457996 167640
rect 458048 167668 458054 167680
rect 537478 167668 537484 167680
rect 458048 167640 537484 167668
rect 458048 167628 458054 167640
rect 537478 167628 537484 167640
rect 537536 167628 537542 167680
rect 457254 167600 457260 167612
rect 451246 167572 457260 167600
rect 457254 167560 457260 167572
rect 457312 167560 457318 167612
rect 445662 167152 445668 167204
rect 445720 167192 445726 167204
rect 446398 167192 446404 167204
rect 445720 167164 446404 167192
rect 445720 167152 445726 167164
rect 446398 167152 446404 167164
rect 446456 167152 446462 167204
rect 384758 167084 384764 167136
rect 384816 167124 384822 167136
rect 393130 167124 393136 167136
rect 384816 167096 393136 167124
rect 384816 167084 384822 167096
rect 393130 167084 393136 167096
rect 393188 167084 393194 167136
rect 430850 167084 430856 167136
rect 430908 167124 430914 167136
rect 449894 167124 449900 167136
rect 430908 167096 449900 167124
rect 430908 167084 430914 167096
rect 449894 167084 449900 167096
rect 449952 167124 449958 167136
rect 450906 167124 450912 167136
rect 449952 167096 450912 167124
rect 449952 167084 449958 167096
rect 450906 167084 450912 167096
rect 450964 167084 450970 167136
rect 383470 167016 383476 167068
rect 383528 167056 383534 167068
rect 434438 167056 434444 167068
rect 383528 167028 434444 167056
rect 383528 167016 383534 167028
rect 434438 167016 434444 167028
rect 434496 167056 434502 167068
rect 449986 167056 449992 167068
rect 434496 167028 449992 167056
rect 434496 167016 434502 167028
rect 449986 167016 449992 167028
rect 450044 167056 450050 167068
rect 450538 167056 450544 167068
rect 450044 167028 450544 167056
rect 450044 167016 450050 167028
rect 450538 167016 450544 167028
rect 450596 167016 450602 167068
rect 536098 166948 536104 167000
rect 536156 166988 536162 167000
rect 580166 166988 580172 167000
rect 536156 166960 580172 166988
rect 536156 166948 536162 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 450906 166336 450912 166388
rect 450964 166376 450970 166388
rect 504358 166376 504364 166388
rect 450964 166348 504364 166376
rect 450964 166336 450970 166348
rect 504358 166336 504364 166348
rect 504416 166336 504422 166388
rect 450538 166268 450544 166320
rect 450596 166308 450602 166320
rect 508498 166308 508504 166320
rect 450596 166280 508504 166308
rect 450596 166268 450602 166280
rect 508498 166268 508504 166280
rect 508556 166268 508562 166320
rect 408034 165724 408040 165776
rect 408092 165764 408098 165776
rect 416222 165764 416228 165776
rect 408092 165736 416228 165764
rect 408092 165724 408098 165736
rect 416222 165724 416228 165736
rect 416280 165724 416286 165776
rect 391566 165656 391572 165708
rect 391624 165696 391630 165708
rect 411898 165696 411904 165708
rect 391624 165668 411904 165696
rect 391624 165656 391630 165668
rect 411898 165656 411904 165668
rect 411956 165656 411962 165708
rect 438026 165656 438032 165708
rect 438084 165696 438090 165708
rect 438762 165696 438768 165708
rect 438084 165668 438768 165696
rect 438084 165656 438090 165668
rect 438762 165656 438768 165668
rect 438820 165696 438826 165708
rect 514754 165696 514760 165708
rect 438820 165668 514760 165696
rect 438820 165656 438826 165668
rect 514754 165656 514760 165668
rect 514812 165656 514818 165708
rect 406654 165588 406660 165640
rect 406712 165628 406718 165640
rect 427078 165628 427084 165640
rect 406712 165600 427084 165628
rect 406712 165588 406718 165600
rect 427078 165588 427084 165600
rect 427136 165588 427142 165640
rect 442718 165588 442724 165640
rect 442776 165628 442782 165640
rect 442902 165628 442908 165640
rect 442776 165600 442908 165628
rect 442776 165588 442782 165600
rect 442902 165588 442908 165600
rect 442960 165628 442966 165640
rect 519170 165628 519176 165640
rect 442960 165600 519176 165628
rect 442960 165588 442966 165600
rect 519170 165588 519176 165600
rect 519228 165588 519234 165640
rect 3786 165520 3792 165572
rect 3844 165560 3850 165572
rect 4890 165560 4896 165572
rect 3844 165532 4896 165560
rect 3844 165520 3850 165532
rect 4890 165520 4896 165532
rect 4948 165520 4954 165572
rect 5258 165520 5264 165572
rect 5316 165560 5322 165572
rect 6270 165560 6276 165572
rect 5316 165532 6276 165560
rect 5316 165520 5322 165532
rect 6270 165520 6276 165532
rect 6328 165520 6334 165572
rect 409874 165452 409880 165504
rect 409932 165492 409938 165504
rect 422202 165492 422208 165504
rect 409932 165464 422208 165492
rect 409932 165452 409938 165464
rect 422202 165452 422208 165464
rect 422260 165452 422266 165504
rect 407666 165384 407672 165436
rect 407724 165424 407730 165436
rect 423122 165424 423128 165436
rect 407724 165396 423128 165424
rect 407724 165384 407730 165396
rect 423122 165384 423128 165396
rect 423180 165384 423186 165436
rect 408494 165316 408500 165368
rect 408552 165356 408558 165368
rect 429286 165356 429292 165368
rect 408552 165328 429292 165356
rect 408552 165316 408558 165328
rect 429286 165316 429292 165328
rect 429344 165316 429350 165368
rect 409506 165248 409512 165300
rect 409564 165288 409570 165300
rect 435358 165288 435364 165300
rect 409564 165260 435364 165288
rect 409564 165248 409570 165260
rect 435358 165248 435364 165260
rect 435416 165248 435422 165300
rect 404170 165180 404176 165232
rect 404228 165220 404234 165232
rect 430850 165220 430856 165232
rect 404228 165192 430856 165220
rect 404228 165180 404234 165192
rect 430850 165180 430856 165192
rect 430908 165180 430914 165232
rect 409230 165112 409236 165164
rect 409288 165152 409294 165164
rect 437980 165152 437986 165164
rect 409288 165124 437986 165152
rect 409288 165112 409294 165124
rect 437980 165112 437986 165124
rect 438038 165112 438044 165164
rect 409322 165044 409328 165096
rect 409380 165084 409386 165096
rect 441660 165084 441666 165096
rect 409380 165056 441666 165084
rect 409380 165044 409386 165056
rect 441660 165044 441666 165056
rect 441718 165084 441724 165096
rect 442718 165084 442724 165096
rect 441718 165056 442724 165084
rect 441718 165044 441724 165056
rect 442718 165044 442724 165056
rect 442776 165044 442782 165096
rect 386046 164976 386052 165028
rect 386104 165016 386110 165028
rect 419718 165016 419724 165028
rect 386104 164988 419724 165016
rect 386104 164976 386110 164988
rect 419718 164976 419724 164988
rect 419776 164976 419782 165028
rect 409414 164908 409420 164960
rect 409472 164948 409478 164960
rect 445202 164948 445208 164960
rect 409472 164920 445208 164948
rect 409472 164908 409478 164920
rect 445202 164908 445208 164920
rect 445260 164908 445266 164960
rect 448330 164908 448336 164960
rect 448388 164948 448394 164960
rect 469858 164948 469864 164960
rect 448388 164920 469864 164948
rect 448388 164908 448394 164920
rect 469858 164908 469864 164920
rect 469916 164908 469922 164960
rect 387702 164840 387708 164892
rect 387760 164880 387766 164892
rect 430758 164880 430764 164892
rect 387760 164852 430764 164880
rect 387760 164840 387766 164852
rect 430758 164840 430764 164852
rect 430816 164840 430822 164892
rect 445662 164840 445668 164892
rect 445720 164880 445726 164892
rect 523770 164880 523776 164892
rect 445720 164852 523776 164880
rect 445720 164840 445726 164852
rect 523770 164840 523776 164852
rect 523828 164840 523834 164892
rect 401594 163548 401600 163600
rect 401652 163588 401658 163600
rect 407666 163588 407672 163600
rect 401652 163560 407672 163588
rect 401652 163548 401658 163560
rect 407666 163548 407672 163560
rect 407724 163548 407730 163600
rect 394510 163412 394516 163464
rect 394568 163452 394574 163464
rect 404446 163452 404452 163464
rect 394568 163424 404452 163452
rect 394568 163412 394574 163424
rect 404446 163412 404452 163424
rect 404504 163412 404510 163464
rect 404354 163208 404360 163260
rect 404412 163248 404418 163260
rect 409874 163248 409880 163260
rect 404412 163220 409880 163248
rect 404412 163208 404418 163220
rect 409874 163208 409880 163220
rect 409932 163208 409938 163260
rect 405550 163140 405556 163192
rect 405608 163180 405614 163192
rect 408494 163180 408500 163192
rect 405608 163152 408500 163180
rect 405608 163140 405614 163152
rect 408494 163140 408500 163152
rect 408552 163140 408558 163192
rect 401410 161440 401416 161492
rect 401468 161480 401474 161492
rect 405550 161480 405556 161492
rect 401468 161452 405556 161480
rect 401468 161440 401474 161452
rect 405550 161440 405556 161452
rect 405608 161440 405614 161492
rect 456794 161236 456800 161288
rect 456852 161276 456858 161288
rect 459002 161276 459008 161288
rect 456852 161248 459008 161276
rect 456852 161236 456858 161248
rect 459002 161236 459008 161248
rect 459060 161236 459066 161288
rect 402422 160080 402428 160132
rect 402480 160120 402486 160132
rect 404354 160120 404360 160132
rect 402480 160092 404360 160120
rect 402480 160080 402486 160092
rect 404354 160080 404360 160092
rect 404412 160080 404418 160132
rect 456794 159944 456800 159996
rect 456852 159984 456858 159996
rect 459094 159984 459100 159996
rect 456852 159956 459100 159984
rect 456852 159944 456858 159956
rect 459094 159944 459100 159956
rect 459152 159944 459158 159996
rect 401594 158760 401600 158772
rect 398852 158732 401600 158760
rect 397178 158652 397184 158704
rect 397236 158692 397242 158704
rect 398852 158692 398880 158732
rect 401594 158720 401600 158732
rect 401652 158720 401658 158772
rect 397236 158664 398880 158692
rect 397236 158652 397242 158664
rect 456794 157020 456800 157072
rect 456852 157060 456858 157072
rect 458910 157060 458916 157072
rect 456852 157032 458916 157060
rect 456852 157020 456858 157032
rect 458910 157020 458916 157032
rect 458968 157020 458974 157072
rect 456794 155320 456800 155372
rect 456852 155360 456858 155372
rect 458726 155360 458732 155372
rect 456852 155332 458732 155360
rect 456852 155320 456858 155332
rect 458726 155320 458732 155332
rect 458784 155320 458790 155372
rect 406838 155252 406844 155304
rect 406896 155292 406902 155304
rect 409506 155292 409512 155304
rect 406896 155264 409512 155292
rect 406896 155252 406902 155264
rect 409506 155252 409512 155264
rect 409564 155252 409570 155304
rect 382274 154504 382280 154556
rect 382332 154544 382338 154556
rect 409414 154544 409420 154556
rect 382332 154516 409420 154544
rect 382332 154504 382338 154516
rect 409414 154504 409420 154516
rect 409472 154504 409478 154556
rect 456794 154096 456800 154148
rect 456852 154136 456858 154148
rect 458634 154136 458640 154148
rect 456852 154108 458640 154136
rect 456852 154096 456858 154108
rect 458634 154096 458640 154108
rect 458692 154096 458698 154148
rect 486418 153824 486424 153876
rect 486476 153864 486482 153876
rect 528554 153864 528560 153876
rect 486476 153836 528560 153864
rect 486476 153824 486482 153836
rect 528554 153824 528560 153836
rect 528612 153824 528618 153876
rect 504358 153144 504364 153196
rect 504416 153184 504422 153196
rect 505462 153184 505468 153196
rect 504416 153156 505468 153184
rect 504416 153144 504422 153156
rect 505462 153144 505468 153156
rect 505520 153144 505526 153196
rect 544378 153144 544384 153196
rect 544436 153184 544442 153196
rect 580166 153184 580172 153196
rect 544436 153156 580172 153184
rect 544436 153144 544442 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 392394 152464 392400 152516
rect 392452 152504 392458 152516
rect 398466 152504 398472 152516
rect 392452 152476 398472 152504
rect 392452 152464 392458 152476
rect 398466 152464 398472 152476
rect 398524 152464 398530 152516
rect 537478 152464 537484 152516
rect 537536 152504 537542 152516
rect 542906 152504 542912 152516
rect 537536 152476 542912 152504
rect 537536 152464 537542 152476
rect 542906 152464 542912 152476
rect 542964 152464 542970 152516
rect 508498 151852 508504 151904
rect 508556 151892 508562 151904
rect 510062 151892 510068 151904
rect 508556 151864 510068 151892
rect 508556 151852 508562 151864
rect 510062 151852 510068 151864
rect 510120 151852 510126 151904
rect 542906 151784 542912 151836
rect 542964 151824 542970 151836
rect 551462 151824 551468 151836
rect 542964 151796 551468 151824
rect 542964 151784 542970 151796
rect 551462 151784 551468 151796
rect 551520 151784 551526 151836
rect 3694 150696 3700 150748
rect 3752 150736 3758 150748
rect 5258 150736 5264 150748
rect 3752 150708 5264 150736
rect 3752 150696 3758 150708
rect 5258 150696 5264 150708
rect 5316 150696 5322 150748
rect 456886 150628 456892 150680
rect 456944 150668 456950 150680
rect 459370 150668 459376 150680
rect 456944 150640 459376 150668
rect 456944 150628 456950 150640
rect 459370 150628 459376 150640
rect 459428 150628 459434 150680
rect 400214 150492 400220 150544
rect 400272 150532 400278 150544
rect 402422 150532 402428 150544
rect 400272 150504 402428 150532
rect 400272 150492 400278 150504
rect 402422 150492 402428 150504
rect 402480 150492 402486 150544
rect 5166 150424 5172 150476
rect 5224 150464 5230 150476
rect 6454 150464 6460 150476
rect 5224 150436 6460 150464
rect 5224 150424 5230 150436
rect 6454 150424 6460 150436
rect 6512 150424 6518 150476
rect 399938 150424 399944 150476
rect 399996 150464 400002 150476
rect 401410 150464 401416 150476
rect 399996 150436 401416 150464
rect 399996 150424 400002 150436
rect 401410 150424 401416 150436
rect 401468 150424 401474 150476
rect 456794 150152 456800 150204
rect 456852 150192 456858 150204
rect 459462 150192 459468 150204
rect 456852 150164 459468 150192
rect 456852 150152 456858 150164
rect 459462 150152 459468 150164
rect 459520 150152 459526 150204
rect 542998 149676 543004 149728
rect 543056 149716 543062 149728
rect 552658 149716 552664 149728
rect 543056 149688 552664 149716
rect 543056 149676 543062 149688
rect 552658 149676 552664 149688
rect 552716 149676 552722 149728
rect 548610 149472 548616 149524
rect 548668 149512 548674 149524
rect 552842 149512 552848 149524
rect 548668 149484 552848 149512
rect 548668 149472 548674 149484
rect 552842 149472 552848 149484
rect 552900 149472 552906 149524
rect 548518 149404 548524 149456
rect 548576 149444 548582 149456
rect 552106 149444 552112 149456
rect 548576 149416 552112 149444
rect 548576 149404 548582 149416
rect 552106 149404 552112 149416
rect 552164 149404 552170 149456
rect 388162 149064 388168 149116
rect 388220 149104 388226 149116
rect 392394 149104 392400 149116
rect 388220 149076 392400 149104
rect 388220 149064 388226 149076
rect 392394 149064 392400 149076
rect 392452 149064 392458 149116
rect 384850 147636 384856 147688
rect 384908 147676 384914 147688
rect 387702 147676 387708 147688
rect 384908 147648 387708 147676
rect 384908 147636 384914 147648
rect 387702 147636 387708 147648
rect 387760 147636 387766 147688
rect 395890 147636 395896 147688
rect 395948 147676 395954 147688
rect 400214 147676 400220 147688
rect 395948 147648 400220 147676
rect 395948 147636 395954 147648
rect 400214 147636 400220 147648
rect 400272 147636 400278 147688
rect 549162 146004 549168 146056
rect 549220 146044 549226 146056
rect 549898 146044 549904 146056
rect 549220 146016 549904 146044
rect 549220 146004 549226 146016
rect 549898 146004 549904 146016
rect 549956 146004 549962 146056
rect 456794 144644 456800 144696
rect 456852 144684 456858 144696
rect 458818 144684 458824 144696
rect 456852 144656 458824 144684
rect 456852 144644 456858 144656
rect 458818 144644 458824 144656
rect 458876 144644 458882 144696
rect 382274 143488 382280 143540
rect 382332 143528 382338 143540
rect 409322 143528 409328 143540
rect 382332 143500 409328 143528
rect 382332 143488 382338 143500
rect 409322 143488 409328 143500
rect 409380 143488 409386 143540
rect 456794 143148 456800 143200
rect 456852 143188 456858 143200
rect 459278 143188 459284 143200
rect 456852 143160 459284 143188
rect 456852 143148 456858 143160
rect 459278 143148 459284 143160
rect 459336 143148 459342 143200
rect 386230 142944 386236 142996
rect 386288 142984 386294 142996
rect 388162 142984 388168 142996
rect 386288 142956 388168 142984
rect 386288 142944 386294 142956
rect 388162 142944 388168 142956
rect 388220 142944 388226 142996
rect 552106 142876 552112 142928
rect 552164 142916 552170 142928
rect 552658 142916 552664 142928
rect 552164 142888 552664 142916
rect 552164 142876 552170 142888
rect 552658 142876 552664 142888
rect 552716 142876 552722 142928
rect 552658 142740 552664 142792
rect 552716 142780 552722 142792
rect 552842 142780 552848 142792
rect 552716 142752 552848 142780
rect 552716 142740 552722 142752
rect 552842 142740 552848 142752
rect 552900 142740 552906 142792
rect 457254 141652 457260 141704
rect 457312 141692 457318 141704
rect 460106 141692 460112 141704
rect 457312 141664 460112 141692
rect 457312 141652 457318 141664
rect 460106 141652 460112 141664
rect 460164 141652 460170 141704
rect 456794 140428 456800 140480
rect 456852 140468 456858 140480
rect 459186 140468 459192 140480
rect 456852 140440 459192 140468
rect 456852 140428 456858 140440
rect 459186 140428 459192 140440
rect 459244 140428 459250 140480
rect 5074 140088 5080 140140
rect 5132 140128 5138 140140
rect 6362 140128 6368 140140
rect 5132 140100 6368 140128
rect 5132 140088 5138 140100
rect 6362 140088 6368 140100
rect 6420 140088 6426 140140
rect 576118 139340 576124 139392
rect 576176 139380 576182 139392
rect 580166 139380 580172 139392
rect 576176 139352 580172 139380
rect 576176 139340 576182 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 457254 138864 457260 138916
rect 457312 138904 457318 138916
rect 460750 138904 460756 138916
rect 457312 138876 460756 138904
rect 457312 138864 457318 138876
rect 460750 138864 460756 138876
rect 460808 138864 460814 138916
rect 3510 138320 3516 138372
rect 3568 138360 3574 138372
rect 5074 138360 5080 138372
rect 3568 138332 5080 138360
rect 3568 138320 3574 138332
rect 5074 138320 5080 138332
rect 5132 138320 5138 138372
rect 394418 137980 394424 138032
rect 394476 138020 394482 138032
rect 395890 138020 395896 138032
rect 394476 137992 395896 138020
rect 394476 137980 394482 137992
rect 395890 137980 395896 137992
rect 395948 137980 395954 138032
rect 457254 137844 457260 137896
rect 457312 137884 457318 137896
rect 460474 137884 460480 137896
rect 457312 137856 460480 137884
rect 457312 137844 457318 137856
rect 460474 137844 460480 137856
rect 460532 137844 460538 137896
rect 390554 137368 390560 137420
rect 390612 137408 390618 137420
rect 394510 137408 394516 137420
rect 390612 137380 394516 137408
rect 390612 137368 390618 137380
rect 394510 137368 394516 137380
rect 394568 137368 394574 137420
rect 384942 133560 384948 133612
rect 385000 133600 385006 133612
rect 390554 133600 390560 133612
rect 385000 133572 390560 133600
rect 385000 133560 385006 133572
rect 390554 133560 390560 133572
rect 390612 133560 390618 133612
rect 457070 132880 457076 132932
rect 457128 132920 457134 132932
rect 460658 132920 460664 132932
rect 457128 132892 460664 132920
rect 457128 132880 457134 132892
rect 460658 132880 460664 132892
rect 460716 132880 460722 132932
rect 382274 132404 382280 132456
rect 382332 132444 382338 132456
rect 409230 132444 409236 132456
rect 382332 132416 409236 132444
rect 382332 132404 382338 132416
rect 409230 132404 409236 132416
rect 409288 132404 409294 132456
rect 382182 131112 382188 131164
rect 382240 131152 382246 131164
rect 384850 131152 384856 131164
rect 382240 131124 384856 131152
rect 382240 131112 382246 131124
rect 384850 131112 384856 131124
rect 384908 131112 384914 131164
rect 457438 128188 457444 128240
rect 457496 128228 457502 128240
rect 460566 128228 460572 128240
rect 457496 128200 460572 128228
rect 457496 128188 457502 128200
rect 460566 128188 460572 128200
rect 460624 128188 460630 128240
rect 405274 127508 405280 127560
rect 405332 127548 405338 127560
rect 406838 127548 406844 127560
rect 405332 127520 406844 127548
rect 405332 127508 405338 127520
rect 406838 127508 406844 127520
rect 406896 127508 406902 127560
rect 558178 126896 558184 126948
rect 558236 126936 558242 126948
rect 580166 126936 580172 126948
rect 558236 126908 580172 126936
rect 558236 126896 558242 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 395890 125468 395896 125520
rect 395948 125508 395954 125520
rect 397178 125508 397184 125520
rect 395948 125480 397184 125508
rect 395948 125468 395954 125480
rect 397178 125468 397184 125480
rect 397236 125468 397242 125520
rect 457346 125196 457352 125248
rect 457404 125236 457410 125248
rect 460382 125236 460388 125248
rect 457404 125208 460388 125236
rect 457404 125196 457410 125208
rect 460382 125196 460388 125208
rect 460440 125196 460446 125248
rect 457070 122544 457076 122596
rect 457128 122584 457134 122596
rect 460290 122584 460296 122596
rect 457128 122556 460296 122584
rect 457128 122544 457134 122556
rect 460290 122544 460296 122556
rect 460348 122544 460354 122596
rect 405274 121496 405280 121508
rect 402946 121468 405280 121496
rect 400214 121388 400220 121440
rect 400272 121428 400278 121440
rect 402946 121428 402974 121468
rect 405274 121456 405280 121468
rect 405332 121456 405338 121508
rect 400272 121400 402974 121428
rect 400272 121388 400278 121400
rect 380618 118872 380624 118924
rect 380676 118912 380682 118924
rect 384942 118912 384948 118924
rect 380676 118884 384948 118912
rect 380676 118872 380682 118884
rect 384942 118872 384948 118884
rect 385000 118872 385006 118924
rect 399938 115988 399944 116000
rect 396092 115960 399944 115988
rect 3970 115880 3976 115932
rect 4028 115920 4034 115932
rect 5166 115920 5172 115932
rect 4028 115892 5172 115920
rect 4028 115880 4034 115892
rect 5166 115880 5172 115892
rect 5224 115880 5230 115932
rect 5350 115880 5356 115932
rect 5408 115920 5414 115932
rect 6546 115920 6552 115932
rect 5408 115892 6552 115920
rect 5408 115880 5414 115892
rect 6546 115880 6552 115892
rect 6604 115880 6610 115932
rect 395982 115880 395988 115932
rect 396040 115920 396046 115932
rect 396092 115920 396120 115960
rect 399938 115948 399944 115960
rect 399996 115948 400002 116000
rect 396040 115892 396120 115920
rect 396040 115880 396046 115892
rect 394510 115540 394516 115592
rect 394568 115580 394574 115592
rect 395890 115580 395896 115592
rect 394568 115552 395896 115580
rect 394568 115540 394574 115552
rect 395890 115540 395896 115552
rect 395948 115540 395954 115592
rect 397362 115200 397368 115252
rect 397420 115240 397426 115252
rect 400122 115240 400128 115252
rect 397420 115212 400128 115240
rect 397420 115200 397426 115212
rect 400122 115200 400128 115212
rect 400180 115200 400186 115252
rect 6178 114588 6184 114640
rect 6236 114628 6242 114640
rect 7742 114628 7748 114640
rect 6236 114600 7748 114628
rect 6236 114588 6242 114600
rect 7742 114588 7748 114600
rect 7800 114588 7806 114640
rect 395982 113200 395988 113212
rect 391952 113172 395988 113200
rect 391658 113092 391664 113144
rect 391716 113132 391722 113144
rect 391952 113132 391980 113172
rect 395982 113160 395988 113172
rect 396040 113160 396046 113212
rect 391716 113104 391980 113132
rect 391716 113092 391722 113104
rect 562318 113092 562324 113144
rect 562376 113132 562382 113144
rect 579798 113132 579804 113144
rect 562376 113104 579804 113132
rect 562376 113092 562382 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 391106 111800 391112 111852
rect 391164 111840 391170 111852
rect 394418 111840 394424 111852
rect 391164 111812 394424 111840
rect 391164 111800 391170 111812
rect 394418 111800 394424 111812
rect 394476 111800 394482 111852
rect 382274 111732 382280 111784
rect 382332 111772 382338 111784
rect 404170 111772 404176 111784
rect 382332 111744 404176 111772
rect 382332 111732 382338 111744
rect 404170 111732 404176 111744
rect 404228 111732 404234 111784
rect 393130 111052 393136 111104
rect 393188 111092 393194 111104
rect 397362 111092 397368 111104
rect 393188 111064 397368 111092
rect 393188 111052 393194 111064
rect 397362 111052 397368 111064
rect 397420 111052 397426 111104
rect 6270 108944 6276 108996
rect 6328 108984 6334 108996
rect 7558 108984 7564 108996
rect 6328 108956 7564 108984
rect 6328 108944 6334 108956
rect 7558 108944 7564 108956
rect 7616 108944 7622 108996
rect 6454 104864 6460 104916
rect 6512 104904 6518 104916
rect 7650 104904 7656 104916
rect 6512 104876 7656 104904
rect 6512 104864 6518 104876
rect 7650 104864 7656 104876
rect 7708 104864 7714 104916
rect 5166 104796 5172 104848
rect 5224 104836 5230 104848
rect 6270 104836 6276 104848
rect 5224 104808 6276 104836
rect 5224 104796 5230 104808
rect 6270 104796 6276 104808
rect 6328 104796 6334 104848
rect 4982 104728 4988 104780
rect 5040 104768 5046 104780
rect 6178 104768 6184 104780
rect 5040 104740 6184 104768
rect 5040 104728 5046 104740
rect 6178 104728 6184 104740
rect 6236 104728 6242 104780
rect 391106 103544 391112 103556
rect 389192 103516 391112 103544
rect 388806 103436 388812 103488
rect 388864 103476 388870 103488
rect 389192 103476 389220 103516
rect 391106 103504 391112 103516
rect 391164 103504 391170 103556
rect 388864 103448 389220 103476
rect 388864 103436 388870 103448
rect 3418 102144 3424 102196
rect 3476 102184 3482 102196
rect 5166 102184 5172 102196
rect 3476 102156 5172 102184
rect 3476 102144 3482 102156
rect 5166 102144 5172 102156
rect 5224 102144 5230 102196
rect 3878 101532 3884 101584
rect 3936 101572 3942 101584
rect 4982 101572 4988 101584
rect 3936 101544 4988 101572
rect 3936 101532 3942 101544
rect 4982 101532 4988 101544
rect 5040 101532 5046 101584
rect 385034 100716 385040 100768
rect 385092 100756 385098 100768
rect 393130 100756 393136 100768
rect 385092 100728 393136 100756
rect 385092 100716 385098 100728
rect 393130 100716 393136 100728
rect 393188 100716 393194 100768
rect 382274 100648 382280 100700
rect 382332 100688 382338 100700
rect 406654 100688 406660 100700
rect 382332 100660 406660 100688
rect 382332 100648 382338 100660
rect 406654 100648 406660 100660
rect 406712 100648 406718 100700
rect 574738 100648 574744 100700
rect 574796 100688 574802 100700
rect 580166 100688 580172 100700
rect 574796 100660 580172 100688
rect 574796 100648 574802 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 391750 99968 391756 100020
rect 391808 100008 391814 100020
rect 394510 100008 394516 100020
rect 391808 99980 394516 100008
rect 391808 99968 391814 99980
rect 394510 99968 394516 99980
rect 394568 99968 394574 100020
rect 385034 99396 385040 99408
rect 383626 99368 385040 99396
rect 383470 99288 383476 99340
rect 383528 99328 383534 99340
rect 383626 99328 383654 99368
rect 385034 99356 385040 99368
rect 385092 99356 385098 99408
rect 383528 99300 383654 99328
rect 383528 99288 383534 99300
rect 3418 96636 3424 96688
rect 3476 96676 3482 96688
rect 20898 96676 20904 96688
rect 3476 96648 20904 96676
rect 3476 96636 3482 96648
rect 20898 96636 20904 96648
rect 20956 96636 20962 96688
rect 6270 96092 6276 96144
rect 6328 96132 6334 96144
rect 8202 96132 8208 96144
rect 6328 96104 8208 96132
rect 6328 96092 6334 96104
rect 8202 96092 8208 96104
rect 8260 96092 8266 96144
rect 5166 91196 5172 91248
rect 5224 91236 5230 91248
rect 6270 91236 6276 91248
rect 5224 91208 6276 91236
rect 5224 91196 5230 91208
rect 6270 91196 6276 91208
rect 6328 91196 6334 91248
rect 380710 91060 380716 91112
rect 380768 91100 380774 91112
rect 383470 91100 383476 91112
rect 380768 91072 383476 91100
rect 380768 91060 380774 91072
rect 383470 91060 383476 91072
rect 383528 91060 383534 91112
rect 6362 90924 6368 90976
rect 6420 90964 6426 90976
rect 7926 90964 7932 90976
rect 6420 90936 7932 90964
rect 6420 90924 6426 90936
rect 7926 90924 7932 90936
rect 7984 90924 7990 90976
rect 3694 90312 3700 90364
rect 3752 90352 3758 90364
rect 10962 90352 10968 90364
rect 3752 90324 10968 90352
rect 3752 90312 3758 90324
rect 10962 90312 10968 90324
rect 11020 90312 11026 90364
rect 3786 89700 3792 89752
rect 3844 89740 3850 89752
rect 5442 89740 5448 89752
rect 3844 89712 5448 89740
rect 3844 89700 3850 89712
rect 5442 89700 5448 89712
rect 5500 89700 5506 89752
rect 382274 89632 382280 89684
rect 382332 89672 382338 89684
rect 409138 89672 409144 89684
rect 382332 89644 409144 89672
rect 382332 89632 382338 89644
rect 409138 89632 409144 89644
rect 409196 89632 409202 89684
rect 8294 88272 8300 88324
rect 8352 88312 8358 88324
rect 11698 88312 11704 88324
rect 8352 88284 11704 88312
rect 8352 88272 8358 88284
rect 11698 88272 11704 88284
rect 11756 88272 11762 88324
rect 381446 87864 381452 87916
rect 381504 87904 381510 87916
rect 384758 87904 384764 87916
rect 381504 87876 384764 87904
rect 381504 87864 381510 87876
rect 384758 87864 384764 87876
rect 384816 87864 384822 87916
rect 383470 87320 383476 87372
rect 383528 87360 383534 87372
rect 386138 87360 386144 87372
rect 383528 87332 386144 87360
rect 383528 87320 383534 87332
rect 386138 87320 386144 87332
rect 386196 87320 386202 87372
rect 555418 86912 555424 86964
rect 555476 86952 555482 86964
rect 580166 86952 580172 86964
rect 555476 86924 580172 86952
rect 555476 86912 555482 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 5534 86572 5540 86624
rect 5592 86612 5598 86624
rect 8018 86612 8024 86624
rect 5592 86584 8024 86612
rect 5592 86572 5598 86584
rect 8018 86572 8024 86584
rect 8076 86572 8082 86624
rect 382826 86232 382832 86284
rect 382884 86272 382890 86284
rect 387610 86272 387616 86284
rect 382884 86244 387616 86272
rect 382884 86232 382890 86244
rect 387610 86232 387616 86244
rect 387668 86232 387674 86284
rect 383562 85552 383568 85604
rect 383620 85592 383626 85604
rect 386230 85592 386236 85604
rect 383620 85564 386236 85592
rect 383620 85552 383626 85564
rect 386230 85552 386236 85564
rect 386288 85552 386294 85604
rect 388806 85592 388812 85604
rect 386432 85564 388812 85592
rect 11054 85484 11060 85536
rect 11112 85524 11118 85536
rect 13722 85524 13728 85536
rect 11112 85496 13728 85524
rect 11112 85484 11118 85496
rect 13722 85484 13728 85496
rect 13780 85484 13786 85536
rect 386138 85484 386144 85536
rect 386196 85524 386202 85536
rect 386432 85524 386460 85564
rect 388806 85552 388812 85564
rect 388864 85552 388870 85604
rect 386196 85496 386460 85524
rect 386196 85484 386202 85496
rect 387610 85484 387616 85536
rect 387668 85524 387674 85536
rect 388714 85524 388720 85536
rect 387668 85496 388720 85524
rect 387668 85484 387674 85496
rect 388714 85484 388720 85496
rect 388772 85484 388778 85536
rect 6546 84260 6552 84312
rect 6604 84300 6610 84312
rect 7834 84300 7840 84312
rect 6604 84272 7840 84300
rect 6604 84260 6610 84272
rect 7834 84260 7840 84272
rect 7892 84260 7898 84312
rect 3326 84192 3332 84244
rect 3384 84232 3390 84244
rect 18598 84232 18604 84244
rect 3384 84204 18604 84232
rect 3384 84192 3390 84204
rect 18598 84192 18604 84204
rect 18656 84192 18662 84244
rect 391658 84232 391664 84244
rect 389192 84204 391664 84232
rect 387794 84124 387800 84176
rect 387852 84164 387858 84176
rect 389192 84164 389220 84204
rect 391658 84192 391664 84204
rect 391716 84192 391722 84244
rect 387852 84136 389220 84164
rect 387852 84124 387858 84136
rect 5074 83172 5080 83224
rect 5132 83212 5138 83224
rect 5994 83212 6000 83224
rect 5132 83184 6000 83212
rect 5132 83172 5138 83184
rect 5994 83172 6000 83184
rect 6052 83172 6058 83224
rect 384758 82832 384764 82884
rect 384816 82872 384822 82884
rect 387610 82872 387616 82884
rect 384816 82844 387616 82872
rect 384816 82832 384822 82844
rect 387610 82832 387616 82844
rect 387668 82832 387674 82884
rect 389450 82832 389456 82884
rect 389508 82872 389514 82884
rect 391750 82872 391756 82884
rect 389508 82844 391756 82872
rect 389508 82832 389514 82844
rect 391750 82832 391756 82844
rect 391808 82832 391814 82884
rect 7742 82084 7748 82136
rect 7800 82124 7806 82136
rect 9122 82124 9128 82136
rect 7800 82096 9128 82124
rect 7800 82084 7806 82096
rect 9122 82084 9128 82096
rect 9180 82084 9186 82136
rect 11698 81404 11704 81456
rect 11756 81444 11762 81456
rect 11756 81416 12480 81444
rect 11756 81404 11762 81416
rect 12452 81376 12480 81416
rect 386230 81404 386236 81456
rect 386288 81444 386294 81456
rect 387794 81444 387800 81456
rect 386288 81416 387800 81444
rect 386288 81404 386294 81416
rect 387794 81404 387800 81416
rect 387852 81404 387858 81456
rect 15838 81376 15844 81388
rect 12452 81348 15844 81376
rect 15838 81336 15844 81348
rect 15896 81336 15902 81388
rect 4982 80044 4988 80096
rect 5040 80084 5046 80096
rect 5040 80056 6914 80084
rect 5040 80044 5046 80056
rect 6886 80016 6914 80056
rect 387610 80044 387616 80096
rect 387668 80084 387674 80096
rect 389450 80084 389456 80096
rect 387668 80056 389456 80084
rect 387668 80044 387674 80056
rect 389450 80044 389456 80056
rect 389508 80044 389514 80096
rect 8386 80016 8392 80028
rect 6886 79988 8392 80016
rect 8386 79976 8392 79988
rect 8444 79976 8450 80028
rect 382274 79908 382280 79960
rect 382332 79948 382338 79960
rect 386046 79948 386052 79960
rect 382332 79920 386052 79948
rect 382332 79908 382338 79920
rect 386046 79908 386052 79920
rect 386104 79908 386110 79960
rect 13722 78684 13728 78736
rect 13780 78724 13786 78736
rect 13780 78696 16574 78724
rect 13780 78684 13786 78696
rect 4890 78616 4896 78668
rect 4948 78656 4954 78668
rect 7742 78656 7748 78668
rect 4948 78628 7748 78656
rect 4948 78616 4954 78628
rect 7742 78616 7748 78628
rect 7800 78616 7806 78668
rect 16546 78656 16574 78696
rect 17218 78656 17224 78668
rect 16546 78628 17224 78656
rect 17218 78616 17224 78628
rect 17276 78616 17282 78668
rect 5994 78548 6000 78600
rect 6052 78588 6058 78600
rect 8938 78588 8944 78600
rect 6052 78560 8944 78588
rect 6052 78548 6058 78560
rect 8938 78548 8944 78560
rect 8996 78548 9002 78600
rect 5534 78480 5540 78532
rect 5592 78520 5598 78532
rect 9030 78520 9036 78532
rect 5592 78492 9036 78520
rect 5592 78480 5598 78492
rect 9030 78480 9036 78492
rect 9088 78480 9094 78532
rect 9030 76440 9036 76492
rect 9088 76480 9094 76492
rect 10962 76480 10968 76492
rect 9088 76452 10968 76480
rect 9088 76440 9094 76452
rect 10962 76440 10968 76452
rect 11020 76440 11026 76492
rect 9122 75828 9128 75880
rect 9180 75868 9186 75880
rect 10318 75868 10324 75880
rect 9180 75840 10324 75868
rect 9180 75828 9186 75840
rect 10318 75828 10324 75840
rect 10376 75828 10382 75880
rect 8386 75760 8392 75812
rect 8444 75800 8450 75812
rect 11698 75800 11704 75812
rect 8444 75772 11704 75800
rect 8444 75760 8450 75772
rect 11698 75760 11704 75772
rect 11756 75760 11762 75812
rect 6270 75148 6276 75200
rect 6328 75188 6334 75200
rect 6914 75188 6920 75200
rect 6328 75160 6920 75188
rect 6328 75148 6334 75160
rect 6914 75148 6920 75160
rect 6972 75148 6978 75200
rect 15838 73176 15844 73228
rect 15896 73216 15902 73228
rect 17310 73216 17316 73228
rect 15896 73188 17316 73216
rect 15896 73176 15902 73188
rect 17310 73176 17316 73188
rect 17368 73176 17374 73228
rect 386046 73176 386052 73228
rect 386104 73216 386110 73228
rect 387610 73216 387616 73228
rect 386104 73188 387616 73216
rect 386104 73176 386110 73188
rect 387610 73176 387616 73188
rect 387668 73176 387674 73228
rect 559558 73108 559564 73160
rect 559616 73148 559622 73160
rect 580166 73148 580172 73160
rect 559616 73120 580172 73148
rect 559616 73108 559622 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 6914 72564 6920 72616
rect 6972 72604 6978 72616
rect 9582 72604 9588 72616
rect 6972 72576 9588 72604
rect 6972 72564 6978 72576
rect 9582 72564 9588 72576
rect 9640 72564 9646 72616
rect 7742 70932 7748 70984
rect 7800 70972 7806 70984
rect 9398 70972 9404 70984
rect 7800 70944 9404 70972
rect 7800 70932 7806 70944
rect 9398 70932 9404 70944
rect 9456 70932 9462 70984
rect 8294 70184 8300 70236
rect 8352 70224 8358 70236
rect 10410 70224 10416 70236
rect 8352 70196 10416 70224
rect 8352 70184 8358 70196
rect 10410 70184 10416 70196
rect 10468 70184 10474 70236
rect 3602 70116 3608 70168
rect 3660 70156 3666 70168
rect 4982 70156 4988 70168
rect 3660 70128 4988 70156
rect 3660 70116 3666 70128
rect 4982 70116 4988 70128
rect 5040 70116 5046 70168
rect 4798 70048 4804 70100
rect 4856 70088 4862 70100
rect 5534 70088 5540 70100
rect 4856 70060 5540 70088
rect 4856 70048 4862 70060
rect 5534 70048 5540 70060
rect 5592 70048 5598 70100
rect 382274 68960 382280 69012
rect 382332 69000 382338 69012
rect 408034 69000 408040 69012
rect 382332 68972 408040 69000
rect 382332 68960 382338 68972
rect 408034 68960 408040 68972
rect 408092 68960 408098 69012
rect 10962 67600 10968 67652
rect 11020 67640 11026 67652
rect 11020 67612 12572 67640
rect 11020 67600 11026 67612
rect 9674 67532 9680 67584
rect 9732 67572 9738 67584
rect 12250 67572 12256 67584
rect 9732 67544 12256 67572
rect 9732 67532 9738 67544
rect 12250 67532 12256 67544
rect 12308 67532 12314 67584
rect 12544 67572 12572 67612
rect 15102 67572 15108 67584
rect 12544 67544 15108 67572
rect 15102 67532 15108 67544
rect 15160 67532 15166 67584
rect 9398 67464 9404 67516
rect 9456 67504 9462 67516
rect 10962 67504 10968 67516
rect 9456 67476 10968 67504
rect 9456 67464 9462 67476
rect 10962 67464 10968 67476
rect 11020 67464 11026 67516
rect 8938 66172 8944 66224
rect 8996 66212 9002 66224
rect 12342 66212 12348 66224
rect 8996 66184 12348 66212
rect 8996 66172 9002 66184
rect 12342 66172 12348 66184
rect 12400 66172 12406 66224
rect 5534 65152 5540 65204
rect 5592 65192 5598 65204
rect 7742 65192 7748 65204
rect 5592 65164 7748 65192
rect 5592 65152 5598 65164
rect 7742 65152 7748 65164
rect 7800 65152 7806 65204
rect 4982 65084 4988 65136
rect 5040 65124 5046 65136
rect 7282 65124 7288 65136
rect 5040 65096 7288 65124
rect 5040 65084 5046 65096
rect 7282 65084 7288 65096
rect 7340 65084 7346 65136
rect 11698 64880 11704 64932
rect 11756 64920 11762 64932
rect 11756 64892 12480 64920
rect 11756 64880 11762 64892
rect 12452 64852 12480 64892
rect 15102 64852 15108 64864
rect 12452 64824 15108 64852
rect 15102 64812 15108 64824
rect 15160 64812 15166 64864
rect 17310 63384 17316 63436
rect 17368 63424 17374 63436
rect 18690 63424 18696 63436
rect 17368 63396 18696 63424
rect 17368 63384 17374 63396
rect 18690 63384 18696 63396
rect 18748 63384 18754 63436
rect 10962 63248 10968 63300
rect 11020 63288 11026 63300
rect 14458 63288 14464 63300
rect 11020 63260 14464 63288
rect 11020 63248 11026 63260
rect 14458 63248 14464 63260
rect 14516 63248 14522 63300
rect 7282 61004 7288 61056
rect 7340 61044 7346 61056
rect 11238 61044 11244 61056
rect 7340 61016 11244 61044
rect 7340 61004 7346 61016
rect 11238 61004 11244 61016
rect 11296 61004 11302 61056
rect 10410 60732 10416 60784
rect 10468 60772 10474 60784
rect 10468 60744 11100 60772
rect 10468 60732 10474 60744
rect 11072 60636 11100 60744
rect 12250 60664 12256 60716
rect 12308 60704 12314 60716
rect 13814 60704 13820 60716
rect 12308 60676 13820 60704
rect 12308 60664 12314 60676
rect 13814 60664 13820 60676
rect 13872 60664 13878 60716
rect 573358 60664 573364 60716
rect 573416 60704 573422 60716
rect 580166 60704 580172 60716
rect 573416 60676 580172 60704
rect 573416 60664 573422 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 13538 60636 13544 60648
rect 11072 60608 13544 60636
rect 13538 60596 13544 60608
rect 13596 60596 13602 60648
rect 12434 59372 12440 59424
rect 12492 59412 12498 59424
rect 12492 59384 14136 59412
rect 12492 59372 12498 59384
rect 14108 59276 14136 59384
rect 15194 59304 15200 59356
rect 15252 59344 15258 59356
rect 17310 59344 17316 59356
rect 15252 59316 17316 59344
rect 15252 59304 15258 59316
rect 17310 59304 17316 59316
rect 17368 59304 17374 59356
rect 17862 59276 17868 59288
rect 14108 59248 17868 59276
rect 17862 59236 17868 59248
rect 17920 59236 17926 59288
rect 13814 59168 13820 59220
rect 13872 59208 13878 59220
rect 17402 59208 17408 59220
rect 13872 59180 17408 59208
rect 13872 59168 13878 59180
rect 17402 59168 17408 59180
rect 17460 59168 17466 59220
rect 15286 59100 15292 59152
rect 15344 59140 15350 59152
rect 18874 59140 18880 59152
rect 15344 59112 18880 59140
rect 15344 59100 15350 59112
rect 18874 59100 18880 59112
rect 18932 59100 18938 59152
rect 8294 57876 8300 57928
rect 8352 57916 8358 57928
rect 13262 57916 13268 57928
rect 8352 57888 13268 57916
rect 8352 57876 8358 57888
rect 13262 57876 13268 57888
rect 13320 57876 13326 57928
rect 17218 57876 17224 57928
rect 17276 57916 17282 57928
rect 18322 57916 18328 57928
rect 17276 57888 18328 57916
rect 17276 57876 17282 57888
rect 18322 57876 18328 57888
rect 18380 57876 18386 57928
rect 382274 57876 382280 57928
rect 382332 57916 382338 57928
rect 391566 57916 391572 57928
rect 382332 57888 391572 57916
rect 382332 57876 382338 57888
rect 391566 57876 391572 57888
rect 391624 57876 391630 57928
rect 6178 56924 6184 56976
rect 6236 56964 6242 56976
rect 8202 56964 8208 56976
rect 6236 56936 8208 56964
rect 6236 56924 6242 56936
rect 8202 56924 8208 56936
rect 8260 56924 8266 56976
rect 11238 56584 11244 56636
rect 11296 56624 11302 56636
rect 11296 56596 13860 56624
rect 11296 56584 11302 56596
rect 7650 56516 7656 56568
rect 7708 56556 7714 56568
rect 8662 56556 8668 56568
rect 7708 56528 8668 56556
rect 7708 56516 7714 56528
rect 8662 56516 8668 56528
rect 8720 56516 8726 56568
rect 13832 56556 13860 56596
rect 16482 56556 16488 56568
rect 13832 56528 16488 56556
rect 16482 56516 16488 56528
rect 16540 56516 16546 56568
rect 7834 56448 7840 56500
rect 7892 56488 7898 56500
rect 10962 56488 10968 56500
rect 7892 56460 10968 56488
rect 7892 56448 7898 56460
rect 10962 56448 10968 56460
rect 11020 56448 11026 56500
rect 7558 56380 7564 56432
rect 7616 56420 7622 56432
rect 10870 56420 10876 56432
rect 7616 56392 10876 56420
rect 7616 56380 7622 56392
rect 10870 56380 10876 56392
rect 10928 56380 10934 56432
rect 13538 55428 13544 55480
rect 13596 55468 13602 55480
rect 18046 55468 18052 55480
rect 13596 55440 18052 55468
rect 13596 55428 13602 55440
rect 18046 55428 18052 55440
rect 18104 55428 18110 55480
rect 14458 54612 14464 54664
rect 14516 54652 14522 54664
rect 15562 54652 15568 54664
rect 14516 54624 15568 54652
rect 14516 54612 14522 54624
rect 15562 54612 15568 54624
rect 15620 54612 15626 54664
rect 17402 54068 17408 54120
rect 17460 54108 17466 54120
rect 19334 54108 19340 54120
rect 17460 54080 19340 54108
rect 17460 54068 17466 54080
rect 19334 54068 19340 54080
rect 19392 54068 19398 54120
rect 10318 53796 10324 53848
rect 10376 53836 10382 53848
rect 10376 53808 11100 53836
rect 10376 53796 10382 53808
rect 11072 53768 11100 53808
rect 15194 53768 15200 53780
rect 11072 53740 15200 53768
rect 15194 53728 15200 53740
rect 15252 53728 15258 53780
rect 11054 53660 11060 53712
rect 11112 53700 11118 53712
rect 13814 53700 13820 53712
rect 11112 53672 13820 53700
rect 11112 53660 11118 53672
rect 13814 53660 13820 53672
rect 13872 53660 13878 53712
rect 17310 53660 17316 53712
rect 17368 53700 17374 53712
rect 19518 53700 19524 53712
rect 17368 53672 19524 53700
rect 17368 53660 17374 53672
rect 19518 53660 19524 53672
rect 19576 53660 19582 53712
rect 538122 53184 538128 53236
rect 538180 53224 538186 53236
rect 551462 53224 551468 53236
rect 538180 53196 551468 53224
rect 538180 53184 538186 53196
rect 551462 53184 551468 53196
rect 551520 53184 551526 53236
rect 8662 53116 8668 53168
rect 8720 53156 8726 53168
rect 20438 53156 20444 53168
rect 8720 53128 20444 53156
rect 8720 53116 8726 53128
rect 20438 53116 20444 53128
rect 20496 53116 20502 53168
rect 7742 53048 7748 53100
rect 7800 53088 7806 53100
rect 20622 53088 20628 53100
rect 7800 53060 20628 53088
rect 7800 53048 7806 53060
rect 20622 53048 20628 53060
rect 20680 53048 20686 53100
rect 540606 53048 540612 53100
rect 540664 53088 540670 53100
rect 554774 53088 554780 53100
rect 540664 53060 554780 53088
rect 540664 53048 540670 53060
rect 554774 53048 554780 53060
rect 554832 53048 554838 53100
rect 13262 52436 13268 52488
rect 13320 52476 13326 52488
rect 13320 52448 16574 52476
rect 13320 52436 13326 52448
rect 10870 52368 10876 52420
rect 10928 52408 10934 52420
rect 12434 52408 12440 52420
rect 10928 52380 12440 52408
rect 10928 52368 10934 52380
rect 12434 52368 12440 52380
rect 12492 52368 12498 52420
rect 16546 52408 16574 52448
rect 19242 52408 19248 52420
rect 16546 52380 19248 52408
rect 19242 52368 19248 52380
rect 19300 52368 19306 52420
rect 19334 52368 19340 52420
rect 19392 52408 19398 52420
rect 20806 52408 20812 52420
rect 19392 52380 20812 52408
rect 19392 52368 19398 52380
rect 20806 52368 20812 52380
rect 20864 52368 20870 52420
rect 18046 52300 18052 52352
rect 18104 52340 18110 52352
rect 20898 52340 20904 52352
rect 18104 52312 20904 52340
rect 18104 52300 18110 52312
rect 20898 52300 20904 52312
rect 20956 52300 20962 52352
rect 15194 52096 15200 52148
rect 15252 52136 15258 52148
rect 20530 52136 20536 52148
rect 15252 52108 20536 52136
rect 15252 52096 15258 52108
rect 20530 52096 20536 52108
rect 20588 52096 20594 52148
rect 3418 52028 3424 52080
rect 3476 52068 3482 52080
rect 460198 52068 460204 52080
rect 3476 52040 460204 52068
rect 3476 52028 3482 52040
rect 460198 52028 460204 52040
rect 460256 52028 460262 52080
rect 3510 51960 3516 52012
rect 3568 52000 3574 52012
rect 455230 52000 455236 52012
rect 3568 51972 455236 52000
rect 3568 51960 3574 51972
rect 455230 51960 455236 51972
rect 455288 51960 455294 52012
rect 16574 51892 16580 51944
rect 16632 51932 16638 51944
rect 382090 51932 382096 51944
rect 16632 51904 382096 51932
rect 16632 51892 16638 51904
rect 382090 51892 382096 51904
rect 382148 51892 382154 51944
rect 18690 51824 18696 51876
rect 18748 51864 18754 51876
rect 383286 51864 383292 51876
rect 18748 51836 383292 51864
rect 18748 51824 18754 51836
rect 383286 51824 383292 51836
rect 383344 51824 383350 51876
rect 18874 51756 18880 51808
rect 18932 51796 18938 51808
rect 383378 51796 383384 51808
rect 18932 51768 383384 51796
rect 18932 51756 18938 51768
rect 383378 51756 383384 51768
rect 383436 51756 383442 51808
rect 15562 51688 15568 51740
rect 15620 51728 15626 51740
rect 20622 51728 20628 51740
rect 15620 51700 20628 51728
rect 15620 51688 15626 51700
rect 20622 51688 20628 51700
rect 20680 51688 20686 51740
rect 20714 51688 20720 51740
rect 20772 51728 20778 51740
rect 383562 51728 383568 51740
rect 20772 51700 383568 51728
rect 20772 51688 20778 51700
rect 383562 51688 383568 51700
rect 383620 51688 383626 51740
rect 18322 51620 18328 51672
rect 18380 51660 18386 51672
rect 380710 51660 380716 51672
rect 18380 51632 380716 51660
rect 18380 51620 18386 51632
rect 380710 51620 380716 51632
rect 380768 51620 380774 51672
rect 19518 51552 19524 51604
rect 19576 51592 19582 51604
rect 381446 51592 381452 51604
rect 19576 51564 381452 51592
rect 19576 51552 19582 51564
rect 381446 51552 381452 51564
rect 381504 51552 381510 51604
rect 382366 51552 382372 51604
rect 382424 51592 382430 51604
rect 384758 51592 384764 51604
rect 382424 51564 384764 51592
rect 382424 51552 382430 51564
rect 384758 51552 384764 51564
rect 384816 51552 384822 51604
rect 20438 51484 20444 51536
rect 20496 51524 20502 51536
rect 20990 51524 20996 51536
rect 20496 51496 20996 51524
rect 20496 51484 20502 51496
rect 20990 51484 20996 51496
rect 21048 51484 21054 51536
rect 378778 51484 378784 51536
rect 378836 51524 378842 51536
rect 384666 51524 384672 51536
rect 378836 51496 384672 51524
rect 378836 51484 378842 51496
rect 384666 51484 384672 51496
rect 384724 51484 384730 51536
rect 382274 51416 382280 51468
rect 382332 51456 382338 51468
rect 386046 51456 386052 51468
rect 382332 51428 386052 51456
rect 382332 51416 382338 51428
rect 386046 51416 386052 51428
rect 386104 51416 386110 51468
rect 378686 51348 378692 51400
rect 378744 51388 378750 51400
rect 386230 51388 386236 51400
rect 378744 51360 386236 51388
rect 378744 51348 378750 51360
rect 386230 51348 386236 51360
rect 386288 51348 386294 51400
rect 377950 51280 377956 51332
rect 378008 51320 378014 51332
rect 382826 51320 382832 51332
rect 378008 51292 382832 51320
rect 378008 51280 378014 51292
rect 382826 51280 382832 51292
rect 382884 51280 382890 51332
rect 378870 51212 378876 51264
rect 378928 51252 378934 51264
rect 386138 51252 386144 51264
rect 378928 51224 386144 51252
rect 378928 51212 378934 51224
rect 386138 51212 386144 51224
rect 386196 51212 386202 51264
rect 21358 51008 21364 51060
rect 21416 51048 21422 51060
rect 455138 51048 455144 51060
rect 21416 51020 455144 51048
rect 21416 51008 21422 51020
rect 455138 51008 455144 51020
rect 455196 51008 455202 51060
rect 8294 50940 8300 50992
rect 8352 50980 8358 50992
rect 377950 50980 377956 50992
rect 8352 50952 377956 50980
rect 8352 50940 8358 50952
rect 377950 50940 377956 50952
rect 378008 50940 378014 50992
rect 17954 50872 17960 50924
rect 18012 50912 18018 50924
rect 382182 50912 382188 50924
rect 18012 50884 382188 50912
rect 18012 50872 18018 50884
rect 382182 50872 382188 50884
rect 382240 50872 382246 50924
rect 20622 50804 20628 50856
rect 20680 50844 20686 50856
rect 383470 50844 383476 50856
rect 20680 50816 383476 50844
rect 20680 50804 20686 50816
rect 383470 50804 383476 50816
rect 383528 50804 383534 50856
rect 19242 50736 19248 50788
rect 19300 50776 19306 50788
rect 378778 50776 378784 50788
rect 19300 50748 378784 50776
rect 19300 50736 19306 50748
rect 378778 50736 378784 50748
rect 378836 50736 378842 50788
rect 20806 50668 20812 50720
rect 20864 50708 20870 50720
rect 380618 50708 380624 50720
rect 20864 50680 380624 50708
rect 20864 50668 20870 50680
rect 380618 50668 380624 50680
rect 380676 50668 380682 50720
rect 20898 50600 20904 50652
rect 20956 50640 20962 50652
rect 380526 50640 380532 50652
rect 20956 50612 380532 50640
rect 20956 50600 20962 50612
rect 380526 50600 380532 50612
rect 380584 50600 380590 50652
rect 65518 50532 65524 50584
rect 65576 50572 65582 50584
rect 401318 50572 401324 50584
rect 65576 50544 401324 50572
rect 65576 50532 65582 50544
rect 401318 50532 401324 50544
rect 401376 50532 401382 50584
rect 20530 50464 20536 50516
rect 20588 50504 20594 50516
rect 33134 50504 33140 50516
rect 20588 50476 33140 50504
rect 20588 50464 20594 50476
rect 33134 50464 33140 50476
rect 33192 50464 33198 50516
rect 62022 50464 62028 50516
rect 62080 50504 62086 50516
rect 403986 50504 403992 50516
rect 62080 50476 403992 50504
rect 62080 50464 62086 50476
rect 403986 50464 403992 50476
rect 404044 50464 404050 50516
rect 20990 50396 20996 50448
rect 21048 50436 21054 50448
rect 42794 50436 42800 50448
rect 21048 50408 42800 50436
rect 21048 50396 21054 50408
rect 42794 50396 42800 50408
rect 42852 50396 42858 50448
rect 58434 50396 58440 50448
rect 58492 50436 58498 50448
rect 404078 50436 404084 50448
rect 58492 50408 404084 50436
rect 58492 50396 58498 50408
rect 404078 50396 404084 50408
rect 404136 50396 404142 50448
rect 13814 50328 13820 50380
rect 13872 50368 13878 50380
rect 44174 50368 44180 50380
rect 13872 50340 44180 50368
rect 13872 50328 13878 50340
rect 44174 50328 44180 50340
rect 44232 50328 44238 50380
rect 54938 50328 54944 50380
rect 54996 50368 55002 50380
rect 403802 50368 403808 50380
rect 54996 50340 403808 50368
rect 54996 50328 55002 50340
rect 403802 50328 403808 50340
rect 403860 50328 403866 50380
rect 70302 50260 70308 50312
rect 70360 50300 70366 50312
rect 387518 50300 387524 50312
rect 70360 50272 387524 50300
rect 70360 50260 70366 50272
rect 387518 50260 387524 50272
rect 387576 50260 387582 50312
rect 93946 50192 93952 50244
rect 94004 50232 94010 50244
rect 395798 50232 395804 50244
rect 94004 50204 395804 50232
rect 94004 50192 94010 50204
rect 395798 50192 395804 50204
rect 395856 50192 395862 50244
rect 115198 50124 115204 50176
rect 115256 50164 115262 50176
rect 395706 50164 395712 50176
rect 115256 50136 395712 50164
rect 115256 50124 115262 50136
rect 395706 50124 395712 50136
rect 395764 50124 395770 50176
rect 12434 49648 12440 49700
rect 12492 49688 12498 49700
rect 378686 49688 378692 49700
rect 12492 49660 378692 49688
rect 12492 49648 12498 49660
rect 378686 49648 378692 49660
rect 378744 49648 378750 49700
rect 33134 49580 33140 49632
rect 33192 49620 33198 49632
rect 382274 49620 382280 49632
rect 33192 49592 382280 49620
rect 33192 49580 33198 49592
rect 382274 49580 382280 49592
rect 382332 49580 382338 49632
rect 44174 49512 44180 49564
rect 44232 49552 44238 49564
rect 382366 49552 382372 49564
rect 44232 49524 382372 49552
rect 44232 49512 44238 49524
rect 382366 49512 382372 49524
rect 382424 49512 382430 49564
rect 42794 49444 42800 49496
rect 42852 49484 42858 49496
rect 378870 49484 378876 49496
rect 42852 49456 378876 49484
rect 42852 49444 42858 49456
rect 378870 49444 378876 49456
rect 378928 49444 378934 49496
rect 101030 48220 101036 48272
rect 101088 48260 101094 48272
rect 395614 48260 395620 48272
rect 101088 48232 395620 48260
rect 101088 48220 101094 48232
rect 395614 48220 395620 48232
rect 395672 48220 395678 48272
rect 87966 48152 87972 48204
rect 88024 48192 88030 48204
rect 384574 48192 384580 48204
rect 88024 48164 384580 48192
rect 88024 48152 88030 48164
rect 384574 48152 384580 48164
rect 384632 48152 384638 48204
rect 97442 48084 97448 48136
rect 97500 48124 97506 48136
rect 395522 48124 395528 48136
rect 97500 48096 395528 48124
rect 97500 48084 97506 48096
rect 395522 48084 395528 48096
rect 395580 48084 395586 48136
rect 90358 48016 90364 48068
rect 90416 48056 90422 48068
rect 398282 48056 398288 48068
rect 90416 48028 398288 48056
rect 90416 48016 90422 48028
rect 398282 48016 398288 48028
rect 398340 48016 398346 48068
rect 86862 47948 86868 48000
rect 86920 47988 86926 48000
rect 398374 47988 398380 48000
rect 86920 47960 398380 47988
rect 86920 47948 86926 47960
rect 398374 47948 398380 47960
rect 398432 47948 398438 48000
rect 83274 47880 83280 47932
rect 83332 47920 83338 47932
rect 398098 47920 398104 47932
rect 83332 47892 398104 47920
rect 83332 47880 83338 47892
rect 398098 47880 398104 47892
rect 398156 47880 398162 47932
rect 79686 47812 79692 47864
rect 79744 47852 79750 47864
rect 401226 47852 401232 47864
rect 79744 47824 401232 47852
rect 79744 47812 79750 47824
rect 401226 47812 401232 47824
rect 401284 47812 401290 47864
rect 76190 47744 76196 47796
rect 76248 47784 76254 47796
rect 401134 47784 401140 47796
rect 76248 47756 401140 47784
rect 76248 47744 76254 47756
rect 401134 47744 401140 47756
rect 401192 47744 401198 47796
rect 72602 47676 72608 47728
rect 72660 47716 72666 47728
rect 401042 47716 401048 47728
rect 72660 47688 401048 47716
rect 72660 47676 72666 47688
rect 401042 47676 401048 47688
rect 401100 47676 401106 47728
rect 69106 47608 69112 47660
rect 69164 47648 69170 47660
rect 400950 47648 400956 47660
rect 69164 47620 400956 47648
rect 69164 47608 69170 47620
rect 400950 47608 400956 47620
rect 401008 47608 401014 47660
rect 12342 47540 12348 47592
rect 12400 47580 12406 47592
rect 398190 47580 398196 47592
rect 12400 47552 398196 47580
rect 12400 47540 12406 47552
rect 398190 47540 398196 47552
rect 398248 47540 398254 47592
rect 104526 47472 104532 47524
rect 104584 47512 104590 47524
rect 395430 47512 395436 47524
rect 104584 47484 395436 47512
rect 104584 47472 104590 47484
rect 395430 47472 395436 47484
rect 395488 47472 395494 47524
rect 110506 47404 110512 47456
rect 110564 47444 110570 47456
rect 399846 47444 399852 47456
rect 110564 47416 399852 47444
rect 110564 47404 110570 47416
rect 399846 47404 399852 47416
rect 399904 47404 399910 47456
rect 569218 46860 569224 46912
rect 569276 46900 569282 46912
rect 580166 46900 580172 46912
rect 569276 46872 580172 46900
rect 569276 46860 569282 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 399754 45540 399760 45552
rect 3476 45512 399760 45540
rect 3476 45500 3482 45512
rect 399754 45500 399760 45512
rect 399812 45500 399818 45552
rect 66714 45432 66720 45484
rect 66772 45472 66778 45484
rect 387426 45472 387432 45484
rect 66772 45444 387432 45472
rect 66772 45432 66778 45444
rect 387426 45432 387432 45444
rect 387484 45432 387490 45484
rect 122282 45364 122288 45416
rect 122340 45404 122346 45416
rect 454954 45404 454960 45416
rect 122340 45376 454960 45404
rect 122340 45364 122346 45376
rect 454954 45364 454960 45376
rect 455012 45364 455018 45416
rect 118786 45296 118792 45348
rect 118844 45336 118850 45348
rect 454862 45336 454868 45348
rect 118844 45308 454868 45336
rect 118844 45296 118850 45308
rect 454862 45296 454868 45308
rect 454920 45296 454926 45348
rect 50154 45228 50160 45280
rect 50212 45268 50218 45280
rect 388622 45268 388628 45280
rect 50212 45240 388628 45268
rect 50212 45228 50218 45240
rect 388622 45228 388628 45240
rect 388680 45228 388686 45280
rect 48958 45160 48964 45212
rect 49016 45200 49022 45212
rect 390278 45200 390284 45212
rect 49016 45172 390284 45200
rect 49016 45160 49022 45172
rect 390278 45160 390284 45172
rect 390336 45160 390342 45212
rect 44266 45092 44272 45144
rect 44324 45132 44330 45144
rect 390186 45132 390192 45144
rect 44324 45104 390192 45132
rect 44324 45092 44330 45104
rect 390186 45092 390192 45104
rect 390244 45092 390250 45144
rect 40678 45024 40684 45076
rect 40736 45064 40742 45076
rect 392946 45064 392952 45076
rect 40736 45036 392952 45064
rect 40736 45024 40742 45036
rect 392946 45024 392952 45036
rect 393004 45024 393010 45076
rect 37182 44956 37188 45008
rect 37240 44996 37246 45008
rect 392762 44996 392768 45008
rect 37240 44968 392768 44996
rect 37240 44956 37246 44968
rect 392762 44956 392768 44968
rect 392820 44956 392826 45008
rect 33594 44888 33600 44940
rect 33652 44928 33658 44940
rect 393038 44928 393044 44940
rect 33652 44900 393044 44928
rect 33652 44888 33658 44900
rect 393038 44888 393044 44900
rect 393096 44888 393102 44940
rect 26510 44820 26516 44872
rect 26568 44860 26574 44872
rect 392854 44860 392860 44872
rect 26568 44832 392860 44860
rect 26568 44820 26574 44832
rect 392854 44820 392860 44832
rect 392912 44820 392918 44872
rect 108114 44752 108120 44804
rect 108172 44792 108178 44804
rect 407942 44792 407948 44804
rect 108172 44764 407948 44792
rect 108172 44752 108178 44764
rect 407942 44752 407948 44764
rect 408000 44752 408006 44804
rect 111610 44684 111616 44736
rect 111668 44724 111674 44736
rect 410518 44724 410524 44736
rect 111668 44696 410524 44724
rect 111668 44684 111674 44696
rect 410518 44684 410524 44696
rect 410576 44684 410582 44736
rect 91554 42712 91560 42764
rect 91612 42752 91618 42764
rect 384390 42752 384396 42764
rect 91612 42724 384396 42752
rect 91612 42712 91618 42724
rect 384390 42712 384396 42724
rect 384448 42712 384454 42764
rect 469858 42712 469864 42764
rect 469916 42752 469922 42764
rect 536834 42752 536840 42764
rect 469916 42724 536840 42752
rect 469916 42712 469922 42724
rect 536834 42712 536840 42724
rect 536892 42712 536898 42764
rect 98638 42644 98644 42696
rect 98696 42684 98702 42696
rect 394326 42684 394332 42696
rect 98696 42656 394332 42684
rect 98696 42644 98702 42656
rect 394326 42644 394332 42656
rect 394384 42644 394390 42696
rect 84470 42576 84476 42628
rect 84528 42616 84534 42628
rect 384482 42616 384488 42628
rect 84528 42588 384488 42616
rect 84528 42576 84534 42588
rect 384482 42576 384488 42588
rect 384540 42576 384546 42628
rect 80882 42508 80888 42560
rect 80940 42548 80946 42560
rect 387242 42548 387248 42560
rect 80940 42520 387248 42548
rect 80940 42508 80946 42520
rect 387242 42508 387248 42520
rect 387300 42508 387306 42560
rect 77386 42440 77392 42492
rect 77444 42480 77450 42492
rect 387150 42480 387156 42492
rect 77444 42452 387156 42480
rect 77444 42440 77450 42452
rect 387150 42440 387156 42452
rect 387208 42440 387214 42492
rect 73798 42372 73804 42424
rect 73856 42412 73862 42424
rect 387058 42412 387064 42424
rect 73856 42384 387064 42412
rect 73856 42372 73862 42384
rect 387058 42372 387064 42384
rect 387116 42372 387122 42424
rect 63218 42304 63224 42356
rect 63276 42344 63282 42356
rect 387334 42344 387340 42356
rect 63276 42316 387340 42344
rect 63276 42304 63282 42316
rect 387334 42304 387340 42316
rect 387392 42304 387398 42356
rect 59630 42236 59636 42288
rect 59688 42276 59694 42288
rect 389910 42276 389916 42288
rect 59688 42248 389916 42276
rect 59688 42236 59694 42248
rect 389910 42236 389916 42248
rect 389968 42236 389974 42288
rect 56042 42168 56048 42220
rect 56100 42208 56106 42220
rect 390002 42208 390008 42220
rect 56100 42180 390008 42208
rect 56100 42168 56106 42180
rect 390002 42168 390008 42180
rect 390060 42168 390066 42220
rect 52546 42100 52552 42152
rect 52604 42140 52610 42152
rect 390094 42140 390100 42152
rect 52604 42112 390100 42140
rect 52604 42100 52610 42112
rect 390094 42100 390100 42112
rect 390152 42100 390158 42152
rect 41874 42032 41880 42084
rect 41932 42072 41938 42084
rect 385954 42072 385960 42084
rect 41932 42044 385960 42072
rect 41932 42032 41938 42044
rect 385954 42032 385960 42044
rect 386012 42032 386018 42084
rect 95142 41964 95148 42016
rect 95200 42004 95206 42016
rect 381998 42004 382004 42016
rect 95200 41976 382004 42004
rect 95200 41964 95206 41976
rect 381998 41964 382004 41976
rect 382056 41964 382062 42016
rect 102226 41896 102232 41948
rect 102284 41936 102290 41948
rect 381906 41936 381912 41948
rect 102284 41908 381912 41936
rect 102284 41896 102290 41908
rect 381906 41896 381912 41908
rect 381964 41896 381970 41948
rect 123478 39992 123484 40044
rect 123536 40032 123542 40044
rect 397086 40032 397092 40044
rect 123536 40004 397092 40032
rect 123536 39992 123542 40004
rect 397086 39992 397092 40004
rect 397144 39992 397150 40044
rect 116394 39924 116400 39976
rect 116452 39964 116458 39976
rect 393958 39964 393964 39976
rect 116452 39936 393964 39964
rect 116452 39924 116458 39936
rect 393958 39924 393964 39936
rect 394016 39924 394022 39976
rect 119890 39856 119896 39908
rect 119948 39896 119954 39908
rect 399478 39896 399484 39908
rect 119948 39868 399484 39896
rect 119948 39856 119954 39868
rect 399478 39856 399484 39868
rect 399536 39856 399542 39908
rect 105722 39788 105728 39840
rect 105780 39828 105786 39840
rect 391474 39828 391480 39840
rect 105780 39800 391480 39828
rect 105780 39788 105786 39800
rect 391474 39788 391480 39800
rect 391532 39788 391538 39840
rect 45462 39720 45468 39772
rect 45520 39760 45526 39772
rect 388530 39760 388536 39772
rect 45520 39732 388536 39760
rect 45520 39720 45526 39732
rect 388530 39720 388536 39732
rect 388588 39720 388594 39772
rect 38378 39652 38384 39704
rect 38436 39692 38442 39704
rect 385770 39692 385776 39704
rect 38436 39664 385776 39692
rect 38436 39652 38442 39664
rect 385770 39652 385776 39664
rect 385828 39652 385834 39704
rect 34790 39584 34796 39636
rect 34848 39624 34854 39636
rect 385678 39624 385684 39636
rect 34848 39596 385684 39624
rect 34848 39584 34854 39596
rect 385678 39584 385684 39596
rect 385736 39584 385742 39636
rect 31294 39516 31300 39568
rect 31352 39556 31358 39568
rect 385862 39556 385868 39568
rect 31352 39528 385868 39556
rect 31352 39516 31358 39528
rect 385862 39516 385868 39528
rect 385920 39516 385926 39568
rect 27706 39448 27712 39500
rect 27764 39488 27770 39500
rect 383102 39488 383108 39500
rect 27764 39460 383108 39488
rect 27764 39448 27770 39460
rect 383102 39448 383108 39460
rect 383160 39448 383166 39500
rect 23014 39380 23020 39432
rect 23072 39420 23078 39432
rect 383194 39420 383200 39432
rect 23072 39392 383200 39420
rect 23072 39380 23078 39392
rect 383194 39380 383200 39392
rect 383252 39380 383258 39432
rect 18230 39312 18236 39364
rect 18288 39352 18294 39364
rect 382918 39352 382924 39364
rect 18288 39324 382924 39352
rect 18288 39312 18294 39324
rect 382918 39312 382924 39324
rect 382976 39312 382982 39364
rect 109310 39244 109316 39296
rect 109368 39284 109374 39296
rect 381814 39284 381820 39296
rect 109368 39256 381820 39284
rect 109368 39244 109374 39256
rect 381814 39244 381820 39256
rect 381872 39244 381878 39296
rect 112806 39176 112812 39228
rect 112864 39216 112870 39228
rect 383010 39216 383016 39228
rect 112864 39188 383016 39216
rect 112864 39176 112870 39188
rect 383010 39176 383016 39188
rect 383068 39176 383074 39228
rect 96246 37204 96252 37256
rect 96304 37244 96310 37256
rect 399662 37244 399668 37256
rect 96304 37216 399668 37244
rect 96304 37204 96310 37216
rect 399662 37204 399668 37216
rect 399720 37204 399726 37256
rect 92750 37136 92756 37188
rect 92808 37176 92814 37188
rect 396902 37176 396908 37188
rect 92808 37148 396908 37176
rect 92808 37136 92814 37148
rect 396902 37136 396908 37148
rect 396960 37136 396966 37188
rect 89162 37068 89168 37120
rect 89220 37108 89226 37120
rect 396994 37108 397000 37120
rect 89220 37080 397000 37108
rect 89220 37068 89226 37080
rect 396994 37068 397000 37080
rect 397052 37068 397058 37120
rect 85666 37000 85672 37052
rect 85724 37040 85730 37052
rect 396810 37040 396816 37052
rect 85724 37012 396816 37040
rect 85724 37000 85730 37012
rect 396810 37000 396816 37012
rect 396868 37000 396874 37052
rect 82078 36932 82084 36984
rect 82136 36972 82142 36984
rect 394142 36972 394148 36984
rect 82136 36944 394148 36972
rect 82136 36932 82142 36944
rect 394142 36932 394148 36944
rect 394200 36932 394206 36984
rect 74994 36864 75000 36916
rect 75052 36904 75058 36916
rect 394234 36904 394240 36916
rect 75052 36876 394240 36904
rect 75052 36864 75058 36876
rect 394234 36864 394240 36876
rect 394292 36864 394298 36916
rect 71498 36796 71504 36848
rect 71556 36836 71562 36848
rect 394050 36836 394056 36848
rect 71556 36808 394056 36836
rect 71556 36796 71562 36808
rect 394050 36796 394056 36808
rect 394108 36796 394114 36848
rect 64322 36728 64328 36780
rect 64380 36768 64386 36780
rect 391382 36768 391388 36780
rect 64380 36740 391388 36768
rect 64380 36728 64386 36740
rect 391382 36728 391388 36740
rect 391440 36728 391446 36780
rect 57238 36660 57244 36712
rect 57296 36700 57302 36712
rect 391198 36700 391204 36712
rect 57296 36672 391204 36700
rect 57296 36660 57302 36672
rect 391198 36660 391204 36672
rect 391256 36660 391262 36712
rect 53742 36592 53748 36644
rect 53800 36632 53806 36644
rect 391290 36632 391296 36644
rect 53800 36604 391296 36632
rect 53800 36592 53806 36604
rect 391290 36592 391296 36604
rect 391348 36592 391354 36644
rect 60826 36524 60832 36576
rect 60884 36564 60890 36576
rect 456242 36564 456248 36576
rect 60884 36536 456248 36564
rect 60884 36524 60890 36536
rect 456242 36524 456248 36536
rect 456300 36524 456306 36576
rect 103330 36456 103336 36508
rect 103388 36496 103394 36508
rect 399570 36496 399576 36508
rect 103388 36468 399576 36496
rect 103388 36456 103394 36468
rect 399570 36456 399576 36468
rect 399628 36456 399634 36508
rect 124674 34076 124680 34128
rect 124732 34116 124738 34128
rect 405090 34116 405096 34128
rect 124732 34088 405096 34116
rect 124732 34076 124738 34088
rect 405090 34076 405096 34088
rect 405148 34076 405154 34128
rect 121086 34008 121092 34060
rect 121144 34048 121150 34060
rect 402330 34048 402336 34060
rect 121144 34020 402336 34048
rect 121144 34008 121150 34020
rect 402330 34008 402336 34020
rect 402388 34008 402394 34060
rect 117590 33940 117596 33992
rect 117648 33980 117654 33992
rect 402238 33980 402244 33992
rect 117648 33952 402244 33980
rect 117648 33940 117654 33952
rect 402238 33940 402244 33952
rect 402296 33940 402302 33992
rect 39574 33872 39580 33924
rect 39632 33912 39638 33924
rect 405182 33912 405188 33924
rect 39632 33884 405188 33912
rect 39632 33872 39638 33884
rect 405182 33872 405188 33884
rect 405240 33872 405246 33924
rect 24210 33804 24216 33856
rect 24268 33844 24274 33856
rect 404998 33844 405004 33856
rect 24268 33816 405004 33844
rect 24268 33804 24274 33816
rect 404998 33804 405004 33816
rect 405056 33804 405062 33856
rect 19426 33736 19432 33788
rect 19484 33776 19490 33788
rect 402514 33776 402520 33788
rect 19484 33748 402520 33776
rect 19484 33736 19490 33748
rect 402514 33736 402520 33748
rect 402572 33736 402578 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 400858 33096 400864 33108
rect 3568 33068 400864 33096
rect 3568 33056 3574 33068
rect 400858 33056 400864 33068
rect 400916 33056 400922 33108
rect 570598 33056 570604 33108
rect 570656 33096 570662 33108
rect 580166 33096 580172 33108
rect 570656 33068 580172 33096
rect 570656 33056 570662 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 403618 20652 403624 20664
rect 3476 20624 403624 20652
rect 3476 20612 3482 20624
rect 403618 20612 403624 20624
rect 403676 20612 403682 20664
rect 571978 20612 571984 20664
rect 572036 20652 572042 20664
rect 579982 20652 579988 20664
rect 572036 20624 579988 20652
rect 572036 20612 572042 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 396718 6848 396724 6860
rect 3476 6820 396724 6848
rect 3476 6808 3482 6820
rect 396718 6808 396724 6820
rect 396776 6808 396782 6860
rect 566458 6808 566464 6860
rect 566516 6848 566522 6860
rect 580166 6848 580172 6860
rect 566516 6820 580172 6848
rect 566516 6808 566522 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 67910 4088 67916 4140
rect 67968 4128 67974 4140
rect 380342 4128 380348 4140
rect 67968 4100 380348 4128
rect 67968 4088 67974 4100
rect 380342 4088 380348 4100
rect 380400 4088 380406 4140
rect 32398 4020 32404 4072
rect 32456 4060 32462 4072
rect 381538 4060 381544 4072
rect 32456 4032 381544 4060
rect 32456 4020 32462 4032
rect 381538 4020 381544 4032
rect 381596 4020 381602 4072
rect 99834 3952 99840 4004
rect 99892 3992 99898 4004
rect 454678 3992 454684 4004
rect 99892 3964 454684 3992
rect 99892 3952 99898 3964
rect 454678 3952 454684 3964
rect 454736 3952 454742 4004
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 380158 3924 380164 3936
rect 14792 3896 380164 3924
rect 14792 3884 14798 3896
rect 380158 3884 380164 3896
rect 380216 3884 380222 3936
rect 13538 3816 13544 3868
rect 13596 3856 13602 3868
rect 384298 3856 384304 3868
rect 13596 3828 384304 3856
rect 13596 3816 13602 3828
rect 384298 3816 384304 3828
rect 384356 3816 384362 3868
rect 21818 3748 21824 3800
rect 21876 3788 21882 3800
rect 392670 3788 392676 3800
rect 21876 3760 392676 3788
rect 21876 3748 21882 3760
rect 392670 3748 392676 3760
rect 392728 3748 392734 3800
rect 17034 3680 17040 3732
rect 17092 3720 17098 3732
rect 395338 3720 395344 3732
rect 17092 3692 395344 3720
rect 17092 3680 17098 3692
rect 395338 3680 395344 3692
rect 395396 3680 395402 3732
rect 28902 3612 28908 3664
rect 28960 3652 28966 3664
rect 407850 3652 407856 3664
rect 28960 3624 407856 3652
rect 28960 3612 28966 3624
rect 407850 3612 407856 3624
rect 407908 3612 407914 3664
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 389818 3584 389824 3596
rect 8812 3556 389824 3584
rect 8812 3544 8818 3556
rect 389818 3544 389824 3556
rect 389876 3544 389882 3596
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 456150 3516 456156 3528
rect 43128 3488 456156 3516
rect 43128 3476 43134 3488
rect 456150 3476 456156 3488
rect 456208 3476 456214 3528
rect 35986 3408 35992 3460
rect 36044 3448 36050 3460
rect 456058 3448 456064 3460
rect 36044 3420 456064 3448
rect 36044 3408 36050 3420
rect 456058 3408 456064 3420
rect 456116 3408 456122 3460
rect 78582 3340 78588 3392
rect 78640 3380 78646 3392
rect 380250 3380 380256 3392
rect 78640 3352 380256 3380
rect 78640 3340 78646 3352
rect 380250 3340 380256 3352
rect 380308 3340 380314 3392
rect 106918 3272 106924 3324
rect 106976 3312 106982 3324
rect 381722 3312 381728 3324
rect 106976 3284 381728 3312
rect 106976 3272 106982 3284
rect 381722 3272 381728 3284
rect 381780 3272 381786 3324
rect 114002 3204 114008 3256
rect 114060 3244 114066 3256
rect 381630 3244 381636 3256
rect 114060 3216 381636 3244
rect 114060 3204 114066 3216
rect 381630 3204 381636 3216
rect 381688 3204 381694 3256
rect 30098 2048 30104 2100
rect 30156 2088 30162 2100
rect 392578 2088 392584 2100
rect 30156 2060 392584 2088
rect 30156 2048 30162 2060
rect 392578 2048 392584 2060
rect 392636 2048 392642 2100
<< via1 >>
rect 397460 700680 397512 700732
rect 418804 700680 418856 700732
rect 444288 700680 444340 700732
rect 478512 700680 478564 700732
rect 364984 700612 365036 700664
rect 446404 700612 446456 700664
rect 332508 700544 332560 700596
rect 445024 700544 445076 700596
rect 218980 700476 219032 700528
rect 416044 700476 416096 700528
rect 444196 700476 444248 700528
rect 494796 700476 494848 700528
rect 235172 700408 235224 700460
rect 446496 700408 446548 700460
rect 170312 700340 170364 700392
rect 449164 700340 449216 700392
rect 137836 700272 137888 700324
rect 445116 700272 445168 700324
rect 527180 700272 527232 700324
rect 543740 700272 543792 700324
rect 3424 683136 3476 683188
rect 446588 683136 446640 683188
rect 570604 683136 570656 683188
rect 579620 683136 579672 683188
rect 448428 679600 448480 679652
rect 462320 679600 462372 679652
rect 3516 670692 3568 670744
rect 446772 670692 446824 670744
rect 573364 670692 573416 670744
rect 580172 670692 580224 670744
rect 348792 670216 348844 670268
rect 446864 670216 446916 670268
rect 283840 670148 283892 670200
rect 445208 670148 445260 670200
rect 154120 670080 154172 670132
rect 446680 670080 446732 670132
rect 89168 670012 89220 670064
rect 413284 670012 413336 670064
rect 72976 669944 73028 669996
rect 418896 669944 418948 669996
rect 267648 668788 267700 668840
rect 445300 668788 445352 668840
rect 23480 668720 23532 668772
rect 380440 668720 380492 668772
rect 20720 668652 20772 668704
rect 378324 668652 378376 668704
rect 20996 668584 21048 668636
rect 378140 668584 378192 668636
rect 21088 668516 21140 668568
rect 380348 668516 380400 668568
rect 20904 668448 20956 668500
rect 380624 668448 380676 668500
rect 18880 668380 18932 668432
rect 378232 668380 378284 668432
rect 20812 668312 20864 668364
rect 381820 668312 381872 668364
rect 19340 668244 19392 668296
rect 381544 668244 381596 668296
rect 18788 668176 18840 668228
rect 380164 668176 380216 668228
rect 17868 668108 17920 668160
rect 381636 668108 381688 668160
rect 7564 668040 7616 668092
rect 381912 668040 381964 668092
rect 3792 667972 3844 668024
rect 447048 667972 447100 668024
rect 3424 667904 3476 667956
rect 446956 667904 447008 667956
rect 378140 667836 378192 667888
rect 380256 667836 380308 667888
rect 19892 667768 19944 667820
rect 23480 667768 23532 667820
rect 378232 667768 378284 667820
rect 381728 667768 381780 667820
rect 19800 667700 19852 667752
rect 20996 667700 21048 667752
rect 378324 667700 378376 667752
rect 380532 667700 380584 667752
rect 18696 667632 18748 667684
rect 21088 667632 21140 667684
rect 21364 667632 21416 667684
rect 420184 667632 420236 667684
rect 3700 667564 3752 667616
rect 418988 667564 419040 667616
rect 18420 666680 18472 666732
rect 20812 666680 20864 666732
rect 17684 666612 17736 666664
rect 19340 666612 19392 666664
rect 20076 666612 20128 666664
rect 20720 666612 20772 666664
rect 19984 666544 20036 666596
rect 20904 666544 20956 666596
rect 16580 665456 16632 665508
rect 19892 665456 19944 665508
rect 13820 665252 13872 665304
rect 17868 665252 17920 665304
rect 10968 665116 11020 665168
rect 17684 665184 17736 665236
rect 18604 664640 18656 664692
rect 19800 664640 19852 664692
rect 11060 663756 11112 663808
rect 16580 663756 16632 663808
rect 15292 663688 15344 663740
rect 18420 663756 18472 663808
rect 17960 662464 18012 662516
rect 20076 662464 20128 662516
rect 8668 662396 8720 662448
rect 10968 662396 11020 662448
rect 13912 662396 13964 662448
rect 18696 662396 18748 662448
rect 14464 661648 14516 661700
rect 18788 661648 18840 661700
rect 11704 660968 11756 661020
rect 15292 661036 15344 661088
rect 15200 660968 15252 661020
rect 18880 661104 18932 661156
rect 18696 661036 18748 661088
rect 19984 661036 20036 661088
rect 382280 661036 382332 661088
rect 403624 661036 403676 661088
rect 5632 660288 5684 660340
rect 7564 660288 7616 660340
rect 5540 659744 5592 659796
rect 8668 659744 8720 659796
rect 9588 659676 9640 659728
rect 13820 659676 13872 659728
rect 8944 658180 8996 658232
rect 11060 658248 11112 658300
rect 14648 657296 14700 657348
rect 15200 657296 15252 657348
rect 10048 656344 10100 656396
rect 13912 656344 13964 656396
rect 7104 656276 7156 656328
rect 9588 656276 9640 656328
rect 460480 655800 460532 655852
rect 460664 655800 460716 655852
rect 3424 655460 3476 655512
rect 5632 655528 5684 655580
rect 15936 655528 15988 655580
rect 17868 655528 17920 655580
rect 4804 654440 4856 654492
rect 5540 654440 5592 654492
rect 8300 652876 8352 652928
rect 14464 652876 14516 652928
rect 5632 652808 5684 652860
rect 8944 652808 8996 652860
rect 5080 652672 5132 652724
rect 7104 652740 7156 652792
rect 9220 652740 9272 652792
rect 11704 652740 11756 652792
rect 17040 652740 17092 652792
rect 18696 652740 18748 652792
rect 3516 651992 3568 652044
rect 10048 651992 10100 652044
rect 12440 651448 12492 651500
rect 14648 651448 14700 651500
rect 13820 651380 13872 651432
rect 15936 651380 15988 651432
rect 382280 651380 382332 651432
rect 396724 651380 396776 651432
rect 5540 650224 5592 650276
rect 9220 650224 9272 650276
rect 3608 649952 3660 650004
rect 5632 650020 5684 650072
rect 4896 649680 4948 649732
rect 8208 649680 8260 649732
rect 8944 648524 8996 648576
rect 12440 648592 12492 648644
rect 15200 648524 15252 648576
rect 18604 648592 18656 648644
rect 11060 646552 11112 646604
rect 13820 646552 13872 646604
rect 13084 645940 13136 645992
rect 17040 645940 17092 645992
rect 12440 645464 12492 645516
rect 15200 645464 15252 645516
rect 460296 643696 460348 643748
rect 460756 643696 460808 643748
rect 4988 643016 5040 643068
rect 8944 643084 8996 643136
rect 8944 640228 8996 640280
rect 11060 640296 11112 640348
rect 9680 637712 9732 637764
rect 12348 637712 12400 637764
rect 6920 636148 6972 636200
rect 9680 636148 9732 636200
rect 10692 632000 10744 632052
rect 13084 632068 13136 632120
rect 7932 631660 7984 631712
rect 8944 631660 8996 631712
rect 3700 630640 3752 630692
rect 6828 630640 6880 630692
rect 577504 630640 577556 630692
rect 580448 630640 580500 630692
rect 382280 629280 382332 629332
rect 395344 629280 395396 629332
rect 5540 628736 5592 628788
rect 7932 628736 7984 628788
rect 4160 626900 4212 626952
rect 5540 626900 5592 626952
rect 8944 625880 8996 625932
rect 10692 625880 10744 625932
rect 382280 619624 382332 619676
rect 399484 619624 399536 619676
rect 3148 619556 3200 619608
rect 20904 619556 20956 619608
rect 7564 617924 7616 617976
rect 8944 617924 8996 617976
rect 571984 616836 572036 616888
rect 580172 616836 580224 616888
rect 457536 610648 457588 610700
rect 457904 610648 457956 610700
rect 382280 608608 382332 608660
rect 393964 608608 394016 608660
rect 460480 602896 460532 602948
rect 460480 602624 460532 602676
rect 6184 601604 6236 601656
rect 7564 601604 7616 601656
rect 460572 600652 460624 600704
rect 461584 600652 461636 600704
rect 457904 600244 457956 600296
rect 462964 600244 463016 600296
rect 457260 600176 457312 600228
rect 463056 600176 463108 600228
rect 457536 599700 457588 599752
rect 464344 599700 464396 599752
rect 457444 599632 457496 599684
rect 467104 599632 467156 599684
rect 518164 599632 518216 599684
rect 543740 599632 543792 599684
rect 460388 599564 460440 599616
rect 503720 599564 503772 599616
rect 515404 599564 515456 599616
rect 580356 599564 580408 599616
rect 457352 598408 457404 598460
rect 468484 598408 468536 598460
rect 457812 598340 457864 598392
rect 471244 598340 471296 598392
rect 459100 598272 459152 598324
rect 502340 598272 502392 598324
rect 460296 598204 460348 598256
rect 495440 598204 495492 598256
rect 496084 598204 496136 598256
rect 540520 598204 540572 598256
rect 382280 597524 382332 597576
rect 406384 597524 406436 597576
rect 457628 596844 457680 596896
rect 467196 596844 467248 596896
rect 459008 596776 459060 596828
rect 496820 596776 496872 596828
rect 457720 595484 457772 595536
rect 468576 595484 468628 595536
rect 460480 595416 460532 595468
rect 500960 595416 501012 595468
rect 458916 592628 458968 592680
rect 494060 592628 494112 592680
rect 459284 591268 459336 591320
rect 503812 591268 503864 591320
rect 459192 589908 459244 589960
rect 499580 589908 499632 589960
rect 3792 587800 3844 587852
rect 6184 587868 6236 587920
rect 382280 587868 382332 587920
rect 392584 587868 392636 587920
rect 3608 578416 3660 578468
rect 5172 578416 5224 578468
rect 382280 576852 382332 576904
rect 419080 576852 419132 576904
rect 518256 576852 518308 576904
rect 579620 576852 579672 576904
rect 381912 573996 381964 574048
rect 384304 573996 384356 574048
rect 381820 572160 381872 572212
rect 383016 572160 383068 572212
rect 3884 565836 3936 565888
rect 5080 565836 5132 565888
rect 382280 565088 382332 565140
rect 407764 565088 407816 565140
rect 515496 563048 515548 563100
rect 580172 563048 580224 563100
rect 383016 559512 383068 559564
rect 387616 559512 387668 559564
rect 384304 556588 384356 556640
rect 385040 556588 385092 556640
rect 382280 556180 382332 556232
rect 391204 556180 391256 556232
rect 385040 554344 385092 554396
rect 387156 554344 387208 554396
rect 3792 553392 3844 553444
rect 4988 553392 5040 553444
rect 380624 553392 380676 553444
rect 383016 553324 383068 553376
rect 387616 552644 387668 552696
rect 389916 552644 389968 552696
rect 382280 545096 382332 545148
rect 389824 545096 389876 545148
rect 389916 543668 389968 543720
rect 394056 543668 394108 543720
rect 380532 543192 380584 543244
rect 381820 543192 381872 543244
rect 381728 537480 381780 537532
rect 389180 537480 389232 537532
rect 460664 537480 460716 537532
rect 498200 537480 498252 537532
rect 518348 536800 518400 536852
rect 580172 536800 580224 536852
rect 383016 536596 383068 536648
rect 384120 536596 384172 536648
rect 389180 535780 389232 535832
rect 391940 535780 391992 535832
rect 382280 534080 382332 534132
rect 387064 534080 387116 534132
rect 391940 534012 391992 534064
rect 394884 534012 394936 534064
rect 381820 533536 381872 533588
rect 383016 533536 383068 533588
rect 384120 532720 384172 532772
rect 389180 532652 389232 532704
rect 394056 531224 394108 531276
rect 396816 531224 396868 531276
rect 389180 529932 389232 529984
rect 394056 529864 394108 529916
rect 394884 529864 394936 529916
rect 397092 529864 397144 529916
rect 381636 529524 381688 529576
rect 385776 529524 385828 529576
rect 3516 525784 3568 525836
rect 4896 525784 4948 525836
rect 382280 524424 382332 524476
rect 385684 524424 385736 524476
rect 458088 522248 458140 522300
rect 467288 522248 467340 522300
rect 397460 521568 397512 521620
rect 402244 521568 402296 521620
rect 482928 520888 482980 520940
rect 531320 520888 531372 520940
rect 461676 520276 461728 520328
rect 488632 520276 488684 520328
rect 460756 519528 460808 519580
rect 493048 519528 493100 519580
rect 457996 518168 458048 518220
rect 469864 518168 469916 518220
rect 387156 518032 387208 518084
rect 391940 518032 391992 518084
rect 394056 517964 394108 518016
rect 394700 517964 394752 518016
rect 450360 517556 450412 517608
rect 491852 517556 491904 517608
rect 450544 517488 450596 517540
rect 514760 517488 514812 517540
rect 489184 517420 489236 517472
rect 450176 516808 450228 516860
rect 480444 516808 480496 516860
rect 450636 516740 450688 516792
rect 494152 516740 494204 516792
rect 383016 516060 383068 516112
rect 384948 516060 385000 516112
rect 391940 516060 391992 516112
rect 395068 516060 395120 516112
rect 494796 515924 494848 515976
rect 498292 515924 498344 515976
rect 396816 514768 396868 514820
rect 400220 514700 400272 514752
rect 514760 514020 514812 514072
rect 547880 514020 547932 514072
rect 382280 513544 382332 513596
rect 384304 513544 384356 513596
rect 395068 513340 395120 513392
rect 399576 513340 399628 513392
rect 506572 512660 506624 512712
rect 543740 512660 543792 512712
rect 494152 512592 494204 512644
rect 538220 512592 538272 512644
rect 519544 510620 519596 510672
rect 580172 510620 580224 510672
rect 385776 510552 385828 510604
rect 387156 510552 387208 510604
rect 394700 510552 394752 510604
rect 397184 510552 397236 510604
rect 400220 510552 400272 510604
rect 402152 510552 402204 510604
rect 385040 510484 385092 510536
rect 388076 510484 388128 510536
rect 498292 509872 498344 509924
rect 540980 509872 541032 509924
rect 397184 509192 397236 509244
rect 403992 509192 404044 509244
rect 492128 508512 492180 508564
rect 534080 508512 534132 508564
rect 3700 507832 3752 507884
rect 4804 507832 4856 507884
rect 494152 505112 494204 505164
rect 531320 505112 531372 505164
rect 388076 504636 388128 504688
rect 389180 504636 389232 504688
rect 402152 503684 402204 503736
rect 404728 503616 404780 503668
rect 382280 502324 382332 502376
rect 410524 502324 410576 502376
rect 389180 502256 389232 502308
rect 392676 502256 392728 502308
rect 403992 502256 404044 502308
rect 405004 502256 405056 502308
rect 387156 500896 387208 500948
rect 389916 500896 389968 500948
rect 404728 500896 404780 500948
rect 406568 500896 406620 500948
rect 450544 500896 450596 500948
rect 472624 500896 472676 500948
rect 494152 500896 494204 500948
rect 464436 497564 464488 497616
rect 485044 497564 485096 497616
rect 454684 497496 454736 497548
rect 486240 497496 486292 497548
rect 453304 497428 453356 497480
rect 489920 497428 489972 497480
rect 399576 497156 399628 497208
rect 400864 497156 400916 497208
rect 461400 494708 461452 494760
rect 461768 494708 461820 494760
rect 382280 492668 382332 492720
rect 411904 492668 411956 492720
rect 405004 492600 405056 492652
rect 406752 492600 406804 492652
rect 481640 490424 481692 490476
rect 482652 490424 482704 490476
rect 380440 489880 380492 489932
rect 383016 489812 383068 489864
rect 392676 488860 392728 488912
rect 395620 488860 395672 488912
rect 395620 485596 395672 485648
rect 400220 485596 400272 485648
rect 400864 485052 400916 485104
rect 406660 485052 406712 485104
rect 402244 484304 402296 484356
rect 403716 484304 403768 484356
rect 406752 484304 406804 484356
rect 407856 484304 407908 484356
rect 382280 481652 382332 481704
rect 414664 481652 414716 481704
rect 400220 480224 400272 480276
rect 403900 480156 403952 480208
rect 380348 478796 380400 478848
rect 381360 478796 381412 478848
rect 389916 477504 389968 477556
rect 394608 477436 394660 477488
rect 403900 476076 403952 476128
rect 406476 476008 406528 476060
rect 380256 473356 380308 473408
rect 394700 473356 394752 473408
rect 382280 473288 382332 473340
rect 401508 473288 401560 473340
rect 381360 470568 381412 470620
rect 382372 470568 382424 470620
rect 419172 470568 419224 470620
rect 514024 470568 514076 470620
rect 579988 470568 580040 470620
rect 384764 470500 384816 470552
rect 382280 469208 382332 469260
rect 385040 469140 385092 469192
rect 384764 468120 384816 468172
rect 387156 468120 387208 468172
rect 401600 467780 401652 467832
rect 403808 467780 403860 467832
rect 494796 466488 494848 466540
rect 528376 466488 528428 466540
rect 385040 466420 385092 466472
rect 406568 466420 406620 466472
rect 388168 466352 388220 466404
rect 454776 466420 454828 466472
rect 525064 466420 525116 466472
rect 408500 466352 408552 466404
rect 511264 465672 511316 465724
rect 580264 465672 580316 465724
rect 464528 465128 464580 465180
rect 554872 465128 554924 465180
rect 458824 465060 458876 465112
rect 558184 465060 558236 465112
rect 406660 464992 406712 465044
rect 407948 464992 408000 465044
rect 388168 463700 388220 463752
rect 408500 463700 408552 463752
rect 391940 463632 391992 463684
rect 407856 463632 407908 463684
rect 409328 463632 409380 463684
rect 412088 463632 412140 463684
rect 391940 461592 391992 461644
rect 400772 461592 400824 461644
rect 449072 461592 449124 461644
rect 487160 461592 487212 461644
rect 383016 460844 383068 460896
rect 384580 460844 384632 460896
rect 400772 460232 400824 460284
rect 404268 460232 404320 460284
rect 449624 460164 449676 460216
rect 488540 460164 488592 460216
rect 382280 459552 382332 459604
rect 400864 459552 400916 459604
rect 404268 458464 404320 458516
rect 405924 458464 405976 458516
rect 468668 458328 468720 458380
rect 474004 458328 474056 458380
rect 478144 458328 478196 458380
rect 456064 458260 456116 458312
rect 482008 458260 482060 458312
rect 384580 458192 384632 458244
rect 403716 458192 403768 458244
rect 387708 458124 387760 458176
rect 409328 458192 409380 458244
rect 410616 458192 410668 458244
rect 457444 458192 457496 458244
rect 490012 458192 490064 458244
rect 494796 458192 494848 458244
rect 407856 458124 407908 458176
rect 449716 457512 449768 457564
rect 481732 457512 481784 457564
rect 449532 457444 449584 457496
rect 481640 457444 481692 457496
rect 405924 456764 405976 456816
rect 570696 456764 570748 456816
rect 580172 456764 580224 456816
rect 410800 456696 410852 456748
rect 449440 456152 449492 456204
rect 480260 456152 480312 456204
rect 407856 456084 407908 456136
rect 411996 456084 412048 456136
rect 449348 456084 449400 456136
rect 483112 456084 483164 456136
rect 449256 456016 449308 456068
rect 491300 456016 491352 456068
rect 403808 453976 403860 454028
rect 406568 453976 406620 454028
rect 387800 452548 387852 452600
rect 389916 452548 389968 452600
rect 382280 449896 382332 449948
rect 399576 449896 399628 449948
rect 387156 449556 387208 449608
rect 390284 449556 390336 449608
rect 389916 448536 389968 448588
rect 391296 448536 391348 448588
rect 407948 448536 408000 448588
rect 410708 448468 410760 448520
rect 410800 448468 410852 448520
rect 413468 448468 413520 448520
rect 447876 447924 447928 447976
rect 458824 447924 458876 447976
rect 447140 447856 447192 447908
rect 447784 447856 447836 447908
rect 464528 447856 464580 447908
rect 449900 447788 449952 447840
rect 450636 447788 450688 447840
rect 468668 447788 468720 447840
rect 437388 447312 437440 447364
rect 447876 447312 447928 447364
rect 448244 447312 448296 447364
rect 432420 447244 432472 447296
rect 447140 447244 447192 447296
rect 427452 447176 427504 447228
rect 446220 447176 446272 447228
rect 390284 447108 390336 447160
rect 422484 447108 422536 447160
rect 449900 447108 449952 447160
rect 395160 447040 395212 447092
rect 410616 445680 410668 445732
rect 411260 445680 411312 445732
rect 429844 445000 429896 445052
rect 445484 445000 445536 445052
rect 442632 444388 442684 444440
rect 446312 444388 446364 444440
rect 395160 444320 395212 444372
rect 402244 444320 402296 444372
rect 411996 442960 412048 443012
rect 413376 442960 413428 443012
rect 411260 441804 411312 441856
rect 413560 441804 413612 441856
rect 391296 440240 391348 440292
rect 392676 440240 392728 440292
rect 406476 440240 406528 440292
rect 409144 440172 409196 440224
rect 413468 439356 413520 439408
rect 415860 439356 415912 439408
rect 406568 439084 406620 439136
rect 408684 439084 408736 439136
rect 413560 437724 413612 437776
rect 414756 437724 414808 437776
rect 410708 436908 410760 436960
rect 411996 436908 412048 436960
rect 408684 436772 408736 436824
rect 410616 436772 410668 436824
rect 415860 436704 415912 436756
rect 418160 436704 418212 436756
rect 418160 434664 418212 434716
rect 420276 434664 420328 434716
rect 414756 431060 414808 431112
rect 416688 431060 416740 431112
rect 411996 430584 412048 430636
rect 414756 430516 414808 430568
rect 464988 429972 465040 430024
rect 474648 429972 474700 430024
rect 466276 429904 466328 429956
rect 477592 429904 477644 429956
rect 479524 429904 479576 429956
rect 489368 429904 489420 429956
rect 466368 429836 466420 429888
rect 480536 429836 480588 429888
rect 485044 429156 485096 429208
rect 486424 429156 486476 429208
rect 490564 429156 490616 429208
rect 492312 429156 492364 429208
rect 402244 429088 402296 429140
rect 404912 429088 404964 429140
rect 409144 428476 409196 428528
rect 411996 428476 412048 428528
rect 416780 427524 416832 427576
rect 419356 427524 419408 427576
rect 463608 427048 463660 427100
rect 471704 427048 471756 427100
rect 412088 426368 412140 426420
rect 413928 426368 413980 426420
rect 410616 424328 410668 424380
rect 416688 424328 416740 424380
rect 413928 423648 413980 423700
rect 404912 423580 404964 423632
rect 407028 423580 407080 423632
rect 415952 423580 416004 423632
rect 536104 423376 536156 423428
rect 545856 423376 545908 423428
rect 537484 423308 537536 423360
rect 547328 423308 547380 423360
rect 533344 423240 533396 423292
rect 544384 423240 544436 423292
rect 544476 423240 544528 423292
rect 553216 423240 553268 423292
rect 523684 423172 523736 423224
rect 532608 423172 532660 423224
rect 540244 423172 540296 423224
rect 551744 423172 551796 423224
rect 518440 423104 518492 423156
rect 528192 423104 528244 423156
rect 538864 423104 538916 423156
rect 550272 423104 550324 423156
rect 512644 423036 512696 423088
rect 556160 423036 556212 423088
rect 512828 422968 512880 423020
rect 557632 422968 557684 423020
rect 512736 422900 512788 422952
rect 559104 422900 559156 422952
rect 522396 422764 522448 422816
rect 529664 422764 529716 422816
rect 519636 422356 519688 422408
rect 525248 422356 525300 422408
rect 515588 421880 515640 421932
rect 520832 421880 520884 421932
rect 547144 421540 547196 421592
rect 554688 421540 554740 421592
rect 416780 420316 416832 420368
rect 419448 420316 419500 420368
rect 518532 420180 518584 420232
rect 541440 420180 541492 420232
rect 419356 419704 419408 419756
rect 421656 419704 421708 419756
rect 415952 419500 416004 419552
rect 420920 419500 420972 419552
rect 382924 418752 382976 418804
rect 439504 418752 439556 418804
rect 407120 418616 407172 418668
rect 408868 418616 408920 418668
rect 413376 418140 413428 418192
rect 417424 418072 417476 418124
rect 420276 418072 420328 418124
rect 424324 418072 424376 418124
rect 424048 417392 424100 417444
rect 443644 417392 443696 417444
rect 408868 416712 408920 416764
rect 410616 416712 410668 416764
rect 414756 416712 414808 416764
rect 421564 416712 421616 416764
rect 421840 416304 421892 416356
rect 422208 416304 422260 416356
rect 423128 416304 423180 416356
rect 423588 416304 423640 416356
rect 392676 416032 392728 416084
rect 398104 416032 398156 416084
rect 381544 414672 381596 414724
rect 386604 414672 386656 414724
rect 419448 413244 419500 413296
rect 428464 413244 428516 413296
rect 420920 412972 420972 413024
rect 423680 412972 423732 413024
rect 522304 411884 522356 411936
rect 580448 411884 580500 411936
rect 398104 411748 398156 411800
rect 398840 411748 398892 411800
rect 424324 411748 424376 411800
rect 425796 411748 425848 411800
rect 421656 411544 421708 411596
rect 424416 411544 424468 411596
rect 386604 410524 386656 410576
rect 403716 410524 403768 410576
rect 410616 409300 410668 409352
rect 412088 409300 412140 409352
rect 423680 408484 423732 408536
rect 428556 408416 428608 408468
rect 425796 408348 425848 408400
rect 427084 408348 427136 408400
rect 382280 407124 382332 407176
rect 435364 407124 435416 407176
rect 461584 406376 461636 406428
rect 473360 406376 473412 406428
rect 398840 405628 398892 405680
rect 401508 405628 401560 405680
rect 380164 404948 380216 405000
rect 389916 404948 389968 405000
rect 421564 404540 421616 404592
rect 424324 404540 424376 404592
rect 401508 401616 401560 401668
rect 405004 401548 405056 401600
rect 412088 400120 412140 400172
rect 415308 400120 415360 400172
rect 382280 396040 382332 396092
rect 436744 396040 436796 396092
rect 417424 394748 417476 394800
rect 415400 394612 415452 394664
rect 417424 394612 417476 394664
rect 421564 394612 421616 394664
rect 411996 391892 412048 391944
rect 414572 391892 414624 391944
rect 424416 390804 424468 390856
rect 425796 390804 425848 390856
rect 414572 389172 414624 389224
rect 417516 389172 417568 389224
rect 403716 388900 403768 388952
rect 406476 388900 406528 388952
rect 427084 387812 427136 387864
rect 429844 387744 429896 387796
rect 471888 387064 471940 387116
rect 490564 387064 490616 387116
rect 382280 386384 382332 386436
rect 443736 386384 443788 386436
rect 389916 385636 389968 385688
rect 398104 385636 398156 385688
rect 468944 385636 468996 385688
rect 485044 385636 485096 385688
rect 515680 385636 515732 385688
rect 547880 385636 547932 385688
rect 470232 384344 470284 384396
rect 479524 384344 479576 384396
rect 447600 384276 447652 384328
rect 454776 384276 454828 384328
rect 467656 384276 467708 384328
rect 483020 384276 483072 384328
rect 519728 384276 519780 384328
rect 542360 384276 542412 384328
rect 468484 383596 468536 383648
rect 477960 383596 478012 383648
rect 467104 383528 467156 383580
rect 479248 383528 479300 383580
rect 469864 383460 469916 383512
rect 481824 383460 481876 383512
rect 462964 383392 463016 383444
rect 476672 383392 476724 383444
rect 471244 383324 471296 383376
rect 486976 383324 487028 383376
rect 468576 383256 468628 383308
rect 485688 383256 485740 383308
rect 467196 383188 467248 383240
rect 483112 383188 483164 383240
rect 463056 383120 463108 383172
rect 480536 383120 480588 383172
rect 424324 383052 424376 383104
rect 425704 383052 425756 383104
rect 467288 383052 467340 383104
rect 484400 383052 484452 383104
rect 448060 382984 448112 383036
rect 456064 382984 456116 383036
rect 464344 382984 464396 383036
rect 488264 382984 488316 383036
rect 494704 382984 494756 383036
rect 506296 382984 506348 383036
rect 450636 382916 450688 382968
rect 554964 382916 555016 382968
rect 405004 382372 405056 382424
rect 408408 382372 408460 382424
rect 442908 382236 442960 382288
rect 450636 382236 450688 382288
rect 452568 382236 452620 382288
rect 453488 382236 453540 382288
rect 455328 382236 455380 382288
rect 456064 382236 456116 382288
rect 450636 381624 450688 381676
rect 457444 381624 457496 381676
rect 447968 381556 448020 381608
rect 461676 381556 461728 381608
rect 448152 381488 448204 381540
rect 496084 381488 496136 381540
rect 514116 381488 514168 381540
rect 539600 381488 539652 381540
rect 428464 381012 428516 381064
rect 431224 381012 431276 381064
rect 428556 380944 428608 380996
rect 429936 380944 429988 380996
rect 447416 380196 447468 380248
rect 454684 380196 454736 380248
rect 447876 380128 447928 380180
rect 464436 380400 464488 380452
rect 515772 380128 515824 380180
rect 535460 380128 535512 380180
rect 543004 380128 543056 380180
rect 561680 380128 561732 380180
rect 448336 379788 448388 379840
rect 453304 379788 453356 379840
rect 449808 379516 449860 379568
rect 564532 379516 564584 379568
rect 398104 379448 398156 379500
rect 403716 379448 403768 379500
rect 512828 379448 512880 379500
rect 543004 379448 543056 379500
rect 570788 378156 570840 378208
rect 579620 378156 579672 378208
rect 512276 378088 512328 378140
rect 547144 378088 547196 378140
rect 512736 377408 512788 377460
rect 536840 377408 536892 377460
rect 406476 376660 406528 376712
rect 411996 376660 412048 376712
rect 403624 376592 403676 376644
rect 447140 376660 447192 376712
rect 417516 376592 417568 376644
rect 420736 376592 420788 376644
rect 513196 376592 513248 376644
rect 540244 376592 540296 376644
rect 408500 376524 408552 376576
rect 412272 376524 412324 376576
rect 513104 376524 513156 376576
rect 538864 376524 538916 376576
rect 513288 376456 513340 376508
rect 544384 376456 544436 376508
rect 512276 375912 512328 375964
rect 515680 375912 515732 375964
rect 382280 375368 382332 375420
rect 439596 375368 439648 375420
rect 395344 375300 395396 375352
rect 447324 375300 447376 375352
rect 512092 375300 512144 375352
rect 537484 375300 537536 375352
rect 396724 375232 396776 375284
rect 447140 375232 447192 375284
rect 513288 375232 513340 375284
rect 536104 375232 536156 375284
rect 439504 375164 439556 375216
rect 447232 375164 447284 375216
rect 512828 375164 512880 375216
rect 533344 375164 533396 375216
rect 393964 373940 394016 373992
rect 447232 373940 447284 373992
rect 513288 373940 513340 373992
rect 519728 373940 519780 373992
rect 399484 373872 399536 373924
rect 447140 373872 447192 373924
rect 513288 373464 513340 373516
rect 518532 373464 518584 373516
rect 512000 373328 512052 373380
rect 514116 373328 514168 373380
rect 517520 373260 517572 373312
rect 538220 373260 538272 373312
rect 429936 373124 429988 373176
rect 430948 373124 431000 373176
rect 412272 372580 412324 372632
rect 415124 372580 415176 372632
rect 392584 372512 392636 372564
rect 447324 372512 447376 372564
rect 513288 372512 513340 372564
rect 517520 372512 517572 372564
rect 406384 372444 406436 372496
rect 447140 372444 447192 372496
rect 513196 372444 513248 372496
rect 534080 372512 534132 372564
rect 419080 372376 419132 372428
rect 447232 372376 447284 372428
rect 421564 371900 421616 371952
rect 422944 371900 422996 371952
rect 512460 371764 512512 371816
rect 515772 371764 515824 371816
rect 417424 371492 417476 371544
rect 418712 371492 418764 371544
rect 425796 371492 425848 371544
rect 427084 371492 427136 371544
rect 389824 371152 389876 371204
rect 447324 371152 447376 371204
rect 513196 371152 513248 371204
rect 529940 371152 529992 371204
rect 391204 371084 391256 371136
rect 447232 371084 447284 371136
rect 513288 371084 513340 371136
rect 523684 371084 523736 371136
rect 407764 371016 407816 371068
rect 447140 371016 447192 371068
rect 513104 371016 513156 371068
rect 522396 371016 522448 371068
rect 418712 370948 418764 371000
rect 420276 370948 420328 371000
rect 420736 370948 420788 371000
rect 423312 370948 423364 371000
rect 385684 369792 385736 369844
rect 447232 369792 447284 369844
rect 513288 369792 513340 369844
rect 525800 369792 525852 369844
rect 387064 369724 387116 369776
rect 447140 369724 447192 369776
rect 513196 369724 513248 369776
rect 523040 369724 523092 369776
rect 430948 369656 431000 369708
rect 432696 369656 432748 369708
rect 513104 369656 513156 369708
rect 518440 369656 518492 369708
rect 403716 369520 403768 369572
rect 409144 369520 409196 369572
rect 513288 369044 513340 369096
rect 519636 369044 519688 369096
rect 423312 368568 423364 368620
rect 424324 368568 424376 368620
rect 384304 368432 384356 368484
rect 447140 368432 447192 368484
rect 512184 368432 512236 368484
rect 521660 368432 521712 368484
rect 410524 368364 410576 368416
rect 447232 368364 447284 368416
rect 411904 368296 411956 368348
rect 447324 368296 447376 368348
rect 415124 368228 415176 368280
rect 420920 368228 420972 368280
rect 512276 367752 512328 367804
rect 515588 367752 515640 367804
rect 513288 367072 513340 367124
rect 547144 367072 547196 367124
rect 414664 367004 414716 367056
rect 447140 367004 447192 367056
rect 419172 366936 419224 366988
rect 447232 366936 447284 366988
rect 513196 366256 513248 366308
rect 518900 366256 518952 366308
rect 513012 365712 513064 365764
rect 547972 365712 548024 365764
rect 383016 365644 383068 365696
rect 447324 365644 447376 365696
rect 399576 365576 399628 365628
rect 447232 365576 447284 365628
rect 400864 365508 400916 365560
rect 447140 365508 447192 365560
rect 420920 364964 420972 365016
rect 425796 364964 425848 365016
rect 512920 364420 512972 364472
rect 548064 364420 548116 364472
rect 431224 364352 431276 364404
rect 432604 364352 432656 364404
rect 513288 364352 513340 364404
rect 549352 364352 549404 364404
rect 572076 364352 572128 364404
rect 580172 364352 580224 364404
rect 383200 364284 383252 364336
rect 447232 364284 447284 364336
rect 383108 364216 383160 364268
rect 447140 364216 447192 364268
rect 512092 363808 512144 363860
rect 514760 363808 514812 363860
rect 382648 363604 382700 363656
rect 443920 363604 443972 363656
rect 513012 363128 513064 363180
rect 514852 363128 514904 363180
rect 420276 362924 420328 362976
rect 421564 362924 421616 362976
rect 513288 362924 513340 362976
rect 550548 362924 550600 362976
rect 435364 362856 435416 362908
rect 447140 362856 447192 362908
rect 436744 362788 436796 362840
rect 447232 362788 447284 362840
rect 443736 362720 443788 362772
rect 447324 362720 447376 362772
rect 513196 362176 513248 362228
rect 549168 362176 549220 362228
rect 512092 361904 512144 361956
rect 514944 361904 514996 361956
rect 513288 361700 513340 361752
rect 523040 361700 523092 361752
rect 512644 361632 512696 361684
rect 517520 361632 517572 361684
rect 439596 361496 439648 361548
rect 447140 361496 447192 361548
rect 443920 361428 443972 361480
rect 447232 361428 447284 361480
rect 512828 360884 512880 360936
rect 550732 360884 550784 360936
rect 513104 360816 513156 360868
rect 409144 360748 409196 360800
rect 411904 360748 411956 360800
rect 429844 360748 429896 360800
rect 431316 360748 431368 360800
rect 551928 360680 551980 360732
rect 550732 360612 550784 360664
rect 551468 360612 551520 360664
rect 513104 360204 513156 360256
rect 520280 360204 520332 360256
rect 549352 360136 549404 360188
rect 557172 360136 557224 360188
rect 517520 360068 517572 360120
rect 550640 360068 550692 360120
rect 547144 360000 547196 360052
rect 568764 360000 568816 360052
rect 550548 359932 550600 359984
rect 553860 359932 553912 359984
rect 514760 359864 514812 359916
rect 555792 359864 555844 359916
rect 547972 359796 548024 359848
rect 567384 359796 567436 359848
rect 425796 359456 425848 359508
rect 427268 359456 427320 359508
rect 444012 358912 444064 358964
rect 447324 358912 447376 358964
rect 439780 358844 439832 358896
rect 447140 358844 447192 358896
rect 433984 358776 434036 358828
rect 447232 358776 447284 358828
rect 513012 358776 513064 358828
rect 523132 358776 523184 358828
rect 425704 358708 425756 358760
rect 427176 358708 427228 358760
rect 551928 358708 551980 358760
rect 559104 358708 559156 358760
rect 424324 358640 424376 358692
rect 426440 358640 426492 358692
rect 514852 358640 514904 358692
rect 552480 358640 552532 358692
rect 548064 358572 548116 358624
rect 562416 358572 562468 358624
rect 549168 358504 549220 358556
rect 560760 358504 560812 358556
rect 518900 358436 518952 358488
rect 565728 358436 565780 358488
rect 551468 358368 551520 358420
rect 564072 358368 564124 358420
rect 513012 357960 513064 358012
rect 520372 357960 520424 358012
rect 512092 357688 512144 357740
rect 514944 357688 514996 357740
rect 440976 357484 441028 357536
rect 447232 357484 447284 357536
rect 435456 357416 435508 357468
rect 447140 357416 447192 357468
rect 513288 357416 513340 357468
rect 523224 357416 523276 357468
rect 443736 356192 443788 356244
rect 447324 356192 447376 356244
rect 512184 356192 512236 356244
rect 514852 356192 514904 356244
rect 439688 356124 439740 356176
rect 447140 356124 447192 356176
rect 436928 356056 436980 356108
rect 447232 356056 447284 356108
rect 512644 356056 512696 356108
rect 516232 356056 516284 356108
rect 512736 354968 512788 355020
rect 517520 354968 517572 355020
rect 426440 354696 426492 354748
rect 513288 354696 513340 354748
rect 523316 354696 523368 354748
rect 430580 354628 430632 354680
rect 432604 354220 432656 354272
rect 434076 354220 434128 354272
rect 512552 354084 512604 354136
rect 517612 354084 517664 354136
rect 411904 353948 411956 354000
rect 423588 353948 423640 354000
rect 513104 353268 513156 353320
rect 518900 353268 518952 353320
rect 512276 352248 512328 352300
rect 520648 352248 520700 352300
rect 513288 351908 513340 351960
rect 523408 351908 523460 351960
rect 430580 351840 430632 351892
rect 434168 351840 434220 351892
rect 512644 351704 512696 351756
rect 516324 351704 516376 351756
rect 513288 351024 513340 351076
rect 520464 351024 520516 351076
rect 423588 350888 423640 350940
rect 431224 350888 431276 350940
rect 512644 350888 512696 350940
rect 516968 350888 517020 350940
rect 422944 350820 422996 350872
rect 425704 350820 425756 350872
rect 513288 350548 513340 350600
rect 517704 350548 517756 350600
rect 421564 350480 421616 350532
rect 423588 350480 423640 350532
rect 424968 350480 425020 350532
rect 447324 350480 447376 350532
rect 431316 350412 431368 350464
rect 433708 350412 433760 350464
rect 426348 350344 426400 350396
rect 447140 350412 447192 350464
rect 427268 350276 427320 350328
rect 428556 350276 428608 350328
rect 426256 350208 426308 350260
rect 447232 350344 447284 350396
rect 513288 349528 513340 349580
rect 518992 349528 519044 349580
rect 512828 349256 512880 349308
rect 520556 349256 520608 349308
rect 512184 349188 512236 349240
rect 515036 349188 515088 349240
rect 427176 349052 427228 349104
rect 428464 349052 428516 349104
rect 423312 348984 423364 349036
rect 447140 349052 447192 349104
rect 443644 348984 443696 349036
rect 447232 348984 447284 349036
rect 513288 348168 513340 348220
rect 520740 348168 520792 348220
rect 513196 347760 513248 347812
rect 521660 347760 521712 347812
rect 422116 347692 422168 347744
rect 447232 347692 447284 347744
rect 422208 347624 422260 347676
rect 447324 347624 447376 347676
rect 428556 347556 428608 347608
rect 429568 347556 429620 347608
rect 423496 347488 423548 347540
rect 447140 347556 447192 347608
rect 512828 346672 512880 346724
rect 519084 346672 519136 346724
rect 513012 346536 513064 346588
rect 521752 346536 521804 346588
rect 427084 346400 427136 346452
rect 512184 346400 512236 346452
rect 513748 346400 513800 346452
rect 430580 346332 430632 346384
rect 433708 346332 433760 346384
rect 435640 346332 435692 346384
rect 513196 345176 513248 345228
rect 519176 345176 519228 345228
rect 407028 345040 407080 345092
rect 447140 345040 447192 345092
rect 513288 345040 513340 345092
rect 521844 345040 521896 345092
rect 446220 344428 446272 344480
rect 447876 344428 447928 344480
rect 513288 344360 513340 344412
rect 520832 344360 520884 344412
rect 423680 344156 423732 344208
rect 426348 344156 426400 344208
rect 512276 343952 512328 344004
rect 515128 343952 515180 344004
rect 425704 343884 425756 343936
rect 427728 343884 427780 343936
rect 512828 343748 512880 343800
rect 521936 343748 521988 343800
rect 382280 343680 382332 343732
rect 386328 343680 386380 343732
rect 382924 343544 382976 343596
rect 447140 343544 447192 343596
rect 426348 343476 426400 343528
rect 429108 343476 429160 343528
rect 411996 342864 412048 342916
rect 418160 342864 418212 342916
rect 512368 342864 512420 342916
rect 515220 342864 515272 342916
rect 513288 342320 513340 342372
rect 519268 342320 519320 342372
rect 428464 342252 428516 342304
rect 434260 342184 434312 342236
rect 386328 341504 386380 341556
rect 402152 341504 402204 341556
rect 512276 341368 512328 341420
rect 513840 341368 513892 341420
rect 512276 341232 512328 341284
rect 519452 341232 519504 341284
rect 435640 341164 435692 341216
rect 438124 341164 438176 341216
rect 513288 340892 513340 340944
rect 522028 340892 522080 340944
rect 427728 340824 427780 340876
rect 430672 340824 430724 340876
rect 430580 340756 430632 340808
rect 432972 340756 433024 340808
rect 418160 340212 418212 340264
rect 432788 340212 432840 340264
rect 413652 340144 413704 340196
rect 449348 340144 449400 340196
rect 513288 339872 513340 339924
rect 517796 339872 517848 339924
rect 513012 339736 513064 339788
rect 518072 339736 518124 339788
rect 512368 339668 512420 339720
rect 515312 339668 515364 339720
rect 512368 339464 512420 339516
rect 514116 339464 514168 339516
rect 429568 339396 429620 339448
rect 433248 339396 433300 339448
rect 449992 339396 450044 339448
rect 450360 339396 450412 339448
rect 450084 339328 450136 339380
rect 450452 339328 450504 339380
rect 449624 339260 449676 339312
rect 450636 339260 450688 339312
rect 447876 339056 447928 339108
rect 450084 339056 450136 339108
rect 450084 338920 450136 338972
rect 450544 338920 450596 338972
rect 383108 338512 383160 338564
rect 447140 338512 447192 338564
rect 429844 338444 429896 338496
rect 450360 338444 450412 338496
rect 425888 338376 425940 338428
rect 450452 338376 450504 338428
rect 513196 338376 513248 338428
rect 517888 338376 517940 338428
rect 417976 338308 418028 338360
rect 450176 338308 450228 338360
rect 414020 338240 414072 338292
rect 450084 338240 450136 338292
rect 512552 338240 512604 338292
rect 515588 338240 515640 338292
rect 410064 338172 410116 338224
rect 449624 338172 449676 338224
rect 513288 338104 513340 338156
rect 522120 338104 522172 338156
rect 434168 338036 434220 338088
rect 437020 338036 437072 338088
rect 420184 337696 420236 337748
rect 439964 337696 440016 337748
rect 418896 337628 418948 337680
rect 442356 337628 442408 337680
rect 416044 337560 416096 337612
rect 440056 337560 440108 337612
rect 418988 337492 419040 337544
rect 445576 337492 445628 337544
rect 413284 337424 413336 337476
rect 439872 337424 439924 337476
rect 418804 337356 418856 337408
rect 449256 337356 449308 337408
rect 512920 337016 512972 337068
rect 516600 337016 516652 337068
rect 430672 336880 430724 336932
rect 432880 336880 432932 336932
rect 382924 336812 382976 336864
rect 447140 336812 447192 336864
rect 383016 336744 383068 336796
rect 447232 336744 447284 336796
rect 513012 336744 513064 336796
rect 522212 336744 522264 336796
rect 402244 336676 402296 336728
rect 442908 336676 442960 336728
rect 447876 336676 447928 336728
rect 429200 336608 429252 336660
rect 431868 336608 431920 336660
rect 513196 335928 513248 335980
rect 517980 335928 518032 335980
rect 442264 335792 442316 335844
rect 447232 335792 447284 335844
rect 443920 335724 443972 335776
rect 447140 335724 447192 335776
rect 513288 335656 513340 335708
rect 519360 335656 519412 335708
rect 512736 335384 512788 335436
rect 516140 335384 516192 335436
rect 431868 335044 431920 335096
rect 434628 335044 434680 335096
rect 439596 334568 439648 334620
rect 447324 334568 447376 334620
rect 434076 334500 434128 334552
rect 435732 334500 435784 334552
rect 513012 334160 513064 334212
rect 516692 334160 516744 334212
rect 433432 334024 433484 334076
rect 434260 333956 434312 334008
rect 435364 334024 435416 334076
rect 436836 334024 436888 334076
rect 447232 334024 447284 334076
rect 512828 334024 512880 334076
rect 516416 334024 516468 334076
rect 436376 333888 436428 333940
rect 447140 333956 447192 334008
rect 437388 333888 437440 333940
rect 512920 332800 512972 332852
rect 516508 332800 516560 332852
rect 513288 332732 513340 332784
rect 519636 332732 519688 332784
rect 440884 332664 440936 332716
rect 447140 332664 447192 332716
rect 432604 332596 432656 332648
rect 447232 332596 447284 332648
rect 512828 332596 512880 332648
rect 523500 332596 523552 332648
rect 433432 331984 433484 332036
rect 439780 331984 439832 332036
rect 434444 331848 434496 331900
rect 444012 331848 444064 331900
rect 513288 331440 513340 331492
rect 519728 331440 519780 331492
rect 443828 331372 443880 331424
rect 447416 331372 447468 331424
rect 443644 331304 443696 331356
rect 447232 331304 447284 331356
rect 432696 331236 432748 331288
rect 439504 331236 439556 331288
rect 447140 331236 447192 331288
rect 512828 331236 512880 331288
rect 516876 331236 516928 331288
rect 435088 331168 435140 331220
rect 436376 331100 436428 331152
rect 438308 331100 438360 331152
rect 432972 330556 433024 330608
rect 436008 330556 436060 330608
rect 436744 330488 436796 330540
rect 447324 330488 447376 330540
rect 434720 329740 434772 329792
rect 438216 329740 438268 329792
rect 446312 329604 446364 329656
rect 448244 329604 448296 329656
rect 431224 329060 431276 329112
rect 435640 329060 435692 329112
rect 512552 328992 512604 329044
rect 514208 328992 514260 329044
rect 512552 328720 512604 328772
rect 513932 328720 513984 328772
rect 442908 328448 442960 328500
rect 447784 328448 447836 328500
rect 448244 328448 448296 328500
rect 513288 328448 513340 328500
rect 523592 328448 523644 328500
rect 432880 328380 432932 328432
rect 433800 328380 433852 328432
rect 435088 328380 435140 328432
rect 437388 328380 437440 328432
rect 513288 327360 513340 327412
rect 520924 327360 520976 327412
rect 438768 327088 438820 327140
rect 448520 327088 448572 327140
rect 435732 327020 435784 327072
rect 437296 327020 437348 327072
rect 437480 327020 437532 327072
rect 439780 327020 439832 327072
rect 447692 327020 447744 327072
rect 450268 327020 450320 327072
rect 438124 325116 438176 325168
rect 440240 325116 440292 325168
rect 434076 324300 434128 324352
rect 440976 324300 441028 324352
rect 437020 323620 437072 323672
rect 440332 323620 440384 323672
rect 433800 323484 433852 323536
rect 436192 323484 436244 323536
rect 436100 322872 436152 322924
rect 442724 322872 442776 322924
rect 435640 322328 435692 322380
rect 440424 322328 440476 322380
rect 433984 322192 434036 322244
rect 443736 322192 443788 322244
rect 511908 322192 511960 322244
rect 580356 322192 580408 322244
rect 438308 321512 438360 321564
rect 438860 321512 438912 321564
rect 439780 321512 439832 321564
rect 440700 321512 440752 321564
rect 511356 320900 511408 320952
rect 580540 320900 580592 320952
rect 509976 320832 510028 320884
rect 580632 320832 580684 320884
rect 437296 320152 437348 320204
rect 442540 320152 442592 320204
rect 440240 320084 440292 320136
rect 441988 320084 442040 320136
rect 442724 320084 442776 320136
rect 445760 320084 445812 320136
rect 449164 319948 449216 320000
rect 461584 319948 461636 320000
rect 572076 319948 572128 320000
rect 446588 319880 446640 319932
rect 462504 319880 462556 319932
rect 468576 319880 468628 319932
rect 470232 319880 470284 319932
rect 570604 319880 570656 319932
rect 432788 319812 432840 319864
rect 451740 319812 451792 319864
rect 451924 319812 451976 319864
rect 474372 319812 474424 319864
rect 485044 319812 485096 319864
rect 570788 319812 570840 319864
rect 451832 319744 451884 319796
rect 461400 319744 461452 319796
rect 469680 319744 469732 319796
rect 518256 319744 518308 319796
rect 436192 319676 436244 319728
rect 451740 319676 451792 319728
rect 451924 319676 451976 319728
rect 484584 319676 484636 319728
rect 437480 319608 437532 319660
rect 446312 319608 446364 319660
rect 446496 319608 446548 319660
rect 451832 319608 451884 319660
rect 469128 319608 469180 319660
rect 514024 319608 514076 319660
rect 440332 319540 440384 319592
rect 484032 319540 484084 319592
rect 445116 319472 445168 319524
rect 471244 319472 471296 319524
rect 500224 319472 500276 319524
rect 580264 319472 580316 319524
rect 438216 319404 438268 319456
rect 446404 319404 446456 319456
rect 481456 319404 481508 319456
rect 579988 319404 580040 319456
rect 447048 319336 447100 319388
rect 483756 319336 483808 319388
rect 446496 319268 446548 319320
rect 460848 319268 460900 319320
rect 433524 319200 433576 319252
rect 435456 319200 435508 319252
rect 446772 319200 446824 319252
rect 438860 319132 438912 319184
rect 479064 319200 479116 319252
rect 485044 319200 485096 319252
rect 461032 319132 461084 319184
rect 484308 319132 484360 319184
rect 472992 319064 473044 319116
rect 461032 318996 461084 319048
rect 471244 318996 471296 319048
rect 482652 318996 482704 319048
rect 442540 318792 442592 318844
rect 445852 318724 445904 318776
rect 446404 318724 446456 318776
rect 463332 318724 463384 318776
rect 478788 318724 478840 318776
rect 481456 318792 481508 318844
rect 480444 318724 480496 318776
rect 489644 318724 489696 318776
rect 458364 318656 458416 318708
rect 580448 318656 580500 318708
rect 445484 318588 445536 318640
rect 460572 318588 460624 318640
rect 469956 318588 470008 318640
rect 577504 318588 577556 318640
rect 444196 318520 444248 318572
rect 460296 318520 460348 318572
rect 470508 318520 470560 318572
rect 516784 318520 516836 318572
rect 441988 318452 442040 318504
rect 444656 318452 444708 318504
rect 449348 318452 449400 318504
rect 471060 318452 471112 318504
rect 480168 318452 480220 318504
rect 522304 318452 522356 318504
rect 468852 318384 468904 318436
rect 509976 318384 510028 318436
rect 469404 318316 469456 318368
rect 511908 318316 511960 318368
rect 445576 318248 445628 318300
rect 462780 318248 462832 318300
rect 479892 318248 479944 318300
rect 518348 318248 518400 318300
rect 446680 318180 446732 318232
rect 472164 318180 472216 318232
rect 479340 318180 479392 318232
rect 458088 318112 458140 318164
rect 462228 318112 462280 318164
rect 478512 318112 478564 318164
rect 479524 318112 479576 318164
rect 480996 318180 481048 318232
rect 481456 318180 481508 318232
rect 487160 318180 487212 318232
rect 488448 318180 488500 318232
rect 489920 318180 489972 318232
rect 491208 318180 491260 318232
rect 494152 318180 494204 318232
rect 494796 318180 494848 318232
rect 498384 318180 498436 318232
rect 543004 318180 543056 318232
rect 500224 318112 500276 318164
rect 503076 318112 503128 318164
rect 548524 318112 548576 318164
rect 440700 318044 440752 318096
rect 444472 318044 444524 318096
rect 461584 318044 461636 318096
rect 445760 317976 445812 318028
rect 473544 317976 473596 318028
rect 445208 317908 445260 317960
rect 471612 317908 471664 317960
rect 477960 318044 478012 318096
rect 478604 318044 478656 318096
rect 484492 318044 484544 318096
rect 485412 318044 485464 318096
rect 485872 318044 485924 318096
rect 486792 318044 486844 318096
rect 487620 318044 487672 318096
rect 488356 318044 488408 318096
rect 490012 318044 490064 318096
rect 490380 318044 490432 318096
rect 494060 318044 494112 318096
rect 494520 318044 494572 318096
rect 497280 318044 497332 318096
rect 548616 318044 548668 318096
rect 477684 317976 477736 318028
rect 478696 317976 478748 318028
rect 481456 317976 481508 318028
rect 476304 317908 476356 317960
rect 477132 317908 477184 317960
rect 477500 317908 477552 317960
rect 480352 317908 480404 317960
rect 481548 317908 481600 317960
rect 484676 317908 484728 317960
rect 485688 317908 485740 317960
rect 485964 317908 486016 317960
rect 486516 317908 486568 317960
rect 487896 317976 487948 318028
rect 488448 317976 488500 318028
rect 518164 317976 518216 318028
rect 488632 317908 488684 317960
rect 489552 317908 489604 317960
rect 489644 317908 489696 317960
rect 515404 317908 515456 317960
rect 456340 317840 456392 317892
rect 461584 317840 461636 317892
rect 462228 317840 462280 317892
rect 580724 317840 580776 317892
rect 446864 317772 446916 317824
rect 471336 317772 471388 317824
rect 479616 317772 479668 317824
rect 511356 317772 511408 317824
rect 445300 317704 445352 317756
rect 482100 317704 482152 317756
rect 486056 317704 486108 317756
rect 487068 317704 487120 317756
rect 490196 317704 490248 317756
rect 490656 317704 490708 317756
rect 491392 317704 491444 317756
rect 492036 317704 492088 317756
rect 492772 317704 492824 317756
rect 493968 317704 494020 317756
rect 444288 317636 444340 317688
rect 470784 317636 470836 317688
rect 485044 317636 485096 317688
rect 486240 317636 486292 317688
rect 490104 317636 490156 317688
rect 490932 317636 490984 317688
rect 491484 317636 491536 317688
rect 492312 317636 492364 317688
rect 471980 317500 472032 317552
rect 474924 317500 474976 317552
rect 460204 317432 460256 317484
rect 465816 317432 465868 317484
rect 472716 317432 472768 317484
rect 475200 317432 475252 317484
rect 446404 317364 446456 317416
rect 447968 317364 448020 317416
rect 459468 317364 459520 317416
rect 571984 317364 572036 317416
rect 459744 317296 459796 317348
rect 573364 317296 573416 317348
rect 458640 317228 458692 317280
rect 570696 317228 570748 317280
rect 458916 317160 458968 317212
rect 519544 317160 519596 317212
rect 459192 317092 459244 317144
rect 515496 317092 515548 317144
rect 445024 317024 445076 317076
rect 481824 317024 481876 317076
rect 440056 316956 440108 317008
rect 471888 316956 471940 317008
rect 444656 316888 444708 316940
rect 473820 316888 473872 316940
rect 439964 316820 440016 316872
rect 473268 316820 473320 316872
rect 481640 316820 481692 316872
rect 485136 316820 485188 316872
rect 446312 316752 446364 316804
rect 474096 316752 474148 316804
rect 494244 316752 494296 316804
rect 495348 316752 495400 316804
rect 450452 316684 450504 316736
rect 451924 316684 451976 316736
rect 439872 316616 439924 316668
rect 472440 316616 472492 316668
rect 440424 316548 440476 316600
rect 463884 316548 463936 316600
rect 445852 316480 445904 316532
rect 463608 316480 463660 316532
rect 444472 316412 444524 316464
rect 463056 316412 463108 316464
rect 456984 316072 457036 316124
rect 457904 316072 457956 316124
rect 457260 316004 457312 316056
rect 457996 316004 458048 316056
rect 442356 315936 442408 315988
rect 481824 315936 481876 315988
rect 498660 315936 498712 315988
rect 499396 315936 499448 315988
rect 501420 315936 501472 315988
rect 502064 315936 502116 315988
rect 450636 315868 450688 315920
rect 452016 315868 452068 315920
rect 450820 315800 450872 315852
rect 453304 315800 453356 315852
rect 448428 315664 448480 315716
rect 480260 315868 480312 315920
rect 497556 315868 497608 315920
rect 498016 315868 498068 315920
rect 500592 315868 500644 315920
rect 500776 315868 500828 315920
rect 501696 315868 501748 315920
rect 502248 315868 502300 315920
rect 449256 315596 449308 315648
rect 480352 315800 480404 315852
rect 455144 315732 455196 315784
rect 476028 315732 476080 315784
rect 500040 315732 500092 315784
rect 500592 315732 500644 315784
rect 454868 315664 454920 315716
rect 510804 315664 510856 315716
rect 456064 315596 456116 315648
rect 512736 315596 512788 315648
rect 456248 315528 456300 315580
rect 512552 315528 512604 315580
rect 454684 315460 454736 315512
rect 512184 315460 512236 315512
rect 454960 315392 455012 315444
rect 513656 315392 513708 315444
rect 448520 315324 448572 315376
rect 471980 315324 472032 315376
rect 478604 315324 478656 315376
rect 538864 315324 538916 315376
rect 455052 315256 455104 315308
rect 516140 315256 516192 315308
rect 456432 315188 456484 315240
rect 456708 315188 456760 315240
rect 457812 315188 457864 315240
rect 461584 315188 461636 315240
rect 463608 315188 463660 315240
rect 464160 315188 464212 315240
rect 473360 315188 473412 315240
rect 486148 315188 486200 315240
rect 455236 315120 455288 315172
rect 465540 315120 465592 315172
rect 434260 315052 434312 315104
rect 436928 315052 436980 315104
rect 456156 314848 456208 314900
rect 456616 314848 456668 314900
rect 462228 314576 462280 314628
rect 464988 314576 465040 314628
rect 479616 314576 479668 314628
rect 481640 314644 481692 314696
rect 481548 314576 481600 314628
rect 484584 314644 484636 314696
rect 467564 314168 467616 314220
rect 467748 314168 467800 314220
rect 460480 314100 460532 314152
rect 491300 314100 491352 314152
rect 440976 314032 441028 314084
rect 475752 314032 475804 314084
rect 499764 314032 499816 314084
rect 550916 314032 550968 314084
rect 459008 313964 459060 314016
rect 495900 313964 495952 314016
rect 496176 313964 496228 314016
rect 550640 313964 550692 314016
rect 455972 313896 456024 313948
rect 566464 313896 566516 313948
rect 466920 313828 466972 313880
rect 467564 313828 467616 313880
rect 468300 313216 468352 313268
rect 580172 313216 580224 313268
rect 472624 313012 472676 313064
rect 474648 313012 474700 313064
rect 465816 312808 465868 312860
rect 473360 312808 473412 312860
rect 460296 312740 460348 312792
rect 488540 312740 488592 312792
rect 499488 312740 499540 312792
rect 460388 312672 460440 312724
rect 488816 312672 488868 312724
rect 501144 312672 501196 312724
rect 501972 312672 502024 312724
rect 502524 312740 502576 312792
rect 549536 312740 549588 312792
rect 550824 312672 550876 312724
rect 458824 312604 458876 312656
rect 492680 312604 492732 312656
rect 498936 312604 498988 312656
rect 550732 312604 550784 312656
rect 456248 312536 456300 312588
rect 518072 312536 518124 312588
rect 460572 311312 460624 311364
rect 465172 311312 465224 311364
rect 461768 311244 461820 311296
rect 463608 311244 463660 311296
rect 500592 311244 500644 311296
rect 551008 311244 551060 311296
rect 458916 311176 458968 311228
rect 494428 311176 494480 311228
rect 501880 311176 501932 311228
rect 552480 311176 552532 311228
rect 456524 311108 456576 311160
rect 558184 311108 558236 311160
rect 477224 310428 477276 310480
rect 481548 310496 481600 310548
rect 443736 310088 443788 310140
rect 448520 310088 448572 310140
rect 459100 309816 459152 309868
rect 495440 309816 495492 309868
rect 501972 309816 502024 309868
rect 552756 309816 552808 309868
rect 452200 309748 452252 309800
rect 463976 309748 464028 309800
rect 477132 309748 477184 309800
rect 562324 309748 562376 309800
rect 502064 308524 502116 308576
rect 552296 308524 552348 308576
rect 497832 308456 497884 308508
rect 549352 308456 549404 308508
rect 456616 308388 456668 308440
rect 569224 308388 569276 308440
rect 457444 307776 457496 307828
rect 462228 307776 462280 307828
rect 465724 307776 465776 307828
rect 472716 307776 472768 307828
rect 433892 307708 433944 307760
rect 439688 307708 439740 307760
rect 483756 307708 483808 307760
rect 485044 307708 485096 307760
rect 488172 307164 488224 307216
rect 529940 307164 529992 307216
rect 496636 307096 496688 307148
rect 549260 307096 549312 307148
rect 478696 307028 478748 307080
rect 544384 307028 544436 307080
rect 473360 306280 473412 306332
rect 477224 306348 477276 306400
rect 458180 306076 458232 306128
rect 461768 306076 461820 306128
rect 438124 306008 438176 306060
rect 460572 306008 460624 306060
rect 474004 306008 474056 306060
rect 484492 306008 484544 306060
rect 406476 305940 406528 305992
rect 485964 305940 486016 305992
rect 383292 305872 383344 305924
rect 443920 305872 443972 305924
rect 477316 305872 477368 305924
rect 570604 305872 570656 305924
rect 403900 305804 403952 305856
rect 511540 305804 511592 305856
rect 403716 305736 403768 305788
rect 511172 305736 511224 305788
rect 380164 305668 380216 305720
rect 512644 305668 512696 305720
rect 380256 305600 380308 305652
rect 512368 305600 512420 305652
rect 438216 304988 438268 305040
rect 440976 304988 441028 305040
rect 488264 304512 488316 304564
rect 531412 304512 531464 304564
rect 410524 304444 410576 304496
rect 514944 304444 514996 304496
rect 382280 304376 382332 304428
rect 442264 304376 442316 304428
rect 448428 304376 448480 304428
rect 458180 304376 458232 304428
rect 467380 304376 467432 304428
rect 573364 304376 573416 304428
rect 407948 304308 408000 304360
rect 516232 304308 516284 304360
rect 381544 304240 381596 304292
rect 512460 304240 512512 304292
rect 481272 303764 481324 303816
rect 483756 303764 483808 303816
rect 472716 303628 472768 303680
rect 475016 303628 475068 303680
rect 401140 303560 401192 303612
rect 510896 303560 510948 303612
rect 404084 303492 404136 303544
rect 514116 303492 514168 303544
rect 403992 303424 404044 303476
rect 515312 303424 515364 303476
rect 403808 303356 403860 303408
rect 515588 303356 515640 303408
rect 401324 303288 401376 303340
rect 513840 303288 513892 303340
rect 401232 303220 401284 303272
rect 513748 303220 513800 303272
rect 398104 303152 398156 303204
rect 510712 303152 510764 303204
rect 401048 303084 401100 303136
rect 515128 303084 515180 303136
rect 400956 303016 401008 303068
rect 515220 303016 515272 303068
rect 381728 302948 381780 303000
rect 512092 302948 512144 303000
rect 381636 302880 381688 302932
rect 512000 302880 512052 302932
rect 456708 302812 456760 302864
rect 555424 302812 555476 302864
rect 400864 302744 400916 302796
rect 465356 302744 465408 302796
rect 440976 302404 441028 302456
rect 443736 302404 443788 302456
rect 446496 302200 446548 302252
rect 448428 302200 448480 302252
rect 478144 302200 478196 302252
rect 479616 302200 479668 302252
rect 3608 302064 3660 302116
rect 4896 302064 4948 302116
rect 477500 301928 477552 301980
rect 481272 301928 481324 301980
rect 457904 301452 457956 301504
rect 536104 301452 536156 301504
rect 395344 300772 395396 300824
rect 510252 300772 510304 300824
rect 395712 300704 395764 300756
rect 509884 300704 509936 300756
rect 398380 300636 398432 300688
rect 515036 300636 515088 300688
rect 392676 300568 392728 300620
rect 510344 300568 510396 300620
rect 395528 300500 395580 300552
rect 513564 300500 513616 300552
rect 398288 300432 398340 300484
rect 517704 300432 517756 300484
rect 395804 300364 395856 300416
rect 516324 300364 516376 300416
rect 392584 300296 392636 300348
rect 514208 300296 514260 300348
rect 395620 300228 395672 300280
rect 517612 300228 517664 300280
rect 395436 300160 395488 300212
rect 517520 300160 517572 300212
rect 392768 300092 392820 300144
rect 516876 300092 516928 300144
rect 448060 300024 448112 300076
rect 546500 300024 546552 300076
rect 477408 299956 477460 300008
rect 559564 299956 559616 300008
rect 461584 299412 461636 299464
rect 580172 299412 580224 299464
rect 435456 299344 435508 299396
rect 438216 299344 438268 299396
rect 470600 298936 470652 298988
rect 473360 298936 473412 298988
rect 475108 298936 475160 298988
rect 477500 298936 477552 298988
rect 387432 298052 387484 298104
rect 510620 298052 510672 298104
rect 390100 297984 390152 298036
rect 516600 297984 516652 298036
rect 390192 297916 390244 297968
rect 516692 297916 516744 297968
rect 390284 297848 390336 297900
rect 517980 297848 518032 297900
rect 390008 297780 390060 297832
rect 517888 297780 517940 297832
rect 389916 297712 389968 297764
rect 517796 297712 517848 297764
rect 387524 297644 387576 297696
rect 519268 297644 519320 297696
rect 387248 297576 387300 297628
rect 519084 297576 519136 297628
rect 387156 297508 387208 297560
rect 519176 297508 519228 297560
rect 387340 297440 387392 297492
rect 519452 297440 519504 297492
rect 387064 297372 387116 297424
rect 520832 297372 520884 297424
rect 452108 297304 452160 297356
rect 457444 297304 457496 297356
rect 457996 297304 458048 297356
rect 533344 297304 533396 297356
rect 457812 296012 457864 296064
rect 537484 296012 537536 296064
rect 380348 295944 380400 295996
rect 512276 295944 512328 295996
rect 394332 295264 394384 295316
rect 513472 295264 513524 295316
rect 393964 295196 394016 295248
rect 513380 295196 513432 295248
rect 399484 295128 399536 295180
rect 520280 295128 520332 295180
rect 382924 295060 382976 295112
rect 508504 295060 508556 295112
rect 384396 294992 384448 295044
rect 516968 294992 517020 295044
rect 381820 294924 381872 294976
rect 514852 294924 514904 294976
rect 384580 294856 384632 294908
rect 518992 294856 519044 294908
rect 384488 294788 384540 294840
rect 520740 294788 520792 294840
rect 381912 294720 381964 294772
rect 518900 294720 518952 294772
rect 383016 294652 383068 294704
rect 520372 294652 520424 294704
rect 382004 294584 382056 294636
rect 520648 294584 520700 294636
rect 478512 294516 478564 294568
rect 540244 294516 540296 294568
rect 457444 294448 457496 294500
rect 492956 294448 493008 294500
rect 444380 294244 444432 294296
rect 446496 294244 446548 294296
rect 399760 293292 399812 293344
rect 485872 293292 485924 293344
rect 488356 293292 488408 293344
rect 531320 293292 531372 293344
rect 440240 293224 440292 293276
rect 444380 293224 444432 293276
rect 467472 293224 467524 293276
rect 576124 293224 576176 293276
rect 471980 292544 472032 292596
rect 475108 292544 475160 292596
rect 476764 292544 476816 292596
rect 478144 292544 478196 292596
rect 397092 292476 397144 292528
rect 514760 292476 514812 292528
rect 383200 292408 383252 292460
rect 510160 292408 510212 292460
rect 388536 292340 388588 292392
rect 516416 292340 516468 292392
rect 385960 292272 386012 292324
rect 516508 292272 516560 292324
rect 391388 292204 391440 292256
rect 522028 292204 522080 292256
rect 388628 292136 388680 292188
rect 519360 292136 519412 292188
rect 383108 292068 383160 292120
rect 513932 292068 513984 292120
rect 391296 292000 391348 292052
rect 522212 292000 522264 292052
rect 391204 291932 391256 291984
rect 522120 291932 522172 291984
rect 385776 291864 385828 291916
rect 519636 291864 519688 291916
rect 385684 291796 385736 291848
rect 519728 291796 519780 291848
rect 467564 291728 467616 291780
rect 574744 291728 574796 291780
rect 396724 291660 396776 291712
rect 486056 291660 486108 291712
rect 466368 290436 466420 290488
rect 571984 290436 572036 290488
rect 468484 290368 468536 290420
rect 470508 290368 470560 290420
rect 405096 289756 405148 289808
rect 523040 289756 523092 289808
rect 402244 289688 402296 289740
rect 523132 289688 523184 289740
rect 399852 289620 399904 289672
rect 523224 289620 523276 289672
rect 396908 289552 396960 289604
rect 520464 289552 520516 289604
rect 397000 289484 397052 289536
rect 520556 289484 520608 289536
rect 399668 289416 399720 289468
rect 523408 289416 523460 289468
rect 399576 289348 399628 289400
rect 523316 289348 523368 289400
rect 396816 289280 396868 289332
rect 521660 289280 521712 289332
rect 394240 289212 394292 289264
rect 521844 289212 521896 289264
rect 394148 289144 394200 289196
rect 521752 289144 521804 289196
rect 394056 289076 394108 289128
rect 521936 289076 521988 289128
rect 405004 289008 405056 289060
rect 520924 289008 520976 289060
rect 432696 288940 432748 288992
rect 435456 288940 435508 288992
rect 479524 288940 479576 288992
rect 580356 288940 580408 288992
rect 467840 288328 467892 288380
rect 471888 288396 471940 288448
rect 467656 287648 467708 287700
rect 580264 287648 580316 287700
rect 436928 286968 436980 287020
rect 440240 287036 440292 287088
rect 403624 286424 403676 286476
rect 476212 286424 476264 286476
rect 407856 286356 407908 286408
rect 523592 286356 523644 286408
rect 405188 286288 405240 286340
rect 523500 286288 523552 286340
rect 449164 285676 449216 285728
rect 452200 285676 452252 285728
rect 461676 285676 461728 285728
rect 465816 285676 465868 285728
rect 466184 285608 466236 285660
rect 467840 285676 467892 285728
rect 471520 285676 471572 285728
rect 474004 285676 474056 285728
rect 469864 284724 469916 284776
rect 472624 284724 472676 284776
rect 466460 284316 466512 284368
rect 468484 284316 468536 284368
rect 436652 283636 436704 283688
rect 461676 283636 461728 283688
rect 457720 283568 457772 283620
rect 494336 283568 494388 283620
rect 439688 282140 439740 282192
rect 472716 282140 472768 282192
rect 464344 282072 464396 282124
rect 466184 282072 466236 282124
rect 382280 281460 382332 281512
rect 439596 281460 439648 281512
rect 406660 280780 406712 280832
rect 436652 280780 436704 280832
rect 467748 280780 467800 280832
rect 543096 280780 543148 280832
rect 457812 279420 457864 279472
rect 494244 279420 494296 279472
rect 458088 278060 458140 278112
rect 466368 278060 466420 278112
rect 488448 278060 488500 278112
rect 530032 278060 530084 278112
rect 459560 277992 459612 278044
rect 471520 277992 471572 278044
rect 500684 277992 500736 278044
rect 551192 277992 551244 278044
rect 400220 276632 400272 276684
rect 406660 276632 406712 276684
rect 457628 276632 457680 276684
rect 492864 276632 492916 276684
rect 445760 276020 445812 276072
rect 449164 276020 449216 276072
rect 458180 275408 458232 275460
rect 464344 275408 464396 275460
rect 460664 275340 460716 275392
rect 490196 275340 490248 275392
rect 380440 275272 380492 275324
rect 512828 275272 512880 275324
rect 435548 275000 435600 275052
rect 440976 275000 441028 275052
rect 482468 274660 482520 274712
rect 484676 274660 484728 274712
rect 452568 274116 452620 274168
rect 458088 274116 458140 274168
rect 460572 273980 460624 274032
rect 488908 273980 488960 274032
rect 431224 273912 431276 273964
rect 438124 273912 438176 273964
rect 457536 273912 457588 273964
rect 490104 273912 490156 273964
rect 497924 273912 497976 273964
rect 549444 273912 549496 273964
rect 452292 273232 452344 273284
rect 459560 273232 459612 273284
rect 499396 272552 499448 272604
rect 549628 272552 549680 272604
rect 420184 272484 420236 272536
rect 435548 272484 435600 272536
rect 458732 272484 458784 272536
rect 494152 272484 494204 272536
rect 498016 272484 498068 272536
rect 552388 272484 552440 272536
rect 463332 271804 463384 271856
rect 469864 271872 469916 271924
rect 472716 271804 472768 271856
rect 476764 271872 476816 271924
rect 449256 271396 449308 271448
rect 452568 271396 452620 271448
rect 433984 271260 434036 271312
rect 436928 271260 436980 271312
rect 502156 271260 502208 271312
rect 549812 271260 549864 271312
rect 453028 271192 453080 271244
rect 458180 271192 458232 271244
rect 459376 271192 459428 271244
rect 492772 271192 492824 271244
rect 497740 271192 497792 271244
rect 552204 271192 552256 271244
rect 458640 271124 458692 271176
rect 494060 271124 494112 271176
rect 496728 271124 496780 271176
rect 552020 271124 552072 271176
rect 443920 271056 443972 271108
rect 446496 271056 446548 271108
rect 382280 270444 382332 270496
rect 436836 270444 436888 270496
rect 397184 270104 397236 270156
rect 400220 270104 400272 270156
rect 473268 270036 473320 270088
rect 482468 270036 482520 270088
rect 460756 269968 460808 270020
rect 491576 269968 491628 270020
rect 502248 269968 502300 270020
rect 549720 269968 549772 270020
rect 460112 269900 460164 269952
rect 491484 269900 491536 269952
rect 505008 269900 505060 269952
rect 554780 269900 554832 269952
rect 459468 269832 459520 269884
rect 493048 269832 493100 269884
rect 500776 269832 500828 269884
rect 551376 269832 551428 269884
rect 452200 269764 452252 269816
rect 463332 269764 463384 269816
rect 468944 269764 468996 269816
rect 580356 269764 580408 269816
rect 451280 268744 451332 268796
rect 453028 268744 453080 268796
rect 456708 268676 456760 268728
rect 472716 268676 472768 268728
rect 449348 268608 449400 268660
rect 465724 268608 465776 268660
rect 443736 268540 443788 268592
rect 473268 268540 473320 268592
rect 457904 268472 457956 268524
rect 487160 268472 487212 268524
rect 503260 268472 503312 268524
rect 552572 268472 552624 268524
rect 459284 268404 459336 268456
rect 491668 268404 491720 268456
rect 500500 268404 500552 268456
rect 551284 268404 551336 268456
rect 440976 268336 441028 268388
rect 445760 268336 445812 268388
rect 459192 268336 459244 268388
rect 491392 268336 491444 268388
rect 499120 268336 499172 268388
rect 551100 268336 551152 268388
rect 3700 266636 3752 266688
rect 5264 266636 5316 266688
rect 413284 266364 413336 266416
rect 420184 266364 420236 266416
rect 427820 266364 427872 266416
rect 431224 266364 431276 266416
rect 453028 266364 453080 266416
rect 456708 266364 456760 266416
rect 448520 264868 448572 264920
rect 453028 264936 453080 264988
rect 383384 264188 383436 264240
rect 443828 264188 443880 264240
rect 449716 263508 449768 263560
rect 456800 263508 456852 263560
rect 447784 263440 447836 263492
rect 451280 263440 451332 263492
rect 438124 262692 438176 262744
rect 443920 262692 443972 262744
rect 445760 260380 445812 260432
rect 448428 260380 448480 260432
rect 382280 259360 382332 259412
rect 435364 259360 435416 259412
rect 425704 258952 425756 259004
rect 427820 258952 427872 259004
rect 429568 258340 429620 258392
rect 433984 258340 434036 258392
rect 449164 258068 449216 258120
rect 452292 258068 452344 258120
rect 424140 257320 424192 257372
rect 432696 257320 432748 257372
rect 437480 257320 437532 257372
rect 449348 257320 449400 257372
rect 424324 255280 424376 255332
rect 429568 255280 429620 255332
rect 446128 255212 446180 255264
rect 449256 255280 449308 255332
rect 409144 254532 409196 254584
rect 424140 254532 424192 254584
rect 441068 254532 441120 254584
rect 445668 254532 445720 254584
rect 3516 253920 3568 253972
rect 5172 253920 5224 253972
rect 394424 253920 394476 253972
rect 397184 253920 397236 253972
rect 435364 252900 435416 252952
rect 437480 252900 437532 252952
rect 426348 251812 426400 251864
rect 438124 251812 438176 251864
rect 418804 250452 418856 250504
rect 425704 250452 425756 250504
rect 443828 250384 443880 250436
rect 446128 250384 446180 250436
rect 382280 249704 382332 249756
rect 432604 249704 432656 249756
rect 411260 249024 411312 249076
rect 426348 249024 426400 249076
rect 447876 249024 447928 249076
rect 457996 249024 458048 249076
rect 436008 248480 436060 248532
rect 439688 248480 439740 248532
rect 422944 246304 422996 246356
rect 435364 246304 435416 246356
rect 3976 245964 4028 246016
rect 5080 245964 5132 246016
rect 405280 245624 405332 245676
rect 411260 245624 411312 245676
rect 446496 245624 446548 245676
rect 447784 245624 447836 245676
rect 537484 245556 537536 245608
rect 580172 245556 580224 245608
rect 390376 245148 390428 245200
rect 394424 245148 394476 245200
rect 429844 244876 429896 244928
rect 436008 244876 436060 244928
rect 420920 244196 420972 244248
rect 424324 244264 424376 244316
rect 445024 243176 445076 243228
rect 446496 243176 446548 243228
rect 443000 240864 443052 240916
rect 449164 240864 449216 240916
rect 419540 239844 419592 239896
rect 420920 239844 420972 239896
rect 395896 239368 395948 239420
rect 413284 239368 413336 239420
rect 382280 238688 382332 238740
rect 440884 238688 440936 238740
rect 417424 237396 417476 237448
rect 419540 237396 419592 237448
rect 420184 235628 420236 235680
rect 422944 235628 422996 235680
rect 434904 235424 434956 235476
rect 443000 235424 443052 235476
rect 383292 235220 383344 235272
rect 390376 235220 390428 235272
rect 453304 234948 453356 235000
rect 457168 234948 457220 235000
rect 450084 234608 450136 234660
rect 452200 234608 452252 234660
rect 416044 233860 416096 233912
rect 418804 233860 418856 233912
rect 540244 233180 540296 233232
rect 580172 233180 580224 233232
rect 449164 232704 449216 232756
rect 452108 232704 452160 232756
rect 427084 232500 427136 232552
rect 434904 232500 434956 232552
rect 447784 231820 447836 231872
rect 450084 231820 450136 231872
rect 435456 230392 435508 230444
rect 443828 230460 443880 230512
rect 422944 229984 422996 230036
rect 429844 229984 429896 230036
rect 397184 229100 397236 229152
rect 405280 229100 405332 229152
rect 387616 227740 387668 227792
rect 395896 227740 395948 227792
rect 382280 227672 382332 227724
rect 436744 227672 436796 227724
rect 411260 226992 411312 227044
rect 416044 226992 416096 227044
rect 421564 224204 421616 224256
rect 427084 224204 427136 224256
rect 438124 224204 438176 224256
rect 441068 224204 441120 224256
rect 416780 223728 416832 223780
rect 420184 223728 420236 223780
rect 444196 223252 444248 223304
rect 449164 223252 449216 223304
rect 452016 222096 452068 222148
rect 457352 222096 457404 222148
rect 433984 220736 434036 220788
rect 435456 220736 435508 220788
rect 408776 220328 408828 220380
rect 411260 220328 411312 220380
rect 411260 220056 411312 220108
rect 416780 220056 416832 220108
rect 435364 219444 435416 219496
rect 444196 219444 444248 219496
rect 442724 218084 442776 218136
rect 445024 218084 445076 218136
rect 417516 216928 417568 216980
rect 422944 216928 422996 216980
rect 440884 216656 440936 216708
rect 442724 216656 442776 216708
rect 3424 215500 3476 215552
rect 5356 215500 5408 215552
rect 406936 215296 406988 215348
rect 411260 215296 411312 215348
rect 413284 215296 413336 215348
rect 417424 215296 417476 215348
rect 384672 214548 384724 214600
rect 397184 214548 397236 214600
rect 399944 213188 399996 213240
rect 408776 213188 408828 213240
rect 3884 212440 3936 212492
rect 4988 212440 5040 212492
rect 402980 212440 403032 212492
rect 406936 212440 406988 212492
rect 436744 212440 436796 212492
rect 438124 212440 438176 212492
rect 425704 211760 425756 211812
rect 440976 211760 441028 211812
rect 443828 211284 443880 211336
rect 447784 211284 447836 211336
rect 383384 207612 383436 207664
rect 399944 207612 399996 207664
rect 451924 207204 451976 207256
rect 456800 207204 456852 207256
rect 382280 206932 382332 206984
rect 439504 206932 439556 206984
rect 533344 206932 533396 206984
rect 579804 206932 579856 206984
rect 393136 206320 393188 206372
rect 402980 206320 403032 206372
rect 395896 206252 395948 206304
rect 409144 206252 409196 206304
rect 411904 205572 411956 205624
rect 413284 205572 413336 205624
rect 432328 202784 432380 202836
rect 435364 202784 435416 202836
rect 422944 201424 422996 201476
rect 425704 201424 425756 201476
rect 438860 201424 438912 201476
rect 440884 201424 440936 201476
rect 408500 199452 408552 199504
rect 421564 199452 421616 199504
rect 384764 199384 384816 199436
rect 395896 199384 395948 199436
rect 402428 199384 402480 199436
rect 417516 199384 417568 199436
rect 432972 198704 433024 198756
rect 433984 198704 434036 198756
rect 433984 197344 434036 197396
rect 436744 197344 436796 197396
rect 429936 196936 429988 196988
rect 432972 196936 433024 196988
rect 400772 196596 400824 196648
rect 408500 196596 408552 196648
rect 436744 195984 436796 196036
rect 438860 195984 438912 196036
rect 382280 195916 382332 195968
rect 443644 195916 443696 195968
rect 429844 193944 429896 193996
rect 432328 193944 432380 193996
rect 410616 193740 410668 193792
rect 411904 193740 411956 193792
rect 538864 193128 538916 193180
rect 580172 193128 580224 193180
rect 398472 192856 398524 192908
rect 400772 192856 400824 192908
rect 440240 189048 440292 189100
rect 443828 189048 443880 189100
rect 4896 188028 4948 188080
rect 6184 188028 6236 188080
rect 3608 187688 3660 187740
rect 4804 187688 4856 187740
rect 407120 187688 407172 187740
rect 410616 187688 410668 187740
rect 416044 187076 416096 187128
rect 422944 187076 422996 187128
rect 439504 186532 439556 186584
rect 443736 186532 443788 186584
rect 390376 186328 390428 186380
rect 393136 186328 393188 186380
rect 382280 186260 382332 186312
rect 447140 186260 447192 186312
rect 382096 186192 382148 186244
rect 384764 186192 384816 186244
rect 447140 185580 447192 185632
rect 448152 185580 448204 185632
rect 536840 185580 536892 185632
rect 428464 185444 428516 185496
rect 429936 185444 429988 185496
rect 405556 183880 405608 183932
rect 407120 183880 407172 183932
rect 432788 183540 432840 183592
rect 433984 183540 434036 183592
rect 438860 183064 438912 183116
rect 440240 183064 440292 183116
rect 397276 182384 397328 182436
rect 402428 182384 402480 182436
rect 397368 182112 397420 182164
rect 405556 182180 405608 182232
rect 431224 182180 431276 182232
rect 432788 182180 432840 182232
rect 435364 182112 435416 182164
rect 436744 182112 436796 182164
rect 436100 179392 436152 179444
rect 438860 179392 438912 179444
rect 543096 179324 543148 179376
rect 580172 179324 580224 179376
rect 401416 178644 401468 178696
rect 416044 178644 416096 178696
rect 393136 175924 393188 175976
rect 397276 175924 397328 175976
rect 426440 175924 426492 175976
rect 428464 175924 428516 175976
rect 430580 175924 430632 175976
rect 436100 175924 436152 175976
rect 422944 175856 422996 175908
rect 429844 175856 429896 175908
rect 382280 175176 382332 175228
rect 447140 175176 447192 175228
rect 447508 175176 447560 175228
rect 447140 174496 447192 174548
rect 532700 174496 532752 174548
rect 395252 173952 395304 174004
rect 397368 173952 397420 174004
rect 423680 173816 423732 173868
rect 426440 173884 426492 173936
rect 380532 173136 380584 173188
rect 390376 173136 390428 173188
rect 429292 172456 429344 172508
rect 431224 172456 431276 172508
rect 393320 172048 393372 172100
rect 395252 172048 395304 172100
rect 429200 171776 429252 171828
rect 430580 171776 430632 171828
rect 422300 169736 422352 169788
rect 423680 169736 423732 169788
rect 388720 169056 388772 169108
rect 393320 169056 393372 169108
rect 449808 169056 449860 169108
rect 452844 169056 452896 169108
rect 386144 168988 386196 169040
rect 401416 168988 401468 169040
rect 423128 168308 423180 168360
rect 429200 168376 429252 168428
rect 449348 168036 449400 168088
rect 456800 168036 456852 168088
rect 457260 167968 457312 168020
rect 482376 167968 482428 168020
rect 430764 167900 430816 167952
rect 439504 167900 439556 167952
rect 456892 167900 456944 167952
rect 457352 167900 457404 167952
rect 487160 167900 487212 167952
rect 419724 167832 419776 167884
rect 458088 167832 458140 167884
rect 416228 167764 416280 167816
rect 456892 167764 456944 167816
rect 491576 167764 491628 167816
rect 404452 167696 404504 167748
rect 422944 167696 422996 167748
rect 427084 167696 427136 167748
rect 450544 167696 450596 167748
rect 500960 167696 501012 167748
rect 411904 167628 411956 167680
rect 456800 167628 456852 167680
rect 457996 167628 458048 167680
rect 537484 167628 537536 167680
rect 457260 167560 457312 167612
rect 445668 167152 445720 167204
rect 446404 167152 446456 167204
rect 384764 167084 384816 167136
rect 393136 167084 393188 167136
rect 430856 167084 430908 167136
rect 449900 167084 449952 167136
rect 450912 167084 450964 167136
rect 383476 167016 383528 167068
rect 434444 167016 434496 167068
rect 449992 167016 450044 167068
rect 450544 167016 450596 167068
rect 536104 166948 536156 167000
rect 580172 166948 580224 167000
rect 450912 166336 450964 166388
rect 504364 166336 504416 166388
rect 450544 166268 450596 166320
rect 508504 166268 508556 166320
rect 408040 165724 408092 165776
rect 416228 165724 416280 165776
rect 391572 165656 391624 165708
rect 411904 165656 411956 165708
rect 438032 165656 438084 165708
rect 438768 165656 438820 165708
rect 514760 165656 514812 165708
rect 406660 165588 406712 165640
rect 427084 165588 427136 165640
rect 442724 165588 442776 165640
rect 442908 165588 442960 165640
rect 519176 165588 519228 165640
rect 3792 165520 3844 165572
rect 4896 165520 4948 165572
rect 5264 165520 5316 165572
rect 6276 165520 6328 165572
rect 409880 165452 409932 165504
rect 422208 165452 422260 165504
rect 407672 165384 407724 165436
rect 423128 165384 423180 165436
rect 408500 165316 408552 165368
rect 429292 165316 429344 165368
rect 409512 165248 409564 165300
rect 435364 165248 435416 165300
rect 404176 165180 404228 165232
rect 430856 165180 430908 165232
rect 409236 165112 409288 165164
rect 437986 165112 438038 165164
rect 409328 165044 409380 165096
rect 441666 165044 441718 165096
rect 442724 165044 442776 165096
rect 386052 164976 386104 165028
rect 419724 164976 419776 165028
rect 409420 164908 409472 164960
rect 445208 164908 445260 164960
rect 448336 164908 448388 164960
rect 469864 164908 469916 164960
rect 387708 164840 387760 164892
rect 430764 164840 430816 164892
rect 445668 164840 445720 164892
rect 523776 164840 523828 164892
rect 401600 163548 401652 163600
rect 407672 163548 407724 163600
rect 394516 163412 394568 163464
rect 404452 163412 404504 163464
rect 404360 163208 404412 163260
rect 409880 163208 409932 163260
rect 405556 163140 405608 163192
rect 408500 163140 408552 163192
rect 401416 161440 401468 161492
rect 405556 161440 405608 161492
rect 456800 161236 456852 161288
rect 459008 161236 459060 161288
rect 402428 160080 402480 160132
rect 404360 160080 404412 160132
rect 456800 159944 456852 159996
rect 459100 159944 459152 159996
rect 397184 158652 397236 158704
rect 401600 158720 401652 158772
rect 456800 157020 456852 157072
rect 458916 157020 458968 157072
rect 456800 155320 456852 155372
rect 458732 155320 458784 155372
rect 406844 155252 406896 155304
rect 409512 155252 409564 155304
rect 382280 154504 382332 154556
rect 409420 154504 409472 154556
rect 456800 154096 456852 154148
rect 458640 154096 458692 154148
rect 486424 153824 486476 153876
rect 528560 153824 528612 153876
rect 504364 153144 504416 153196
rect 505468 153144 505520 153196
rect 544384 153144 544436 153196
rect 580172 153144 580224 153196
rect 392400 152464 392452 152516
rect 398472 152464 398524 152516
rect 537484 152464 537536 152516
rect 542912 152464 542964 152516
rect 508504 151852 508556 151904
rect 510068 151852 510120 151904
rect 542912 151784 542964 151836
rect 551468 151784 551520 151836
rect 3700 150696 3752 150748
rect 5264 150696 5316 150748
rect 456892 150628 456944 150680
rect 459376 150628 459428 150680
rect 400220 150492 400272 150544
rect 402428 150492 402480 150544
rect 5172 150424 5224 150476
rect 6460 150424 6512 150476
rect 399944 150424 399996 150476
rect 401416 150424 401468 150476
rect 456800 150152 456852 150204
rect 459468 150152 459520 150204
rect 543004 149676 543056 149728
rect 552664 149676 552716 149728
rect 548616 149472 548668 149524
rect 552848 149472 552900 149524
rect 548524 149404 548576 149456
rect 552112 149404 552164 149456
rect 388168 149064 388220 149116
rect 392400 149064 392452 149116
rect 384856 147636 384908 147688
rect 387708 147636 387760 147688
rect 395896 147636 395948 147688
rect 400220 147636 400272 147688
rect 549168 146004 549220 146056
rect 549904 146004 549956 146056
rect 456800 144644 456852 144696
rect 458824 144644 458876 144696
rect 382280 143488 382332 143540
rect 409328 143488 409380 143540
rect 456800 143148 456852 143200
rect 459284 143148 459336 143200
rect 386236 142944 386288 142996
rect 388168 142944 388220 142996
rect 552112 142876 552164 142928
rect 552664 142876 552716 142928
rect 552664 142740 552716 142792
rect 552848 142740 552900 142792
rect 457260 141652 457312 141704
rect 460112 141652 460164 141704
rect 456800 140428 456852 140480
rect 459192 140428 459244 140480
rect 5080 140088 5132 140140
rect 6368 140088 6420 140140
rect 576124 139340 576176 139392
rect 580172 139340 580224 139392
rect 457260 138864 457312 138916
rect 460756 138864 460808 138916
rect 3516 138320 3568 138372
rect 5080 138320 5132 138372
rect 394424 137980 394476 138032
rect 395896 137980 395948 138032
rect 457260 137844 457312 137896
rect 460480 137844 460532 137896
rect 390560 137368 390612 137420
rect 394516 137368 394568 137420
rect 384948 133560 385000 133612
rect 390560 133560 390612 133612
rect 457076 132880 457128 132932
rect 460664 132880 460716 132932
rect 382280 132404 382332 132456
rect 409236 132404 409288 132456
rect 382188 131112 382240 131164
rect 384856 131112 384908 131164
rect 457444 128188 457496 128240
rect 460572 128188 460624 128240
rect 405280 127508 405332 127560
rect 406844 127508 406896 127560
rect 558184 126896 558236 126948
rect 580172 126896 580224 126948
rect 395896 125468 395948 125520
rect 397184 125468 397236 125520
rect 457352 125196 457404 125248
rect 460388 125196 460440 125248
rect 457076 122544 457128 122596
rect 460296 122544 460348 122596
rect 400220 121388 400272 121440
rect 405280 121456 405332 121508
rect 380624 118872 380676 118924
rect 384948 118872 385000 118924
rect 3976 115880 4028 115932
rect 5172 115880 5224 115932
rect 5356 115880 5408 115932
rect 6552 115880 6604 115932
rect 395988 115880 396040 115932
rect 399944 115948 399996 116000
rect 394516 115540 394568 115592
rect 395896 115540 395948 115592
rect 397368 115200 397420 115252
rect 400128 115200 400180 115252
rect 6184 114588 6236 114640
rect 7748 114588 7800 114640
rect 391664 113092 391716 113144
rect 395988 113160 396040 113212
rect 562324 113092 562376 113144
rect 579804 113092 579856 113144
rect 391112 111800 391164 111852
rect 394424 111800 394476 111852
rect 382280 111732 382332 111784
rect 404176 111732 404228 111784
rect 393136 111052 393188 111104
rect 397368 111052 397420 111104
rect 6276 108944 6328 108996
rect 7564 108944 7616 108996
rect 6460 104864 6512 104916
rect 7656 104864 7708 104916
rect 5172 104796 5224 104848
rect 6276 104796 6328 104848
rect 4988 104728 5040 104780
rect 6184 104728 6236 104780
rect 388812 103436 388864 103488
rect 391112 103504 391164 103556
rect 3424 102144 3476 102196
rect 5172 102144 5224 102196
rect 3884 101532 3936 101584
rect 4988 101532 5040 101584
rect 385040 100716 385092 100768
rect 393136 100716 393188 100768
rect 382280 100648 382332 100700
rect 406660 100648 406712 100700
rect 574744 100648 574796 100700
rect 580172 100648 580224 100700
rect 391756 99968 391808 100020
rect 394516 99968 394568 100020
rect 383476 99288 383528 99340
rect 385040 99356 385092 99408
rect 3424 96636 3476 96688
rect 20904 96636 20956 96688
rect 6276 96092 6328 96144
rect 8208 96092 8260 96144
rect 5172 91196 5224 91248
rect 6276 91196 6328 91248
rect 380716 91060 380768 91112
rect 383476 91060 383528 91112
rect 6368 90924 6420 90976
rect 7932 90924 7984 90976
rect 3700 90312 3752 90364
rect 10968 90312 11020 90364
rect 3792 89700 3844 89752
rect 5448 89700 5500 89752
rect 382280 89632 382332 89684
rect 409144 89632 409196 89684
rect 8300 88272 8352 88324
rect 11704 88272 11756 88324
rect 381452 87864 381504 87916
rect 384764 87864 384816 87916
rect 383476 87320 383528 87372
rect 386144 87320 386196 87372
rect 555424 86912 555476 86964
rect 580172 86912 580224 86964
rect 5540 86572 5592 86624
rect 8024 86572 8076 86624
rect 382832 86232 382884 86284
rect 387616 86232 387668 86284
rect 383568 85552 383620 85604
rect 386236 85552 386288 85604
rect 11060 85484 11112 85536
rect 13728 85484 13780 85536
rect 386144 85484 386196 85536
rect 388812 85552 388864 85604
rect 387616 85484 387668 85536
rect 388720 85484 388772 85536
rect 6552 84260 6604 84312
rect 7840 84260 7892 84312
rect 3332 84192 3384 84244
rect 18604 84192 18656 84244
rect 387800 84124 387852 84176
rect 391664 84192 391716 84244
rect 5080 83172 5132 83224
rect 6000 83172 6052 83224
rect 384764 82832 384816 82884
rect 387616 82832 387668 82884
rect 389456 82832 389508 82884
rect 391756 82832 391808 82884
rect 7748 82084 7800 82136
rect 9128 82084 9180 82136
rect 11704 81404 11756 81456
rect 386236 81404 386288 81456
rect 387800 81404 387852 81456
rect 15844 81336 15896 81388
rect 4988 80044 5040 80096
rect 387616 80044 387668 80096
rect 389456 80044 389508 80096
rect 8392 79976 8444 80028
rect 382280 79908 382332 79960
rect 386052 79908 386104 79960
rect 13728 78684 13780 78736
rect 4896 78616 4948 78668
rect 7748 78616 7800 78668
rect 17224 78616 17276 78668
rect 6000 78548 6052 78600
rect 8944 78548 8996 78600
rect 5540 78480 5592 78532
rect 9036 78480 9088 78532
rect 9036 76440 9088 76492
rect 10968 76440 11020 76492
rect 9128 75828 9180 75880
rect 10324 75828 10376 75880
rect 8392 75760 8444 75812
rect 11704 75760 11756 75812
rect 6276 75148 6328 75200
rect 6920 75148 6972 75200
rect 15844 73176 15896 73228
rect 17316 73176 17368 73228
rect 386052 73176 386104 73228
rect 387616 73176 387668 73228
rect 559564 73108 559616 73160
rect 580172 73108 580224 73160
rect 6920 72564 6972 72616
rect 9588 72564 9640 72616
rect 7748 70932 7800 70984
rect 9404 70932 9456 70984
rect 8300 70184 8352 70236
rect 10416 70184 10468 70236
rect 3608 70116 3660 70168
rect 4988 70116 5040 70168
rect 4804 70048 4856 70100
rect 5540 70048 5592 70100
rect 382280 68960 382332 69012
rect 408040 68960 408092 69012
rect 10968 67600 11020 67652
rect 9680 67532 9732 67584
rect 12256 67532 12308 67584
rect 15108 67532 15160 67584
rect 9404 67464 9456 67516
rect 10968 67464 11020 67516
rect 8944 66172 8996 66224
rect 12348 66172 12400 66224
rect 5540 65152 5592 65204
rect 7748 65152 7800 65204
rect 4988 65084 5040 65136
rect 7288 65084 7340 65136
rect 11704 64880 11756 64932
rect 15108 64812 15160 64864
rect 17316 63384 17368 63436
rect 18696 63384 18748 63436
rect 10968 63248 11020 63300
rect 14464 63248 14516 63300
rect 7288 61004 7340 61056
rect 11244 61004 11296 61056
rect 10416 60732 10468 60784
rect 12256 60664 12308 60716
rect 13820 60664 13872 60716
rect 573364 60664 573416 60716
rect 580172 60664 580224 60716
rect 13544 60596 13596 60648
rect 12440 59372 12492 59424
rect 15200 59304 15252 59356
rect 17316 59304 17368 59356
rect 17868 59236 17920 59288
rect 13820 59168 13872 59220
rect 17408 59168 17460 59220
rect 15292 59100 15344 59152
rect 18880 59100 18932 59152
rect 8300 57876 8352 57928
rect 13268 57876 13320 57928
rect 17224 57876 17276 57928
rect 18328 57876 18380 57928
rect 382280 57876 382332 57928
rect 391572 57876 391624 57928
rect 6184 56924 6236 56976
rect 8208 56924 8260 56976
rect 11244 56584 11296 56636
rect 7656 56516 7708 56568
rect 8668 56516 8720 56568
rect 16488 56516 16540 56568
rect 7840 56448 7892 56500
rect 10968 56448 11020 56500
rect 7564 56380 7616 56432
rect 10876 56380 10928 56432
rect 13544 55428 13596 55480
rect 18052 55428 18104 55480
rect 14464 54612 14516 54664
rect 15568 54612 15620 54664
rect 17408 54068 17460 54120
rect 19340 54068 19392 54120
rect 10324 53796 10376 53848
rect 15200 53728 15252 53780
rect 11060 53660 11112 53712
rect 13820 53660 13872 53712
rect 17316 53660 17368 53712
rect 19524 53660 19576 53712
rect 538128 53184 538180 53236
rect 551468 53184 551520 53236
rect 8668 53116 8720 53168
rect 20444 53116 20496 53168
rect 7748 53048 7800 53100
rect 20628 53048 20680 53100
rect 540612 53048 540664 53100
rect 554780 53048 554832 53100
rect 13268 52436 13320 52488
rect 10876 52368 10928 52420
rect 12440 52368 12492 52420
rect 19248 52368 19300 52420
rect 19340 52368 19392 52420
rect 20812 52368 20864 52420
rect 18052 52300 18104 52352
rect 20904 52300 20956 52352
rect 15200 52096 15252 52148
rect 20536 52096 20588 52148
rect 3424 52028 3476 52080
rect 460204 52028 460256 52080
rect 3516 51960 3568 52012
rect 455236 51960 455288 52012
rect 16580 51892 16632 51944
rect 382096 51892 382148 51944
rect 18696 51824 18748 51876
rect 383292 51824 383344 51876
rect 18880 51756 18932 51808
rect 383384 51756 383436 51808
rect 15568 51688 15620 51740
rect 20628 51688 20680 51740
rect 20720 51688 20772 51740
rect 383568 51688 383620 51740
rect 18328 51620 18380 51672
rect 380716 51620 380768 51672
rect 19524 51552 19576 51604
rect 381452 51552 381504 51604
rect 382372 51552 382424 51604
rect 384764 51552 384816 51604
rect 20444 51484 20496 51536
rect 20996 51484 21048 51536
rect 378784 51484 378836 51536
rect 384672 51484 384724 51536
rect 382280 51416 382332 51468
rect 386052 51416 386104 51468
rect 378692 51348 378744 51400
rect 386236 51348 386288 51400
rect 377956 51280 378008 51332
rect 382832 51280 382884 51332
rect 378876 51212 378928 51264
rect 386144 51212 386196 51264
rect 21364 51008 21416 51060
rect 455144 51008 455196 51060
rect 8300 50940 8352 50992
rect 377956 50940 378008 50992
rect 17960 50872 18012 50924
rect 382188 50872 382240 50924
rect 20628 50804 20680 50856
rect 383476 50804 383528 50856
rect 19248 50736 19300 50788
rect 378784 50736 378836 50788
rect 20812 50668 20864 50720
rect 380624 50668 380676 50720
rect 20904 50600 20956 50652
rect 380532 50600 380584 50652
rect 65524 50532 65576 50584
rect 401324 50532 401376 50584
rect 20536 50464 20588 50516
rect 33140 50464 33192 50516
rect 62028 50464 62080 50516
rect 403992 50464 404044 50516
rect 20996 50396 21048 50448
rect 42800 50396 42852 50448
rect 58440 50396 58492 50448
rect 404084 50396 404136 50448
rect 13820 50328 13872 50380
rect 44180 50328 44232 50380
rect 54944 50328 54996 50380
rect 403808 50328 403860 50380
rect 70308 50260 70360 50312
rect 387524 50260 387576 50312
rect 93952 50192 94004 50244
rect 395804 50192 395856 50244
rect 115204 50124 115256 50176
rect 395712 50124 395764 50176
rect 12440 49648 12492 49700
rect 378692 49648 378744 49700
rect 33140 49580 33192 49632
rect 382280 49580 382332 49632
rect 44180 49512 44232 49564
rect 382372 49512 382424 49564
rect 42800 49444 42852 49496
rect 378876 49444 378928 49496
rect 101036 48220 101088 48272
rect 395620 48220 395672 48272
rect 87972 48152 88024 48204
rect 384580 48152 384632 48204
rect 97448 48084 97500 48136
rect 395528 48084 395580 48136
rect 90364 48016 90416 48068
rect 398288 48016 398340 48068
rect 86868 47948 86920 48000
rect 398380 47948 398432 48000
rect 83280 47880 83332 47932
rect 398104 47880 398156 47932
rect 79692 47812 79744 47864
rect 401232 47812 401284 47864
rect 76196 47744 76248 47796
rect 401140 47744 401192 47796
rect 72608 47676 72660 47728
rect 401048 47676 401100 47728
rect 69112 47608 69164 47660
rect 400956 47608 401008 47660
rect 12348 47540 12400 47592
rect 398196 47540 398248 47592
rect 104532 47472 104584 47524
rect 395436 47472 395488 47524
rect 110512 47404 110564 47456
rect 399852 47404 399904 47456
rect 569224 46860 569276 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 399760 45500 399812 45552
rect 66720 45432 66772 45484
rect 387432 45432 387484 45484
rect 122288 45364 122340 45416
rect 454960 45364 455012 45416
rect 118792 45296 118844 45348
rect 454868 45296 454920 45348
rect 50160 45228 50212 45280
rect 388628 45228 388680 45280
rect 48964 45160 49016 45212
rect 390284 45160 390336 45212
rect 44272 45092 44324 45144
rect 390192 45092 390244 45144
rect 40684 45024 40736 45076
rect 392952 45024 393004 45076
rect 37188 44956 37240 45008
rect 392768 44956 392820 45008
rect 33600 44888 33652 44940
rect 393044 44888 393096 44940
rect 26516 44820 26568 44872
rect 392860 44820 392912 44872
rect 108120 44752 108172 44804
rect 407948 44752 408000 44804
rect 111616 44684 111668 44736
rect 410524 44684 410576 44736
rect 91560 42712 91612 42764
rect 384396 42712 384448 42764
rect 469864 42712 469916 42764
rect 536840 42712 536892 42764
rect 98644 42644 98696 42696
rect 394332 42644 394384 42696
rect 84476 42576 84528 42628
rect 384488 42576 384540 42628
rect 80888 42508 80940 42560
rect 387248 42508 387300 42560
rect 77392 42440 77444 42492
rect 387156 42440 387208 42492
rect 73804 42372 73856 42424
rect 387064 42372 387116 42424
rect 63224 42304 63276 42356
rect 387340 42304 387392 42356
rect 59636 42236 59688 42288
rect 389916 42236 389968 42288
rect 56048 42168 56100 42220
rect 390008 42168 390060 42220
rect 52552 42100 52604 42152
rect 390100 42100 390152 42152
rect 41880 42032 41932 42084
rect 385960 42032 386012 42084
rect 95148 41964 95200 42016
rect 382004 41964 382056 42016
rect 102232 41896 102284 41948
rect 381912 41896 381964 41948
rect 123484 39992 123536 40044
rect 397092 39992 397144 40044
rect 116400 39924 116452 39976
rect 393964 39924 394016 39976
rect 119896 39856 119948 39908
rect 399484 39856 399536 39908
rect 105728 39788 105780 39840
rect 391480 39788 391532 39840
rect 45468 39720 45520 39772
rect 388536 39720 388588 39772
rect 38384 39652 38436 39704
rect 385776 39652 385828 39704
rect 34796 39584 34848 39636
rect 385684 39584 385736 39636
rect 31300 39516 31352 39568
rect 385868 39516 385920 39568
rect 27712 39448 27764 39500
rect 383108 39448 383160 39500
rect 23020 39380 23072 39432
rect 383200 39380 383252 39432
rect 18236 39312 18288 39364
rect 382924 39312 382976 39364
rect 109316 39244 109368 39296
rect 381820 39244 381872 39296
rect 112812 39176 112864 39228
rect 383016 39176 383068 39228
rect 96252 37204 96304 37256
rect 399668 37204 399720 37256
rect 92756 37136 92808 37188
rect 396908 37136 396960 37188
rect 89168 37068 89220 37120
rect 397000 37068 397052 37120
rect 85672 37000 85724 37052
rect 396816 37000 396868 37052
rect 82084 36932 82136 36984
rect 394148 36932 394200 36984
rect 75000 36864 75052 36916
rect 394240 36864 394292 36916
rect 71504 36796 71556 36848
rect 394056 36796 394108 36848
rect 64328 36728 64380 36780
rect 391388 36728 391440 36780
rect 57244 36660 57296 36712
rect 391204 36660 391256 36712
rect 53748 36592 53800 36644
rect 391296 36592 391348 36644
rect 60832 36524 60884 36576
rect 456248 36524 456300 36576
rect 103336 36456 103388 36508
rect 399576 36456 399628 36508
rect 124680 34076 124732 34128
rect 405096 34076 405148 34128
rect 121092 34008 121144 34060
rect 402336 34008 402388 34060
rect 117596 33940 117648 33992
rect 402244 33940 402296 33992
rect 39580 33872 39632 33924
rect 405188 33872 405240 33924
rect 24216 33804 24268 33856
rect 405004 33804 405056 33856
rect 19432 33736 19484 33788
rect 402520 33736 402572 33788
rect 3516 33056 3568 33108
rect 400864 33056 400916 33108
rect 570604 33056 570656 33108
rect 580172 33056 580224 33108
rect 3424 20612 3476 20664
rect 403624 20612 403676 20664
rect 571984 20612 572036 20664
rect 579988 20612 580040 20664
rect 3424 6808 3476 6860
rect 396724 6808 396776 6860
rect 566464 6808 566516 6860
rect 580172 6808 580224 6860
rect 67916 4088 67968 4140
rect 380348 4088 380400 4140
rect 32404 4020 32456 4072
rect 381544 4020 381596 4072
rect 99840 3952 99892 4004
rect 454684 3952 454736 4004
rect 14740 3884 14792 3936
rect 380164 3884 380216 3936
rect 13544 3816 13596 3868
rect 384304 3816 384356 3868
rect 21824 3748 21876 3800
rect 392676 3748 392728 3800
rect 17040 3680 17092 3732
rect 395344 3680 395396 3732
rect 28908 3612 28960 3664
rect 407856 3612 407908 3664
rect 8760 3544 8812 3596
rect 389824 3544 389876 3596
rect 43076 3476 43128 3528
rect 456156 3476 456208 3528
rect 35992 3408 36044 3460
rect 456064 3408 456116 3460
rect 78588 3340 78640 3392
rect 380256 3340 380308 3392
rect 106924 3272 106976 3324
rect 381728 3272 381780 3324
rect 114008 3204 114060 3256
rect 381636 3204 381688 3256
rect 30104 2048 30156 2100
rect 392584 2048 392636 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 8128 668545 8156 703520
rect 23480 668772 23532 668778
rect 23480 668714 23532 668720
rect 20720 668704 20772 668710
rect 20720 668646 20772 668652
rect 8114 668536 8170 668545
rect 8114 668471 8170 668480
rect 18880 668432 18932 668438
rect 18880 668374 18932 668380
rect 18788 668228 18840 668234
rect 18788 668170 18840 668176
rect 17868 668160 17920 668166
rect 17868 668102 17920 668108
rect 7564 668092 7616 668098
rect 7564 668034 7616 668040
rect 3792 668024 3844 668030
rect 3792 667966 3844 667972
rect 3424 667956 3476 667962
rect 3424 667898 3476 667904
rect 3436 658209 3464 667898
rect 3700 667616 3752 667622
rect 3700 667558 3752 667564
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3424 655512 3476 655518
rect 3424 655454 3476 655460
rect 3148 619608 3200 619614
rect 3148 619550 3200 619556
rect 3160 619177 3188 619550
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3436 501809 3464 655454
rect 3516 652044 3568 652050
rect 3516 651986 3568 651992
rect 3528 527921 3556 651986
rect 3608 650004 3660 650010
rect 3608 649946 3660 649952
rect 3620 580009 3648 649946
rect 3712 632097 3740 667558
rect 3698 632088 3754 632097
rect 3698 632023 3754 632032
rect 3700 630692 3752 630698
rect 3700 630634 3752 630640
rect 3606 580000 3662 580009
rect 3606 579935 3662 579944
rect 3608 578468 3660 578474
rect 3608 578410 3660 578416
rect 3514 527912 3570 527921
rect 3514 527847 3570 527856
rect 3516 525836 3568 525842
rect 3516 525778 3568 525784
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 3528 423609 3556 525778
rect 3620 462641 3648 578410
rect 3712 514865 3740 630634
rect 3804 606121 3832 667966
rect 7576 660346 7604 668034
rect 17684 666664 17736 666670
rect 17684 666606 17736 666612
rect 16580 665508 16632 665514
rect 16580 665450 16632 665456
rect 13820 665304 13872 665310
rect 13820 665246 13872 665252
rect 10968 665168 11020 665174
rect 10968 665110 11020 665116
rect 10980 662454 11008 665110
rect 11060 663808 11112 663814
rect 11060 663750 11112 663756
rect 8668 662448 8720 662454
rect 8668 662390 8720 662396
rect 10968 662448 11020 662454
rect 10968 662390 11020 662396
rect 5632 660340 5684 660346
rect 5632 660282 5684 660288
rect 7564 660340 7616 660346
rect 7564 660282 7616 660288
rect 5540 659796 5592 659802
rect 5540 659738 5592 659744
rect 5552 654498 5580 659738
rect 5644 655586 5672 660282
rect 8680 659802 8708 662390
rect 8668 659796 8720 659802
rect 8668 659738 8720 659744
rect 9588 659728 9640 659734
rect 9588 659670 9640 659676
rect 8944 658232 8996 658238
rect 8944 658174 8996 658180
rect 7104 656328 7156 656334
rect 7104 656270 7156 656276
rect 5632 655580 5684 655586
rect 5632 655522 5684 655528
rect 4804 654492 4856 654498
rect 4804 654434 4856 654440
rect 5540 654492 5592 654498
rect 5540 654434 5592 654440
rect 4160 626952 4212 626958
rect 4160 626894 4212 626900
rect 4172 622418 4200 626894
rect 3988 622390 4200 622418
rect 3790 606112 3846 606121
rect 3790 606047 3846 606056
rect 3792 587852 3844 587858
rect 3792 587794 3844 587800
rect 3804 566953 3832 587794
rect 3790 566944 3846 566953
rect 3790 566879 3846 566888
rect 3884 565888 3936 565894
rect 3884 565830 3936 565836
rect 3792 553444 3844 553450
rect 3792 553386 3844 553392
rect 3698 514856 3754 514865
rect 3698 514791 3754 514800
rect 3700 507884 3752 507890
rect 3700 507826 3752 507832
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3712 410553 3740 507826
rect 3804 449585 3832 553386
rect 3896 475697 3924 565830
rect 3988 553897 4016 622390
rect 3974 553888 4030 553897
rect 3974 553823 4030 553832
rect 4816 507890 4844 654434
rect 5632 652860 5684 652866
rect 5632 652802 5684 652808
rect 5080 652724 5132 652730
rect 5080 652666 5132 652672
rect 4896 649732 4948 649738
rect 4896 649674 4948 649680
rect 4908 525842 4936 649674
rect 4988 643068 5040 643074
rect 4988 643010 5040 643016
rect 5000 553450 5028 643010
rect 5092 565894 5120 652666
rect 5540 650276 5592 650282
rect 5540 650218 5592 650224
rect 5552 644474 5580 650218
rect 5644 650078 5672 652802
rect 7116 652798 7144 656270
rect 8300 652928 8352 652934
rect 8300 652870 8352 652876
rect 7104 652792 7156 652798
rect 7104 652734 7156 652740
rect 8312 651386 8340 652870
rect 8956 652866 8984 658174
rect 9600 656334 9628 659670
rect 11072 658306 11100 663750
rect 11704 661020 11756 661026
rect 11704 660962 11756 660968
rect 11060 658300 11112 658306
rect 11060 658242 11112 658248
rect 10048 656396 10100 656402
rect 10048 656338 10100 656344
rect 9588 656328 9640 656334
rect 9588 656270 9640 656276
rect 8944 652860 8996 652866
rect 8944 652802 8996 652808
rect 9220 652792 9272 652798
rect 9220 652734 9272 652740
rect 8220 651358 8340 651386
rect 5632 650072 5684 650078
rect 5632 650014 5684 650020
rect 8220 649738 8248 651358
rect 9232 650282 9260 652734
rect 10060 652050 10088 656338
rect 11716 652798 11744 660962
rect 13832 659734 13860 665246
rect 16592 663814 16620 665450
rect 17696 665242 17724 666606
rect 17880 665310 17908 668102
rect 18696 667684 18748 667690
rect 18696 667626 18748 667632
rect 18420 666732 18472 666738
rect 18420 666674 18472 666680
rect 17868 665304 17920 665310
rect 17868 665246 17920 665252
rect 17684 665236 17736 665242
rect 17684 665178 17736 665184
rect 18432 663814 18460 666674
rect 18604 664692 18656 664698
rect 18604 664634 18656 664640
rect 16580 663808 16632 663814
rect 16580 663750 16632 663756
rect 18420 663808 18472 663814
rect 18420 663750 18472 663756
rect 15292 663740 15344 663746
rect 15292 663682 15344 663688
rect 13912 662448 13964 662454
rect 13912 662390 13964 662396
rect 13820 659728 13872 659734
rect 13820 659670 13872 659676
rect 13924 656402 13952 662390
rect 14464 661700 14516 661706
rect 14464 661642 14516 661648
rect 13912 656396 13964 656402
rect 13912 656338 13964 656344
rect 14476 652934 14504 661642
rect 15304 661094 15332 663682
rect 17960 662516 18012 662522
rect 17960 662458 18012 662464
rect 15292 661088 15344 661094
rect 15292 661030 15344 661036
rect 15200 661020 15252 661026
rect 15200 660962 15252 660968
rect 15212 657354 15240 660962
rect 14648 657348 14700 657354
rect 14648 657290 14700 657296
rect 15200 657348 15252 657354
rect 15200 657290 15252 657296
rect 14464 652928 14516 652934
rect 14464 652870 14516 652876
rect 11704 652792 11756 652798
rect 11704 652734 11756 652740
rect 10048 652044 10100 652050
rect 10048 651986 10100 651992
rect 14660 651506 14688 657290
rect 17972 656962 18000 662458
rect 17880 656934 18000 656962
rect 17880 655586 17908 656934
rect 15936 655580 15988 655586
rect 15936 655522 15988 655528
rect 17868 655580 17920 655586
rect 17868 655522 17920 655528
rect 12440 651500 12492 651506
rect 12440 651442 12492 651448
rect 14648 651500 14700 651506
rect 14648 651442 14700 651448
rect 9220 650276 9272 650282
rect 9220 650218 9272 650224
rect 8208 649732 8260 649738
rect 8208 649674 8260 649680
rect 12452 648650 12480 651442
rect 15948 651438 15976 655522
rect 17040 652792 17092 652798
rect 17040 652734 17092 652740
rect 13820 651432 13872 651438
rect 13820 651374 13872 651380
rect 15936 651432 15988 651438
rect 15936 651374 15988 651380
rect 12440 648644 12492 648650
rect 12440 648586 12492 648592
rect 8944 648576 8996 648582
rect 8944 648518 8996 648524
rect 5184 644446 5580 644474
rect 5184 578474 5212 644446
rect 8956 643142 8984 648518
rect 13832 646610 13860 651374
rect 15200 648576 15252 648582
rect 15200 648518 15252 648524
rect 11060 646604 11112 646610
rect 11060 646546 11112 646552
rect 13820 646604 13872 646610
rect 13820 646546 13872 646552
rect 8944 643136 8996 643142
rect 8944 643078 8996 643084
rect 11072 640354 11100 646546
rect 13084 645992 13136 645998
rect 13084 645934 13136 645940
rect 12440 645516 12492 645522
rect 12440 645458 12492 645464
rect 12452 641730 12480 645458
rect 12360 641702 12480 641730
rect 11060 640348 11112 640354
rect 11060 640290 11112 640296
rect 8944 640280 8996 640286
rect 8944 640222 8996 640228
rect 6920 636200 6972 636206
rect 6920 636142 6972 636148
rect 6932 632074 6960 636142
rect 6840 632046 6960 632074
rect 6840 630698 6868 632046
rect 8956 631718 8984 640222
rect 12360 637770 12388 641702
rect 9680 637764 9732 637770
rect 9680 637706 9732 637712
rect 12348 637764 12400 637770
rect 12348 637706 12400 637712
rect 9692 636206 9720 637706
rect 9680 636200 9732 636206
rect 9680 636142 9732 636148
rect 13096 632126 13124 645934
rect 15212 645522 15240 648518
rect 17052 645998 17080 652734
rect 18616 648650 18644 664634
rect 18708 662454 18736 667626
rect 18696 662448 18748 662454
rect 18696 662390 18748 662396
rect 18800 661706 18828 668170
rect 18788 661700 18840 661706
rect 18788 661642 18840 661648
rect 18892 661162 18920 668374
rect 19340 668296 19392 668302
rect 19340 668238 19392 668244
rect 19352 666670 19380 668238
rect 19892 667820 19944 667826
rect 19892 667762 19944 667768
rect 19800 667752 19852 667758
rect 19800 667694 19852 667700
rect 19340 666664 19392 666670
rect 19340 666606 19392 666612
rect 19812 664698 19840 667694
rect 19904 665514 19932 667762
rect 20732 666670 20760 668646
rect 20996 668636 21048 668642
rect 20996 668578 21048 668584
rect 20904 668500 20956 668506
rect 20904 668442 20956 668448
rect 20812 668364 20864 668370
rect 20812 668306 20864 668312
rect 20824 666738 20852 668306
rect 20812 666732 20864 666738
rect 20812 666674 20864 666680
rect 20076 666664 20128 666670
rect 20076 666606 20128 666612
rect 20720 666664 20772 666670
rect 20720 666606 20772 666612
rect 19984 666596 20036 666602
rect 19984 666538 20036 666544
rect 19892 665508 19944 665514
rect 19892 665450 19944 665456
rect 19800 664692 19852 664698
rect 19800 664634 19852 664640
rect 18880 661156 18932 661162
rect 18880 661098 18932 661104
rect 19996 661094 20024 666538
rect 20088 662522 20116 666606
rect 20916 666602 20944 668442
rect 21008 667758 21036 668578
rect 21088 668568 21140 668574
rect 21088 668510 21140 668516
rect 20996 667752 21048 667758
rect 20996 667694 21048 667700
rect 21100 667690 21128 668510
rect 23492 667826 23520 668714
rect 24320 668681 24348 703520
rect 40512 700369 40540 703520
rect 40498 700360 40554 700369
rect 40498 700295 40554 700304
rect 72988 670002 73016 703520
rect 89180 670070 89208 703520
rect 105464 700505 105492 703520
rect 105450 700496 105506 700505
rect 105450 700431 105506 700440
rect 137848 700330 137876 703520
rect 137836 700324 137888 700330
rect 137836 700266 137888 700272
rect 154132 670138 154160 703520
rect 170324 700398 170352 703520
rect 170312 700392 170364 700398
rect 170312 700334 170364 700340
rect 202800 671401 202828 703520
rect 218992 700534 219020 703520
rect 218980 700528 219032 700534
rect 218980 700470 219032 700476
rect 235184 700466 235212 703520
rect 235172 700460 235224 700466
rect 235172 700402 235224 700408
rect 202786 671392 202842 671401
rect 202786 671327 202842 671336
rect 154120 670132 154172 670138
rect 154120 670074 154172 670080
rect 89168 670064 89220 670070
rect 89168 670006 89220 670012
rect 72976 669996 73028 670002
rect 72976 669938 73028 669944
rect 267660 668846 267688 703520
rect 283852 670206 283880 703520
rect 300136 700641 300164 703520
rect 300122 700632 300178 700641
rect 332520 700602 332548 703520
rect 300122 700567 300178 700576
rect 332508 700596 332560 700602
rect 332508 700538 332560 700544
rect 348804 670274 348832 703520
rect 364996 700670 365024 703520
rect 397472 700738 397500 703520
rect 397460 700732 397512 700738
rect 397460 700674 397512 700680
rect 364984 700664 365036 700670
rect 364984 700606 365036 700612
rect 348792 670268 348844 670274
rect 348792 670210 348844 670216
rect 283840 670200 283892 670206
rect 283840 670142 283892 670148
rect 413284 670064 413336 670070
rect 413284 670006 413336 670012
rect 267648 668840 267700 668846
rect 267648 668782 267700 668788
rect 380440 668772 380492 668778
rect 380440 668714 380492 668720
rect 378324 668704 378376 668710
rect 24306 668672 24362 668681
rect 378324 668646 378376 668652
rect 24306 668607 24362 668616
rect 378140 668636 378192 668642
rect 378140 668578 378192 668584
rect 378152 667894 378180 668578
rect 378232 668432 378284 668438
rect 378232 668374 378284 668380
rect 378140 667888 378192 667894
rect 378140 667830 378192 667836
rect 378244 667826 378272 668374
rect 23480 667820 23532 667826
rect 23480 667762 23532 667768
rect 378232 667820 378284 667826
rect 378232 667762 378284 667768
rect 378336 667758 378364 668646
rect 380348 668568 380400 668574
rect 380348 668510 380400 668516
rect 380164 668228 380216 668234
rect 380164 668170 380216 668176
rect 378324 667752 378376 667758
rect 378324 667694 378376 667700
rect 21088 667684 21140 667690
rect 21088 667626 21140 667632
rect 21364 667684 21416 667690
rect 21364 667626 21416 667632
rect 20904 666596 20956 666602
rect 20904 666538 20956 666544
rect 20076 662516 20128 662522
rect 20076 662458 20128 662464
rect 18696 661088 18748 661094
rect 18696 661030 18748 661036
rect 19984 661088 20036 661094
rect 19984 661030 20036 661036
rect 18708 652798 18736 661030
rect 18696 652792 18748 652798
rect 18696 652734 18748 652740
rect 18604 648644 18656 648650
rect 18604 648586 18656 648592
rect 17040 645992 17092 645998
rect 17040 645934 17092 645940
rect 15200 645516 15252 645522
rect 15200 645458 15252 645464
rect 13084 632120 13136 632126
rect 13084 632062 13136 632068
rect 10692 632052 10744 632058
rect 10692 631994 10744 632000
rect 7932 631712 7984 631718
rect 7932 631654 7984 631660
rect 8944 631712 8996 631718
rect 8944 631654 8996 631660
rect 6828 630692 6880 630698
rect 6828 630634 6880 630640
rect 7944 628794 7972 631654
rect 5540 628788 5592 628794
rect 5540 628730 5592 628736
rect 7932 628788 7984 628794
rect 7932 628730 7984 628736
rect 5552 626958 5580 628730
rect 5540 626952 5592 626958
rect 5540 626894 5592 626900
rect 10704 625938 10732 631994
rect 8944 625932 8996 625938
rect 8944 625874 8996 625880
rect 10692 625932 10744 625938
rect 10692 625874 10744 625880
rect 8956 617982 8984 625874
rect 21376 625154 21404 667626
rect 20916 625126 21404 625154
rect 20916 619614 20944 625126
rect 20904 619608 20956 619614
rect 20904 619550 20956 619556
rect 7564 617976 7616 617982
rect 7564 617918 7616 617924
rect 8944 617976 8996 617982
rect 8944 617918 8996 617924
rect 7576 601662 7604 617918
rect 6184 601656 6236 601662
rect 6184 601598 6236 601604
rect 7564 601656 7616 601662
rect 7564 601598 7616 601604
rect 6196 587926 6224 601598
rect 6184 587920 6236 587926
rect 6184 587862 6236 587868
rect 5172 578468 5224 578474
rect 5172 578410 5224 578416
rect 5080 565888 5132 565894
rect 5080 565830 5132 565836
rect 4988 553444 5040 553450
rect 4988 553386 5040 553392
rect 4896 525836 4948 525842
rect 4896 525778 4948 525784
rect 4804 507884 4856 507890
rect 4804 507826 4856 507832
rect 3882 475688 3938 475697
rect 3882 475623 3938 475632
rect 3790 449576 3846 449585
rect 3790 449511 3846 449520
rect 3698 410544 3754 410553
rect 3698 410479 3754 410488
rect 380176 405006 380204 668170
rect 380256 667888 380308 667894
rect 380256 667830 380308 667836
rect 380268 473414 380296 667830
rect 380360 478854 380388 668510
rect 380452 489938 380480 668714
rect 380624 668500 380676 668506
rect 380624 668442 380676 668448
rect 380532 667752 380584 667758
rect 380532 667694 380584 667700
rect 380544 543250 380572 667694
rect 380636 553450 380664 668442
rect 381820 668364 381872 668370
rect 381820 668306 381872 668312
rect 381544 668296 381596 668302
rect 381544 668238 381596 668244
rect 380624 553444 380676 553450
rect 380624 553386 380676 553392
rect 380532 543244 380584 543250
rect 380532 543186 380584 543192
rect 380440 489932 380492 489938
rect 380440 489874 380492 489880
rect 380348 478848 380400 478854
rect 380348 478790 380400 478796
rect 381360 478848 381412 478854
rect 381360 478790 381412 478796
rect 380256 473408 380308 473414
rect 380256 473350 380308 473356
rect 381372 470626 381400 478790
rect 381360 470620 381412 470626
rect 381360 470562 381412 470568
rect 381556 414730 381584 668238
rect 381636 668160 381688 668166
rect 381636 668102 381688 668108
rect 381648 529582 381676 668102
rect 381728 667820 381780 667826
rect 381728 667762 381780 667768
rect 381740 537538 381768 667762
rect 381832 572218 381860 668306
rect 381912 668092 381964 668098
rect 381912 668034 381964 668040
rect 381924 574054 381952 668034
rect 382278 662416 382334 662425
rect 382278 662351 382334 662360
rect 382292 661094 382320 662351
rect 382280 661088 382332 661094
rect 382280 661030 382332 661036
rect 403624 661088 403676 661094
rect 403624 661030 403676 661036
rect 382278 651808 382334 651817
rect 382278 651743 382334 651752
rect 382292 651438 382320 651743
rect 382280 651432 382332 651438
rect 382280 651374 382332 651380
rect 396724 651432 396776 651438
rect 396724 651374 396776 651380
rect 382922 641200 382978 641209
rect 382922 641135 382978 641144
rect 382278 630592 382334 630601
rect 382278 630527 382334 630536
rect 382292 629338 382320 630527
rect 382280 629332 382332 629338
rect 382280 629274 382332 629280
rect 382278 619984 382334 619993
rect 382278 619919 382334 619928
rect 382292 619682 382320 619919
rect 382280 619676 382332 619682
rect 382280 619618 382332 619624
rect 382278 609376 382334 609385
rect 382278 609311 382334 609320
rect 382292 608666 382320 609311
rect 382280 608660 382332 608666
rect 382280 608602 382332 608608
rect 382278 598768 382334 598777
rect 382278 598703 382334 598712
rect 382292 597582 382320 598703
rect 382280 597576 382332 597582
rect 382280 597518 382332 597524
rect 382278 588160 382334 588169
rect 382278 588095 382334 588104
rect 382292 587926 382320 588095
rect 382280 587920 382332 587926
rect 382280 587862 382332 587868
rect 382278 577552 382334 577561
rect 382278 577487 382334 577496
rect 382292 576910 382320 577487
rect 382280 576904 382332 576910
rect 382280 576846 382332 576852
rect 381912 574048 381964 574054
rect 381912 573990 381964 573996
rect 381820 572212 381872 572218
rect 381820 572154 381872 572160
rect 382278 566944 382334 566953
rect 382278 566879 382334 566888
rect 382292 565146 382320 566879
rect 382280 565140 382332 565146
rect 382280 565082 382332 565088
rect 382278 556336 382334 556345
rect 382278 556271 382334 556280
rect 382292 556238 382320 556271
rect 382280 556232 382332 556238
rect 382280 556174 382332 556180
rect 382278 545728 382334 545737
rect 382278 545663 382334 545672
rect 382292 545154 382320 545663
rect 382280 545148 382332 545154
rect 382280 545090 382332 545096
rect 381820 543244 381872 543250
rect 381820 543186 381872 543192
rect 381728 537532 381780 537538
rect 381728 537474 381780 537480
rect 381832 533594 381860 543186
rect 382278 535120 382334 535129
rect 382278 535055 382334 535064
rect 382292 534138 382320 535055
rect 382280 534132 382332 534138
rect 382280 534074 382332 534080
rect 381820 533588 381872 533594
rect 381820 533530 381872 533536
rect 381636 529576 381688 529582
rect 381636 529518 381688 529524
rect 382278 524512 382334 524521
rect 382278 524447 382280 524456
rect 382332 524447 382334 524456
rect 382280 524418 382332 524424
rect 382278 513904 382334 513913
rect 382278 513839 382334 513848
rect 382292 513602 382320 513839
rect 382280 513596 382332 513602
rect 382280 513538 382332 513544
rect 382278 503296 382334 503305
rect 382278 503231 382334 503240
rect 382292 502382 382320 503231
rect 382280 502376 382332 502382
rect 382280 502318 382332 502324
rect 382280 492720 382332 492726
rect 382278 492688 382280 492697
rect 382332 492688 382334 492697
rect 382278 492623 382334 492632
rect 382278 482080 382334 482089
rect 382278 482015 382334 482024
rect 382292 481710 382320 482015
rect 382280 481704 382332 481710
rect 382280 481646 382332 481652
rect 382280 473340 382332 473346
rect 382280 473282 382332 473288
rect 382292 469266 382320 473282
rect 382370 471472 382426 471481
rect 382370 471407 382426 471416
rect 382384 470626 382412 471407
rect 382372 470620 382424 470626
rect 382372 470562 382424 470568
rect 382280 469260 382332 469266
rect 382280 469202 382332 469208
rect 382278 460864 382334 460873
rect 382278 460799 382334 460808
rect 382292 459610 382320 460799
rect 382280 459604 382332 459610
rect 382280 459546 382332 459552
rect 382278 450256 382334 450265
rect 382278 450191 382334 450200
rect 382292 449954 382320 450191
rect 382280 449948 382332 449954
rect 382280 449890 382332 449896
rect 382936 418810 382964 641135
rect 395344 629332 395396 629338
rect 395344 629274 395396 629280
rect 393964 608660 394016 608666
rect 393964 608602 394016 608608
rect 392584 587920 392636 587926
rect 392584 587862 392636 587868
rect 384304 574048 384356 574054
rect 384304 573990 384356 573996
rect 383016 572212 383068 572218
rect 383016 572154 383068 572160
rect 383028 559570 383056 572154
rect 383016 559564 383068 559570
rect 383016 559506 383068 559512
rect 384316 556646 384344 573990
rect 387616 559564 387668 559570
rect 387616 559506 387668 559512
rect 384304 556640 384356 556646
rect 384304 556582 384356 556588
rect 385040 556640 385092 556646
rect 385040 556582 385092 556588
rect 385052 554402 385080 556582
rect 385040 554396 385092 554402
rect 385040 554338 385092 554344
rect 387156 554396 387208 554402
rect 387156 554338 387208 554344
rect 383016 553376 383068 553382
rect 383016 553318 383068 553324
rect 383028 536654 383056 553318
rect 383016 536648 383068 536654
rect 383016 536590 383068 536596
rect 384120 536648 384172 536654
rect 384120 536590 384172 536596
rect 383016 533588 383068 533594
rect 383016 533530 383068 533536
rect 383028 516118 383056 533530
rect 384132 532778 384160 536590
rect 387064 534132 387116 534138
rect 387064 534074 387116 534080
rect 384120 532772 384172 532778
rect 384120 532714 384172 532720
rect 385776 529576 385828 529582
rect 385776 529518 385828 529524
rect 385684 524476 385736 524482
rect 385684 524418 385736 524424
rect 383016 516112 383068 516118
rect 383016 516054 383068 516060
rect 384948 516112 385000 516118
rect 384948 516054 385000 516060
rect 384304 513596 384356 513602
rect 384304 513538 384356 513544
rect 383016 489864 383068 489870
rect 383016 489806 383068 489812
rect 383028 460902 383056 489806
rect 383016 460896 383068 460902
rect 383016 460838 383068 460844
rect 383014 439648 383070 439657
rect 383014 439583 383070 439592
rect 382924 418804 382976 418810
rect 382924 418746 382976 418752
rect 381544 414724 381596 414730
rect 381544 414666 381596 414672
rect 382278 407824 382334 407833
rect 382278 407759 382334 407768
rect 382292 407182 382320 407759
rect 382280 407176 382332 407182
rect 382280 407118 382332 407124
rect 380164 405000 380216 405006
rect 380164 404942 380216 404948
rect 3514 397488 3570 397497
rect 3514 397423 3570 397432
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 215558 3464 371311
rect 3528 253978 3556 397423
rect 382278 397216 382334 397225
rect 382278 397151 382334 397160
rect 382292 396098 382320 397151
rect 382280 396092 382332 396098
rect 382280 396034 382332 396040
rect 382278 386608 382334 386617
rect 382278 386543 382334 386552
rect 382292 386442 382320 386543
rect 382280 386436 382332 386442
rect 382280 386378 382332 386384
rect 382278 376000 382334 376009
rect 382278 375935 382334 375944
rect 382292 375426 382320 375935
rect 382280 375420 382332 375426
rect 382280 375362 382332 375368
rect 383028 365702 383056 439583
rect 383106 429040 383162 429049
rect 383106 428975 383162 428984
rect 383016 365696 383068 365702
rect 383016 365638 383068 365644
rect 382646 365392 382702 365401
rect 382646 365327 382702 365336
rect 382660 363662 382688 365327
rect 383120 364274 383148 428975
rect 383198 418432 383254 418441
rect 383198 418367 383254 418376
rect 383212 364342 383240 418367
rect 384316 368490 384344 513538
rect 384960 513346 384988 516054
rect 384960 513318 385080 513346
rect 385052 510542 385080 513318
rect 385040 510536 385092 510542
rect 385040 510478 385092 510484
rect 384764 470552 384816 470558
rect 384764 470494 384816 470500
rect 384776 468178 384804 470494
rect 385040 469192 385092 469198
rect 385040 469134 385092 469140
rect 384764 468172 384816 468178
rect 384764 468114 384816 468120
rect 385052 466478 385080 469134
rect 385040 466472 385092 466478
rect 385040 466414 385092 466420
rect 384580 460896 384632 460902
rect 384580 460838 384632 460844
rect 384592 458250 384620 460838
rect 384580 458244 384632 458250
rect 384580 458186 384632 458192
rect 385696 369850 385724 524418
rect 385788 510610 385816 529518
rect 385776 510604 385828 510610
rect 385776 510546 385828 510552
rect 386604 414724 386656 414730
rect 386604 414666 386656 414672
rect 386616 410582 386644 414666
rect 386604 410576 386656 410582
rect 386604 410518 386656 410524
rect 385684 369844 385736 369850
rect 385684 369786 385736 369792
rect 387076 369782 387104 534074
rect 387168 518090 387196 554338
rect 387628 552702 387656 559506
rect 391204 556232 391256 556238
rect 391204 556174 391256 556180
rect 387616 552696 387668 552702
rect 387616 552638 387668 552644
rect 389916 552696 389968 552702
rect 389916 552638 389968 552644
rect 389824 545148 389876 545154
rect 389824 545090 389876 545096
rect 389180 537532 389232 537538
rect 389180 537474 389232 537480
rect 389192 535838 389220 537474
rect 389180 535832 389232 535838
rect 389180 535774 389232 535780
rect 389180 532704 389232 532710
rect 389180 532646 389232 532652
rect 389192 529990 389220 532646
rect 389180 529984 389232 529990
rect 389180 529926 389232 529932
rect 387156 518084 387208 518090
rect 387156 518026 387208 518032
rect 387156 510604 387208 510610
rect 387156 510546 387208 510552
rect 387168 500954 387196 510546
rect 388076 510536 388128 510542
rect 388076 510478 388128 510484
rect 388088 504694 388116 510478
rect 388076 504688 388128 504694
rect 388076 504630 388128 504636
rect 389180 504688 389232 504694
rect 389180 504630 389232 504636
rect 389192 502314 389220 504630
rect 389180 502308 389232 502314
rect 389180 502250 389232 502256
rect 387156 500948 387208 500954
rect 387156 500890 387208 500896
rect 387156 468172 387208 468178
rect 387156 468114 387208 468120
rect 387168 449614 387196 468114
rect 388168 466404 388220 466410
rect 388168 466346 388220 466352
rect 388180 463758 388208 466346
rect 388168 463752 388220 463758
rect 388168 463694 388220 463700
rect 387708 458176 387760 458182
rect 387708 458118 387760 458124
rect 387720 455410 387748 458118
rect 387720 455382 387840 455410
rect 387812 452606 387840 455382
rect 387800 452600 387852 452606
rect 387800 452542 387852 452548
rect 387156 449608 387208 449614
rect 387156 449550 387208 449556
rect 389836 371210 389864 545090
rect 389928 543726 389956 552638
rect 389916 543720 389968 543726
rect 389916 543662 389968 543668
rect 389916 500948 389968 500954
rect 389916 500890 389968 500896
rect 389928 477562 389956 500890
rect 389916 477556 389968 477562
rect 389916 477498 389968 477504
rect 389916 452600 389968 452606
rect 389916 452542 389968 452548
rect 389928 448594 389956 452542
rect 390284 449608 390336 449614
rect 390284 449550 390336 449556
rect 389916 448588 389968 448594
rect 389916 448530 389968 448536
rect 390296 447166 390324 449550
rect 390284 447160 390336 447166
rect 390284 447102 390336 447108
rect 389916 405000 389968 405006
rect 389916 404942 389968 404948
rect 389928 385694 389956 404942
rect 389916 385688 389968 385694
rect 389916 385630 389968 385636
rect 389824 371204 389876 371210
rect 389824 371146 389876 371152
rect 391216 371142 391244 556174
rect 391940 535832 391992 535838
rect 391940 535774 391992 535780
rect 391952 534070 391980 535774
rect 391940 534064 391992 534070
rect 391940 534006 391992 534012
rect 391940 518084 391992 518090
rect 391940 518026 391992 518032
rect 391952 516118 391980 518026
rect 391940 516112 391992 516118
rect 391940 516054 391992 516060
rect 391940 463684 391992 463690
rect 391940 463626 391992 463632
rect 391952 461650 391980 463626
rect 391940 461644 391992 461650
rect 391940 461586 391992 461592
rect 391296 448588 391348 448594
rect 391296 448530 391348 448536
rect 391308 440298 391336 448530
rect 391296 440292 391348 440298
rect 391296 440234 391348 440240
rect 392596 372570 392624 587862
rect 392676 502308 392728 502314
rect 392676 502250 392728 502256
rect 392688 488918 392716 502250
rect 392676 488912 392728 488918
rect 392676 488854 392728 488860
rect 392676 440292 392728 440298
rect 392676 440234 392728 440240
rect 392688 416090 392716 440234
rect 392676 416084 392728 416090
rect 392676 416026 392728 416032
rect 393976 373998 394004 608602
rect 394056 543720 394108 543726
rect 394056 543662 394108 543668
rect 394068 531282 394096 543662
rect 394884 534064 394936 534070
rect 394884 534006 394936 534012
rect 394056 531276 394108 531282
rect 394056 531218 394108 531224
rect 394896 529922 394924 534006
rect 394056 529916 394108 529922
rect 394056 529858 394108 529864
rect 394884 529916 394936 529922
rect 394884 529858 394936 529864
rect 394068 518022 394096 529858
rect 394056 518016 394108 518022
rect 394056 517958 394108 517964
rect 394700 518016 394752 518022
rect 394700 517958 394752 517964
rect 394712 510610 394740 517958
rect 395068 516112 395120 516118
rect 395068 516054 395120 516060
rect 395080 513398 395108 516054
rect 395068 513392 395120 513398
rect 395068 513334 395120 513340
rect 394700 510604 394752 510610
rect 394700 510546 394752 510552
rect 394608 477488 394660 477494
rect 394608 477430 394660 477436
rect 394620 476082 394648 477430
rect 394620 476054 394740 476082
rect 394712 473414 394740 476054
rect 394700 473408 394752 473414
rect 394700 473350 394752 473356
rect 395160 447092 395212 447098
rect 395160 447034 395212 447040
rect 395172 444378 395200 447034
rect 395160 444372 395212 444378
rect 395160 444314 395212 444320
rect 395356 375358 395384 629274
rect 395620 488912 395672 488918
rect 395620 488854 395672 488860
rect 395632 485654 395660 488854
rect 395620 485648 395672 485654
rect 395620 485590 395672 485596
rect 395344 375352 395396 375358
rect 395344 375294 395396 375300
rect 396736 375290 396764 651374
rect 399484 619676 399536 619682
rect 399484 619618 399536 619624
rect 396816 531276 396868 531282
rect 396816 531218 396868 531224
rect 396828 514826 396856 531218
rect 397092 529916 397144 529922
rect 397092 529858 397144 529864
rect 397104 524498 397132 529858
rect 397104 524470 397500 524498
rect 397472 521626 397500 524470
rect 397460 521620 397512 521626
rect 397460 521562 397512 521568
rect 396816 514820 396868 514826
rect 396816 514762 396868 514768
rect 397184 510604 397236 510610
rect 397184 510546 397236 510552
rect 397196 509250 397224 510546
rect 397184 509244 397236 509250
rect 397184 509186 397236 509192
rect 398104 416084 398156 416090
rect 398104 416026 398156 416032
rect 398116 411806 398144 416026
rect 398104 411800 398156 411806
rect 398104 411742 398156 411748
rect 398840 411800 398892 411806
rect 398840 411742 398892 411748
rect 398852 405686 398880 411742
rect 398840 405680 398892 405686
rect 398840 405622 398892 405628
rect 398104 385688 398156 385694
rect 398104 385630 398156 385636
rect 398116 379506 398144 385630
rect 398104 379500 398156 379506
rect 398104 379442 398156 379448
rect 396724 375284 396776 375290
rect 396724 375226 396776 375232
rect 393964 373992 394016 373998
rect 393964 373934 394016 373940
rect 399496 373930 399524 619618
rect 402244 521620 402296 521626
rect 402244 521562 402296 521568
rect 400220 514752 400272 514758
rect 400220 514694 400272 514700
rect 399576 513392 399628 513398
rect 399576 513334 399628 513340
rect 399588 497214 399616 513334
rect 400232 510610 400260 514694
rect 400220 510604 400272 510610
rect 400220 510546 400272 510552
rect 402152 510604 402204 510610
rect 402152 510546 402204 510552
rect 402164 503742 402192 510546
rect 402152 503736 402204 503742
rect 402152 503678 402204 503684
rect 399576 497208 399628 497214
rect 399576 497150 399628 497156
rect 400864 497208 400916 497214
rect 400864 497150 400916 497156
rect 400220 485648 400272 485654
rect 400220 485590 400272 485596
rect 400232 480282 400260 485590
rect 400876 485110 400904 497150
rect 400864 485104 400916 485110
rect 400864 485046 400916 485052
rect 402256 484362 402284 521562
rect 402244 484356 402296 484362
rect 402244 484298 402296 484304
rect 400220 480276 400272 480282
rect 400220 480218 400272 480224
rect 401508 473340 401560 473346
rect 401508 473282 401560 473288
rect 401520 470594 401548 473282
rect 401520 470566 401640 470594
rect 401612 467838 401640 470566
rect 401600 467832 401652 467838
rect 401600 467774 401652 467780
rect 400772 461644 400824 461650
rect 400772 461586 400824 461592
rect 400784 460290 400812 461586
rect 400772 460284 400824 460290
rect 400772 460226 400824 460232
rect 400864 459604 400916 459610
rect 400864 459546 400916 459552
rect 399576 449948 399628 449954
rect 399576 449890 399628 449896
rect 399484 373924 399536 373930
rect 399484 373866 399536 373872
rect 392584 372564 392636 372570
rect 392584 372506 392636 372512
rect 391204 371136 391256 371142
rect 391204 371078 391256 371084
rect 387064 369776 387116 369782
rect 387064 369718 387116 369724
rect 384304 368484 384356 368490
rect 384304 368426 384356 368432
rect 399588 365634 399616 449890
rect 399576 365628 399628 365634
rect 399576 365570 399628 365576
rect 400876 365566 400904 459546
rect 402244 444372 402296 444378
rect 402244 444314 402296 444320
rect 402256 429146 402284 444314
rect 402244 429140 402296 429146
rect 402244 429082 402296 429088
rect 401508 405680 401560 405686
rect 401508 405622 401560 405628
rect 401520 401674 401548 405622
rect 401508 401668 401560 401674
rect 401508 401610 401560 401616
rect 403636 376650 403664 661030
rect 406384 597576 406436 597582
rect 406384 597518 406436 597524
rect 403992 509244 404044 509250
rect 403992 509186 404044 509192
rect 404004 502314 404032 509186
rect 404728 503668 404780 503674
rect 404728 503610 404780 503616
rect 403992 502308 404044 502314
rect 403992 502250 404044 502256
rect 404740 500954 404768 503610
rect 405004 502308 405056 502314
rect 405004 502250 405056 502256
rect 404728 500948 404780 500954
rect 404728 500890 404780 500896
rect 405016 492658 405044 502250
rect 405004 492652 405056 492658
rect 405004 492594 405056 492600
rect 403716 484356 403768 484362
rect 403716 484298 403768 484304
rect 403728 458250 403756 484298
rect 403900 480208 403952 480214
rect 403900 480150 403952 480156
rect 403912 476134 403940 480150
rect 403900 476128 403952 476134
rect 403900 476070 403952 476076
rect 403808 467832 403860 467838
rect 403808 467774 403860 467780
rect 403716 458244 403768 458250
rect 403716 458186 403768 458192
rect 403820 454034 403848 467774
rect 404268 460284 404320 460290
rect 404268 460226 404320 460232
rect 404280 458522 404308 460226
rect 404268 458516 404320 458522
rect 404268 458458 404320 458464
rect 405924 458516 405976 458522
rect 405924 458458 405976 458464
rect 405936 456822 405964 458458
rect 405924 456816 405976 456822
rect 405924 456758 405976 456764
rect 403808 454028 403860 454034
rect 403808 453970 403860 453976
rect 404912 429140 404964 429146
rect 404912 429082 404964 429088
rect 404924 423638 404952 429082
rect 404912 423632 404964 423638
rect 404912 423574 404964 423580
rect 403716 410576 403768 410582
rect 403716 410518 403768 410524
rect 403728 388958 403756 410518
rect 405004 401600 405056 401606
rect 405004 401542 405056 401548
rect 403716 388952 403768 388958
rect 403716 388894 403768 388900
rect 405016 382430 405044 401542
rect 405004 382424 405056 382430
rect 405004 382366 405056 382372
rect 403716 379500 403768 379506
rect 403716 379442 403768 379448
rect 403624 376644 403676 376650
rect 403624 376586 403676 376592
rect 403728 369578 403756 379442
rect 406396 372502 406424 597518
rect 407764 565140 407816 565146
rect 407764 565082 407816 565088
rect 406568 500948 406620 500954
rect 406568 500890 406620 500896
rect 406476 476060 406528 476066
rect 406476 476002 406528 476008
rect 406488 440298 406516 476002
rect 406580 466478 406608 500890
rect 406752 492652 406804 492658
rect 406752 492594 406804 492600
rect 406660 485104 406712 485110
rect 406660 485046 406712 485052
rect 406568 466472 406620 466478
rect 406568 466414 406620 466420
rect 406672 465050 406700 485046
rect 406764 484362 406792 492594
rect 406752 484356 406804 484362
rect 406752 484298 406804 484304
rect 406660 465044 406712 465050
rect 406660 464986 406712 464992
rect 406568 454028 406620 454034
rect 406568 453970 406620 453976
rect 406476 440292 406528 440298
rect 406476 440234 406528 440240
rect 406580 439142 406608 453970
rect 406568 439136 406620 439142
rect 406568 439078 406620 439084
rect 407028 423632 407080 423638
rect 407028 423574 407080 423580
rect 407040 422294 407068 423574
rect 407040 422266 407160 422294
rect 407132 418674 407160 422266
rect 407120 418668 407172 418674
rect 407120 418610 407172 418616
rect 406476 388952 406528 388958
rect 406476 388894 406528 388900
rect 406488 376718 406516 388894
rect 406476 376712 406528 376718
rect 406476 376654 406528 376660
rect 406384 372496 406436 372502
rect 406384 372438 406436 372444
rect 407776 371074 407804 565082
rect 410524 502376 410576 502382
rect 410524 502318 410576 502324
rect 407856 484356 407908 484362
rect 407856 484298 407908 484304
rect 407868 463690 407896 484298
rect 408500 466404 408552 466410
rect 408500 466346 408552 466352
rect 407948 465044 408000 465050
rect 407948 464986 408000 464992
rect 407856 463684 407908 463690
rect 407856 463626 407908 463632
rect 407856 458176 407908 458182
rect 407856 458118 407908 458124
rect 407868 456142 407896 458118
rect 407856 456136 407908 456142
rect 407856 456078 407908 456084
rect 407960 448594 407988 464986
rect 408512 463758 408540 466346
rect 408500 463752 408552 463758
rect 408500 463694 408552 463700
rect 409328 463684 409380 463690
rect 409328 463626 409380 463632
rect 409340 458250 409368 463626
rect 409328 458244 409380 458250
rect 409328 458186 409380 458192
rect 407948 448588 408000 448594
rect 407948 448530 408000 448536
rect 409144 440224 409196 440230
rect 409144 440166 409196 440172
rect 408684 439136 408736 439142
rect 408684 439078 408736 439084
rect 408696 436830 408724 439078
rect 408684 436824 408736 436830
rect 408684 436766 408736 436772
rect 409156 428534 409184 440166
rect 409144 428528 409196 428534
rect 409144 428470 409196 428476
rect 408868 418668 408920 418674
rect 408868 418610 408920 418616
rect 408880 416770 408908 418610
rect 408868 416764 408920 416770
rect 408868 416706 408920 416712
rect 408408 382424 408460 382430
rect 408408 382366 408460 382372
rect 408420 378026 408448 382366
rect 408420 377998 408540 378026
rect 408512 376582 408540 377998
rect 408500 376576 408552 376582
rect 408500 376518 408552 376524
rect 407764 371068 407816 371074
rect 407764 371010 407816 371016
rect 403716 369572 403768 369578
rect 403716 369514 403768 369520
rect 409144 369572 409196 369578
rect 409144 369514 409196 369520
rect 400864 365560 400916 365566
rect 400864 365502 400916 365508
rect 383200 364336 383252 364342
rect 383200 364278 383252 364284
rect 383108 364268 383160 364274
rect 383108 364210 383160 364216
rect 382648 363656 382700 363662
rect 382648 363598 382700 363604
rect 409156 360806 409184 369514
rect 410536 368422 410564 502318
rect 411904 492720 411956 492726
rect 411904 492662 411956 492668
rect 410616 458244 410668 458250
rect 410616 458186 410668 458192
rect 410628 445738 410656 458186
rect 410800 456748 410852 456754
rect 410800 456690 410852 456696
rect 410812 448526 410840 456690
rect 410708 448520 410760 448526
rect 410708 448462 410760 448468
rect 410800 448520 410852 448526
rect 410800 448462 410852 448468
rect 410616 445732 410668 445738
rect 410616 445674 410668 445680
rect 410720 436966 410748 448462
rect 411260 445732 411312 445738
rect 411260 445674 411312 445680
rect 411272 441862 411300 445674
rect 411260 441856 411312 441862
rect 411260 441798 411312 441804
rect 410708 436960 410760 436966
rect 410708 436902 410760 436908
rect 410616 436824 410668 436830
rect 410616 436766 410668 436772
rect 410628 424386 410656 436766
rect 410616 424380 410668 424386
rect 410616 424322 410668 424328
rect 410616 416764 410668 416770
rect 410616 416706 410668 416712
rect 410628 409358 410656 416706
rect 410616 409352 410668 409358
rect 410616 409294 410668 409300
rect 410524 368416 410576 368422
rect 410524 368358 410576 368364
rect 411916 368354 411944 492662
rect 412088 463684 412140 463690
rect 412088 463626 412140 463632
rect 411996 456136 412048 456142
rect 411996 456078 412048 456084
rect 412008 443018 412036 456078
rect 411996 443012 412048 443018
rect 411996 442954 412048 442960
rect 411996 436960 412048 436966
rect 411996 436902 412048 436908
rect 412008 430642 412036 436902
rect 411996 430636 412048 430642
rect 411996 430578 412048 430584
rect 411996 428528 412048 428534
rect 411996 428470 412048 428476
rect 412008 391950 412036 428470
rect 412100 426426 412128 463626
rect 412088 426420 412140 426426
rect 412088 426362 412140 426368
rect 412088 409352 412140 409358
rect 412088 409294 412140 409300
rect 412100 400178 412128 409294
rect 412088 400172 412140 400178
rect 412088 400114 412140 400120
rect 411996 391944 412048 391950
rect 411996 391886 412048 391892
rect 411996 376712 412048 376718
rect 411996 376654 412048 376660
rect 411904 368348 411956 368354
rect 411904 368290 411956 368296
rect 409144 360800 409196 360806
rect 409144 360742 409196 360748
rect 411904 360800 411956 360806
rect 411904 360742 411956 360748
rect 3606 358456 3662 358465
rect 3606 358391 3662 358400
rect 3620 302122 3648 358391
rect 382922 354784 382978 354793
rect 382922 354719 382978 354728
rect 3698 345400 3754 345409
rect 3698 345335 3754 345344
rect 3608 302116 3660 302122
rect 3608 302058 3660 302064
rect 3606 293176 3662 293185
rect 3606 293111 3662 293120
rect 3516 253972 3568 253978
rect 3516 253914 3568 253920
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3424 215552 3476 215558
rect 3424 215494 3476 215500
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3436 102202 3464 214911
rect 3528 138378 3556 241023
rect 3620 187746 3648 293111
rect 3712 266694 3740 345335
rect 382278 344176 382334 344185
rect 382278 344111 382334 344120
rect 382292 343738 382320 344111
rect 382280 343732 382332 343738
rect 382280 343674 382332 343680
rect 382936 343602 382964 354719
rect 411916 354006 411944 360742
rect 411904 354000 411956 354006
rect 411904 353942 411956 353948
rect 407028 345092 407080 345098
rect 407028 345034 407080 345040
rect 386328 343732 386380 343738
rect 386328 343674 386380 343680
rect 382924 343596 382976 343602
rect 382924 343538 382976 343544
rect 386340 341562 386368 343674
rect 386328 341556 386380 341562
rect 386328 341498 386380 341504
rect 402152 341556 402204 341562
rect 402152 341498 402204 341504
rect 383108 338564 383160 338570
rect 383108 338506 383160 338512
rect 382924 336864 382976 336870
rect 382924 336806 382976 336812
rect 3974 319288 4030 319297
rect 3974 319223 4030 319232
rect 3882 306232 3938 306241
rect 3882 306167 3938 306176
rect 3790 267200 3846 267209
rect 3790 267135 3846 267144
rect 3700 266688 3752 266694
rect 3700 266630 3752 266636
rect 3698 254144 3754 254153
rect 3698 254079 3754 254088
rect 3608 187740 3660 187746
rect 3608 187682 3660 187688
rect 3712 150754 3740 254079
rect 3804 165578 3832 267135
rect 3896 212498 3924 306167
rect 3988 246022 4016 319223
rect 382936 312361 382964 336806
rect 383016 336796 383068 336802
rect 383016 336738 383068 336744
rect 383028 322969 383056 336738
rect 383120 333577 383148 338506
rect 402164 336954 402192 341498
rect 407040 337090 407068 345034
rect 412008 342922 412036 376654
rect 412272 376576 412324 376582
rect 412272 376518 412324 376524
rect 412284 372638 412312 376518
rect 412272 372632 412324 372638
rect 412272 372574 412324 372580
rect 411996 342916 412048 342922
rect 411996 342858 412048 342864
rect 410064 338224 410116 338230
rect 410064 338166 410116 338172
rect 406488 337062 407068 337090
rect 406488 336954 406516 337062
rect 402164 336940 402284 336954
rect 402178 336926 402284 336940
rect 406134 336926 406516 336954
rect 410076 336940 410104 338166
rect 413296 337482 413324 670006
rect 413468 448520 413520 448526
rect 413468 448462 413520 448468
rect 413376 443012 413428 443018
rect 413376 442954 413428 442960
rect 413388 418198 413416 442954
rect 413480 439414 413508 448462
rect 413560 441856 413612 441862
rect 413560 441798 413612 441804
rect 413468 439408 413520 439414
rect 413468 439350 413520 439356
rect 413572 437782 413600 441798
rect 413560 437776 413612 437782
rect 413560 437718 413612 437724
rect 413376 418192 413428 418198
rect 413376 418134 413428 418140
rect 413664 340202 413692 703520
rect 418804 700732 418856 700738
rect 418804 700674 418856 700680
rect 416044 700528 416096 700534
rect 416044 700470 416096 700476
rect 414664 481704 414716 481710
rect 414664 481646 414716 481652
rect 413928 426420 413980 426426
rect 413928 426362 413980 426368
rect 413940 423706 413968 426362
rect 413928 423700 413980 423706
rect 413928 423642 413980 423648
rect 414572 391944 414624 391950
rect 414572 391886 414624 391892
rect 414584 389230 414612 391886
rect 414572 389224 414624 389230
rect 414572 389166 414624 389172
rect 414676 367062 414704 481646
rect 415860 439408 415912 439414
rect 415860 439350 415912 439356
rect 414756 437776 414808 437782
rect 414756 437718 414808 437724
rect 414768 431118 414796 437718
rect 415872 436762 415900 439350
rect 415860 436756 415912 436762
rect 415860 436698 415912 436704
rect 414756 431112 414808 431118
rect 414756 431054 414808 431060
rect 414756 430568 414808 430574
rect 414756 430510 414808 430516
rect 414768 416770 414796 430510
rect 415952 423632 416004 423638
rect 415952 423574 416004 423580
rect 415964 419558 415992 423574
rect 415952 419552 416004 419558
rect 415952 419494 416004 419500
rect 414756 416764 414808 416770
rect 414756 416706 414808 416712
rect 415308 400172 415360 400178
rect 415308 400114 415360 400120
rect 415320 398834 415348 400114
rect 415320 398806 415440 398834
rect 415412 394670 415440 398806
rect 415400 394664 415452 394670
rect 415400 394606 415452 394612
rect 415124 372632 415176 372638
rect 415124 372574 415176 372580
rect 415136 368286 415164 372574
rect 415124 368280 415176 368286
rect 415124 368222 415176 368228
rect 414664 367056 414716 367062
rect 414664 366998 414716 367004
rect 413652 340196 413704 340202
rect 413652 340138 413704 340144
rect 414020 338292 414072 338298
rect 414020 338234 414072 338240
rect 413284 337476 413336 337482
rect 413284 337418 413336 337424
rect 414032 336940 414060 338234
rect 416056 337618 416084 700470
rect 418160 436756 418212 436762
rect 418160 436698 418212 436704
rect 418172 434722 418200 436698
rect 418160 434716 418212 434722
rect 418160 434658 418212 434664
rect 416688 431112 416740 431118
rect 416688 431054 416740 431060
rect 416700 430522 416728 431054
rect 416700 430494 416820 430522
rect 416792 427582 416820 430494
rect 416780 427576 416832 427582
rect 416780 427518 416832 427524
rect 416688 424380 416740 424386
rect 416688 424322 416740 424328
rect 416700 422294 416728 424322
rect 416700 422266 416820 422294
rect 416792 420374 416820 422266
rect 416780 420368 416832 420374
rect 416780 420310 416832 420316
rect 417424 418124 417476 418130
rect 417424 418066 417476 418072
rect 417436 394806 417464 418066
rect 417424 394800 417476 394806
rect 417424 394742 417476 394748
rect 417424 394664 417476 394670
rect 417424 394606 417476 394612
rect 417436 371550 417464 394606
rect 417516 389224 417568 389230
rect 417516 389166 417568 389172
rect 417528 376650 417556 389166
rect 417516 376644 417568 376650
rect 417516 376586 417568 376592
rect 417424 371544 417476 371550
rect 417424 371486 417476 371492
rect 418712 371544 418764 371550
rect 418712 371486 418764 371492
rect 418724 371006 418752 371486
rect 418712 371000 418764 371006
rect 418712 370942 418764 370948
rect 418160 342916 418212 342922
rect 418160 342858 418212 342864
rect 418172 340270 418200 342858
rect 418160 340264 418212 340270
rect 418160 340206 418212 340212
rect 417976 338360 418028 338366
rect 417976 338302 418028 338308
rect 416044 337612 416096 337618
rect 416044 337554 416096 337560
rect 417988 336940 418016 338302
rect 418816 337414 418844 700674
rect 418896 669996 418948 670002
rect 418896 669938 418948 669944
rect 418908 337686 418936 669938
rect 420184 667684 420236 667690
rect 420184 667626 420236 667632
rect 418988 667616 419040 667622
rect 418988 667558 419040 667564
rect 418896 337680 418948 337686
rect 418896 337622 418948 337628
rect 419000 337550 419028 667558
rect 419080 576904 419132 576910
rect 419080 576846 419132 576852
rect 419092 372434 419120 576846
rect 419172 470620 419224 470626
rect 419172 470562 419224 470568
rect 419080 372428 419132 372434
rect 419080 372370 419132 372376
rect 419184 366994 419212 470562
rect 419356 427576 419408 427582
rect 419356 427518 419408 427524
rect 419368 419762 419396 427518
rect 419448 420368 419500 420374
rect 419448 420310 419500 420316
rect 419356 419756 419408 419762
rect 419356 419698 419408 419704
rect 419460 413302 419488 420310
rect 419448 413296 419500 413302
rect 419448 413238 419500 413244
rect 419172 366988 419224 366994
rect 419172 366930 419224 366936
rect 420196 337754 420224 667626
rect 427452 447228 427504 447234
rect 427452 447170 427504 447176
rect 422484 447160 422536 447166
rect 422484 447102 422536 447108
rect 422496 444924 422524 447102
rect 427464 444924 427492 447170
rect 429856 445058 429884 703520
rect 444288 700732 444340 700738
rect 444288 700674 444340 700680
rect 444196 700528 444248 700534
rect 444196 700470 444248 700476
rect 437388 447364 437440 447370
rect 437388 447306 437440 447312
rect 432420 447296 432472 447302
rect 432420 447238 432472 447244
rect 429844 445052 429896 445058
rect 429844 444994 429896 445000
rect 432432 444924 432460 447238
rect 437400 444924 437428 447306
rect 442632 444440 442684 444446
rect 442382 444388 442632 444394
rect 442382 444382 442684 444388
rect 442382 444366 442672 444382
rect 420276 434716 420328 434722
rect 420276 434658 420328 434664
rect 420288 418130 420316 434658
rect 421498 420022 421880 420050
rect 421656 419756 421708 419762
rect 421656 419698 421708 419704
rect 420920 419552 420972 419558
rect 420920 419494 420972 419500
rect 420276 418124 420328 418130
rect 420276 418066 420328 418072
rect 420932 413030 420960 419494
rect 421564 416764 421616 416770
rect 421564 416706 421616 416712
rect 420920 413024 420972 413030
rect 420920 412966 420972 412972
rect 421576 404598 421604 416706
rect 421668 411602 421696 419698
rect 421852 416362 421880 420022
rect 421840 416356 421892 416362
rect 421840 416298 421892 416304
rect 421656 411596 421708 411602
rect 421656 411538 421708 411544
rect 421564 404592 421616 404598
rect 421564 404534 421616 404540
rect 421564 394664 421616 394670
rect 421564 394606 421616 394612
rect 420736 376644 420788 376650
rect 420736 376586 420788 376592
rect 420748 371006 420776 376586
rect 421576 371958 421604 394606
rect 421564 371952 421616 371958
rect 421564 371894 421616 371900
rect 420276 371000 420328 371006
rect 420276 370942 420328 370948
rect 420736 371000 420788 371006
rect 420736 370942 420788 370948
rect 420288 362982 420316 370942
rect 420920 368280 420972 368286
rect 420920 368222 420972 368228
rect 420932 365022 420960 368222
rect 420920 365016 420972 365022
rect 420920 364958 420972 364964
rect 420276 362976 420328 362982
rect 420276 362918 420328 362924
rect 421564 362976 421616 362982
rect 421564 362918 421616 362924
rect 421576 350538 421604 362918
rect 421564 350532 421616 350538
rect 421564 350474 421616 350480
rect 422128 347750 422156 420036
rect 422786 420022 423168 420050
rect 423430 420022 423536 420050
rect 423140 416362 423168 420022
rect 422208 416356 422260 416362
rect 422208 416298 422260 416304
rect 423128 416356 423180 416362
rect 423128 416298 423180 416304
rect 422116 347744 422168 347750
rect 422116 347686 422168 347692
rect 422220 347682 422248 416298
rect 422944 371952 422996 371958
rect 422944 371894 422996 371900
rect 422956 350878 422984 371894
rect 423312 371000 423364 371006
rect 423312 370942 423364 370948
rect 423324 368626 423352 370942
rect 423312 368620 423364 368626
rect 423312 368562 423364 368568
rect 423508 354226 423536 420022
rect 424060 417450 424088 420036
rect 424718 420022 425008 420050
rect 425362 420022 425928 420050
rect 426006 420022 426388 420050
rect 424324 418124 424376 418130
rect 424324 418066 424376 418072
rect 424048 417444 424100 417450
rect 424048 417386 424100 417392
rect 423588 416356 423640 416362
rect 423588 416298 423640 416304
rect 423324 354198 423536 354226
rect 422944 350872 422996 350878
rect 422944 350814 422996 350820
rect 423324 349042 423352 354198
rect 423600 354090 423628 416298
rect 423680 413024 423732 413030
rect 423680 412966 423732 412972
rect 423692 408542 423720 412966
rect 424336 411806 424364 418066
rect 424324 411800 424376 411806
rect 424324 411742 424376 411748
rect 424416 411596 424468 411602
rect 424416 411538 424468 411544
rect 423680 408536 423732 408542
rect 423680 408478 423732 408484
rect 424324 404592 424376 404598
rect 424324 404534 424376 404540
rect 424336 383110 424364 404534
rect 424428 390862 424456 411538
rect 424416 390856 424468 390862
rect 424416 390798 424468 390804
rect 424324 383104 424376 383110
rect 424324 383046 424376 383052
rect 424324 368620 424376 368626
rect 424324 368562 424376 368568
rect 424336 358698 424364 368562
rect 424324 358692 424376 358698
rect 424324 358634 424376 358640
rect 423508 354062 423628 354090
rect 423312 349036 423364 349042
rect 423312 348978 423364 348984
rect 422208 347676 422260 347682
rect 422208 347618 422260 347624
rect 423508 347546 423536 354062
rect 423588 354000 423640 354006
rect 423588 353942 423640 353948
rect 423600 350946 423628 353942
rect 423588 350940 423640 350946
rect 423588 350882 423640 350888
rect 424980 350538 425008 420022
rect 425900 412634 425928 420022
rect 425900 412606 426296 412634
rect 425796 411800 425848 411806
rect 425796 411742 425848 411748
rect 425808 408406 425836 411742
rect 425796 408400 425848 408406
rect 425796 408342 425848 408348
rect 425796 390856 425848 390862
rect 425796 390798 425848 390804
rect 425704 383104 425756 383110
rect 425704 383046 425756 383052
rect 425716 358766 425744 383046
rect 425808 371550 425836 390798
rect 425796 371544 425848 371550
rect 425796 371486 425848 371492
rect 425796 365016 425848 365022
rect 425796 364958 425848 364964
rect 425808 359514 425836 364958
rect 425796 359508 425848 359514
rect 425796 359450 425848 359456
rect 425704 358760 425756 358766
rect 425704 358702 425756 358708
rect 425704 350872 425756 350878
rect 425704 350814 425756 350820
rect 423588 350532 423640 350538
rect 423588 350474 423640 350480
rect 424968 350532 425020 350538
rect 424968 350474 425020 350480
rect 423496 347540 423548 347546
rect 423496 347482 423548 347488
rect 423600 345014 423628 350474
rect 423600 344986 423720 345014
rect 423692 344214 423720 344986
rect 423680 344208 423732 344214
rect 423680 344150 423732 344156
rect 425716 343942 425744 350814
rect 426268 350266 426296 412606
rect 426360 350402 426388 420022
rect 439504 418804 439556 418810
rect 439504 418746 439556 418752
rect 428464 413296 428516 413302
rect 428464 413238 428516 413244
rect 427084 408400 427136 408406
rect 427084 408342 427136 408348
rect 427096 387870 427124 408342
rect 427084 387864 427136 387870
rect 427084 387806 427136 387812
rect 428476 381070 428504 413238
rect 428556 408468 428608 408474
rect 428556 408410 428608 408416
rect 428464 381064 428516 381070
rect 428464 381006 428516 381012
rect 428568 381002 428596 408410
rect 435364 407176 435416 407182
rect 435364 407118 435416 407124
rect 429844 387796 429896 387802
rect 429844 387738 429896 387744
rect 428556 380996 428608 381002
rect 428556 380938 428608 380944
rect 427084 371544 427136 371550
rect 427084 371486 427136 371492
rect 426440 358692 426492 358698
rect 426440 358634 426492 358640
rect 426452 354754 426480 358634
rect 426440 354748 426492 354754
rect 426440 354690 426492 354696
rect 426348 350396 426400 350402
rect 426348 350338 426400 350344
rect 426256 350260 426308 350266
rect 426256 350202 426308 350208
rect 427096 346458 427124 371486
rect 429856 360806 429884 387738
rect 431224 381064 431276 381070
rect 431224 381006 431276 381012
rect 429936 380996 429988 381002
rect 429936 380938 429988 380944
rect 429948 373182 429976 380938
rect 429936 373176 429988 373182
rect 429936 373118 429988 373124
rect 430948 373176 431000 373182
rect 430948 373118 431000 373124
rect 430960 369714 430988 373118
rect 430948 369708 431000 369714
rect 430948 369650 431000 369656
rect 431236 364410 431264 381006
rect 432696 369708 432748 369714
rect 432696 369650 432748 369656
rect 431224 364404 431276 364410
rect 431224 364346 431276 364352
rect 432604 364404 432656 364410
rect 432604 364346 432656 364352
rect 429844 360800 429896 360806
rect 429844 360742 429896 360748
rect 431316 360800 431368 360806
rect 431316 360742 431368 360748
rect 427268 359508 427320 359514
rect 427268 359450 427320 359456
rect 427176 358760 427228 358766
rect 427176 358702 427228 358708
rect 427188 349110 427216 358702
rect 427280 350334 427308 359450
rect 430580 354680 430632 354686
rect 430580 354622 430632 354628
rect 430592 351898 430620 354622
rect 430580 351892 430632 351898
rect 430580 351834 430632 351840
rect 431224 350940 431276 350946
rect 431224 350882 431276 350888
rect 427268 350328 427320 350334
rect 427268 350270 427320 350276
rect 428556 350328 428608 350334
rect 428556 350270 428608 350276
rect 427176 349104 427228 349110
rect 427176 349046 427228 349052
rect 428464 349104 428516 349110
rect 428464 349046 428516 349052
rect 427084 346452 427136 346458
rect 427084 346394 427136 346400
rect 426348 344208 426400 344214
rect 426348 344150 426400 344156
rect 425704 343936 425756 343942
rect 425704 343878 425756 343884
rect 426360 343534 426388 344150
rect 427728 343936 427780 343942
rect 427728 343878 427780 343884
rect 426348 343528 426400 343534
rect 426348 343470 426400 343476
rect 427740 340882 427768 343878
rect 428476 342310 428504 349046
rect 428568 347614 428596 350270
rect 428556 347608 428608 347614
rect 428556 347550 428608 347556
rect 429568 347608 429620 347614
rect 429568 347550 429620 347556
rect 429108 343528 429160 343534
rect 429108 343470 429160 343476
rect 428464 342304 428516 342310
rect 428464 342246 428516 342252
rect 427728 340876 427780 340882
rect 427728 340818 427780 340824
rect 429120 339402 429148 343470
rect 429580 339454 429608 347550
rect 430580 346384 430632 346390
rect 430580 346326 430632 346332
rect 430592 340814 430620 346326
rect 430672 340876 430724 340882
rect 430672 340818 430724 340824
rect 430580 340808 430632 340814
rect 430580 340750 430632 340756
rect 429568 339448 429620 339454
rect 429120 339374 429240 339402
rect 429568 339390 429620 339396
rect 425888 338428 425940 338434
rect 425888 338370 425940 338376
rect 420184 337748 420236 337754
rect 420184 337690 420236 337696
rect 418988 337544 419040 337550
rect 418988 337486 419040 337492
rect 418804 337408 418856 337414
rect 418804 337350 418856 337356
rect 425900 336940 425928 338370
rect 402256 336734 402284 336926
rect 422206 336832 422262 336841
rect 421958 336790 422206 336818
rect 422206 336767 422262 336776
rect 402244 336728 402296 336734
rect 402244 336670 402296 336676
rect 429212 336666 429240 339374
rect 429844 338496 429896 338502
rect 429844 338438 429896 338444
rect 429856 336940 429884 338438
rect 430684 336938 430712 340818
rect 430672 336932 430724 336938
rect 430672 336874 430724 336880
rect 429200 336660 429252 336666
rect 429200 336602 429252 336608
rect 383106 333568 383162 333577
rect 383106 333503 383162 333512
rect 431236 329118 431264 350882
rect 431328 350470 431356 360742
rect 432616 354278 432644 364346
rect 432604 354272 432656 354278
rect 432604 354214 432656 354220
rect 431316 350464 431368 350470
rect 431316 350406 431368 350412
rect 431868 336660 431920 336666
rect 431868 336602 431920 336608
rect 431880 335102 431908 336602
rect 431868 335096 431920 335102
rect 431868 335038 431920 335044
rect 432604 332648 432656 332654
rect 432604 332590 432656 332596
rect 431224 329112 431276 329118
rect 431224 329054 431276 329060
rect 383014 322960 383070 322969
rect 383014 322895 383070 322904
rect 382922 312352 382978 312361
rect 382922 312287 382978 312296
rect 406476 305992 406528 305998
rect 406476 305934 406528 305940
rect 406750 305960 406806 305969
rect 383292 305924 383344 305930
rect 383292 305866 383344 305872
rect 380164 305720 380216 305726
rect 380164 305662 380216 305668
rect 4896 302116 4948 302122
rect 4896 302058 4948 302064
rect 3976 246016 4028 246022
rect 3976 245958 4028 245964
rect 3884 212492 3936 212498
rect 3884 212434 3936 212440
rect 3882 201920 3938 201929
rect 3882 201855 3938 201864
rect 3792 165572 3844 165578
rect 3792 165514 3844 165520
rect 3790 162888 3846 162897
rect 3790 162823 3846 162832
rect 3700 150748 3752 150754
rect 3700 150690 3752 150696
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 3516 138372 3568 138378
rect 3516 138314 3568 138320
rect 3514 110664 3570 110673
rect 3514 110599 3570 110608
rect 3424 102196 3476 102202
rect 3424 102138 3476 102144
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3436 96694 3464 97543
rect 3424 96688 3476 96694
rect 3424 96630 3476 96636
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3344 84250 3372 84623
rect 3332 84244 3384 84250
rect 3332 84186 3384 84192
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3436 52086 3464 71567
rect 3424 52080 3476 52086
rect 3424 52022 3476 52028
rect 3528 52018 3556 110599
rect 3620 70174 3648 149767
rect 3698 136776 3754 136785
rect 3698 136711 3754 136720
rect 3712 90370 3740 136711
rect 3700 90364 3752 90370
rect 3700 90306 3752 90312
rect 3804 89758 3832 162823
rect 3896 101590 3924 201855
rect 3974 188864 4030 188873
rect 3974 188799 4030 188808
rect 3988 115938 4016 188799
rect 4908 188086 4936 302058
rect 5264 266688 5316 266694
rect 5264 266630 5316 266636
rect 5172 253972 5224 253978
rect 5172 253914 5224 253920
rect 5080 246016 5132 246022
rect 5080 245958 5132 245964
rect 4988 212492 5040 212498
rect 4988 212434 5040 212440
rect 4896 188080 4948 188086
rect 4896 188022 4948 188028
rect 4804 187740 4856 187746
rect 4804 187682 4856 187688
rect 3976 115932 4028 115938
rect 3976 115874 4028 115880
rect 3884 101584 3936 101590
rect 3884 101526 3936 101532
rect 3792 89752 3844 89758
rect 3792 89694 3844 89700
rect 3608 70168 3660 70174
rect 3608 70110 3660 70116
rect 4816 70106 4844 187682
rect 4896 165572 4948 165578
rect 4896 165514 4948 165520
rect 4908 78674 4936 165514
rect 5000 104786 5028 212434
rect 5092 140146 5120 245958
rect 5184 150482 5212 253914
rect 5276 165578 5304 266630
rect 5356 215552 5408 215558
rect 5356 215494 5408 215500
rect 5264 165572 5316 165578
rect 5264 165514 5316 165520
rect 5264 150748 5316 150754
rect 5264 150690 5316 150696
rect 5172 150476 5224 150482
rect 5172 150418 5224 150424
rect 5080 140140 5132 140146
rect 5080 140082 5132 140088
rect 5080 138372 5132 138378
rect 5080 138314 5132 138320
rect 4988 104780 5040 104786
rect 4988 104722 5040 104728
rect 4988 101584 5040 101590
rect 4988 101526 5040 101532
rect 5000 80102 5028 101526
rect 5092 83230 5120 138314
rect 5172 115932 5224 115938
rect 5172 115874 5224 115880
rect 5184 104854 5212 115874
rect 5172 104848 5224 104854
rect 5172 104790 5224 104796
rect 5172 102196 5224 102202
rect 5172 102138 5224 102144
rect 5184 91254 5212 102138
rect 5172 91248 5224 91254
rect 5172 91190 5224 91196
rect 5276 90250 5304 150690
rect 5368 115938 5396 215494
rect 6184 188080 6236 188086
rect 6184 188022 6236 188028
rect 5356 115932 5408 115938
rect 5356 115874 5408 115880
rect 6196 114646 6224 188022
rect 6276 165572 6328 165578
rect 6276 165514 6328 165520
rect 6184 114640 6236 114646
rect 6184 114582 6236 114588
rect 6288 109002 6316 165514
rect 6460 150476 6512 150482
rect 6460 150418 6512 150424
rect 6368 140140 6420 140146
rect 6368 140082 6420 140088
rect 6276 108996 6328 109002
rect 6276 108938 6328 108944
rect 6276 104848 6328 104854
rect 6276 104790 6328 104796
rect 6184 104780 6236 104786
rect 6184 104722 6236 104728
rect 5276 90222 5580 90250
rect 5448 89752 5500 89758
rect 5448 89694 5500 89700
rect 5460 86442 5488 89694
rect 5552 86630 5580 90222
rect 5540 86624 5592 86630
rect 5540 86566 5592 86572
rect 5460 86414 5580 86442
rect 5080 83224 5132 83230
rect 5080 83166 5132 83172
rect 4988 80096 5040 80102
rect 4988 80038 5040 80044
rect 4896 78668 4948 78674
rect 4896 78610 4948 78616
rect 5552 78538 5580 86414
rect 6000 83224 6052 83230
rect 6000 83166 6052 83172
rect 6012 78606 6040 83166
rect 6000 78600 6052 78606
rect 6000 78542 6052 78548
rect 5540 78532 5592 78538
rect 5540 78474 5592 78480
rect 4988 70168 5040 70174
rect 4988 70110 5040 70116
rect 4804 70100 4856 70106
rect 4804 70042 4856 70048
rect 5000 65142 5028 70110
rect 5540 70100 5592 70106
rect 5540 70042 5592 70048
rect 5552 65210 5580 70042
rect 5540 65204 5592 65210
rect 5540 65146 5592 65152
rect 4988 65136 5040 65142
rect 4988 65078 5040 65084
rect 3606 58576 3662 58585
rect 3606 58511 3662 58520
rect 3620 52057 3648 58511
rect 6196 56982 6224 104722
rect 6288 96150 6316 104790
rect 6276 96144 6328 96150
rect 6276 96086 6328 96092
rect 6276 91248 6328 91254
rect 6276 91190 6328 91196
rect 6288 75206 6316 91190
rect 6380 90982 6408 140082
rect 6472 104922 6500 150418
rect 6552 115932 6604 115938
rect 6552 115874 6604 115880
rect 6460 104916 6512 104922
rect 6460 104858 6512 104864
rect 6368 90976 6420 90982
rect 6368 90918 6420 90924
rect 6564 84318 6592 115874
rect 7748 114640 7800 114646
rect 7748 114582 7800 114588
rect 7564 108996 7616 109002
rect 7564 108938 7616 108944
rect 6552 84312 6604 84318
rect 6552 84254 6604 84260
rect 6276 75200 6328 75206
rect 6276 75142 6328 75148
rect 6920 75200 6972 75206
rect 6920 75142 6972 75148
rect 6932 72622 6960 75142
rect 6920 72616 6972 72622
rect 6920 72558 6972 72564
rect 7288 65136 7340 65142
rect 7288 65078 7340 65084
rect 7300 61062 7328 65078
rect 7288 61056 7340 61062
rect 7288 60998 7340 61004
rect 6184 56976 6236 56982
rect 6184 56918 6236 56924
rect 7576 56438 7604 108938
rect 7656 104916 7708 104922
rect 7656 104858 7708 104864
rect 7668 56574 7696 104858
rect 7760 82142 7788 114582
rect 20904 96688 20956 96694
rect 20904 96630 20956 96636
rect 8208 96144 8260 96150
rect 8208 96086 8260 96092
rect 7932 90976 7984 90982
rect 7932 90918 7984 90924
rect 7840 84312 7892 84318
rect 7840 84254 7892 84260
rect 7748 82136 7800 82142
rect 7748 82078 7800 82084
rect 7748 78668 7800 78674
rect 7748 78610 7800 78616
rect 7760 70990 7788 78610
rect 7748 70984 7800 70990
rect 7748 70926 7800 70932
rect 7748 65204 7800 65210
rect 7748 65146 7800 65152
rect 7656 56568 7708 56574
rect 7656 56510 7708 56516
rect 7564 56432 7616 56438
rect 7564 56374 7616 56380
rect 7760 53106 7788 65146
rect 7852 56506 7880 84254
rect 7944 60738 7972 90918
rect 8220 89842 8248 96086
rect 20916 93854 20944 96630
rect 20916 93826 21404 93854
rect 10968 90364 11020 90370
rect 10968 90306 11020 90312
rect 8220 89814 8340 89842
rect 8312 88330 8340 89814
rect 8300 88324 8352 88330
rect 8300 88266 8352 88272
rect 10980 88210 11008 90306
rect 11704 88324 11756 88330
rect 11704 88266 11756 88272
rect 10980 88182 11100 88210
rect 8024 86624 8076 86630
rect 8024 86566 8076 86572
rect 8036 77194 8064 86566
rect 11072 85542 11100 88182
rect 11060 85536 11112 85542
rect 11060 85478 11112 85484
rect 9128 82136 9180 82142
rect 9128 82078 9180 82084
rect 8392 80028 8444 80034
rect 8392 79970 8444 79976
rect 8036 77166 8340 77194
rect 8312 70242 8340 77166
rect 8404 75818 8432 79970
rect 8944 78600 8996 78606
rect 8944 78542 8996 78548
rect 8392 75812 8444 75818
rect 8392 75754 8444 75760
rect 8300 70236 8352 70242
rect 8300 70178 8352 70184
rect 8956 66230 8984 78542
rect 9036 78532 9088 78538
rect 9036 78474 9088 78480
rect 9048 76498 9076 78474
rect 9036 76492 9088 76498
rect 9036 76434 9088 76440
rect 9140 75886 9168 82078
rect 11716 81462 11744 88266
rect 13728 85536 13780 85542
rect 13728 85478 13780 85484
rect 11704 81456 11756 81462
rect 11704 81398 11756 81404
rect 13740 78742 13768 85478
rect 18604 84244 18656 84250
rect 18604 84186 18656 84192
rect 15844 81388 15896 81394
rect 15844 81330 15896 81336
rect 13728 78736 13780 78742
rect 13728 78678 13780 78684
rect 10968 76492 11020 76498
rect 10968 76434 11020 76440
rect 9128 75880 9180 75886
rect 9128 75822 9180 75828
rect 10324 75880 10376 75886
rect 10324 75822 10376 75828
rect 9588 72616 9640 72622
rect 9588 72558 9640 72564
rect 9404 70984 9456 70990
rect 9404 70926 9456 70932
rect 9416 67522 9444 70926
rect 9600 70394 9628 72558
rect 9600 70366 9720 70394
rect 9692 67590 9720 70366
rect 9680 67584 9732 67590
rect 9680 67526 9732 67532
rect 9404 67516 9456 67522
rect 9404 67458 9456 67464
rect 8944 66224 8996 66230
rect 8944 66166 8996 66172
rect 7944 60710 8340 60738
rect 8312 57934 8340 60710
rect 8300 57928 8352 57934
rect 8300 57870 8352 57876
rect 8208 56976 8260 56982
rect 8208 56918 8260 56924
rect 7840 56500 7892 56506
rect 7840 56442 7892 56448
rect 8220 53122 8248 56918
rect 8668 56568 8720 56574
rect 8668 56510 8720 56516
rect 8680 53174 8708 56510
rect 10336 53854 10364 75822
rect 10416 70236 10468 70242
rect 10416 70178 10468 70184
rect 10428 60790 10456 70178
rect 10980 67658 11008 76434
rect 11704 75812 11756 75818
rect 11704 75754 11756 75760
rect 10968 67652 11020 67658
rect 10968 67594 11020 67600
rect 10968 67516 11020 67522
rect 10968 67458 11020 67464
rect 10980 63306 11008 67458
rect 11716 64938 11744 75754
rect 15856 73234 15884 81330
rect 17224 78668 17276 78674
rect 17224 78610 17276 78616
rect 15844 73228 15896 73234
rect 15844 73170 15896 73176
rect 12256 67584 12308 67590
rect 12256 67526 12308 67532
rect 15108 67584 15160 67590
rect 15108 67526 15160 67532
rect 11704 64932 11756 64938
rect 11704 64874 11756 64880
rect 10968 63300 11020 63306
rect 10968 63242 11020 63248
rect 11244 61056 11296 61062
rect 11244 60998 11296 61004
rect 10416 60784 10468 60790
rect 10416 60726 10468 60732
rect 11256 56642 11284 60998
rect 12268 60722 12296 67526
rect 12348 66224 12400 66230
rect 12348 66166 12400 66172
rect 12360 62098 12388 66166
rect 15120 64954 15148 67526
rect 15120 64926 15240 64954
rect 15212 64874 15240 64926
rect 15108 64864 15160 64870
rect 15212 64846 15332 64874
rect 15108 64806 15160 64812
rect 14464 63300 14516 63306
rect 14464 63242 14516 63248
rect 12360 62070 12480 62098
rect 12256 60716 12308 60722
rect 12256 60658 12308 60664
rect 12452 59430 12480 62070
rect 13820 60716 13872 60722
rect 13820 60658 13872 60664
rect 13544 60648 13596 60654
rect 13544 60590 13596 60596
rect 12440 59424 12492 59430
rect 12440 59366 12492 59372
rect 13268 57928 13320 57934
rect 13268 57870 13320 57876
rect 11244 56636 11296 56642
rect 11244 56578 11296 56584
rect 10968 56500 11020 56506
rect 10968 56442 11020 56448
rect 10876 56432 10928 56438
rect 10876 56374 10928 56380
rect 10324 53848 10376 53854
rect 10324 53790 10376 53796
rect 8668 53168 8720 53174
rect 7748 53100 7800 53106
rect 8220 53094 8340 53122
rect 8668 53110 8720 53116
rect 7748 53042 7800 53048
rect 3606 52048 3662 52057
rect 3516 52012 3568 52018
rect 3606 51983 3662 51992
rect 3516 51954 3568 51960
rect 8312 50998 8340 53094
rect 10888 52426 10916 56374
rect 10980 55214 11008 56442
rect 10980 55186 11100 55214
rect 11072 53718 11100 55186
rect 11060 53712 11112 53718
rect 11060 53654 11112 53660
rect 13280 52494 13308 57870
rect 13556 55486 13584 60590
rect 13832 59226 13860 60658
rect 13820 59220 13872 59226
rect 13820 59162 13872 59168
rect 13544 55480 13596 55486
rect 13544 55422 13596 55428
rect 14476 54670 14504 63242
rect 15120 62098 15148 64806
rect 15120 62070 15240 62098
rect 15212 59362 15240 62070
rect 15200 59356 15252 59362
rect 15200 59298 15252 59304
rect 15304 59158 15332 64846
rect 15292 59152 15344 59158
rect 15292 59094 15344 59100
rect 17236 57934 17264 78610
rect 17316 73228 17368 73234
rect 17316 73170 17368 73176
rect 17328 63442 17356 73170
rect 17316 63436 17368 63442
rect 17316 63378 17368 63384
rect 17316 59356 17368 59362
rect 17316 59298 17368 59304
rect 17224 57928 17276 57934
rect 17224 57870 17276 57876
rect 16488 56568 16540 56574
rect 16488 56510 16540 56516
rect 16500 55162 16528 56510
rect 16500 55134 16620 55162
rect 14464 54664 14516 54670
rect 14464 54606 14516 54612
rect 15568 54664 15620 54670
rect 15568 54606 15620 54612
rect 15200 53780 15252 53786
rect 15200 53722 15252 53728
rect 13820 53712 13872 53718
rect 13820 53654 13872 53660
rect 13268 52488 13320 52494
rect 13268 52430 13320 52436
rect 10876 52420 10928 52426
rect 10876 52362 10928 52368
rect 12440 52420 12492 52426
rect 12440 52362 12492 52368
rect 8300 50992 8352 50998
rect 8300 50934 8352 50940
rect 7654 50552 7710 50561
rect 7654 50487 7710 50496
rect 2870 50416 2926 50425
rect 2870 50351 2926 50360
rect 1674 3632 1730 3641
rect 1674 3567 1730 3576
rect 570 3360 626 3369
rect 570 3295 626 3304
rect 584 480 612 3295
rect 1688 480 1716 3567
rect 2884 480 2912 50351
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 5262 4040 5318 4049
rect 5262 3975 5318 3984
rect 4066 3496 4122 3505
rect 4066 3431 4122 3440
rect 4080 480 4108 3431
rect 5276 480 5304 3975
rect 6458 3768 6514 3777
rect 6458 3703 6514 3712
rect 6472 480 6500 3703
rect 7668 480 7696 50487
rect 12452 49706 12480 52362
rect 13832 50386 13860 53654
rect 15212 52154 15240 53722
rect 15200 52148 15252 52154
rect 15200 52090 15252 52096
rect 15580 51746 15608 54606
rect 16592 51950 16620 55134
rect 17328 53718 17356 59298
rect 17868 59288 17920 59294
rect 17868 59230 17920 59236
rect 17408 59220 17460 59226
rect 17408 59162 17460 59168
rect 17420 54126 17448 59162
rect 17880 57882 17908 59230
rect 18328 57928 18380 57934
rect 17880 57854 18000 57882
rect 18328 57870 18380 57876
rect 17408 54120 17460 54126
rect 17408 54062 17460 54068
rect 17316 53712 17368 53718
rect 17316 53654 17368 53660
rect 16580 51944 16632 51950
rect 16580 51886 16632 51892
rect 15568 51740 15620 51746
rect 15568 51682 15620 51688
rect 17972 50930 18000 57854
rect 18052 55480 18104 55486
rect 18052 55422 18104 55428
rect 18064 52358 18092 55422
rect 18052 52352 18104 52358
rect 18052 52294 18104 52300
rect 18340 51678 18368 57870
rect 18616 51921 18644 84186
rect 18696 63436 18748 63442
rect 18696 63378 18748 63384
rect 18602 51912 18658 51921
rect 18708 51882 18736 63378
rect 18880 59152 18932 59158
rect 18880 59094 18932 59100
rect 18602 51847 18658 51856
rect 18696 51876 18748 51882
rect 18696 51818 18748 51824
rect 18892 51814 18920 59094
rect 19340 54120 19392 54126
rect 19340 54062 19392 54068
rect 19352 52426 19380 54062
rect 19524 53712 19576 53718
rect 19524 53654 19576 53660
rect 19248 52420 19300 52426
rect 19248 52362 19300 52368
rect 19340 52420 19392 52426
rect 19340 52362 19392 52368
rect 18880 51808 18932 51814
rect 18880 51750 18932 51756
rect 18328 51672 18380 51678
rect 18328 51614 18380 51620
rect 17960 50924 18012 50930
rect 17960 50866 18012 50872
rect 19260 50794 19288 52362
rect 19536 51610 19564 53654
rect 20444 53168 20496 53174
rect 20444 53110 20496 53116
rect 19524 51604 19576 51610
rect 19524 51546 19576 51552
rect 20456 51542 20484 53110
rect 20628 53100 20680 53106
rect 20628 53042 20680 53048
rect 20536 52148 20588 52154
rect 20536 52090 20588 52096
rect 20444 51536 20496 51542
rect 20444 51478 20496 51484
rect 19248 50788 19300 50794
rect 19248 50730 19300 50736
rect 20548 50522 20576 52090
rect 20640 51898 20668 53042
rect 20812 52420 20864 52426
rect 20812 52362 20864 52368
rect 20640 51870 20760 51898
rect 20732 51746 20760 51870
rect 20628 51740 20680 51746
rect 20628 51682 20680 51688
rect 20720 51740 20772 51746
rect 20720 51682 20772 51688
rect 20640 50862 20668 51682
rect 20628 50856 20680 50862
rect 20628 50798 20680 50804
rect 20824 50726 20852 52362
rect 20904 52352 20956 52358
rect 20904 52294 20956 52300
rect 20812 50720 20864 50726
rect 20812 50662 20864 50668
rect 20916 50658 20944 52294
rect 20996 51536 21048 51542
rect 20996 51478 21048 51484
rect 20904 50652 20956 50658
rect 20904 50594 20956 50600
rect 20536 50516 20588 50522
rect 20536 50458 20588 50464
rect 21008 50454 21036 51478
rect 21376 51066 21404 93826
rect 378784 51536 378836 51542
rect 378784 51478 378836 51484
rect 378692 51400 378744 51406
rect 378692 51342 378744 51348
rect 377956 51332 378008 51338
rect 377956 51274 378008 51280
rect 21364 51060 21416 51066
rect 21364 51002 21416 51008
rect 377968 50998 377996 51274
rect 377956 50992 378008 50998
rect 377956 50934 378008 50940
rect 51354 50824 51410 50833
rect 51354 50759 51410 50768
rect 47858 50688 47914 50697
rect 47858 50623 47914 50632
rect 33140 50516 33192 50522
rect 33140 50458 33192 50464
rect 20996 50448 21048 50454
rect 20996 50390 21048 50396
rect 13820 50380 13872 50386
rect 13820 50322 13872 50328
rect 12440 49700 12492 49706
rect 12440 49642 12492 49648
rect 33152 49638 33180 50458
rect 42800 50448 42852 50454
rect 42800 50390 42852 50396
rect 33140 49632 33192 49638
rect 33140 49574 33192 49580
rect 42812 49502 42840 50390
rect 44180 50380 44232 50386
rect 44180 50322 44232 50328
rect 44192 49570 44220 50322
rect 46662 50280 46718 50289
rect 46662 50215 46718 50224
rect 44180 49564 44232 49570
rect 44180 49506 44232 49512
rect 42800 49496 42852 49502
rect 42800 49438 42852 49444
rect 12348 47592 12400 47598
rect 12348 47534 12400 47540
rect 9954 3904 10010 3913
rect 9954 3839 10010 3848
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 480 8800 3538
rect 9968 480 9996 3839
rect 12360 480 12388 47534
rect 44272 45144 44324 45150
rect 44272 45086 44324 45092
rect 40684 45076 40736 45082
rect 40684 45018 40736 45024
rect 37188 45008 37240 45014
rect 37188 44950 37240 44956
rect 33600 44940 33652 44946
rect 33600 44882 33652 44888
rect 26516 44872 26568 44878
rect 26516 44814 26568 44820
rect 23020 39432 23072 39438
rect 23020 39374 23072 39380
rect 18236 39364 18288 39370
rect 18236 39306 18288 39312
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 13544 3868 13596 3874
rect 13544 3810 13596 3816
rect 13556 480 13584 3810
rect 14752 480 14780 3878
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 17052 480 17080 3674
rect 18248 480 18276 39306
rect 19432 33788 19484 33794
rect 19432 33730 19484 33736
rect 19444 480 19472 33730
rect 21824 3800 21876 3806
rect 21824 3742 21876 3748
rect 21836 480 21864 3742
rect 23032 480 23060 39374
rect 24216 33856 24268 33862
rect 24216 33798 24268 33804
rect 24228 480 24256 33798
rect 26528 480 26556 44814
rect 31300 39568 31352 39574
rect 31300 39510 31352 39516
rect 27712 39500 27764 39506
rect 27712 39442 27764 39448
rect 27724 480 27752 39442
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 28920 480 28948 3606
rect 30104 2100 30156 2106
rect 30104 2042 30156 2048
rect 30116 480 30144 2042
rect 31312 480 31340 39510
rect 32404 4072 32456 4078
rect 32404 4014 32456 4020
rect 32416 480 32444 4014
rect 33612 480 33640 44882
rect 34796 39636 34848 39642
rect 34796 39578 34848 39584
rect 34808 480 34836 39578
rect 35992 3460 36044 3466
rect 35992 3402 36044 3408
rect 36004 480 36032 3402
rect 37200 480 37228 44950
rect 38384 39704 38436 39710
rect 38384 39646 38436 39652
rect 38396 480 38424 39646
rect 39580 33924 39632 33930
rect 39580 33866 39632 33872
rect 39592 480 39620 33866
rect 40696 480 40724 45018
rect 41880 42084 41932 42090
rect 41880 42026 41932 42032
rect 41892 480 41920 42026
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 43088 480 43116 3470
rect 44284 480 44312 45086
rect 45468 39772 45520 39778
rect 45468 39714 45520 39720
rect 45480 480 45508 39714
rect 46676 480 46704 50215
rect 47872 480 47900 50623
rect 50160 45280 50212 45286
rect 50160 45222 50212 45228
rect 48964 45212 49016 45218
rect 48964 45154 49016 45160
rect 48976 480 49004 45154
rect 50172 480 50200 45222
rect 51368 480 51396 50759
rect 65524 50584 65576 50590
rect 65524 50526 65576 50532
rect 62028 50516 62080 50522
rect 62028 50458 62080 50464
rect 58440 50448 58492 50454
rect 58440 50390 58492 50396
rect 54944 50380 54996 50386
rect 54944 50322 54996 50328
rect 52552 42152 52604 42158
rect 52552 42094 52604 42100
rect 52564 480 52592 42094
rect 53748 36644 53800 36650
rect 53748 36586 53800 36592
rect 53760 480 53788 36586
rect 54956 480 54984 50322
rect 56048 42220 56100 42226
rect 56048 42162 56100 42168
rect 56060 480 56088 42162
rect 57244 36712 57296 36718
rect 57244 36654 57296 36660
rect 57256 480 57284 36654
rect 58452 480 58480 50390
rect 59636 42288 59688 42294
rect 59636 42230 59688 42236
rect 59648 480 59676 42230
rect 60832 36576 60884 36582
rect 60832 36518 60884 36524
rect 60844 480 60872 36518
rect 62040 480 62068 50458
rect 63224 42356 63276 42362
rect 63224 42298 63276 42304
rect 63236 480 63264 42298
rect 64328 36780 64380 36786
rect 64328 36722 64380 36728
rect 64340 480 64368 36722
rect 65536 480 65564 50526
rect 70308 50312 70360 50318
rect 70308 50254 70360 50260
rect 69112 47660 69164 47666
rect 69112 47602 69164 47608
rect 66720 45484 66772 45490
rect 66720 45426 66772 45432
rect 66732 480 66760 45426
rect 67916 4140 67968 4146
rect 67916 4082 67968 4088
rect 67928 480 67956 4082
rect 69124 480 69152 47602
rect 70320 480 70348 50254
rect 93952 50244 94004 50250
rect 93952 50186 94004 50192
rect 87972 48204 88024 48210
rect 87972 48146 88024 48152
rect 86868 48000 86920 48006
rect 86868 47942 86920 47948
rect 83280 47932 83332 47938
rect 83280 47874 83332 47880
rect 79692 47864 79744 47870
rect 79692 47806 79744 47812
rect 76196 47796 76248 47802
rect 76196 47738 76248 47744
rect 72608 47728 72660 47734
rect 72608 47670 72660 47676
rect 71504 36848 71556 36854
rect 71504 36790 71556 36796
rect 71516 480 71544 36790
rect 72620 480 72648 47670
rect 73804 42424 73856 42430
rect 73804 42366 73856 42372
rect 73816 480 73844 42366
rect 75000 36916 75052 36922
rect 75000 36858 75052 36864
rect 75012 480 75040 36858
rect 76208 480 76236 47738
rect 77392 42492 77444 42498
rect 77392 42434 77444 42440
rect 77404 480 77432 42434
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 78600 480 78628 3334
rect 79704 480 79732 47806
rect 80888 42560 80940 42566
rect 80888 42502 80940 42508
rect 80900 480 80928 42502
rect 82084 36984 82136 36990
rect 82084 36926 82136 36932
rect 82096 480 82124 36926
rect 83292 480 83320 47874
rect 84476 42628 84528 42634
rect 84476 42570 84528 42576
rect 84488 480 84516 42570
rect 85672 37052 85724 37058
rect 85672 36994 85724 37000
rect 85684 480 85712 36994
rect 86880 480 86908 47942
rect 87984 480 88012 48146
rect 90364 48068 90416 48074
rect 90364 48010 90416 48016
rect 89168 37120 89220 37126
rect 89168 37062 89220 37068
rect 89180 480 89208 37062
rect 90376 480 90404 48010
rect 91560 42764 91612 42770
rect 91560 42706 91612 42712
rect 91572 480 91600 42706
rect 92756 37188 92808 37194
rect 92756 37130 92808 37136
rect 92768 480 92796 37130
rect 93964 480 93992 50186
rect 115204 50176 115256 50182
rect 115204 50118 115256 50124
rect 101036 48272 101088 48278
rect 101036 48214 101088 48220
rect 97448 48136 97500 48142
rect 97448 48078 97500 48084
rect 95148 42016 95200 42022
rect 95148 41958 95200 41964
rect 95160 480 95188 41958
rect 96252 37256 96304 37262
rect 96252 37198 96304 37204
rect 96264 480 96292 37198
rect 97460 480 97488 48078
rect 98644 42696 98696 42702
rect 98644 42638 98696 42644
rect 98656 480 98684 42638
rect 99840 4004 99892 4010
rect 99840 3946 99892 3952
rect 99852 480 99880 3946
rect 101048 480 101076 48214
rect 104532 47524 104584 47530
rect 104532 47466 104584 47472
rect 102232 41948 102284 41954
rect 102232 41890 102284 41896
rect 102244 480 102272 41890
rect 103336 36508 103388 36514
rect 103336 36450 103388 36456
rect 103348 480 103376 36450
rect 104544 480 104572 47466
rect 110512 47456 110564 47462
rect 110512 47398 110564 47404
rect 108120 44804 108172 44810
rect 108120 44746 108172 44752
rect 105728 39840 105780 39846
rect 105728 39782 105780 39788
rect 105740 480 105768 39782
rect 106924 3324 106976 3330
rect 106924 3266 106976 3272
rect 106936 480 106964 3266
rect 108132 480 108160 44746
rect 109316 39296 109368 39302
rect 109316 39238 109368 39244
rect 109328 480 109356 39238
rect 110524 480 110552 47398
rect 111616 44736 111668 44742
rect 111616 44678 111668 44684
rect 111628 480 111656 44678
rect 112812 39228 112864 39234
rect 112812 39170 112864 39176
rect 112824 480 112852 39170
rect 114008 3256 114060 3262
rect 114008 3198 114060 3204
rect 114020 480 114048 3198
rect 115216 480 115244 50118
rect 378704 49706 378732 51342
rect 378796 50794 378824 51478
rect 378876 51264 378928 51270
rect 378876 51206 378928 51212
rect 378784 50788 378836 50794
rect 378784 50730 378836 50736
rect 378692 49700 378744 49706
rect 378692 49642 378744 49648
rect 378888 49502 378916 51206
rect 378876 49496 378928 49502
rect 378876 49438 378928 49444
rect 122288 45416 122340 45422
rect 122288 45358 122340 45364
rect 118792 45348 118844 45354
rect 118792 45290 118844 45296
rect 116400 39976 116452 39982
rect 116400 39918 116452 39924
rect 116412 480 116440 39918
rect 117596 33992 117648 33998
rect 117596 33934 117648 33940
rect 117608 480 117636 33934
rect 118804 480 118832 45290
rect 119896 39908 119948 39914
rect 119896 39850 119948 39856
rect 119908 480 119936 39850
rect 121092 34060 121144 34066
rect 121092 34002 121144 34008
rect 121104 480 121132 34002
rect 122300 480 122328 45358
rect 123484 40044 123536 40050
rect 123484 39986 123536 39992
rect 123496 480 123524 39986
rect 124680 34128 124732 34134
rect 124680 34070 124732 34076
rect 124692 480 124720 34070
rect 380176 3942 380204 305662
rect 380256 305652 380308 305658
rect 380256 305594 380308 305600
rect 380164 3936 380216 3942
rect 380164 3878 380216 3884
rect 380268 3398 380296 305594
rect 382280 304428 382332 304434
rect 382280 304370 382332 304376
rect 381544 304292 381596 304298
rect 381544 304234 381596 304240
rect 380348 295996 380400 296002
rect 380348 295938 380400 295944
rect 380360 4146 380388 295938
rect 380440 275324 380492 275330
rect 380440 275266 380492 275272
rect 380348 4140 380400 4146
rect 380348 4082 380400 4088
rect 380452 4049 380480 275266
rect 380532 173188 380584 173194
rect 380532 173130 380584 173136
rect 380544 50658 380572 173130
rect 380624 118924 380676 118930
rect 380624 118866 380676 118872
rect 380636 50726 380664 118866
rect 380716 91112 380768 91118
rect 380716 91054 380768 91060
rect 380728 51678 380756 91054
rect 381452 87916 381504 87922
rect 381452 87858 381504 87864
rect 380716 51672 380768 51678
rect 380716 51614 380768 51620
rect 381464 51610 381492 87858
rect 381452 51604 381504 51610
rect 381452 51546 381504 51552
rect 380624 50720 380676 50726
rect 380624 50662 380676 50668
rect 380532 50652 380584 50658
rect 380532 50594 380584 50600
rect 381556 4078 381584 304234
rect 381728 303000 381780 303006
rect 381728 302942 381780 302948
rect 381636 302932 381688 302938
rect 381636 302874 381688 302880
rect 381544 4072 381596 4078
rect 380438 4040 380494 4049
rect 381544 4014 381596 4020
rect 380438 3975 380494 3984
rect 380256 3392 380308 3398
rect 380256 3334 380308 3340
rect 381648 3262 381676 302874
rect 381740 3330 381768 302942
rect 382292 301753 382320 304370
rect 382278 301744 382334 301753
rect 382278 301679 382334 301688
rect 382924 295112 382976 295118
rect 382924 295054 382976 295060
rect 381820 294976 381872 294982
rect 381820 294918 381872 294924
rect 381832 39302 381860 294918
rect 381912 294772 381964 294778
rect 381912 294714 381964 294720
rect 381924 41954 381952 294714
rect 382004 294636 382056 294642
rect 382004 294578 382056 294584
rect 382016 42022 382044 294578
rect 382280 281512 382332 281518
rect 382280 281454 382332 281460
rect 382292 280537 382320 281454
rect 382278 280528 382334 280537
rect 382278 280463 382334 280472
rect 382280 270496 382332 270502
rect 382280 270438 382332 270444
rect 382292 269929 382320 270438
rect 382278 269920 382334 269929
rect 382278 269855 382334 269864
rect 382280 259412 382332 259418
rect 382280 259354 382332 259360
rect 382292 259321 382320 259354
rect 382278 259312 382334 259321
rect 382278 259247 382334 259256
rect 382280 249756 382332 249762
rect 382280 249698 382332 249704
rect 382292 248713 382320 249698
rect 382278 248704 382334 248713
rect 382278 248639 382334 248648
rect 382280 238740 382332 238746
rect 382280 238682 382332 238688
rect 382292 238105 382320 238682
rect 382278 238096 382334 238105
rect 382278 238031 382334 238040
rect 382280 227724 382332 227730
rect 382280 227666 382332 227672
rect 382292 227497 382320 227666
rect 382278 227488 382334 227497
rect 382278 227423 382334 227432
rect 382280 206984 382332 206990
rect 382280 206926 382332 206932
rect 382292 206281 382320 206926
rect 382278 206272 382334 206281
rect 382278 206207 382334 206216
rect 382280 195968 382332 195974
rect 382280 195910 382332 195916
rect 382292 195673 382320 195910
rect 382278 195664 382334 195673
rect 382278 195599 382334 195608
rect 382280 186312 382332 186318
rect 382280 186254 382332 186260
rect 382096 186244 382148 186250
rect 382096 186186 382148 186192
rect 382108 51950 382136 186186
rect 382292 185065 382320 186254
rect 382278 185056 382334 185065
rect 382278 184991 382334 185000
rect 382280 175228 382332 175234
rect 382280 175170 382332 175176
rect 382292 174457 382320 175170
rect 382278 174448 382334 174457
rect 382278 174383 382334 174392
rect 382280 154556 382332 154562
rect 382280 154498 382332 154504
rect 382292 153241 382320 154498
rect 382278 153232 382334 153241
rect 382278 153167 382334 153176
rect 382280 143540 382332 143546
rect 382280 143482 382332 143488
rect 382292 142633 382320 143482
rect 382278 142624 382334 142633
rect 382278 142559 382334 142568
rect 382280 132456 382332 132462
rect 382280 132398 382332 132404
rect 382292 132025 382320 132398
rect 382278 132016 382334 132025
rect 382278 131951 382334 131960
rect 382188 131164 382240 131170
rect 382188 131106 382240 131112
rect 382096 51944 382148 51950
rect 382096 51886 382148 51892
rect 382200 50930 382228 131106
rect 382280 111784 382332 111790
rect 382280 111726 382332 111732
rect 382292 110809 382320 111726
rect 382278 110800 382334 110809
rect 382278 110735 382334 110744
rect 382280 100700 382332 100706
rect 382280 100642 382332 100648
rect 382292 100201 382320 100642
rect 382278 100192 382334 100201
rect 382278 100127 382334 100136
rect 382280 89684 382332 89690
rect 382280 89626 382332 89632
rect 382292 89593 382320 89626
rect 382278 89584 382334 89593
rect 382278 89519 382334 89528
rect 382832 86284 382884 86290
rect 382832 86226 382884 86232
rect 382280 79960 382332 79966
rect 382280 79902 382332 79908
rect 382292 78985 382320 79902
rect 382278 78976 382334 78985
rect 382278 78911 382334 78920
rect 382280 69012 382332 69018
rect 382280 68954 382332 68960
rect 382292 68377 382320 68954
rect 382278 68368 382334 68377
rect 382278 68303 382334 68312
rect 382280 57928 382332 57934
rect 382280 57870 382332 57876
rect 382292 57769 382320 57870
rect 382278 57760 382334 57769
rect 382278 57695 382334 57704
rect 382372 51604 382424 51610
rect 382372 51546 382424 51552
rect 382280 51468 382332 51474
rect 382280 51410 382332 51416
rect 382188 50924 382240 50930
rect 382188 50866 382240 50872
rect 382292 49638 382320 51410
rect 382280 49632 382332 49638
rect 382280 49574 382332 49580
rect 382384 49570 382412 51546
rect 382844 51338 382872 86226
rect 382832 51332 382884 51338
rect 382832 51274 382884 51280
rect 382372 49564 382424 49570
rect 382372 49506 382424 49512
rect 382004 42016 382056 42022
rect 382004 41958 382056 41964
rect 381912 41948 381964 41954
rect 381912 41890 381964 41896
rect 382936 39370 382964 295054
rect 383016 294704 383068 294710
rect 383016 294646 383068 294652
rect 382924 39364 382976 39370
rect 382924 39306 382976 39312
rect 381820 39296 381872 39302
rect 381820 39238 381872 39244
rect 383028 39234 383056 294646
rect 383200 292460 383252 292466
rect 383200 292402 383252 292408
rect 383108 292120 383160 292126
rect 383108 292062 383160 292068
rect 383120 39506 383148 292062
rect 383108 39500 383160 39506
rect 383108 39442 383160 39448
rect 383212 39438 383240 292402
rect 383304 291145 383332 305866
rect 403900 305856 403952 305862
rect 403900 305798 403952 305804
rect 406382 305824 406438 305833
rect 403716 305788 403768 305794
rect 403716 305730 403768 305736
rect 401140 303612 401192 303618
rect 401140 303554 401192 303560
rect 398104 303204 398156 303210
rect 398104 303146 398156 303152
rect 395344 300824 395396 300830
rect 395344 300766 395396 300772
rect 392676 300620 392728 300626
rect 392676 300562 392728 300568
rect 392584 300348 392636 300354
rect 392584 300290 392636 300296
rect 387432 298104 387484 298110
rect 387432 298046 387484 298052
rect 387248 297628 387300 297634
rect 387248 297570 387300 297576
rect 387156 297560 387208 297566
rect 387156 297502 387208 297508
rect 387064 297424 387116 297430
rect 387064 297366 387116 297372
rect 384396 295044 384448 295050
rect 384396 294986 384448 294992
rect 384302 294536 384358 294545
rect 384302 294471 384358 294480
rect 383290 291136 383346 291145
rect 383290 291071 383346 291080
rect 383384 264240 383436 264246
rect 383384 264182 383436 264188
rect 383292 235272 383344 235278
rect 383292 235214 383344 235220
rect 383304 51882 383332 235214
rect 383396 216889 383424 264182
rect 383382 216880 383438 216889
rect 383382 216815 383438 216824
rect 383384 207664 383436 207670
rect 383384 207606 383436 207612
rect 383292 51876 383344 51882
rect 383292 51818 383344 51824
rect 383396 51814 383424 207606
rect 383476 167068 383528 167074
rect 383476 167010 383528 167016
rect 383488 121417 383516 167010
rect 383474 121408 383530 121417
rect 383474 121343 383530 121352
rect 383476 99340 383528 99346
rect 383476 99282 383528 99288
rect 383488 91118 383516 99282
rect 383476 91112 383528 91118
rect 383476 91054 383528 91060
rect 383476 87372 383528 87378
rect 383476 87314 383528 87320
rect 383384 51808 383436 51814
rect 383384 51750 383436 51756
rect 383488 50862 383516 87314
rect 383568 85604 383620 85610
rect 383568 85546 383620 85552
rect 383580 51746 383608 85546
rect 383568 51740 383620 51746
rect 383568 51682 383620 51688
rect 383476 50856 383528 50862
rect 383476 50798 383528 50804
rect 383200 39432 383252 39438
rect 383200 39374 383252 39380
rect 383016 39228 383068 39234
rect 383016 39170 383068 39176
rect 384316 3874 384344 294471
rect 384408 42770 384436 294986
rect 384580 294908 384632 294914
rect 384580 294850 384632 294856
rect 384488 294840 384540 294846
rect 384488 294782 384540 294788
rect 384396 42764 384448 42770
rect 384396 42706 384448 42712
rect 384500 42634 384528 294782
rect 384592 48210 384620 294850
rect 385960 292324 386012 292330
rect 385960 292266 386012 292272
rect 385776 291916 385828 291922
rect 385776 291858 385828 291864
rect 385684 291848 385736 291854
rect 385684 291790 385736 291796
rect 384672 214600 384724 214606
rect 384672 214542 384724 214548
rect 384684 51542 384712 214542
rect 384764 199436 384816 199442
rect 384764 199378 384816 199384
rect 384776 186250 384804 199378
rect 384764 186244 384816 186250
rect 384764 186186 384816 186192
rect 384764 167136 384816 167142
rect 384764 167078 384816 167084
rect 384776 87922 384804 167078
rect 384856 147688 384908 147694
rect 384856 147630 384908 147636
rect 384868 131170 384896 147630
rect 384948 133612 385000 133618
rect 384948 133554 385000 133560
rect 384856 131164 384908 131170
rect 384856 131106 384908 131112
rect 384960 118930 384988 133554
rect 384948 118924 385000 118930
rect 384948 118866 385000 118872
rect 385040 100768 385092 100774
rect 385040 100710 385092 100716
rect 385052 99414 385080 100710
rect 385040 99408 385092 99414
rect 385040 99350 385092 99356
rect 384764 87916 384816 87922
rect 384764 87858 384816 87864
rect 384764 82884 384816 82890
rect 384764 82826 384816 82832
rect 384776 51610 384804 82826
rect 384764 51604 384816 51610
rect 384764 51546 384816 51552
rect 384672 51536 384724 51542
rect 384672 51478 384724 51484
rect 384580 48204 384632 48210
rect 384580 48146 384632 48152
rect 384488 42628 384540 42634
rect 384488 42570 384540 42576
rect 385696 39642 385724 291790
rect 385788 39710 385816 291858
rect 385866 291816 385922 291825
rect 385866 291751 385922 291760
rect 385776 39704 385828 39710
rect 385776 39646 385828 39652
rect 385684 39636 385736 39642
rect 385684 39578 385736 39584
rect 385880 39574 385908 291751
rect 385972 42090 386000 292266
rect 386144 169040 386196 169046
rect 386144 168982 386196 168988
rect 386052 165028 386104 165034
rect 386052 164970 386104 164976
rect 386064 79966 386092 164970
rect 386156 87378 386184 168982
rect 386236 142996 386288 143002
rect 386236 142938 386288 142944
rect 386144 87372 386196 87378
rect 386144 87314 386196 87320
rect 386248 85610 386276 142938
rect 386236 85604 386288 85610
rect 386236 85546 386288 85552
rect 386144 85536 386196 85542
rect 386144 85478 386196 85484
rect 386052 79960 386104 79966
rect 386052 79902 386104 79908
rect 386052 73228 386104 73234
rect 386052 73170 386104 73176
rect 386064 51474 386092 73170
rect 386052 51468 386104 51474
rect 386052 51410 386104 51416
rect 386156 51270 386184 85478
rect 386236 81456 386288 81462
rect 386236 81398 386288 81404
rect 386248 51406 386276 81398
rect 386236 51400 386288 51406
rect 386236 51342 386288 51348
rect 386144 51264 386196 51270
rect 386144 51206 386196 51212
rect 387076 42430 387104 297366
rect 387168 42498 387196 297502
rect 387260 42566 387288 297570
rect 387340 297492 387392 297498
rect 387340 297434 387392 297440
rect 387248 42560 387300 42566
rect 387248 42502 387300 42508
rect 387156 42492 387208 42498
rect 387156 42434 387208 42440
rect 387064 42424 387116 42430
rect 387064 42366 387116 42372
rect 387352 42362 387380 297434
rect 387444 45490 387472 298046
rect 390100 298036 390152 298042
rect 390100 297978 390152 297984
rect 390008 297832 390060 297838
rect 390008 297774 390060 297780
rect 389916 297764 389968 297770
rect 389916 297706 389968 297712
rect 387524 297696 387576 297702
rect 387524 297638 387576 297644
rect 387536 50318 387564 297638
rect 389822 297528 389878 297537
rect 389822 297463 389878 297472
rect 388536 292392 388588 292398
rect 388536 292334 388588 292340
rect 388442 291952 388498 291961
rect 388442 291887 388498 291896
rect 387616 227792 387668 227798
rect 387616 227734 387668 227740
rect 387628 86290 387656 227734
rect 387708 164892 387760 164898
rect 387708 164834 387760 164840
rect 387720 147694 387748 164834
rect 388168 149116 388220 149122
rect 388168 149058 388220 149064
rect 387708 147688 387760 147694
rect 387708 147630 387760 147636
rect 388180 143002 388208 149058
rect 388168 142996 388220 143002
rect 388168 142938 388220 142944
rect 387616 86284 387668 86290
rect 387616 86226 387668 86232
rect 387616 85536 387668 85542
rect 387616 85478 387668 85484
rect 387628 82890 387656 85478
rect 387800 84176 387852 84182
rect 387800 84118 387852 84124
rect 387616 82884 387668 82890
rect 387616 82826 387668 82832
rect 387812 81462 387840 84118
rect 387800 81456 387852 81462
rect 387800 81398 387852 81404
rect 387616 80096 387668 80102
rect 387616 80038 387668 80044
rect 387628 73234 387656 80038
rect 387616 73228 387668 73234
rect 387616 73170 387668 73176
rect 387524 50312 387576 50318
rect 387524 50254 387576 50260
rect 387432 45484 387484 45490
rect 387432 45426 387484 45432
rect 387340 42356 387392 42362
rect 387340 42298 387392 42304
rect 385960 42084 386012 42090
rect 385960 42026 386012 42032
rect 385868 39568 385920 39574
rect 385868 39510 385920 39516
rect 388456 3913 388484 291887
rect 388548 39778 388576 292334
rect 388628 292188 388680 292194
rect 388628 292130 388680 292136
rect 388640 45286 388668 292130
rect 388720 169108 388772 169114
rect 388720 169050 388772 169056
rect 388732 85542 388760 169050
rect 388812 103488 388864 103494
rect 388812 103430 388864 103436
rect 388824 85610 388852 103430
rect 388812 85604 388864 85610
rect 388812 85546 388864 85552
rect 388720 85536 388772 85542
rect 388720 85478 388772 85484
rect 389456 82884 389508 82890
rect 389456 82826 389508 82832
rect 389468 80102 389496 82826
rect 389456 80096 389508 80102
rect 389456 80038 389508 80044
rect 388628 45280 388680 45286
rect 388628 45222 388680 45228
rect 388536 39772 388588 39778
rect 388536 39714 388588 39720
rect 388442 3904 388498 3913
rect 384304 3868 384356 3874
rect 388442 3839 388498 3848
rect 384304 3810 384356 3816
rect 389836 3602 389864 297463
rect 389928 42294 389956 297706
rect 389916 42288 389968 42294
rect 389916 42230 389968 42236
rect 390020 42226 390048 297774
rect 390008 42220 390060 42226
rect 390008 42162 390060 42168
rect 390112 42158 390140 297978
rect 390192 297968 390244 297974
rect 390192 297910 390244 297916
rect 390204 45150 390232 297910
rect 390284 297900 390336 297906
rect 390284 297842 390336 297848
rect 390296 45218 390324 297842
rect 391478 294672 391534 294681
rect 391478 294607 391534 294616
rect 391388 292256 391440 292262
rect 391388 292198 391440 292204
rect 391296 292052 391348 292058
rect 391296 291994 391348 292000
rect 391204 291984 391256 291990
rect 391204 291926 391256 291932
rect 390376 245200 390428 245206
rect 390376 245142 390428 245148
rect 390388 235278 390416 245142
rect 390376 235272 390428 235278
rect 390376 235214 390428 235220
rect 390376 186380 390428 186386
rect 390376 186322 390428 186328
rect 390388 173194 390416 186322
rect 390376 173188 390428 173194
rect 390376 173130 390428 173136
rect 390560 137420 390612 137426
rect 390560 137362 390612 137368
rect 390572 133618 390600 137362
rect 390560 133612 390612 133618
rect 390560 133554 390612 133560
rect 391112 111852 391164 111858
rect 391112 111794 391164 111800
rect 391124 103562 391152 111794
rect 391112 103556 391164 103562
rect 391112 103498 391164 103504
rect 390284 45212 390336 45218
rect 390284 45154 390336 45160
rect 390192 45144 390244 45150
rect 390192 45086 390244 45092
rect 390100 42152 390152 42158
rect 390100 42094 390152 42100
rect 391216 36718 391244 291926
rect 391204 36712 391256 36718
rect 391204 36654 391256 36660
rect 391308 36650 391336 291994
rect 391400 36786 391428 292198
rect 391492 39846 391520 294607
rect 391572 165708 391624 165714
rect 391572 165650 391624 165656
rect 391584 57934 391612 165650
rect 392400 152516 392452 152522
rect 392400 152458 392452 152464
rect 392412 149122 392440 152458
rect 392400 149116 392452 149122
rect 392400 149058 392452 149064
rect 391664 113144 391716 113150
rect 391664 113086 391716 113092
rect 391676 84250 391704 113086
rect 391756 100020 391808 100026
rect 391756 99962 391808 99968
rect 391664 84244 391716 84250
rect 391664 84186 391716 84192
rect 391768 82890 391796 99962
rect 391756 82884 391808 82890
rect 391756 82826 391808 82832
rect 391572 57928 391624 57934
rect 391572 57870 391624 57876
rect 391480 39840 391532 39846
rect 391480 39782 391532 39788
rect 391388 36780 391440 36786
rect 391388 36722 391440 36728
rect 391296 36644 391348 36650
rect 391296 36586 391348 36592
rect 389824 3596 389876 3602
rect 389824 3538 389876 3544
rect 381728 3324 381780 3330
rect 381728 3266 381780 3272
rect 381636 3256 381688 3262
rect 381636 3198 381688 3204
rect 392596 2106 392624 300290
rect 392688 3806 392716 300562
rect 393042 300248 393098 300257
rect 393042 300183 393098 300192
rect 392768 300144 392820 300150
rect 392768 300086 392820 300092
rect 392858 300112 392914 300121
rect 392780 45014 392808 300086
rect 392858 300047 392914 300056
rect 392768 45008 392820 45014
rect 392768 44950 392820 44956
rect 392872 44878 392900 300047
rect 392950 297392 393006 297401
rect 392950 297327 393006 297336
rect 392964 45082 392992 297327
rect 392952 45076 393004 45082
rect 392952 45018 393004 45024
rect 393056 44946 393084 300183
rect 394332 295316 394384 295322
rect 394332 295258 394384 295264
rect 393964 295248 394016 295254
rect 393964 295190 394016 295196
rect 393136 206372 393188 206378
rect 393136 206314 393188 206320
rect 393148 186386 393176 206314
rect 393136 186380 393188 186386
rect 393136 186322 393188 186328
rect 393136 175976 393188 175982
rect 393136 175918 393188 175924
rect 393148 167142 393176 175918
rect 393320 172100 393372 172106
rect 393320 172042 393372 172048
rect 393332 169114 393360 172042
rect 393320 169108 393372 169114
rect 393320 169050 393372 169056
rect 393136 167136 393188 167142
rect 393136 167078 393188 167084
rect 393136 111104 393188 111110
rect 393136 111046 393188 111052
rect 393148 100774 393176 111046
rect 393136 100768 393188 100774
rect 393136 100710 393188 100716
rect 393044 44940 393096 44946
rect 393044 44882 393096 44888
rect 392860 44872 392912 44878
rect 392860 44814 392912 44820
rect 393976 39982 394004 295190
rect 394240 289264 394292 289270
rect 394240 289206 394292 289212
rect 394148 289196 394200 289202
rect 394148 289138 394200 289144
rect 394056 289128 394108 289134
rect 394056 289070 394108 289076
rect 393964 39976 394016 39982
rect 393964 39918 394016 39924
rect 394068 36854 394096 289070
rect 394160 36990 394188 289138
rect 394148 36984 394200 36990
rect 394148 36926 394200 36932
rect 394252 36922 394280 289206
rect 394344 42702 394372 295258
rect 394424 253972 394476 253978
rect 394424 253914 394476 253920
rect 394436 245206 394464 253914
rect 394424 245200 394476 245206
rect 394424 245142 394476 245148
rect 395252 174004 395304 174010
rect 395252 173946 395304 173952
rect 395264 172106 395292 173946
rect 395252 172100 395304 172106
rect 395252 172042 395304 172048
rect 394516 163464 394568 163470
rect 394516 163406 394568 163412
rect 394424 138032 394476 138038
rect 394424 137974 394476 137980
rect 394436 111858 394464 137974
rect 394528 137426 394556 163406
rect 394516 137420 394568 137426
rect 394516 137362 394568 137368
rect 394516 115592 394568 115598
rect 394516 115534 394568 115540
rect 394424 111852 394476 111858
rect 394424 111794 394476 111800
rect 394528 100026 394556 115534
rect 394516 100020 394568 100026
rect 394516 99962 394568 99968
rect 394332 42696 394384 42702
rect 394332 42638 394384 42644
rect 394240 36916 394292 36922
rect 394240 36858 394292 36864
rect 394056 36848 394108 36854
rect 394056 36790 394108 36796
rect 392676 3800 392728 3806
rect 392676 3742 392728 3748
rect 395356 3738 395384 300766
rect 395712 300756 395764 300762
rect 395712 300698 395764 300704
rect 395528 300552 395580 300558
rect 395528 300494 395580 300500
rect 395436 300212 395488 300218
rect 395436 300154 395488 300160
rect 395448 47530 395476 300154
rect 395540 48142 395568 300494
rect 395620 300280 395672 300286
rect 395620 300222 395672 300228
rect 395632 48278 395660 300222
rect 395724 50182 395752 300698
rect 395804 300416 395856 300422
rect 395804 300358 395856 300364
rect 395816 50250 395844 300358
rect 397092 292528 397144 292534
rect 397092 292470 397144 292476
rect 396724 291712 396776 291718
rect 396724 291654 396776 291660
rect 395896 239420 395948 239426
rect 395896 239362 395948 239368
rect 395908 227798 395936 239362
rect 395896 227792 395948 227798
rect 395896 227734 395948 227740
rect 395896 206304 395948 206310
rect 395896 206246 395948 206252
rect 395908 199442 395936 206246
rect 395896 199436 395948 199442
rect 395896 199378 395948 199384
rect 395896 147688 395948 147694
rect 395896 147630 395948 147636
rect 395908 138038 395936 147630
rect 395896 138032 395948 138038
rect 395896 137974 395948 137980
rect 395896 125520 395948 125526
rect 395896 125462 395948 125468
rect 395908 115598 395936 125462
rect 395988 115932 396040 115938
rect 395988 115874 396040 115880
rect 395896 115592 395948 115598
rect 395896 115534 395948 115540
rect 396000 113218 396028 115874
rect 395988 113212 396040 113218
rect 395988 113154 396040 113160
rect 395804 50244 395856 50250
rect 395804 50186 395856 50192
rect 395712 50176 395764 50182
rect 395712 50118 395764 50124
rect 395620 48272 395672 48278
rect 395620 48214 395672 48220
rect 395528 48136 395580 48142
rect 395528 48078 395580 48084
rect 395436 47524 395488 47530
rect 395436 47466 395488 47472
rect 396736 6866 396764 291654
rect 396908 289604 396960 289610
rect 396908 289546 396960 289552
rect 396816 289332 396868 289338
rect 396816 289274 396868 289280
rect 396828 37058 396856 289274
rect 396920 37194 396948 289546
rect 397000 289536 397052 289542
rect 397000 289478 397052 289484
rect 396908 37188 396960 37194
rect 396908 37130 396960 37136
rect 397012 37126 397040 289478
rect 397104 40050 397132 292470
rect 397184 270156 397236 270162
rect 397184 270098 397236 270104
rect 397196 253978 397224 270098
rect 397184 253972 397236 253978
rect 397184 253914 397236 253920
rect 397184 229152 397236 229158
rect 397184 229094 397236 229100
rect 397196 214606 397224 229094
rect 397184 214600 397236 214606
rect 397184 214542 397236 214548
rect 397276 182436 397328 182442
rect 397276 182378 397328 182384
rect 397288 175982 397316 182378
rect 397368 182164 397420 182170
rect 397368 182106 397420 182112
rect 397276 175976 397328 175982
rect 397276 175918 397328 175924
rect 397380 174010 397408 182106
rect 397368 174004 397420 174010
rect 397368 173946 397420 173952
rect 397184 158704 397236 158710
rect 397184 158646 397236 158652
rect 397196 125526 397224 158646
rect 397184 125520 397236 125526
rect 397184 125462 397236 125468
rect 397368 115252 397420 115258
rect 397368 115194 397420 115200
rect 397380 111110 397408 115194
rect 397368 111104 397420 111110
rect 397368 111046 397420 111052
rect 398116 47938 398144 303146
rect 401048 303136 401100 303142
rect 401048 303078 401100 303084
rect 400956 303068 401008 303074
rect 400956 303010 401008 303016
rect 398194 302832 398250 302841
rect 398194 302767 398250 302776
rect 400864 302796 400916 302802
rect 398104 47932 398156 47938
rect 398104 47874 398156 47880
rect 398208 47598 398236 302767
rect 400864 302738 400916 302744
rect 398380 300688 398432 300694
rect 398380 300630 398432 300636
rect 398288 300484 398340 300490
rect 398288 300426 398340 300432
rect 398300 48074 398328 300426
rect 398288 48068 398340 48074
rect 398288 48010 398340 48016
rect 398392 48006 398420 300630
rect 399484 295180 399536 295186
rect 399484 295122 399536 295128
rect 398472 192908 398524 192914
rect 398472 192850 398524 192856
rect 398484 152522 398512 192850
rect 398472 152516 398524 152522
rect 398472 152458 398524 152464
rect 398380 48000 398432 48006
rect 398380 47942 398432 47948
rect 398196 47592 398248 47598
rect 398196 47534 398248 47540
rect 397092 40044 397144 40050
rect 397092 39986 397144 39992
rect 399496 39914 399524 295122
rect 399760 293344 399812 293350
rect 399760 293286 399812 293292
rect 399668 289468 399720 289474
rect 399668 289410 399720 289416
rect 399576 289400 399628 289406
rect 399576 289342 399628 289348
rect 399484 39908 399536 39914
rect 399484 39850 399536 39856
rect 397000 37120 397052 37126
rect 397000 37062 397052 37068
rect 396816 37052 396868 37058
rect 396816 36994 396868 37000
rect 399588 36514 399616 289342
rect 399680 37262 399708 289410
rect 399772 45558 399800 293286
rect 399852 289672 399904 289678
rect 399852 289614 399904 289620
rect 399864 47462 399892 289614
rect 400220 276684 400272 276690
rect 400220 276626 400272 276632
rect 400232 270162 400260 276626
rect 400220 270156 400272 270162
rect 400220 270098 400272 270104
rect 399944 213240 399996 213246
rect 399944 213182 399996 213188
rect 399956 207670 399984 213182
rect 399944 207664 399996 207670
rect 399944 207606 399996 207612
rect 400772 196648 400824 196654
rect 400772 196590 400824 196596
rect 400784 192914 400812 196590
rect 400772 192908 400824 192914
rect 400772 192850 400824 192856
rect 400220 150544 400272 150550
rect 400220 150486 400272 150492
rect 399944 150476 399996 150482
rect 399944 150418 399996 150424
rect 399956 116006 399984 150418
rect 400232 147694 400260 150486
rect 400220 147688 400272 147694
rect 400220 147630 400272 147636
rect 400220 121440 400272 121446
rect 400220 121382 400272 121388
rect 400232 118810 400260 121382
rect 400140 118782 400260 118810
rect 399944 116000 399996 116006
rect 399944 115942 399996 115948
rect 400140 115258 400168 118782
rect 400128 115252 400180 115258
rect 400128 115194 400180 115200
rect 399852 47456 399904 47462
rect 399852 47398 399904 47404
rect 399760 45552 399812 45558
rect 399760 45494 399812 45500
rect 399668 37256 399720 37262
rect 399668 37198 399720 37204
rect 399576 36508 399628 36514
rect 399576 36450 399628 36456
rect 400876 33114 400904 302738
rect 400968 47666 400996 303010
rect 401060 47734 401088 303078
rect 401152 47802 401180 303554
rect 401324 303340 401376 303346
rect 401324 303282 401376 303288
rect 401232 303272 401284 303278
rect 401232 303214 401284 303220
rect 401244 47870 401272 303214
rect 401336 50590 401364 303282
rect 402244 289740 402296 289746
rect 402244 289682 402296 289688
rect 401416 178696 401468 178702
rect 401416 178638 401468 178644
rect 401428 169046 401456 178638
rect 401416 169040 401468 169046
rect 401416 168982 401468 168988
rect 401600 163600 401652 163606
rect 401600 163542 401652 163548
rect 401416 161492 401468 161498
rect 401416 161434 401468 161440
rect 401428 150482 401456 161434
rect 401612 158778 401640 163542
rect 401600 158772 401652 158778
rect 401600 158714 401652 158720
rect 401416 150476 401468 150482
rect 401416 150418 401468 150424
rect 401324 50584 401376 50590
rect 401324 50526 401376 50532
rect 401232 47864 401284 47870
rect 401232 47806 401284 47812
rect 401140 47796 401192 47802
rect 401140 47738 401192 47744
rect 401048 47728 401100 47734
rect 401048 47670 401100 47676
rect 400956 47660 401008 47666
rect 400956 47602 401008 47608
rect 402256 33998 402284 289682
rect 402334 289232 402390 289241
rect 402334 289167 402390 289176
rect 402348 34066 402376 289167
rect 402518 289096 402574 289105
rect 402518 289031 402574 289040
rect 402428 199436 402480 199442
rect 402428 199378 402480 199384
rect 402440 182442 402468 199378
rect 402428 182436 402480 182442
rect 402428 182378 402480 182384
rect 402428 160132 402480 160138
rect 402428 160074 402480 160080
rect 402440 150550 402468 160074
rect 402428 150544 402480 150550
rect 402428 150486 402480 150492
rect 402336 34060 402388 34066
rect 402336 34002 402388 34008
rect 402244 33992 402296 33998
rect 402244 33934 402296 33940
rect 402532 33794 402560 289031
rect 403624 286476 403676 286482
rect 403624 286418 403676 286424
rect 402980 212492 403032 212498
rect 402980 212434 403032 212440
rect 402992 206378 403020 212434
rect 402980 206372 403032 206378
rect 402980 206314 403032 206320
rect 402520 33788 402572 33794
rect 402520 33730 402572 33736
rect 400864 33108 400916 33114
rect 400864 33050 400916 33056
rect 403636 20670 403664 286418
rect 403728 50833 403756 305730
rect 403808 303408 403860 303414
rect 403808 303350 403860 303356
rect 403714 50824 403770 50833
rect 403714 50759 403770 50768
rect 403820 50386 403848 303350
rect 403912 50697 403940 305798
rect 406382 305759 406438 305768
rect 404084 303544 404136 303550
rect 404084 303486 404136 303492
rect 403992 303476 404044 303482
rect 403992 303418 404044 303424
rect 403898 50688 403954 50697
rect 403898 50623 403954 50632
rect 404004 50522 404032 303418
rect 403992 50516 404044 50522
rect 403992 50458 404044 50464
rect 404096 50454 404124 303486
rect 405096 289808 405148 289814
rect 405096 289750 405148 289756
rect 405004 289060 405056 289066
rect 405004 289002 405056 289008
rect 404452 167748 404504 167754
rect 404452 167690 404504 167696
rect 404176 165232 404228 165238
rect 404176 165174 404228 165180
rect 404188 111790 404216 165174
rect 404464 163470 404492 167690
rect 404452 163464 404504 163470
rect 404452 163406 404504 163412
rect 404360 163260 404412 163266
rect 404360 163202 404412 163208
rect 404372 160138 404400 163202
rect 404360 160132 404412 160138
rect 404360 160074 404412 160080
rect 404176 111784 404228 111790
rect 404176 111726 404228 111732
rect 404084 50448 404136 50454
rect 404084 50390 404136 50396
rect 403808 50380 403860 50386
rect 403808 50322 403860 50328
rect 405016 33862 405044 289002
rect 405108 34134 405136 289750
rect 405188 286340 405240 286346
rect 405188 286282 405240 286288
rect 405096 34128 405148 34134
rect 405096 34070 405148 34076
rect 405200 33930 405228 286282
rect 405280 245676 405332 245682
rect 405280 245618 405332 245624
rect 405292 229158 405320 245618
rect 405280 229152 405332 229158
rect 405280 229094 405332 229100
rect 405556 183932 405608 183938
rect 405556 183874 405608 183880
rect 405568 182238 405596 183874
rect 405556 182232 405608 182238
rect 405556 182174 405608 182180
rect 405556 163192 405608 163198
rect 405556 163134 405608 163140
rect 405568 161498 405596 163134
rect 405556 161492 405608 161498
rect 405556 161434 405608 161440
rect 405280 127560 405332 127566
rect 405280 127502 405332 127508
rect 405292 121514 405320 127502
rect 405280 121508 405332 121514
rect 405280 121450 405332 121456
rect 405188 33924 405240 33930
rect 405188 33866 405240 33872
rect 405004 33856 405056 33862
rect 405004 33798 405056 33804
rect 403624 20664 403676 20670
rect 403624 20606 403676 20612
rect 396724 6860 396776 6866
rect 396724 6802 396776 6808
rect 395344 3732 395396 3738
rect 395344 3674 395396 3680
rect 406396 3641 406424 305759
rect 406488 51921 406516 305934
rect 406750 305895 406806 305904
rect 406566 305688 406622 305697
rect 406566 305623 406622 305632
rect 406474 51912 406530 51921
rect 406474 51847 406530 51856
rect 406580 50425 406608 305623
rect 406660 280832 406712 280838
rect 406660 280774 406712 280780
rect 406672 276690 406700 280774
rect 406660 276684 406712 276690
rect 406660 276626 406712 276632
rect 406660 165640 406712 165646
rect 406660 165582 406712 165588
rect 406672 100706 406700 165582
rect 406660 100700 406712 100706
rect 406660 100642 406712 100648
rect 406764 50561 406792 305895
rect 410524 304496 410576 304502
rect 410524 304438 410576 304444
rect 407948 304360 408000 304366
rect 407948 304302 408000 304308
rect 407856 286408 407908 286414
rect 407762 286376 407818 286385
rect 407856 286350 407908 286356
rect 407762 286311 407818 286320
rect 406936 215348 406988 215354
rect 406936 215290 406988 215296
rect 406948 212498 406976 215290
rect 406936 212492 406988 212498
rect 406936 212434 406988 212440
rect 407120 187740 407172 187746
rect 407120 187682 407172 187688
rect 407132 183938 407160 187682
rect 407120 183932 407172 183938
rect 407120 183874 407172 183880
rect 407672 165436 407724 165442
rect 407672 165378 407724 165384
rect 407684 163606 407712 165378
rect 407672 163600 407724 163606
rect 407672 163542 407724 163548
rect 406844 155304 406896 155310
rect 406844 155246 406896 155252
rect 406856 127566 406884 155246
rect 406844 127560 406896 127566
rect 406844 127502 406896 127508
rect 406750 50552 406806 50561
rect 406750 50487 406806 50496
rect 406566 50416 406622 50425
rect 406566 50351 406622 50360
rect 407776 3777 407804 286311
rect 407762 3768 407818 3777
rect 407762 3703 407818 3712
rect 407868 3670 407896 286350
rect 407960 44810 407988 304302
rect 409144 254584 409196 254590
rect 409144 254526 409196 254532
rect 408776 220380 408828 220386
rect 408776 220322 408828 220328
rect 408788 213246 408816 220322
rect 408776 213240 408828 213246
rect 408776 213182 408828 213188
rect 409156 206310 409184 254526
rect 409144 206304 409196 206310
rect 409144 206246 409196 206252
rect 408500 199504 408552 199510
rect 408500 199446 408552 199452
rect 408512 196654 408540 199446
rect 408500 196648 408552 196654
rect 408500 196590 408552 196596
rect 408040 165776 408092 165782
rect 408040 165718 408092 165724
rect 408052 69018 408080 165718
rect 409880 165504 409932 165510
rect 409880 165446 409932 165452
rect 408500 165368 408552 165374
rect 408500 165310 408552 165316
rect 408512 163198 408540 165310
rect 409512 165300 409564 165306
rect 409512 165242 409564 165248
rect 409236 165164 409288 165170
rect 409236 165106 409288 165112
rect 409142 163432 409198 163441
rect 409142 163367 409198 163376
rect 408500 163192 408552 163198
rect 408500 163134 408552 163140
rect 409156 89690 409184 163367
rect 409248 132462 409276 165106
rect 409328 165096 409380 165102
rect 409328 165038 409380 165044
rect 409340 143546 409368 165038
rect 409420 164960 409472 164966
rect 409420 164902 409472 164908
rect 409432 154562 409460 164902
rect 409524 155310 409552 165242
rect 409892 163266 409920 165446
rect 409880 163260 409932 163266
rect 409880 163202 409932 163208
rect 409512 155304 409564 155310
rect 409512 155246 409564 155252
rect 409420 154556 409472 154562
rect 409420 154498 409472 154504
rect 409328 143540 409380 143546
rect 409328 143482 409380 143488
rect 409236 132456 409288 132462
rect 409236 132398 409288 132404
rect 409144 89684 409196 89690
rect 409144 89626 409196 89632
rect 408040 69012 408092 69018
rect 408040 68954 408092 68960
rect 407948 44804 408000 44810
rect 407948 44746 408000 44752
rect 410536 44742 410564 304438
rect 431224 273964 431276 273970
rect 431224 273906 431276 273912
rect 420184 272536 420236 272542
rect 420184 272478 420236 272484
rect 420196 266422 420224 272478
rect 431236 266422 431264 273906
rect 413284 266416 413336 266422
rect 413284 266358 413336 266364
rect 420184 266416 420236 266422
rect 420184 266358 420236 266364
rect 427820 266416 427872 266422
rect 427820 266358 427872 266364
rect 431224 266416 431276 266422
rect 431224 266358 431276 266364
rect 411260 249076 411312 249082
rect 411260 249018 411312 249024
rect 411272 245682 411300 249018
rect 411260 245676 411312 245682
rect 411260 245618 411312 245624
rect 413296 239426 413324 266358
rect 427832 259010 427860 266358
rect 425704 259004 425756 259010
rect 425704 258946 425756 258952
rect 427820 259004 427872 259010
rect 427820 258946 427872 258952
rect 424140 257372 424192 257378
rect 424140 257314 424192 257320
rect 424152 254590 424180 257314
rect 424324 255332 424376 255338
rect 424324 255274 424376 255280
rect 424140 254584 424192 254590
rect 424140 254526 424192 254532
rect 418804 250504 418856 250510
rect 418804 250446 418856 250452
rect 413284 239420 413336 239426
rect 413284 239362 413336 239368
rect 417424 237448 417476 237454
rect 417424 237390 417476 237396
rect 416044 233912 416096 233918
rect 416044 233854 416096 233860
rect 416056 227050 416084 233854
rect 411260 227044 411312 227050
rect 411260 226986 411312 226992
rect 416044 227044 416096 227050
rect 416044 226986 416096 226992
rect 411272 220386 411300 226986
rect 416780 223780 416832 223786
rect 416780 223722 416832 223728
rect 411260 220380 411312 220386
rect 411260 220322 411312 220328
rect 416792 220114 416820 223722
rect 411260 220108 411312 220114
rect 411260 220050 411312 220056
rect 416780 220108 416832 220114
rect 416780 220050 416832 220056
rect 411272 215354 411300 220050
rect 417436 215354 417464 237390
rect 418816 233918 418844 250446
rect 422944 246356 422996 246362
rect 422944 246298 422996 246304
rect 420920 244248 420972 244254
rect 420920 244190 420972 244196
rect 420932 239902 420960 244190
rect 419540 239896 419592 239902
rect 419540 239838 419592 239844
rect 420920 239896 420972 239902
rect 420920 239838 420972 239844
rect 419552 237454 419580 239838
rect 419540 237448 419592 237454
rect 419540 237390 419592 237396
rect 422956 235686 422984 246298
rect 424336 244322 424364 255274
rect 425716 250510 425744 258946
rect 429568 258392 429620 258398
rect 429568 258334 429620 258340
rect 429580 255338 429608 258334
rect 429568 255332 429620 255338
rect 429568 255274 429620 255280
rect 426348 251864 426400 251870
rect 426348 251806 426400 251812
rect 425704 250504 425756 250510
rect 425704 250446 425756 250452
rect 426360 249082 426388 251806
rect 432616 249762 432644 332590
rect 432708 331294 432736 369650
rect 435376 362914 435404 407118
rect 436744 396092 436796 396098
rect 436744 396034 436796 396040
rect 435364 362908 435416 362914
rect 435364 362850 435416 362856
rect 436756 362846 436784 396034
rect 439516 375222 439544 418746
rect 443644 417444 443696 417450
rect 443644 417386 443696 417392
rect 442908 382288 442960 382294
rect 442908 382230 442960 382236
rect 439596 375420 439648 375426
rect 439596 375362 439648 375368
rect 439504 375216 439556 375222
rect 439504 375158 439556 375164
rect 436744 362840 436796 362846
rect 436744 362782 436796 362788
rect 439608 361554 439636 375362
rect 439596 361548 439648 361554
rect 439596 361490 439648 361496
rect 439780 358896 439832 358902
rect 439780 358838 439832 358844
rect 433984 358828 434036 358834
rect 433984 358770 434036 358776
rect 433708 350464 433760 350470
rect 433708 350406 433760 350412
rect 433720 346390 433748 350406
rect 433708 346384 433760 346390
rect 433708 346326 433760 346332
rect 432972 340808 433024 340814
rect 432972 340750 433024 340756
rect 432788 340264 432840 340270
rect 432788 340206 432840 340212
rect 432696 331288 432748 331294
rect 432696 331230 432748 331236
rect 432800 319870 432828 340206
rect 432880 336932 432932 336938
rect 432880 336874 432932 336880
rect 432892 328438 432920 336874
rect 432984 330614 433012 340750
rect 433248 339448 433300 339454
rect 433248 339390 433300 339396
rect 433260 335354 433288 339390
rect 433260 335326 433472 335354
rect 433444 334082 433472 335326
rect 433996 334801 434024 358770
rect 435456 357468 435508 357474
rect 435456 357410 435508 357416
rect 434076 354272 434128 354278
rect 434076 354214 434128 354220
rect 433982 334792 434038 334801
rect 433982 334727 434038 334736
rect 434088 334558 434116 354214
rect 434168 351892 434220 351898
rect 434168 351834 434220 351840
rect 434180 338094 434208 351834
rect 434260 342236 434312 342242
rect 434260 342178 434312 342184
rect 434168 338088 434220 338094
rect 434168 338030 434220 338036
rect 434076 334552 434128 334558
rect 434076 334494 434128 334500
rect 433432 334076 433484 334082
rect 433432 334018 433484 334024
rect 434272 334014 434300 342178
rect 434628 335096 434680 335102
rect 434628 335038 434680 335044
rect 434260 334008 434312 334014
rect 434260 333950 434312 333956
rect 434640 332466 434668 335038
rect 435364 334076 435416 334082
rect 435364 334018 435416 334024
rect 434640 332438 434760 332466
rect 433432 332036 433484 332042
rect 433432 331978 433484 331984
rect 433444 330857 433472 331978
rect 434444 331900 434496 331906
rect 434444 331842 434496 331848
rect 433430 330848 433486 330857
rect 433430 330783 433486 330792
rect 432972 330608 433024 330614
rect 432972 330550 433024 330556
rect 432880 328432 432932 328438
rect 432880 328374 432932 328380
rect 433800 328432 433852 328438
rect 433800 328374 433852 328380
rect 433812 323542 433840 328374
rect 434456 326913 434484 331842
rect 434732 329798 434760 332438
rect 435088 331220 435140 331226
rect 435088 331162 435140 331168
rect 434720 329792 434772 329798
rect 434720 329734 434772 329740
rect 435100 328438 435128 331162
rect 435088 328432 435140 328438
rect 435088 328374 435140 328380
rect 434442 326904 434498 326913
rect 434442 326839 434498 326848
rect 434076 324352 434128 324358
rect 434076 324294 434128 324300
rect 433800 323536 433852 323542
rect 433800 323478 433852 323484
rect 434088 322969 434116 324294
rect 434074 322960 434130 322969
rect 434074 322895 434130 322904
rect 433984 322244 434036 322250
rect 433984 322186 434036 322192
rect 432788 319864 432840 319870
rect 432788 319806 432840 319812
rect 433524 319252 433576 319258
rect 433524 319194 433576 319200
rect 433536 319025 433564 319194
rect 433522 319016 433578 319025
rect 433522 318951 433578 318960
rect 433996 311137 434024 322186
rect 434260 315104 434312 315110
rect 434258 315072 434260 315081
rect 434312 315072 434314 315081
rect 434258 315007 434314 315016
rect 433982 311128 434038 311137
rect 433982 311063 434038 311072
rect 433892 307760 433944 307766
rect 433892 307702 433944 307708
rect 433904 307193 433932 307702
rect 433890 307184 433946 307193
rect 433890 307119 433946 307128
rect 432696 288992 432748 288998
rect 432696 288934 432748 288940
rect 432708 257378 432736 288934
rect 433984 271312 434036 271318
rect 433984 271254 434036 271260
rect 433996 258398 434024 271254
rect 435376 259418 435404 334018
rect 435468 319258 435496 357410
rect 439688 356176 439740 356182
rect 439688 356118 439740 356124
rect 436928 356108 436980 356114
rect 436928 356050 436980 356056
rect 435640 346384 435692 346390
rect 435640 346326 435692 346332
rect 435652 341222 435680 346326
rect 435640 341216 435692 341222
rect 435640 341158 435692 341164
rect 435732 334552 435784 334558
rect 435732 334494 435784 334500
rect 435640 329112 435692 329118
rect 435640 329054 435692 329060
rect 435652 322386 435680 329054
rect 435744 327078 435772 334494
rect 436836 334076 436888 334082
rect 436836 334018 436888 334024
rect 436376 333940 436428 333946
rect 436376 333882 436428 333888
rect 436388 331158 436416 333882
rect 436376 331152 436428 331158
rect 436376 331094 436428 331100
rect 436008 330608 436060 330614
rect 436008 330550 436060 330556
rect 436020 328386 436048 330550
rect 436744 330540 436796 330546
rect 436744 330482 436796 330488
rect 436020 328358 436140 328386
rect 435732 327072 435784 327078
rect 435732 327014 435784 327020
rect 436112 322930 436140 328358
rect 436192 323536 436244 323542
rect 436192 323478 436244 323484
rect 436100 322924 436152 322930
rect 436100 322866 436152 322872
rect 435640 322380 435692 322386
rect 435640 322322 435692 322328
rect 436204 319734 436232 323478
rect 436192 319728 436244 319734
rect 436192 319670 436244 319676
rect 435456 319252 435508 319258
rect 435456 319194 435508 319200
rect 435456 299396 435508 299402
rect 435456 299338 435508 299344
rect 435468 288998 435496 299338
rect 435456 288992 435508 288998
rect 435456 288934 435508 288940
rect 436652 283688 436704 283694
rect 436652 283630 436704 283636
rect 436664 280838 436692 283630
rect 436652 280832 436704 280838
rect 436652 280774 436704 280780
rect 435548 275052 435600 275058
rect 435548 274994 435600 275000
rect 435560 272542 435588 274994
rect 435548 272536 435600 272542
rect 435548 272478 435600 272484
rect 435364 259412 435416 259418
rect 435364 259354 435416 259360
rect 433984 258392 434036 258398
rect 433984 258334 434036 258340
rect 432696 257372 432748 257378
rect 432696 257314 432748 257320
rect 435364 252952 435416 252958
rect 435364 252894 435416 252900
rect 432604 249756 432656 249762
rect 432604 249698 432656 249704
rect 426348 249076 426400 249082
rect 426348 249018 426400 249024
rect 435376 246362 435404 252894
rect 436008 248532 436060 248538
rect 436008 248474 436060 248480
rect 435364 246356 435416 246362
rect 435364 246298 435416 246304
rect 436020 244934 436048 248474
rect 429844 244928 429896 244934
rect 429844 244870 429896 244876
rect 436008 244928 436060 244934
rect 436008 244870 436060 244876
rect 424324 244316 424376 244322
rect 424324 244258 424376 244264
rect 420184 235680 420236 235686
rect 420184 235622 420236 235628
rect 422944 235680 422996 235686
rect 422944 235622 422996 235628
rect 418804 233912 418856 233918
rect 418804 233854 418856 233860
rect 420196 223786 420224 235622
rect 427084 232552 427136 232558
rect 427084 232494 427136 232500
rect 422944 230036 422996 230042
rect 422944 229978 422996 229984
rect 421564 224256 421616 224262
rect 421564 224198 421616 224204
rect 420184 223780 420236 223786
rect 420184 223722 420236 223728
rect 417516 216980 417568 216986
rect 417516 216922 417568 216928
rect 411260 215348 411312 215354
rect 411260 215290 411312 215296
rect 413284 215348 413336 215354
rect 413284 215290 413336 215296
rect 417424 215348 417476 215354
rect 417424 215290 417476 215296
rect 413296 205630 413324 215290
rect 411904 205624 411956 205630
rect 411904 205566 411956 205572
rect 413284 205624 413336 205630
rect 413284 205566 413336 205572
rect 411916 193798 411944 205566
rect 417528 199442 417556 216922
rect 421576 199510 421604 224198
rect 422956 216986 422984 229978
rect 427096 224262 427124 232494
rect 429856 230042 429884 244870
rect 434904 235476 434956 235482
rect 434904 235418 434956 235424
rect 434916 232558 434944 235418
rect 434904 232552 434956 232558
rect 434904 232494 434956 232500
rect 435456 230444 435508 230450
rect 435456 230386 435508 230392
rect 429844 230036 429896 230042
rect 429844 229978 429896 229984
rect 427084 224256 427136 224262
rect 427084 224198 427136 224204
rect 435468 220794 435496 230386
rect 436756 227730 436784 330482
rect 436848 270502 436876 334018
rect 436940 315110 436968 356050
rect 438124 341216 438176 341222
rect 438124 341158 438176 341164
rect 437020 338088 437072 338094
rect 437020 338030 437072 338036
rect 437032 323678 437060 338030
rect 437388 333940 437440 333946
rect 437388 333882 437440 333888
rect 437400 332466 437428 333882
rect 437400 332438 437520 332466
rect 437388 328432 437440 328438
rect 437388 328374 437440 328380
rect 437296 327072 437348 327078
rect 437296 327014 437348 327020
rect 437020 323672 437072 323678
rect 437020 323614 437072 323620
rect 437308 320210 437336 327014
rect 437400 325694 437428 328374
rect 437492 327078 437520 332438
rect 437480 327072 437532 327078
rect 437480 327014 437532 327020
rect 437400 325666 437520 325694
rect 437296 320204 437348 320210
rect 437296 320146 437348 320152
rect 437492 319666 437520 325666
rect 438136 325174 438164 341158
rect 439596 334620 439648 334626
rect 439596 334562 439648 334568
rect 439504 331288 439556 331294
rect 439504 331230 439556 331236
rect 438308 331152 438360 331158
rect 438308 331094 438360 331100
rect 438216 329792 438268 329798
rect 438216 329734 438268 329740
rect 438124 325168 438176 325174
rect 438124 325110 438176 325116
rect 437480 319660 437532 319666
rect 437480 319602 437532 319608
rect 438228 319462 438256 329734
rect 438320 321570 438348 331094
rect 438768 327140 438820 327146
rect 438768 327082 438820 327088
rect 438308 321564 438360 321570
rect 438308 321506 438360 321512
rect 438216 319456 438268 319462
rect 438216 319398 438268 319404
rect 436928 315104 436980 315110
rect 436928 315046 436980 315052
rect 438124 306060 438176 306066
rect 438124 306002 438176 306008
rect 436928 287020 436980 287026
rect 436928 286962 436980 286968
rect 436940 271318 436968 286962
rect 438136 273970 438164 306002
rect 438216 305040 438268 305046
rect 438216 304982 438268 304988
rect 438228 299402 438256 304982
rect 438216 299396 438268 299402
rect 438216 299338 438268 299344
rect 438124 273964 438176 273970
rect 438124 273906 438176 273912
rect 436928 271312 436980 271318
rect 436928 271254 436980 271260
rect 436836 270496 436888 270502
rect 436836 270438 436888 270444
rect 438124 262744 438176 262750
rect 438124 262686 438176 262692
rect 437480 257372 437532 257378
rect 437480 257314 437532 257320
rect 437492 252958 437520 257314
rect 437480 252952 437532 252958
rect 437480 252894 437532 252900
rect 438136 251870 438164 262686
rect 438124 251864 438176 251870
rect 438124 251806 438176 251812
rect 436744 227724 436796 227730
rect 436744 227666 436796 227672
rect 438124 224256 438176 224262
rect 438124 224198 438176 224204
rect 433984 220788 434036 220794
rect 433984 220730 434036 220736
rect 435456 220788 435508 220794
rect 435456 220730 435508 220736
rect 422944 216980 422996 216986
rect 422944 216922 422996 216928
rect 425704 211812 425756 211818
rect 425704 211754 425756 211760
rect 425716 201482 425744 211754
rect 432328 202836 432380 202842
rect 432328 202778 432380 202784
rect 422944 201476 422996 201482
rect 422944 201418 422996 201424
rect 425704 201476 425756 201482
rect 425704 201418 425756 201424
rect 421564 199504 421616 199510
rect 421564 199446 421616 199452
rect 417516 199436 417568 199442
rect 417516 199378 417568 199384
rect 410616 193792 410668 193798
rect 410616 193734 410668 193740
rect 411904 193792 411956 193798
rect 411904 193734 411956 193740
rect 410628 187746 410656 193734
rect 410616 187740 410668 187746
rect 410616 187682 410668 187688
rect 422956 187134 422984 201418
rect 429936 196988 429988 196994
rect 429936 196930 429988 196936
rect 429844 193996 429896 194002
rect 429844 193938 429896 193944
rect 416044 187128 416096 187134
rect 416044 187070 416096 187076
rect 422944 187128 422996 187134
rect 422944 187070 422996 187076
rect 416056 178702 416084 187070
rect 428464 185496 428516 185502
rect 428464 185438 428516 185444
rect 416044 178696 416096 178702
rect 416044 178638 416096 178644
rect 428476 175982 428504 185438
rect 426440 175976 426492 175982
rect 426440 175918 426492 175924
rect 428464 175976 428516 175982
rect 428464 175918 428516 175924
rect 422944 175908 422996 175914
rect 422944 175850 422996 175856
rect 422300 169788 422352 169794
rect 422300 169730 422352 169736
rect 419724 167884 419776 167890
rect 419724 167826 419776 167832
rect 416228 167816 416280 167822
rect 416228 167758 416280 167764
rect 411904 167680 411956 167686
rect 411904 167622 411956 167628
rect 411916 165714 411944 167622
rect 416240 165782 416268 167758
rect 416228 165776 416280 165782
rect 416228 165718 416280 165724
rect 411904 165708 411956 165714
rect 411904 165650 411956 165656
rect 411916 164914 411944 165650
rect 416240 164914 416268 165718
rect 419736 165034 419764 167826
rect 422312 165730 422340 169730
rect 422956 167754 422984 175850
rect 426452 173942 426480 175918
rect 429856 175914 429884 193938
rect 429948 185502 429976 196930
rect 432340 194002 432368 202778
rect 433996 198762 434024 220730
rect 435364 219496 435416 219502
rect 435364 219438 435416 219444
rect 435376 202842 435404 219438
rect 438136 212498 438164 224198
rect 436744 212492 436796 212498
rect 436744 212434 436796 212440
rect 438124 212492 438176 212498
rect 438124 212434 438176 212440
rect 435364 202836 435416 202842
rect 435364 202778 435416 202784
rect 432972 198756 433024 198762
rect 432972 198698 433024 198704
rect 433984 198756 434036 198762
rect 433984 198698 434036 198704
rect 432984 196994 433012 198698
rect 436756 197402 436784 212434
rect 433984 197396 434036 197402
rect 433984 197338 434036 197344
rect 436744 197396 436796 197402
rect 436744 197338 436796 197344
rect 432972 196988 433024 196994
rect 432972 196930 433024 196936
rect 432328 193996 432380 194002
rect 432328 193938 432380 193944
rect 429936 185496 429988 185502
rect 429936 185438 429988 185444
rect 433996 183598 434024 197338
rect 436744 196036 436796 196042
rect 436744 195978 436796 195984
rect 432788 183592 432840 183598
rect 432788 183534 432840 183540
rect 433984 183592 434036 183598
rect 433984 183534 434036 183540
rect 432800 182238 432828 183534
rect 431224 182232 431276 182238
rect 431224 182174 431276 182180
rect 432788 182232 432840 182238
rect 432788 182174 432840 182180
rect 430580 175976 430632 175982
rect 430580 175918 430632 175924
rect 429844 175908 429896 175914
rect 429844 175850 429896 175856
rect 426440 173936 426492 173942
rect 426440 173878 426492 173884
rect 423680 173868 423732 173874
rect 423680 173810 423732 173816
rect 423692 169794 423720 173810
rect 429292 172508 429344 172514
rect 429292 172450 429344 172456
rect 429200 171828 429252 171834
rect 429200 171770 429252 171776
rect 423680 169788 423732 169794
rect 423680 169730 423732 169736
rect 429212 168434 429240 171770
rect 429200 168428 429252 168434
rect 429200 168370 429252 168376
rect 423128 168360 423180 168366
rect 423128 168302 423180 168308
rect 422944 167748 422996 167754
rect 422944 167690 422996 167696
rect 422220 165702 422340 165730
rect 422220 165510 422248 165702
rect 422208 165504 422260 165510
rect 422208 165446 422260 165452
rect 423140 165442 423168 168302
rect 427084 167748 427136 167754
rect 427084 167690 427136 167696
rect 427096 165646 427124 167690
rect 427084 165640 427136 165646
rect 427084 165582 427136 165588
rect 423128 165436 423180 165442
rect 423128 165378 423180 165384
rect 419724 165028 419776 165034
rect 419724 164970 419776 164976
rect 411916 164886 412252 164914
rect 415932 164886 416268 164914
rect 419736 164778 419764 164970
rect 427096 164778 427124 165582
rect 429304 165374 429332 172450
rect 430592 171834 430620 175918
rect 431236 172514 431264 182174
rect 436756 182170 436784 195978
rect 435364 182164 435416 182170
rect 435364 182106 435416 182112
rect 436744 182164 436796 182170
rect 436744 182106 436796 182112
rect 431224 172508 431276 172514
rect 431224 172450 431276 172456
rect 430580 171828 430632 171834
rect 430580 171770 430632 171776
rect 430764 167952 430816 167958
rect 430764 167894 430816 167900
rect 429292 165368 429344 165374
rect 429292 165310 429344 165316
rect 430776 164898 430804 167894
rect 430856 167136 430908 167142
rect 430856 167078 430908 167084
rect 430868 165238 430896 167078
rect 434444 167068 434496 167074
rect 434444 167010 434496 167016
rect 430856 165232 430908 165238
rect 430856 165174 430908 165180
rect 430764 164892 430816 164898
rect 430764 164834 430816 164840
rect 419612 164750 419764 164778
rect 426972 164750 427124 164778
rect 430868 164642 430896 165174
rect 434456 164642 434484 167010
rect 435376 165306 435404 182106
rect 436100 179444 436152 179450
rect 436100 179386 436152 179392
rect 436112 175982 436140 179386
rect 436100 175976 436152 175982
rect 436100 175918 436152 175924
rect 438780 165714 438808 327082
rect 438860 321564 438912 321570
rect 438860 321506 438912 321512
rect 438872 319190 438900 321506
rect 438860 319184 438912 319190
rect 438860 319126 438912 319132
rect 439516 206990 439544 331230
rect 439608 281518 439636 334562
rect 439700 307766 439728 356118
rect 439792 332042 439820 358838
rect 440976 357536 441028 357542
rect 440976 357478 441028 357484
rect 439964 337748 440016 337754
rect 439964 337690 440016 337696
rect 439872 337476 439924 337482
rect 439872 337418 439924 337424
rect 439780 332036 439832 332042
rect 439780 331978 439832 331984
rect 439780 327072 439832 327078
rect 439780 327014 439832 327020
rect 439792 321570 439820 327014
rect 439780 321564 439832 321570
rect 439780 321506 439832 321512
rect 439884 316674 439912 337418
rect 439976 316878 440004 337690
rect 440056 337612 440108 337618
rect 440056 337554 440108 337560
rect 440068 317014 440096 337554
rect 440884 332716 440936 332722
rect 440884 332658 440936 332664
rect 440240 325168 440292 325174
rect 440240 325110 440292 325116
rect 440252 320142 440280 325110
rect 440332 323672 440384 323678
rect 440332 323614 440384 323620
rect 440240 320136 440292 320142
rect 440240 320078 440292 320084
rect 440344 319598 440372 323614
rect 440424 322380 440476 322386
rect 440424 322322 440476 322328
rect 440332 319592 440384 319598
rect 440332 319534 440384 319540
rect 440056 317008 440108 317014
rect 440056 316950 440108 316956
rect 439964 316872 440016 316878
rect 439964 316814 440016 316820
rect 439872 316668 439924 316674
rect 439872 316610 439924 316616
rect 440436 316606 440464 322322
rect 440700 321564 440752 321570
rect 440700 321506 440752 321512
rect 440712 318102 440740 321506
rect 440700 318096 440752 318102
rect 440700 318038 440752 318044
rect 440424 316600 440476 316606
rect 440424 316542 440476 316548
rect 439688 307760 439740 307766
rect 439688 307702 439740 307708
rect 440240 293276 440292 293282
rect 440240 293218 440292 293224
rect 440252 287094 440280 293218
rect 440240 287088 440292 287094
rect 440240 287030 440292 287036
rect 439688 282192 439740 282198
rect 439688 282134 439740 282140
rect 439596 281512 439648 281518
rect 439596 281454 439648 281460
rect 439700 248538 439728 282134
rect 439688 248532 439740 248538
rect 439688 248474 439740 248480
rect 440896 238746 440924 332658
rect 440988 324358 441016 357478
rect 442356 337680 442408 337686
rect 442356 337622 442408 337628
rect 442264 335844 442316 335850
rect 442264 335786 442316 335792
rect 440976 324352 441028 324358
rect 440976 324294 441028 324300
rect 441988 320136 442040 320142
rect 441988 320078 442040 320084
rect 442000 318510 442028 320078
rect 441988 318504 442040 318510
rect 441988 318446 442040 318452
rect 440976 314084 441028 314090
rect 440976 314026 441028 314032
rect 440988 305046 441016 314026
rect 440976 305040 441028 305046
rect 440976 304982 441028 304988
rect 442276 304434 442304 335786
rect 442368 315994 442396 337622
rect 442920 336734 442948 382230
rect 443656 349042 443684 417386
rect 443736 386436 443788 386442
rect 443736 386378 443788 386384
rect 443748 362778 443776 386378
rect 443920 363656 443972 363662
rect 443920 363598 443972 363604
rect 443736 362772 443788 362778
rect 443736 362714 443788 362720
rect 443932 361486 443960 363598
rect 443920 361480 443972 361486
rect 443920 361422 443972 361428
rect 444012 358964 444064 358970
rect 444012 358906 444064 358912
rect 443736 356244 443788 356250
rect 443736 356186 443788 356192
rect 443644 349036 443696 349042
rect 443644 348978 443696 348984
rect 442908 336728 442960 336734
rect 442908 336670 442960 336676
rect 443644 331356 443696 331362
rect 443644 331298 443696 331304
rect 442908 328500 442960 328506
rect 442908 328442 442960 328448
rect 442724 322924 442776 322930
rect 442724 322866 442776 322872
rect 442540 320204 442592 320210
rect 442540 320146 442592 320152
rect 442552 318850 442580 320146
rect 442736 320142 442764 322866
rect 442724 320136 442776 320142
rect 442724 320078 442776 320084
rect 442540 318844 442592 318850
rect 442540 318786 442592 318792
rect 442356 315988 442408 315994
rect 442356 315930 442408 315936
rect 442264 304428 442316 304434
rect 442264 304370 442316 304376
rect 440976 302456 441028 302462
rect 440976 302398 441028 302404
rect 440988 275058 441016 302398
rect 440976 275052 441028 275058
rect 440976 274994 441028 275000
rect 440976 268388 441028 268394
rect 440976 268330 441028 268336
rect 440884 238740 440936 238746
rect 440884 238682 440936 238688
rect 440884 216708 440936 216714
rect 440884 216650 440936 216656
rect 439504 206984 439556 206990
rect 439504 206926 439556 206932
rect 440896 201482 440924 216650
rect 440988 211818 441016 268330
rect 441068 254584 441120 254590
rect 441068 254526 441120 254532
rect 441080 224262 441108 254526
rect 441068 224256 441120 224262
rect 441068 224198 441120 224204
rect 442724 218136 442776 218142
rect 442724 218078 442776 218084
rect 442736 216714 442764 218078
rect 442724 216708 442776 216714
rect 442724 216650 442776 216656
rect 440976 211812 441028 211818
rect 440976 211754 441028 211760
rect 438860 201476 438912 201482
rect 438860 201418 438912 201424
rect 440884 201476 440936 201482
rect 440884 201418 440936 201424
rect 438872 196042 438900 201418
rect 438860 196036 438912 196042
rect 438860 195978 438912 195984
rect 440240 189100 440292 189106
rect 440240 189042 440292 189048
rect 439504 186584 439556 186590
rect 439504 186526 439556 186532
rect 438860 183116 438912 183122
rect 438860 183058 438912 183064
rect 438872 179450 438900 183058
rect 438860 179444 438912 179450
rect 438860 179386 438912 179392
rect 439516 167958 439544 186526
rect 440252 183122 440280 189042
rect 440240 183116 440292 183122
rect 440240 183058 440292 183064
rect 439504 167952 439556 167958
rect 439504 167894 439556 167900
rect 438032 165708 438084 165714
rect 438032 165650 438084 165656
rect 438768 165708 438820 165714
rect 438768 165650 438820 165656
rect 435364 165300 435416 165306
rect 435364 165242 435416 165248
rect 438044 165186 438072 165650
rect 442920 165646 442948 328442
rect 443000 240916 443052 240922
rect 443000 240858 443052 240864
rect 443012 235482 443040 240858
rect 443000 235476 443052 235482
rect 443000 235418 443052 235424
rect 443656 195974 443684 331298
rect 443748 322250 443776 356186
rect 443920 335776 443972 335782
rect 443920 335718 443972 335724
rect 443828 331424 443880 331430
rect 443828 331366 443880 331372
rect 443736 322244 443788 322250
rect 443736 322186 443788 322192
rect 443736 310140 443788 310146
rect 443736 310082 443788 310088
rect 443748 302462 443776 310082
rect 443736 302456 443788 302462
rect 443736 302398 443788 302404
rect 443736 268592 443788 268598
rect 443736 268534 443788 268540
rect 443644 195968 443696 195974
rect 443644 195910 443696 195916
rect 443748 186590 443776 268534
rect 443840 264246 443868 331366
rect 443932 305930 443960 335718
rect 444024 331906 444052 358906
rect 444012 331900 444064 331906
rect 444012 331842 444064 331848
rect 444208 318578 444236 700470
rect 444196 318572 444248 318578
rect 444196 318514 444248 318520
rect 444300 317694 444328 700674
rect 446404 700664 446456 700670
rect 446404 700606 446456 700612
rect 445024 700596 445076 700602
rect 445024 700538 445076 700544
rect 444656 318504 444708 318510
rect 444656 318446 444708 318452
rect 444472 318096 444524 318102
rect 444472 318038 444524 318044
rect 444288 317688 444340 317694
rect 444288 317630 444340 317636
rect 444484 316470 444512 318038
rect 444668 316946 444696 318446
rect 445036 317082 445064 700538
rect 445116 700324 445168 700330
rect 445116 700266 445168 700272
rect 445128 319530 445156 700266
rect 445208 670200 445260 670206
rect 445208 670142 445260 670148
rect 445116 319524 445168 319530
rect 445116 319466 445168 319472
rect 445220 317966 445248 670142
rect 445300 668840 445352 668846
rect 445300 668782 445352 668788
rect 445208 317960 445260 317966
rect 445208 317902 445260 317908
rect 445312 317762 445340 668782
rect 445390 668536 445446 668545
rect 445390 668471 445446 668480
rect 445404 318753 445432 668471
rect 446220 447228 446272 447234
rect 446220 447170 446272 447176
rect 445484 445052 445536 445058
rect 445484 444994 445536 445000
rect 445390 318744 445446 318753
rect 445390 318679 445446 318688
rect 445496 318646 445524 444994
rect 446232 344486 446260 447170
rect 446312 444440 446364 444446
rect 446312 444382 446364 444388
rect 446220 344480 446272 344486
rect 446220 344422 446272 344428
rect 445576 337544 445628 337550
rect 445576 337486 445628 337492
rect 445484 318640 445536 318646
rect 445484 318582 445536 318588
rect 445588 318306 445616 337486
rect 446324 329662 446352 444382
rect 446312 329656 446364 329662
rect 446312 329598 446364 329604
rect 445760 320136 445812 320142
rect 445760 320078 445812 320084
rect 445576 318300 445628 318306
rect 445576 318242 445628 318248
rect 445772 318034 445800 320078
rect 446312 319660 446364 319666
rect 446312 319602 446364 319608
rect 445852 318776 445904 318782
rect 445852 318718 445904 318724
rect 445760 318028 445812 318034
rect 445760 317970 445812 317976
rect 445300 317756 445352 317762
rect 445300 317698 445352 317704
rect 445024 317076 445076 317082
rect 445024 317018 445076 317024
rect 444656 316940 444708 316946
rect 444656 316882 444708 316888
rect 445864 316538 445892 318718
rect 446324 316810 446352 319602
rect 446416 319546 446444 700606
rect 446496 700460 446548 700466
rect 446496 700402 446548 700408
rect 446508 319666 446536 700402
rect 449164 700392 449216 700398
rect 449164 700334 449216 700340
rect 446588 683188 446640 683194
rect 446588 683130 446640 683136
rect 446600 319938 446628 683130
rect 448428 679652 448480 679658
rect 448428 679594 448480 679600
rect 446772 670744 446824 670750
rect 446772 670686 446824 670692
rect 446680 670132 446732 670138
rect 446680 670074 446732 670080
rect 446588 319932 446640 319938
rect 446588 319874 446640 319880
rect 446496 319660 446548 319666
rect 446496 319602 446548 319608
rect 446416 319518 446536 319546
rect 446404 319456 446456 319462
rect 446404 319398 446456 319404
rect 446416 318782 446444 319398
rect 446508 319326 446536 319518
rect 446496 319320 446548 319326
rect 446496 319262 446548 319268
rect 446404 318776 446456 318782
rect 446404 318718 446456 318724
rect 446692 318238 446720 670074
rect 446784 319258 446812 670686
rect 446864 670268 446916 670274
rect 446864 670210 446916 670216
rect 446772 319252 446824 319258
rect 446772 319194 446824 319200
rect 446680 318232 446732 318238
rect 446680 318174 446732 318180
rect 446876 317830 446904 670210
rect 447048 668024 447100 668030
rect 447048 667966 447100 667972
rect 446956 667956 447008 667962
rect 446956 667898 447008 667904
rect 446968 318617 446996 667898
rect 447060 319394 447088 667966
rect 447876 447976 447928 447982
rect 447876 447918 447928 447924
rect 447140 447908 447192 447914
rect 447140 447850 447192 447856
rect 447784 447908 447836 447914
rect 447784 447850 447836 447856
rect 447152 447302 447180 447850
rect 447140 447296 447192 447302
rect 447140 447238 447192 447244
rect 447600 384328 447652 384334
rect 447600 384270 447652 384276
rect 447416 380248 447468 380254
rect 447416 380190 447468 380196
rect 447140 376712 447192 376718
rect 447140 376654 447192 376660
rect 447152 375873 447180 376654
rect 447138 375864 447194 375873
rect 447138 375799 447194 375808
rect 447324 375352 447376 375358
rect 447138 375320 447194 375329
rect 447324 375294 447376 375300
rect 447138 375255 447140 375264
rect 447192 375255 447194 375264
rect 447140 375226 447192 375232
rect 447232 375216 447284 375222
rect 447232 375158 447284 375164
rect 447244 374785 447272 375158
rect 447230 374776 447286 374785
rect 447230 374711 447286 374720
rect 447336 374241 447364 375294
rect 447322 374232 447378 374241
rect 447322 374167 447378 374176
rect 447232 373992 447284 373998
rect 447232 373934 447284 373940
rect 447140 373924 447192 373930
rect 447140 373866 447192 373872
rect 447152 373697 447180 373866
rect 447138 373688 447194 373697
rect 447138 373623 447194 373632
rect 447244 373153 447272 373934
rect 447230 373144 447286 373153
rect 447230 373079 447286 373088
rect 447138 372600 447194 372609
rect 447138 372535 447194 372544
rect 447324 372564 447376 372570
rect 447152 372502 447180 372535
rect 447324 372506 447376 372512
rect 447140 372496 447192 372502
rect 447140 372438 447192 372444
rect 447232 372428 447284 372434
rect 447232 372370 447284 372376
rect 447244 371521 447272 372370
rect 447336 372065 447364 372506
rect 447322 372056 447378 372065
rect 447322 371991 447378 372000
rect 447230 371512 447286 371521
rect 447230 371447 447286 371456
rect 447324 371204 447376 371210
rect 447324 371146 447376 371152
rect 447232 371136 447284 371142
rect 447232 371078 447284 371084
rect 447140 371068 447192 371074
rect 447140 371010 447192 371016
rect 447152 370977 447180 371010
rect 447138 370968 447194 370977
rect 447138 370903 447194 370912
rect 447244 370433 447272 371078
rect 447230 370424 447286 370433
rect 447230 370359 447286 370368
rect 447336 369889 447364 371146
rect 447322 369880 447378 369889
rect 447232 369844 447284 369850
rect 447322 369815 447378 369824
rect 447232 369786 447284 369792
rect 447140 369776 447192 369782
rect 447140 369718 447192 369724
rect 447152 369345 447180 369718
rect 447138 369336 447194 369345
rect 447138 369271 447194 369280
rect 447244 368801 447272 369786
rect 447230 368792 447286 368801
rect 447230 368727 447286 368736
rect 447140 368484 447192 368490
rect 447140 368426 447192 368432
rect 447152 368257 447180 368426
rect 447232 368416 447284 368422
rect 447232 368358 447284 368364
rect 447138 368248 447194 368257
rect 447138 368183 447194 368192
rect 447244 367713 447272 368358
rect 447324 368348 447376 368354
rect 447324 368290 447376 368296
rect 447230 367704 447286 367713
rect 447230 367639 447286 367648
rect 447336 367169 447364 368290
rect 447322 367160 447378 367169
rect 447322 367095 447378 367104
rect 447140 367056 447192 367062
rect 447140 366998 447192 367004
rect 447152 366625 447180 366998
rect 447232 366988 447284 366994
rect 447232 366930 447284 366936
rect 447138 366616 447194 366625
rect 447138 366551 447194 366560
rect 447244 366081 447272 366930
rect 447230 366072 447286 366081
rect 447230 366007 447286 366016
rect 447324 365696 447376 365702
rect 447324 365638 447376 365644
rect 447232 365628 447284 365634
rect 447232 365570 447284 365576
rect 447140 365560 447192 365566
rect 447138 365528 447140 365537
rect 447192 365528 447194 365537
rect 447138 365463 447194 365472
rect 447244 364993 447272 365570
rect 447230 364984 447286 364993
rect 447230 364919 447286 364928
rect 447336 364449 447364 365638
rect 447322 364440 447378 364449
rect 447322 364375 447378 364384
rect 447232 364336 447284 364342
rect 447232 364278 447284 364284
rect 447140 364268 447192 364274
rect 447140 364210 447192 364216
rect 447152 363905 447180 364210
rect 447138 363896 447194 363905
rect 447138 363831 447194 363840
rect 447244 363361 447272 364278
rect 447230 363352 447286 363361
rect 447230 363287 447286 363296
rect 447140 362908 447192 362914
rect 447140 362850 447192 362856
rect 447152 362817 447180 362850
rect 447232 362840 447284 362846
rect 447138 362808 447194 362817
rect 447232 362782 447284 362788
rect 447138 362743 447194 362752
rect 447244 362273 447272 362782
rect 447324 362772 447376 362778
rect 447324 362714 447376 362720
rect 447230 362264 447286 362273
rect 447230 362199 447286 362208
rect 447336 361729 447364 362714
rect 447322 361720 447378 361729
rect 447322 361655 447378 361664
rect 447140 361548 447192 361554
rect 447140 361490 447192 361496
rect 447152 361185 447180 361490
rect 447232 361480 447284 361486
rect 447232 361422 447284 361428
rect 447138 361176 447194 361185
rect 447138 361111 447194 361120
rect 447244 360641 447272 361422
rect 447230 360632 447286 360641
rect 447230 360567 447286 360576
rect 447230 360088 447286 360097
rect 447230 360023 447286 360032
rect 447138 359544 447194 359553
rect 447138 359479 447194 359488
rect 447152 358902 447180 359479
rect 447140 358896 447192 358902
rect 447140 358838 447192 358844
rect 447244 358834 447272 360023
rect 447322 359000 447378 359009
rect 447322 358935 447324 358944
rect 447376 358935 447378 358944
rect 447324 358906 447376 358912
rect 447232 358828 447284 358834
rect 447232 358770 447284 358776
rect 447230 358456 447286 358465
rect 447230 358391 447286 358400
rect 447138 357912 447194 357921
rect 447138 357847 447194 357856
rect 447152 357474 447180 357847
rect 447244 357542 447272 358391
rect 447232 357536 447284 357542
rect 447232 357478 447284 357484
rect 447140 357468 447192 357474
rect 447140 357410 447192 357416
rect 447230 357368 447286 357377
rect 447230 357303 447286 357312
rect 447138 356280 447194 356289
rect 447138 356215 447194 356224
rect 447152 356182 447180 356215
rect 447140 356176 447192 356182
rect 447140 356118 447192 356124
rect 447244 356114 447272 357303
rect 447322 356824 447378 356833
rect 447322 356759 447378 356768
rect 447336 356250 447364 356759
rect 447324 356244 447376 356250
rect 447324 356186 447376 356192
rect 447232 356108 447284 356114
rect 447232 356050 447284 356056
rect 447428 353569 447456 380190
rect 447414 353560 447470 353569
rect 447414 353495 447470 353504
rect 447324 350532 447376 350538
rect 447324 350474 447376 350480
rect 447140 350464 447192 350470
rect 447140 350406 447192 350412
rect 447152 350305 447180 350406
rect 447232 350396 447284 350402
rect 447232 350338 447284 350344
rect 447138 350296 447194 350305
rect 447138 350231 447194 350240
rect 447244 349761 447272 350338
rect 447230 349752 447286 349761
rect 447230 349687 447286 349696
rect 447336 349217 447364 350474
rect 447322 349208 447378 349217
rect 447322 349143 447378 349152
rect 447140 349104 447192 349110
rect 447140 349046 447192 349052
rect 447152 348129 447180 349046
rect 447232 349036 447284 349042
rect 447232 348978 447284 348984
rect 447244 348673 447272 348978
rect 447230 348664 447286 348673
rect 447230 348599 447286 348608
rect 447138 348120 447194 348129
rect 447138 348055 447194 348064
rect 447232 347744 447284 347750
rect 447232 347686 447284 347692
rect 447140 347608 447192 347614
rect 447138 347576 447140 347585
rect 447192 347576 447194 347585
rect 447138 347511 447194 347520
rect 447244 347041 447272 347686
rect 447324 347676 447376 347682
rect 447324 347618 447376 347624
rect 447230 347032 447286 347041
rect 447230 346967 447286 346976
rect 447336 346497 447364 347618
rect 447322 346488 447378 346497
rect 447322 346423 447378 346432
rect 447138 345400 447194 345409
rect 447138 345335 447194 345344
rect 447152 345098 447180 345335
rect 447140 345092 447192 345098
rect 447140 345034 447192 345040
rect 447140 343596 447192 343602
rect 447140 343538 447192 343544
rect 447152 342689 447180 343538
rect 447138 342680 447194 342689
rect 447138 342615 447194 342624
rect 447612 342145 447640 384270
rect 447598 342136 447654 342145
rect 447598 342071 447654 342080
rect 447140 338564 447192 338570
rect 447140 338506 447192 338512
rect 447152 338337 447180 338506
rect 447138 338328 447194 338337
rect 447138 338263 447194 338272
rect 447690 338056 447746 338065
rect 447690 337991 447746 338000
rect 447230 337784 447286 337793
rect 447230 337719 447286 337728
rect 447138 337240 447194 337249
rect 447138 337175 447194 337184
rect 447152 336870 447180 337175
rect 447140 336864 447192 336870
rect 447140 336806 447192 336812
rect 447244 336802 447272 337719
rect 447704 336841 447732 337991
rect 447690 336832 447746 336841
rect 447232 336796 447284 336802
rect 447690 336767 447746 336776
rect 447232 336738 447284 336744
rect 447230 336696 447286 336705
rect 447230 336631 447286 336640
rect 447138 336152 447194 336161
rect 447138 336087 447194 336096
rect 447152 335782 447180 336087
rect 447244 335850 447272 336631
rect 447232 335844 447284 335850
rect 447232 335786 447284 335792
rect 447140 335776 447192 335782
rect 447140 335718 447192 335724
rect 447322 335608 447378 335617
rect 447322 335543 447378 335552
rect 447230 335064 447286 335073
rect 447230 334999 447286 335008
rect 447138 334520 447194 334529
rect 447138 334455 447194 334464
rect 447152 334014 447180 334455
rect 447244 334082 447272 334999
rect 447336 334626 447364 335543
rect 447324 334620 447376 334626
rect 447324 334562 447376 334568
rect 447232 334076 447284 334082
rect 447232 334018 447284 334024
rect 447140 334008 447192 334014
rect 447140 333950 447192 333956
rect 447230 333976 447286 333985
rect 447230 333911 447286 333920
rect 447138 333432 447194 333441
rect 447138 333367 447194 333376
rect 447152 332722 447180 333367
rect 447140 332716 447192 332722
rect 447140 332658 447192 332664
rect 447244 332654 447272 333911
rect 447322 332888 447378 332897
rect 447322 332823 447378 332832
rect 447232 332648 447284 332654
rect 447232 332590 447284 332596
rect 447138 331800 447194 331809
rect 447138 331735 447194 331744
rect 447152 331294 447180 331735
rect 447232 331356 447284 331362
rect 447232 331298 447284 331304
rect 447140 331288 447192 331294
rect 447244 331265 447272 331298
rect 447140 331230 447192 331236
rect 447230 331256 447286 331265
rect 447230 331191 447286 331200
rect 447336 330546 447364 332823
rect 447414 332344 447470 332353
rect 447414 332279 447470 332288
rect 447428 331430 447456 332279
rect 447416 331424 447468 331430
rect 447416 331366 447468 331372
rect 447324 330540 447376 330546
rect 447324 330482 447376 330488
rect 447506 330168 447562 330177
rect 447506 330103 447562 330112
rect 447048 319388 447100 319394
rect 447048 319330 447100 319336
rect 446954 318608 447010 318617
rect 446954 318543 447010 318552
rect 446864 317824 446916 317830
rect 446864 317766 446916 317772
rect 446404 317416 446456 317422
rect 446404 317358 446456 317364
rect 446312 316804 446364 316810
rect 446312 316746 446364 316752
rect 445852 316532 445904 316538
rect 445852 316474 445904 316480
rect 444472 316464 444524 316470
rect 444472 316406 444524 316412
rect 443920 305924 443972 305930
rect 443920 305866 443972 305872
rect 444380 294296 444432 294302
rect 444380 294238 444432 294244
rect 444392 293282 444420 294238
rect 444380 293276 444432 293282
rect 444380 293218 444432 293224
rect 445760 276072 445812 276078
rect 445760 276014 445812 276020
rect 443920 271108 443972 271114
rect 443920 271050 443972 271056
rect 443828 264240 443880 264246
rect 443828 264182 443880 264188
rect 443932 262750 443960 271050
rect 445772 268394 445800 276014
rect 445760 268388 445812 268394
rect 445760 268330 445812 268336
rect 443920 262744 443972 262750
rect 443920 262686 443972 262692
rect 445760 260432 445812 260438
rect 445760 260374 445812 260380
rect 445772 258074 445800 260374
rect 445680 258046 445800 258074
rect 445680 254590 445708 258046
rect 446128 255264 446180 255270
rect 446128 255206 446180 255212
rect 445668 254584 445720 254590
rect 445668 254526 445720 254532
rect 446140 250442 446168 255206
rect 443828 250436 443880 250442
rect 443828 250378 443880 250384
rect 446128 250436 446180 250442
rect 446128 250378 446180 250384
rect 443840 230518 443868 250378
rect 445024 243228 445076 243234
rect 445024 243170 445076 243176
rect 443828 230512 443880 230518
rect 443828 230454 443880 230460
rect 444196 223304 444248 223310
rect 444196 223246 444248 223252
rect 444208 219502 444236 223246
rect 444196 219496 444248 219502
rect 444196 219438 444248 219444
rect 445036 218142 445064 243170
rect 445024 218136 445076 218142
rect 445024 218078 445076 218084
rect 443828 211336 443880 211342
rect 443828 211278 443880 211284
rect 443840 189106 443868 211278
rect 443828 189100 443880 189106
rect 443828 189042 443880 189048
rect 443736 186584 443788 186590
rect 443736 186526 443788 186532
rect 446416 167210 446444 317358
rect 446496 302252 446548 302258
rect 446496 302194 446548 302200
rect 446508 294302 446536 302194
rect 446496 294296 446548 294302
rect 446496 294238 446548 294244
rect 446494 276720 446550 276729
rect 446494 276655 446550 276664
rect 446508 271114 446536 276655
rect 446496 271108 446548 271114
rect 446496 271050 446548 271056
rect 446496 245676 446548 245682
rect 446496 245618 446548 245624
rect 446508 243234 446536 245618
rect 446496 243228 446548 243234
rect 446496 243170 446548 243176
rect 447140 186312 447192 186318
rect 447140 186254 447192 186260
rect 447152 185638 447180 186254
rect 447140 185632 447192 185638
rect 447140 185574 447192 185580
rect 447520 175234 447548 330103
rect 447704 327078 447732 336767
rect 447796 328506 447824 447850
rect 447888 447370 447916 447918
rect 447876 447364 447928 447370
rect 447876 447306 447928 447312
rect 448244 447364 448296 447370
rect 448244 447306 448296 447312
rect 448060 383036 448112 383042
rect 448060 382978 448112 382984
rect 447968 381608 448020 381614
rect 447968 381550 448020 381556
rect 447876 380180 447928 380186
rect 447876 380122 447928 380128
rect 447888 353025 447916 380122
rect 447874 353016 447930 353025
rect 447874 352951 447930 352960
rect 447876 344480 447928 344486
rect 447876 344422 447928 344428
rect 447888 340513 447916 344422
rect 447980 344321 448008 381550
rect 447966 344312 448022 344321
rect 447966 344247 448022 344256
rect 448072 343777 448100 382978
rect 448152 381540 448204 381546
rect 448152 381482 448204 381488
rect 448058 343768 448114 343777
rect 448058 343703 448114 343712
rect 448164 341601 448192 381482
rect 448150 341592 448206 341601
rect 448150 341527 448206 341536
rect 448058 341048 448114 341057
rect 448058 340983 448114 340992
rect 447874 340504 447930 340513
rect 447874 340439 447930 340448
rect 447876 339108 447928 339114
rect 447876 339050 447928 339056
rect 447888 336734 447916 339050
rect 447876 336728 447928 336734
rect 447876 336670 447928 336676
rect 447784 328500 447836 328506
rect 447784 328442 447836 328448
rect 447692 327072 447744 327078
rect 447692 327014 447744 327020
rect 447784 263492 447836 263498
rect 447784 263434 447836 263440
rect 447796 245682 447824 263434
rect 447888 249082 447916 336670
rect 447966 329760 448022 329769
rect 447966 329695 448022 329704
rect 447980 329089 448008 329695
rect 447966 329080 448022 329089
rect 447966 329015 448022 329024
rect 447980 317422 448008 329015
rect 447968 317416 448020 317422
rect 447968 317358 448020 317364
rect 448072 300082 448100 340983
rect 448150 330712 448206 330721
rect 448150 330647 448206 330656
rect 448060 300076 448112 300082
rect 448060 300018 448112 300024
rect 447876 249076 447928 249082
rect 447876 249018 447928 249024
rect 447784 245676 447836 245682
rect 447784 245618 447836 245624
rect 447784 231872 447836 231878
rect 447784 231814 447836 231820
rect 447796 211342 447824 231814
rect 447784 211336 447836 211342
rect 447784 211278 447836 211284
rect 448164 185638 448192 330647
rect 448256 329769 448284 447306
rect 448336 379840 448388 379846
rect 448336 379782 448388 379788
rect 448348 355201 448376 379782
rect 448334 355192 448390 355201
rect 448334 355127 448390 355136
rect 448334 345944 448390 345953
rect 448334 345879 448390 345888
rect 448242 329760 448298 329769
rect 448242 329695 448298 329704
rect 448244 329656 448296 329662
rect 448242 329624 448244 329633
rect 448296 329624 448298 329633
rect 448242 329559 448298 329568
rect 448242 328536 448298 328545
rect 448242 328471 448244 328480
rect 448296 328471 448298 328480
rect 448244 328442 448296 328448
rect 448152 185632 448204 185638
rect 448152 185574 448204 185580
rect 447140 175228 447192 175234
rect 447140 175170 447192 175176
rect 447508 175228 447560 175234
rect 447508 175170 447560 175176
rect 447152 174554 447180 175170
rect 447140 174548 447192 174554
rect 447140 174490 447192 174496
rect 445668 167204 445720 167210
rect 445668 167146 445720 167152
rect 446404 167204 446456 167210
rect 446404 167146 446456 167152
rect 442724 165640 442776 165646
rect 442724 165582 442776 165588
rect 442908 165640 442960 165646
rect 442908 165582 442960 165588
rect 437998 165170 438072 165186
rect 437986 165164 438072 165170
rect 438038 165158 438072 165164
rect 437986 165106 438038 165112
rect 437998 164900 438026 165106
rect 442736 165102 442764 165582
rect 441666 165096 441718 165102
rect 441666 165038 441718 165044
rect 442724 165096 442776 165102
rect 442724 165038 442776 165044
rect 441678 164900 441706 165038
rect 445208 164960 445260 164966
rect 445680 164914 445708 167146
rect 448348 164966 448376 345879
rect 448440 315722 448468 679594
rect 449072 461644 449124 461650
rect 449072 461586 449124 461592
rect 449084 354113 449112 461586
rect 449070 354104 449126 354113
rect 449070 354039 449126 354048
rect 448518 327992 448574 328001
rect 448518 327927 448574 327936
rect 448532 327146 448560 327927
rect 448520 327140 448572 327146
rect 448520 327082 448572 327088
rect 449176 320006 449204 700334
rect 462332 679658 462360 703520
rect 478524 700738 478552 703520
rect 478512 700732 478564 700738
rect 478512 700674 478564 700680
rect 494808 700534 494836 703520
rect 494796 700528 494848 700534
rect 494796 700470 494848 700476
rect 527192 700330 527220 703520
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 543476 699825 543504 703520
rect 543740 700324 543792 700330
rect 543740 700266 543792 700272
rect 543462 699816 543518 699825
rect 543462 699751 543518 699760
rect 462320 679652 462372 679658
rect 462320 679594 462372 679600
rect 458730 678600 458786 678609
rect 458730 678535 458786 678544
rect 457902 632904 457958 632913
rect 457902 632839 457958 632848
rect 457810 630048 457866 630057
rect 457810 629983 457866 629992
rect 457718 627192 457774 627201
rect 457718 627127 457774 627136
rect 457626 621480 457682 621489
rect 457626 621415 457682 621424
rect 457534 615768 457590 615777
rect 457534 615703 457590 615712
rect 457548 615494 457576 615703
rect 457272 615466 457576 615494
rect 457272 600234 457300 615466
rect 457442 612912 457498 612921
rect 457442 612847 457498 612856
rect 457350 610056 457406 610065
rect 457350 609991 457406 610000
rect 457260 600228 457312 600234
rect 457260 600170 457312 600176
rect 457364 598466 457392 609991
rect 457456 599690 457484 612847
rect 457536 610700 457588 610706
rect 457536 610642 457588 610648
rect 457548 599758 457576 610642
rect 457536 599752 457588 599758
rect 457536 599694 457588 599700
rect 457444 599684 457496 599690
rect 457444 599626 457496 599632
rect 457352 598460 457404 598466
rect 457352 598402 457404 598408
rect 457640 596902 457668 621415
rect 457628 596896 457680 596902
rect 457628 596838 457680 596844
rect 457732 595542 457760 627127
rect 457824 598398 457852 629983
rect 457916 610706 457944 632839
rect 458086 624336 458142 624345
rect 458086 624271 458142 624280
rect 457994 618624 458050 618633
rect 457994 618559 458050 618568
rect 457904 610700 457956 610706
rect 457904 610642 457956 610648
rect 457902 607200 457958 607209
rect 457902 607135 457958 607144
rect 457916 600302 457944 607135
rect 457904 600296 457956 600302
rect 457904 600238 457956 600244
rect 457812 598392 457864 598398
rect 457812 598334 457864 598340
rect 457720 595536 457772 595542
rect 457720 595478 457772 595484
rect 458008 518226 458036 618559
rect 458100 522306 458128 624271
rect 458744 599593 458772 678535
rect 459282 670032 459338 670041
rect 459282 669967 459338 669976
rect 459098 664320 459154 664329
rect 459098 664255 459154 664264
rect 459006 652896 459062 652905
rect 459006 652831 459062 652840
rect 458914 647184 458970 647193
rect 458914 647119 458970 647128
rect 458822 641472 458878 641481
rect 458822 641407 458878 641416
rect 458730 599584 458786 599593
rect 458730 599519 458786 599528
rect 458836 596873 458864 641407
rect 458822 596864 458878 596873
rect 458822 596799 458878 596808
rect 458928 592686 458956 647119
rect 459020 596834 459048 652831
rect 459112 598330 459140 664255
rect 459190 658608 459246 658617
rect 459190 658543 459246 658552
rect 459100 598324 459152 598330
rect 459100 598266 459152 598272
rect 459008 596828 459060 596834
rect 459008 596770 459060 596776
rect 458916 592680 458968 592686
rect 458916 592622 458968 592628
rect 459204 589966 459232 658543
rect 459296 591326 459324 669967
rect 460570 666632 460626 666641
rect 460570 666567 460626 666576
rect 460386 661056 460442 661065
rect 460386 660991 460442 661000
rect 460400 654134 460428 660991
rect 460478 655888 460534 655897
rect 460478 655823 460480 655832
rect 460532 655823 460534 655832
rect 460480 655794 460532 655800
rect 460400 654106 460520 654134
rect 460386 650176 460442 650185
rect 460386 650111 460442 650120
rect 460294 643784 460350 643793
rect 460294 643719 460296 643728
rect 460348 643719 460350 643728
rect 460296 643690 460348 643696
rect 459466 638616 459522 638625
rect 459466 638551 459522 638560
rect 459374 604344 459430 604353
rect 459374 604279 459430 604288
rect 459388 594017 459416 604279
rect 459374 594008 459430 594017
rect 459374 593943 459430 593952
rect 459284 591320 459336 591326
rect 459284 591262 459336 591268
rect 459192 589960 459244 589966
rect 459192 589902 459244 589908
rect 458088 522300 458140 522306
rect 458088 522242 458140 522248
rect 457996 518220 458048 518226
rect 457996 518162 458048 518168
rect 459480 518129 459508 638551
rect 460400 605834 460428 650111
rect 460308 605806 460428 605834
rect 460308 598262 460336 605806
rect 460492 602954 460520 654106
rect 460480 602948 460532 602954
rect 460480 602890 460532 602896
rect 460584 602834 460612 666567
rect 460664 655852 460716 655858
rect 460664 655794 460716 655800
rect 460400 602806 460612 602834
rect 460400 599622 460428 602806
rect 460480 602676 460532 602682
rect 460480 602618 460532 602624
rect 460388 599616 460440 599622
rect 460388 599558 460440 599564
rect 460296 598256 460348 598262
rect 460296 598198 460348 598204
rect 460492 595474 460520 602618
rect 460570 600944 460626 600953
rect 460570 600879 460626 600888
rect 460584 600710 460612 600879
rect 460572 600704 460624 600710
rect 460572 600646 460624 600652
rect 460480 595468 460532 595474
rect 460480 595410 460532 595416
rect 460676 537538 460704 655794
rect 460756 643748 460808 643754
rect 460756 643690 460808 643696
rect 460664 537532 460716 537538
rect 460664 537474 460716 537480
rect 460768 519586 460796 643690
rect 461584 600704 461636 600710
rect 461584 600646 461636 600652
rect 460756 519580 460808 519586
rect 460756 519522 460808 519528
rect 459466 518120 459522 518129
rect 459466 518055 459522 518064
rect 450360 517608 450412 517614
rect 450360 517550 450412 517556
rect 450176 516860 450228 516866
rect 450176 516802 450228 516808
rect 449990 512408 450046 512417
rect 449990 512343 450046 512352
rect 449624 460216 449676 460222
rect 449624 460158 449676 460164
rect 449532 457496 449584 457502
rect 449532 457438 449584 457444
rect 449440 456204 449492 456210
rect 449440 456146 449492 456152
rect 449348 456136 449400 456142
rect 449348 456078 449400 456084
rect 449256 456068 449308 456074
rect 449256 456010 449308 456016
rect 449268 355745 449296 456010
rect 449254 355736 449310 355745
rect 449254 355671 449310 355680
rect 449360 352481 449388 456078
rect 449346 352472 449402 352481
rect 449346 352407 449402 352416
rect 449452 350849 449480 456146
rect 449544 351937 449572 457438
rect 449636 354657 449664 460158
rect 449716 457564 449768 457570
rect 449716 457506 449768 457512
rect 449622 354648 449678 354657
rect 449622 354583 449678 354592
rect 449530 351928 449586 351937
rect 449530 351863 449586 351872
rect 449728 351393 449756 457506
rect 449900 447840 449952 447846
rect 449900 447782 449952 447788
rect 449912 447166 449940 447782
rect 449900 447160 449952 447166
rect 449900 447102 449952 447108
rect 449808 379568 449860 379574
rect 449808 379510 449860 379516
rect 449714 351384 449770 351393
rect 449714 351319 449770 351328
rect 449438 350840 449494 350849
rect 449438 350775 449494 350784
rect 449714 344856 449770 344865
rect 449714 344791 449770 344800
rect 449348 340196 449400 340202
rect 449348 340138 449400 340144
rect 449256 337408 449308 337414
rect 449256 337350 449308 337356
rect 449164 320000 449216 320006
rect 449164 319942 449216 319948
rect 448428 315716 448480 315722
rect 448428 315658 448480 315664
rect 449268 315654 449296 337350
rect 449360 318510 449388 340138
rect 449624 339312 449676 339318
rect 449624 339254 449676 339260
rect 449636 338230 449664 339254
rect 449624 338224 449676 338230
rect 449624 338166 449676 338172
rect 449636 324193 449664 338166
rect 449622 324184 449678 324193
rect 449622 324119 449678 324128
rect 449348 318504 449400 318510
rect 449348 318446 449400 318452
rect 449256 315648 449308 315654
rect 449256 315590 449308 315596
rect 448520 315376 448572 315382
rect 448520 315318 448572 315324
rect 448532 310146 448560 315318
rect 448520 310140 448572 310146
rect 448520 310082 448572 310088
rect 448428 304428 448480 304434
rect 448428 304370 448480 304376
rect 448440 302258 448468 304370
rect 448428 302252 448480 302258
rect 448428 302194 448480 302200
rect 449164 285728 449216 285734
rect 449164 285670 449216 285676
rect 449176 276078 449204 285670
rect 449164 276072 449216 276078
rect 449164 276014 449216 276020
rect 449256 271448 449308 271454
rect 449256 271390 449308 271396
rect 448520 264920 448572 264926
rect 448520 264862 448572 264868
rect 448532 262290 448560 264862
rect 448440 262262 448560 262290
rect 448440 260438 448468 262262
rect 448428 260432 448480 260438
rect 448428 260374 448480 260380
rect 449164 258120 449216 258126
rect 449164 258062 449216 258068
rect 449176 240922 449204 258062
rect 449268 255338 449296 271390
rect 449348 268660 449400 268666
rect 449348 268602 449400 268608
rect 449360 257378 449388 268602
rect 449728 263566 449756 344791
rect 449820 343233 449848 379510
rect 449806 343224 449862 343233
rect 449806 343159 449862 343168
rect 449806 339960 449862 339969
rect 449806 339895 449862 339904
rect 449716 263560 449768 263566
rect 449716 263502 449768 263508
rect 449348 257372 449400 257378
rect 449348 257314 449400 257320
rect 449256 255332 449308 255338
rect 449256 255274 449308 255280
rect 449164 240916 449216 240922
rect 449164 240858 449216 240864
rect 449164 232756 449216 232762
rect 449164 232698 449216 232704
rect 449176 223310 449204 232698
rect 449164 223304 449216 223310
rect 449164 223246 449216 223252
rect 449820 169114 449848 339895
rect 450004 339454 450032 512343
rect 450082 510232 450138 510241
rect 450082 510167 450138 510176
rect 449992 339448 450044 339454
rect 449992 339390 450044 339396
rect 450096 339386 450124 510167
rect 450188 505481 450216 516802
rect 450372 510241 450400 517550
rect 450544 517540 450596 517546
rect 450544 517482 450596 517488
rect 450450 517032 450506 517041
rect 450450 516967 450506 516976
rect 450464 512417 450492 516967
rect 450556 514729 450584 517482
rect 450636 516792 450688 516798
rect 450636 516734 450688 516740
rect 450542 514720 450598 514729
rect 450542 514655 450598 514664
rect 450450 512408 450506 512417
rect 450450 512343 450506 512352
rect 450358 510232 450414 510241
rect 450358 510167 450414 510176
rect 450266 507648 450322 507657
rect 450648 507634 450676 516734
rect 450322 507606 450676 507634
rect 450266 507583 450322 507592
rect 450174 505472 450230 505481
rect 450174 505407 450230 505416
rect 450084 339380 450136 339386
rect 450084 339322 450136 339328
rect 450082 339144 450138 339153
rect 450082 339079 450084 339088
rect 450136 339079 450138 339088
rect 450084 339050 450136 339056
rect 450084 338972 450136 338978
rect 450084 338914 450136 338920
rect 450096 338298 450124 338914
rect 450188 338366 450216 505407
rect 450176 338360 450228 338366
rect 450176 338302 450228 338308
rect 450084 338292 450136 338298
rect 450084 338234 450136 338240
rect 449990 327176 450046 327185
rect 449990 327111 450046 327120
rect 449898 326632 449954 326641
rect 449898 326567 449954 326576
rect 449808 169108 449860 169114
rect 449808 169050 449860 169056
rect 449348 168088 449400 168094
rect 449348 168030 449400 168036
rect 445260 164908 445708 164914
rect 445208 164902 445708 164908
rect 448336 164960 448388 164966
rect 449360 164914 449388 168030
rect 449912 167142 449940 326567
rect 449900 167136 449952 167142
rect 449900 167078 449952 167084
rect 450004 167074 450032 327111
rect 450096 325009 450124 338234
rect 450188 325553 450216 338302
rect 450280 338065 450308 507583
rect 450542 503296 450598 503305
rect 450542 503231 450598 503240
rect 450556 500954 450584 503231
rect 450544 500948 450596 500954
rect 450544 500890 450596 500896
rect 450360 339448 450412 339454
rect 450360 339390 450412 339396
rect 450372 338502 450400 339390
rect 450452 339380 450504 339386
rect 450452 339322 450504 339328
rect 450360 338496 450412 338502
rect 450360 338438 450412 338444
rect 450266 338056 450322 338065
rect 450266 337991 450322 338000
rect 450268 327072 450320 327078
rect 450268 327014 450320 327020
rect 450280 326097 450308 327014
rect 450372 326641 450400 338438
rect 450464 338434 450492 339322
rect 450556 338978 450584 500890
rect 450754 500126 451228 500154
rect 452226 500126 452608 500154
rect 451200 496890 451228 500126
rect 451200 496862 451320 496890
rect 450636 447840 450688 447846
rect 450636 447782 450688 447788
rect 450648 382974 450676 447782
rect 451292 402974 451320 496862
rect 451292 402946 451872 402974
rect 450636 382968 450688 382974
rect 450636 382910 450688 382916
rect 450648 382294 450676 382910
rect 450636 382288 450688 382294
rect 450636 382230 450688 382236
rect 450636 381676 450688 381682
rect 450636 381618 450688 381624
rect 450648 339318 450676 381618
rect 451844 379930 451872 402946
rect 452580 382294 452608 500126
rect 453304 497480 453356 497486
rect 453304 497422 453356 497428
rect 452568 382288 452620 382294
rect 452568 382230 452620 382236
rect 451844 379902 452226 379930
rect 453316 379846 453344 497422
rect 453684 496890 453712 500140
rect 455170 500126 455368 500154
rect 454684 497548 454736 497554
rect 454684 497490 454736 497496
rect 453684 496862 454080 496890
rect 454052 402974 454080 496862
rect 454052 402946 454448 402974
rect 453488 382288 453540 382294
rect 453488 382230 453540 382236
rect 453500 379916 453528 382230
rect 454420 379930 454448 402946
rect 454696 380254 454724 497490
rect 454776 466472 454828 466478
rect 454776 466414 454828 466420
rect 454788 384334 454816 466414
rect 454776 384328 454828 384334
rect 454776 384270 454828 384276
rect 455340 382294 455368 500126
rect 456628 499574 456656 500140
rect 456628 499546 456748 499574
rect 456064 458312 456116 458318
rect 456064 458254 456116 458260
rect 456076 383042 456104 458254
rect 456720 383654 456748 499546
rect 457444 458244 457496 458250
rect 457444 458186 457496 458192
rect 456720 383626 457024 383654
rect 456064 383036 456116 383042
rect 456064 382978 456116 382984
rect 455328 382288 455380 382294
rect 455328 382230 455380 382236
rect 456064 382288 456116 382294
rect 456064 382230 456116 382236
rect 454684 380248 454736 380254
rect 454684 380190 454736 380196
rect 454420 379902 454802 379930
rect 456076 379916 456104 382230
rect 456996 379930 457024 383626
rect 457456 381682 457484 458186
rect 458100 431954 458128 500140
rect 459586 500126 460244 500154
rect 461058 500126 461440 500154
rect 458824 465112 458876 465118
rect 458824 465054 458876 465060
rect 458836 447982 458864 465054
rect 458824 447976 458876 447982
rect 458824 447918 458876 447924
rect 458100 431926 458220 431954
rect 458192 402974 458220 431926
rect 458192 402946 458312 402974
rect 457444 381676 457496 381682
rect 457444 381618 457496 381624
rect 458284 379930 458312 402946
rect 460216 379930 460244 500126
rect 461412 494766 461440 500126
rect 461400 494760 461452 494766
rect 461400 494702 461452 494708
rect 461596 406434 461624 600646
rect 462964 600296 463016 600302
rect 462964 600238 463016 600244
rect 461676 520328 461728 520334
rect 461676 520270 461728 520276
rect 461584 406428 461636 406434
rect 461584 406370 461636 406376
rect 461688 381614 461716 520270
rect 461768 494760 461820 494766
rect 461768 494702 461820 494708
rect 461676 381608 461728 381614
rect 461676 381550 461728 381556
rect 461780 379930 461808 494702
rect 462976 383450 463004 600238
rect 463056 600228 463108 600234
rect 463056 600170 463108 600176
rect 462964 383444 463016 383450
rect 462964 383386 463016 383392
rect 463068 383178 463096 600170
rect 464370 600086 464476 600114
rect 464344 599752 464396 599758
rect 464344 599694 464396 599700
rect 463608 427100 463660 427106
rect 463608 427042 463660 427048
rect 463620 383654 463648 427042
rect 463160 383626 463648 383654
rect 463056 383172 463108 383178
rect 463056 383114 463108 383120
rect 463160 380610 463188 383626
rect 464356 383042 464384 599694
rect 464448 501129 464476 600086
rect 472636 600086 472834 600114
rect 480456 600086 481298 600114
rect 489196 600086 489762 600114
rect 498226 600086 498332 600114
rect 467104 599684 467156 599690
rect 467104 599626 467156 599632
rect 464434 501120 464490 501129
rect 464434 501055 464490 501064
rect 464436 497616 464488 497622
rect 464436 497558 464488 497564
rect 464344 383036 464396 383042
rect 464344 382978 464396 382984
rect 462976 380582 463188 380610
rect 462976 379930 463004 380582
rect 464448 380458 464476 497558
rect 464528 465180 464580 465186
rect 464528 465122 464580 465128
rect 464540 447914 464568 465122
rect 464528 447908 464580 447914
rect 464528 447850 464580 447856
rect 464988 430024 465040 430030
rect 464988 429966 465040 429972
rect 465000 383654 465028 429966
rect 466276 429956 466328 429962
rect 466276 429898 466328 429904
rect 466288 383654 466316 429898
rect 466368 429888 466420 429894
rect 466368 429830 466420 429836
rect 464540 383626 465028 383654
rect 465552 383626 466316 383654
rect 464436 380452 464488 380458
rect 464436 380394 464488 380400
rect 464540 380338 464568 383626
rect 464264 380310 464568 380338
rect 464264 379930 464292 380310
rect 465552 379930 465580 383626
rect 456996 379902 457378 379930
rect 458284 379902 458666 379930
rect 459954 379902 460244 379930
rect 461242 379902 461808 379930
rect 462530 379902 463004 379930
rect 463818 379902 464292 379930
rect 465106 379902 465580 379930
rect 466380 379916 466408 429830
rect 467116 383586 467144 599626
rect 468484 598460 468536 598466
rect 468484 598402 468536 598408
rect 467196 596896 467248 596902
rect 467196 596838 467248 596844
rect 467104 383580 467156 383586
rect 467104 383522 467156 383528
rect 467208 383246 467236 596838
rect 467288 522300 467340 522306
rect 467288 522242 467340 522248
rect 467196 383240 467248 383246
rect 467196 383182 467248 383188
rect 467300 383110 467328 522242
rect 467656 384328 467708 384334
rect 467656 384270 467708 384276
rect 467288 383104 467340 383110
rect 467288 383046 467340 383052
rect 467668 379916 467696 384270
rect 468496 383654 468524 598402
rect 471244 598392 471296 598398
rect 471244 598334 471296 598340
rect 468576 595536 468628 595542
rect 468576 595478 468628 595484
rect 468484 383648 468536 383654
rect 468484 383590 468536 383596
rect 468588 383314 468616 595478
rect 469864 518220 469916 518226
rect 469864 518162 469916 518168
rect 468668 458380 468720 458386
rect 468668 458322 468720 458328
rect 468680 447846 468708 458322
rect 468668 447840 468720 447846
rect 468668 447782 468720 447788
rect 468944 385688 468996 385694
rect 468944 385630 468996 385636
rect 468576 383308 468628 383314
rect 468576 383250 468628 383256
rect 468956 379916 468984 385630
rect 469876 383518 469904 518162
rect 470232 384396 470284 384402
rect 470232 384338 470284 384344
rect 469864 383512 469916 383518
rect 469864 383454 469916 383460
rect 470244 379916 470272 384338
rect 471256 383382 471284 598334
rect 472636 500954 472664 600086
rect 480456 516905 480484 600086
rect 482928 520940 482980 520946
rect 482928 520882 482980 520888
rect 482742 517576 482798 517585
rect 482940 517562 482968 520882
rect 488632 520328 488684 520334
rect 488632 520270 488684 520276
rect 488644 517970 488672 520270
rect 488644 517942 488980 517970
rect 482798 517534 483000 517562
rect 482742 517511 482798 517520
rect 489196 517478 489224 600086
rect 495440 598256 495492 598262
rect 495440 598198 495492 598204
rect 496084 598256 496136 598262
rect 496084 598198 496136 598204
rect 494060 592680 494112 592686
rect 494060 592622 494112 592628
rect 493048 519580 493100 519586
rect 493048 519522 493100 519528
rect 491852 517608 491904 517614
rect 491852 517550 491904 517556
rect 489184 517472 489236 517478
rect 489184 517414 489236 517420
rect 480442 516896 480498 516905
rect 480442 516831 480444 516840
rect 480496 516831 480498 516840
rect 480444 516802 480496 516808
rect 491864 516633 491892 517550
rect 492126 516896 492182 516905
rect 492126 516831 492182 516840
rect 491850 516624 491906 516633
rect 491850 516559 491906 516568
rect 492140 508949 492168 516831
rect 492126 508940 492182 508949
rect 492126 508875 492182 508884
rect 492140 508570 492168 508875
rect 492128 508564 492180 508570
rect 492128 508506 492180 508512
rect 472624 500948 472676 500954
rect 472624 500890 472676 500896
rect 480272 500126 480608 500154
rect 481744 500126 481804 500154
rect 482664 500126 483000 500154
rect 483124 500126 484196 500154
rect 485056 500126 485392 500154
rect 486252 500126 486588 500154
rect 487172 500126 487784 500154
rect 488552 500126 488980 500154
rect 489932 500126 490176 500154
rect 491312 500126 491372 500154
rect 478142 467120 478198 467129
rect 478142 467055 478198 467064
rect 478156 458386 478184 467055
rect 474004 458380 474056 458386
rect 474004 458322 474056 458328
rect 478144 458380 478196 458386
rect 478144 458322 478196 458328
rect 474016 455940 474044 458322
rect 480272 456210 480300 500126
rect 481640 490476 481692 490482
rect 481640 490418 481692 490424
rect 481652 457502 481680 490418
rect 481744 457570 481772 500126
rect 482664 490482 482692 500126
rect 482652 490476 482704 490482
rect 482652 490418 482704 490424
rect 482008 458312 482060 458318
rect 482008 458254 482060 458260
rect 481732 457564 481784 457570
rect 481732 457506 481784 457512
rect 481640 457496 481692 457502
rect 481640 457438 481692 457444
rect 480260 456204 480312 456210
rect 480260 456146 480312 456152
rect 482020 455940 482048 458254
rect 483124 456142 483152 500126
rect 485056 497622 485084 500126
rect 485044 497616 485096 497622
rect 485044 497558 485096 497564
rect 486252 497554 486280 500126
rect 486240 497548 486292 497554
rect 486240 497490 486292 497496
rect 487172 461650 487200 500126
rect 487160 461644 487212 461650
rect 487160 461586 487212 461592
rect 488552 460222 488580 500126
rect 489932 497486 489960 500126
rect 489920 497480 489972 497486
rect 489920 497422 489972 497428
rect 488540 460216 488592 460222
rect 488540 460158 488592 460164
rect 490012 458244 490064 458250
rect 490012 458186 490064 458192
rect 483112 456136 483164 456142
rect 483112 456078 483164 456084
rect 490024 455940 490052 458186
rect 491312 456074 491340 500126
rect 491300 456068 491352 456074
rect 491300 456010 491352 456016
rect 471716 427106 471744 432140
rect 474660 430030 474688 432140
rect 474648 430024 474700 430030
rect 474648 429966 474700 429972
rect 477604 429962 477632 432140
rect 477592 429956 477644 429962
rect 477592 429898 477644 429904
rect 479524 429956 479576 429962
rect 479524 429898 479576 429904
rect 471704 427100 471756 427106
rect 471704 427042 471756 427048
rect 473360 406428 473412 406434
rect 473360 406370 473412 406376
rect 473372 402974 473400 406370
rect 473372 402946 473768 402974
rect 471888 387116 471940 387122
rect 471888 387058 471940 387064
rect 471244 383376 471296 383382
rect 471244 383318 471296 383324
rect 471900 379930 471928 387058
rect 472806 382392 472862 382401
rect 472806 382327 472862 382336
rect 471546 379902 471928 379930
rect 472820 379916 472848 382327
rect 473740 379930 473768 402946
rect 479536 384402 479564 429898
rect 480548 429894 480576 432140
rect 483032 432126 483506 432154
rect 480536 429888 480588 429894
rect 480536 429830 480588 429836
rect 479524 384396 479576 384402
rect 479524 384338 479576 384344
rect 483032 384334 483060 432126
rect 486436 429214 486464 432140
rect 489380 429962 489408 432140
rect 489368 429956 489420 429962
rect 489368 429898 489420 429904
rect 492324 429214 492352 432140
rect 485044 429208 485096 429214
rect 485044 429150 485096 429156
rect 486424 429208 486476 429214
rect 486424 429150 486476 429156
rect 490564 429208 490616 429214
rect 490564 429150 490616 429156
rect 492312 429208 492364 429214
rect 492312 429150 492364 429156
rect 485056 385694 485084 429150
rect 489182 391232 489238 391241
rect 489182 391167 489238 391176
rect 485044 385688 485096 385694
rect 485044 385630 485096 385636
rect 483020 384328 483072 384334
rect 483020 384270 483072 384276
rect 477960 383648 478012 383654
rect 477960 383590 478012 383596
rect 476672 383444 476724 383450
rect 476672 383386 476724 383392
rect 475382 382392 475438 382401
rect 475382 382327 475438 382336
rect 473740 379902 474122 379930
rect 475396 379916 475424 382327
rect 476684 379916 476712 383386
rect 477972 379916 478000 383590
rect 479248 383580 479300 383586
rect 479248 383522 479300 383528
rect 479260 379916 479288 383522
rect 481824 383512 481876 383518
rect 481824 383454 481876 383460
rect 480536 383172 480588 383178
rect 480536 383114 480588 383120
rect 480548 379916 480576 383114
rect 481836 379916 481864 383454
rect 486976 383376 487028 383382
rect 486976 383318 487028 383324
rect 485688 383308 485740 383314
rect 485688 383250 485740 383256
rect 483112 383240 483164 383246
rect 483112 383182 483164 383188
rect 483124 379916 483152 383182
rect 484400 383104 484452 383110
rect 484400 383046 484452 383052
rect 484412 379916 484440 383046
rect 485700 379916 485728 383250
rect 486988 379916 487016 383318
rect 488264 383036 488316 383042
rect 488264 382978 488316 382984
rect 488276 379916 488304 382978
rect 489196 379930 489224 391167
rect 490576 387122 490604 429150
rect 490564 387116 490616 387122
rect 490564 387058 490616 387064
rect 490838 382392 490894 382401
rect 490838 382327 490894 382336
rect 492126 382392 492182 382401
rect 492126 382327 492182 382336
rect 489196 379902 489578 379930
rect 490852 379916 490880 382327
rect 492140 379916 492168 382327
rect 493060 379930 493088 519522
rect 494072 402974 494100 592622
rect 494702 520976 494758 520985
rect 494702 520911 494758 520920
rect 494152 516792 494204 516798
rect 494152 516734 494204 516740
rect 494164 512650 494192 516734
rect 494152 512644 494204 512650
rect 494152 512586 494204 512592
rect 494164 512553 494192 512586
rect 494150 512544 494206 512553
rect 494150 512479 494206 512488
rect 494150 505200 494206 505209
rect 494150 505135 494152 505144
rect 494204 505135 494206 505144
rect 494152 505106 494204 505112
rect 494164 500954 494192 505106
rect 494152 500948 494204 500954
rect 494152 500890 494204 500896
rect 494072 402946 494376 402974
rect 494348 379930 494376 402946
rect 494716 383042 494744 520911
rect 494796 515976 494848 515982
rect 494794 515944 494796 515953
rect 494848 515944 494850 515953
rect 494794 515879 494850 515888
rect 494794 501256 494850 501265
rect 494794 501191 494850 501200
rect 494808 466546 494836 501191
rect 494796 466540 494848 466546
rect 494796 466482 494848 466488
rect 494808 458250 494836 466482
rect 494796 458244 494848 458250
rect 494796 458186 494848 458192
rect 495452 402974 495480 598198
rect 495452 402946 495664 402974
rect 494704 383036 494756 383042
rect 494704 382978 494756 382984
rect 495636 379930 495664 402946
rect 496096 381546 496124 598198
rect 496820 596828 496872 596834
rect 496820 596770 496872 596776
rect 496832 402974 496860 596770
rect 498200 537532 498252 537538
rect 498200 537474 498252 537480
rect 496832 402946 496952 402974
rect 496084 381540 496136 381546
rect 496084 381482 496136 381488
rect 496924 379930 496952 402946
rect 498212 379930 498240 537474
rect 498304 515982 498332 600086
rect 506584 600086 506690 600114
rect 514772 600086 515154 600114
rect 523618 600086 523724 600114
rect 503720 599616 503772 599622
rect 503720 599558 503772 599564
rect 502340 598324 502392 598330
rect 502340 598266 502392 598272
rect 500960 595468 501012 595474
rect 500960 595410 501012 595416
rect 499580 589960 499632 589966
rect 499580 589902 499632 589908
rect 498292 515976 498344 515982
rect 498292 515918 498344 515924
rect 498304 509930 498332 515918
rect 498292 509924 498344 509930
rect 498292 509866 498344 509872
rect 499592 379930 499620 589902
rect 500972 379930 501000 595410
rect 502352 379930 502380 598266
rect 493060 379902 493442 379930
rect 494348 379902 494730 379930
rect 495636 379902 496018 379930
rect 496924 379902 497306 379930
rect 498212 379902 498594 379930
rect 499592 379902 499882 379930
rect 500972 379902 501170 379930
rect 502352 379902 502458 379930
rect 503732 379916 503760 599558
rect 503812 591320 503864 591326
rect 503812 591262 503864 591268
rect 503824 402974 503852 591262
rect 506478 537432 506534 537441
rect 506478 537367 506534 537376
rect 506492 402974 506520 537367
rect 506584 517041 506612 600086
rect 514772 517546 514800 600086
rect 518164 599684 518216 599690
rect 518164 599626 518216 599632
rect 515404 599616 515456 599622
rect 515404 599558 515456 599564
rect 514760 517540 514812 517546
rect 514760 517482 514812 517488
rect 506570 517032 506626 517041
rect 506570 516967 506626 516976
rect 506584 512718 506612 516967
rect 514772 514078 514800 517482
rect 514760 514072 514812 514078
rect 514760 514014 514812 514020
rect 506572 512712 506624 512718
rect 506572 512654 506624 512660
rect 514024 470620 514076 470626
rect 514024 470562 514076 470568
rect 511264 465724 511316 465730
rect 511264 465666 511316 465672
rect 503824 402946 504680 402974
rect 506492 402946 507256 402974
rect 504652 379930 504680 402946
rect 506296 383036 506348 383042
rect 506296 382978 506348 382984
rect 504652 379902 505034 379930
rect 506308 379916 506336 382978
rect 507228 379930 507256 402946
rect 507228 379902 507610 379930
rect 453304 379840 453356 379846
rect 453304 379782 453356 379788
rect 510986 361176 511042 361185
rect 510986 361111 511042 361120
rect 510802 360360 510858 360369
rect 510802 360295 510858 360304
rect 510066 359136 510122 359145
rect 510066 359071 510122 359080
rect 510080 354674 510108 359071
rect 509896 354646 510108 354674
rect 450636 339312 450688 339318
rect 450636 339254 450688 339260
rect 450544 338972 450596 338978
rect 450544 338914 450596 338920
rect 450452 338428 450504 338434
rect 450452 338370 450504 338376
rect 450464 331214 450492 338370
rect 450464 331186 450584 331214
rect 450358 326632 450414 326641
rect 450358 326567 450414 326576
rect 450556 326097 450584 331186
rect 450266 326088 450322 326097
rect 450266 326023 450322 326032
rect 450542 326088 450598 326097
rect 450542 326023 450598 326032
rect 450174 325544 450230 325553
rect 450174 325479 450230 325488
rect 450082 325000 450138 325009
rect 450082 324935 450138 324944
rect 450450 323912 450506 323921
rect 450450 323847 450506 323856
rect 450464 316742 450492 323847
rect 450452 316736 450504 316742
rect 450452 316678 450504 316684
rect 450084 234660 450136 234666
rect 450084 234602 450136 234608
rect 450096 231878 450124 234602
rect 450084 231872 450136 231878
rect 450084 231814 450136 231820
rect 450556 167754 450584 326023
rect 450634 325544 450690 325553
rect 450690 325502 450860 325530
rect 450634 325479 450690 325488
rect 450634 325000 450690 325009
rect 450634 324935 450690 324944
rect 450648 315926 450676 324935
rect 450636 315920 450688 315926
rect 450636 315862 450688 315868
rect 450832 315858 450860 325502
rect 464434 320376 464490 320385
rect 464434 320311 464490 320320
rect 460018 320104 460074 320113
rect 451752 319926 451964 319954
rect 451752 319870 451780 319926
rect 451936 319870 451964 319926
rect 451740 319864 451792 319870
rect 451740 319806 451792 319812
rect 451924 319864 451976 319870
rect 451924 319806 451976 319812
rect 455938 319818 455966 320076
rect 451832 319796 451884 319802
rect 455938 319790 456012 319818
rect 451832 319738 451884 319744
rect 451740 319728 451792 319734
rect 451740 319670 451792 319676
rect 451752 319546 451780 319670
rect 451844 319666 451872 319738
rect 451924 319728 451976 319734
rect 451924 319670 451976 319676
rect 451832 319660 451884 319666
rect 451832 319602 451884 319608
rect 451936 319546 451964 319670
rect 451752 319518 451964 319546
rect 451924 316736 451976 316742
rect 451924 316678 451976 316684
rect 450820 315852 450872 315858
rect 450820 315794 450872 315800
rect 451280 268796 451332 268802
rect 451280 268738 451332 268744
rect 451292 263498 451320 268738
rect 451280 263492 451332 263498
rect 451280 263434 451332 263440
rect 451936 207262 451964 316678
rect 452016 315920 452068 315926
rect 452016 315862 452068 315868
rect 452028 222154 452056 315862
rect 453304 315852 453356 315858
rect 453304 315794 453356 315800
rect 452200 309800 452252 309806
rect 452200 309742 452252 309748
rect 452108 297356 452160 297362
rect 452108 297298 452160 297304
rect 452120 232762 452148 297298
rect 452212 285734 452240 309742
rect 452200 285728 452252 285734
rect 452200 285670 452252 285676
rect 452568 274168 452620 274174
rect 452568 274110 452620 274116
rect 452292 273284 452344 273290
rect 452292 273226 452344 273232
rect 452200 269816 452252 269822
rect 452200 269758 452252 269764
rect 452212 234666 452240 269758
rect 452304 258126 452332 273226
rect 452580 271454 452608 274110
rect 452568 271448 452620 271454
rect 452568 271390 452620 271396
rect 453028 271244 453080 271250
rect 453028 271186 453080 271192
rect 453040 268802 453068 271186
rect 453028 268796 453080 268802
rect 453028 268738 453080 268744
rect 453028 266416 453080 266422
rect 453028 266358 453080 266364
rect 453040 264994 453068 266358
rect 453028 264988 453080 264994
rect 453028 264930 453080 264936
rect 452292 258120 452344 258126
rect 452292 258062 452344 258068
rect 453316 235006 453344 315794
rect 455144 315784 455196 315790
rect 455144 315726 455196 315732
rect 454868 315716 454920 315722
rect 454868 315658 454920 315664
rect 454684 315512 454736 315518
rect 454684 315454 454736 315460
rect 453304 235000 453356 235006
rect 453304 234942 453356 234948
rect 452200 234660 452252 234666
rect 452200 234602 452252 234608
rect 452108 232756 452160 232762
rect 452108 232698 452160 232704
rect 452016 222148 452068 222154
rect 452016 222090 452068 222096
rect 451924 207256 451976 207262
rect 451924 207198 451976 207204
rect 452844 169108 452896 169114
rect 452844 169050 452896 169056
rect 450544 167748 450596 167754
rect 450544 167690 450596 167696
rect 450912 167136 450964 167142
rect 450912 167078 450964 167084
rect 449992 167068 450044 167074
rect 449992 167010 450044 167016
rect 450544 167068 450596 167074
rect 450544 167010 450596 167016
rect 450556 166326 450584 167010
rect 450924 166394 450952 167078
rect 450912 166388 450964 166394
rect 450912 166330 450964 166336
rect 450544 166320 450596 166326
rect 450544 166262 450596 166268
rect 448336 164902 448388 164908
rect 445220 164898 445708 164902
rect 445220 164892 445720 164898
rect 445220 164886 445668 164892
rect 449052 164886 449388 164914
rect 445668 164834 445720 164840
rect 452856 164642 452884 169050
rect 430652 164614 430896 164642
rect 434332 164614 434484 164642
rect 452732 164614 452884 164642
rect 423264 164384 423320 164393
rect 423264 164319 423320 164328
rect 410524 44736 410576 44742
rect 410524 44678 410576 44684
rect 454696 4010 454724 315454
rect 454774 315344 454830 315353
rect 454774 315279 454830 315288
rect 454684 4004 454736 4010
rect 454684 3946 454736 3952
rect 407856 3664 407908 3670
rect 406382 3632 406438 3641
rect 407856 3606 407908 3612
rect 406382 3567 406438 3576
rect 454788 3505 454816 315279
rect 454880 45354 454908 315658
rect 454960 315444 455012 315450
rect 454960 315386 455012 315392
rect 454972 45422 455000 315386
rect 455052 315308 455104 315314
rect 455052 315250 455104 315256
rect 455064 50289 455092 315250
rect 455156 51066 455184 315726
rect 455236 315172 455288 315178
rect 455236 315114 455288 315120
rect 455248 52018 455276 315114
rect 455984 313954 456012 319790
rect 456064 315648 456116 315654
rect 456064 315590 456116 315596
rect 455972 313948 456024 313954
rect 455972 313890 456024 313896
rect 455236 52012 455288 52018
rect 455236 51954 455288 51960
rect 455144 51060 455196 51066
rect 455144 51002 455196 51008
rect 455050 50280 455106 50289
rect 455050 50215 455106 50224
rect 454960 45416 455012 45422
rect 454960 45358 455012 45364
rect 454868 45348 454920 45354
rect 454868 45290 454920 45296
rect 454774 3496 454830 3505
rect 456076 3466 456104 315590
rect 456168 314906 456196 320076
rect 456340 317892 456392 317898
rect 456340 317834 456392 317840
rect 456248 315580 456300 315586
rect 456248 315522 456300 315528
rect 456156 314900 456208 314906
rect 456156 314842 456208 314848
rect 456260 313698 456288 315522
rect 456168 313670 456288 313698
rect 456168 3534 456196 313670
rect 456248 312588 456300 312594
rect 456248 312530 456300 312536
rect 456260 36582 456288 312530
rect 456352 52057 456380 317834
rect 456444 315246 456472 320076
rect 456720 316010 456748 320076
rect 456996 316130 457024 320076
rect 456984 316124 457036 316130
rect 456984 316066 457036 316072
rect 457272 316062 457300 320076
rect 456536 315982 456748 316010
rect 457260 316056 457312 316062
rect 457260 315998 457312 316004
rect 456432 315240 456484 315246
rect 456432 315182 456484 315188
rect 456536 311166 456564 315982
rect 456708 315240 456760 315246
rect 456708 315182 456760 315188
rect 456616 314900 456668 314906
rect 456616 314842 456668 314848
rect 456524 311160 456576 311166
rect 456524 311102 456576 311108
rect 456628 308446 456656 314842
rect 456616 308440 456668 308446
rect 456616 308382 456668 308388
rect 456720 302870 456748 315182
rect 457548 311894 457576 320076
rect 457824 315246 457852 320076
rect 458100 318170 458128 320076
rect 458376 318714 458404 320076
rect 458364 318708 458416 318714
rect 458364 318650 458416 318656
rect 458088 318164 458140 318170
rect 458088 318106 458140 318112
rect 458652 317286 458680 320076
rect 458640 317280 458692 317286
rect 458640 317222 458692 317228
rect 458928 317218 458956 320076
rect 458916 317212 458968 317218
rect 458916 317154 458968 317160
rect 459204 317150 459232 320076
rect 459480 317422 459508 320076
rect 459468 317416 459520 317422
rect 459468 317358 459520 317364
rect 459756 317354 459784 320076
rect 460018 320039 460074 320048
rect 460308 318578 460336 320076
rect 460584 318646 460612 320076
rect 460860 319326 460888 320076
rect 461136 319841 461164 320076
rect 461122 319832 461178 319841
rect 461412 319802 461440 320076
rect 461584 320000 461636 320006
rect 461688 319954 461716 320076
rect 461636 319948 461716 319954
rect 461584 319942 461716 319948
rect 461596 319926 461716 319942
rect 461122 319767 461178 319776
rect 461400 319796 461452 319802
rect 461400 319738 461452 319744
rect 461964 319569 461992 320076
rect 462134 319968 462190 319977
rect 462240 319954 462268 320076
rect 462190 319926 462268 319954
rect 462516 319938 462544 320076
rect 462504 319932 462556 319938
rect 462134 319903 462190 319912
rect 462504 319874 462556 319880
rect 461950 319560 462006 319569
rect 461950 319495 462006 319504
rect 460848 319320 460900 319326
rect 460848 319262 460900 319268
rect 461032 319184 461084 319190
rect 461032 319126 461084 319132
rect 461044 319054 461072 319126
rect 461032 319048 461084 319054
rect 461032 318990 461084 318996
rect 460572 318640 460624 318646
rect 460572 318582 460624 318588
rect 460296 318572 460348 318578
rect 460296 318514 460348 318520
rect 462792 318306 462820 320076
rect 462780 318300 462832 318306
rect 462780 318242 462832 318248
rect 462228 318164 462280 318170
rect 462228 318106 462280 318112
rect 461584 318096 461636 318102
rect 461584 318038 461636 318044
rect 461596 317898 461624 318038
rect 462240 317898 462268 318106
rect 461584 317892 461636 317898
rect 461584 317834 461636 317840
rect 462228 317892 462280 317898
rect 462228 317834 462280 317840
rect 460204 317484 460256 317490
rect 460204 317426 460256 317432
rect 459744 317348 459796 317354
rect 459744 317290 459796 317296
rect 459192 317144 459244 317150
rect 459192 317086 459244 317092
rect 457904 316124 457956 316130
rect 457904 316066 457956 316072
rect 457812 315240 457864 315246
rect 457812 315182 457864 315188
rect 457548 311866 457852 311894
rect 457444 307828 457496 307834
rect 457444 307770 457496 307776
rect 456708 302864 456760 302870
rect 456708 302806 456760 302812
rect 457456 297362 457484 307770
rect 457444 297356 457496 297362
rect 457444 297298 457496 297304
rect 457824 296070 457852 311866
rect 457916 301510 457944 316066
rect 457996 316056 458048 316062
rect 457996 315998 458048 316004
rect 457904 301504 457956 301510
rect 457904 301446 457956 301452
rect 458008 297362 458036 315998
rect 459008 314016 459060 314022
rect 459008 313958 459060 313964
rect 458824 312656 458876 312662
rect 458824 312598 458876 312604
rect 458180 306128 458232 306134
rect 458180 306070 458232 306076
rect 458192 304434 458220 306070
rect 458180 304428 458232 304434
rect 458180 304370 458232 304376
rect 457996 297356 458048 297362
rect 457996 297298 458048 297304
rect 457812 296064 457864 296070
rect 457812 296006 457864 296012
rect 457444 294500 457496 294506
rect 457444 294442 457496 294448
rect 456708 268728 456760 268734
rect 456708 268670 456760 268676
rect 456720 266422 456748 268670
rect 456708 266416 456760 266422
rect 456708 266358 456760 266364
rect 456800 263560 456852 263566
rect 456800 263502 456852 263508
rect 456812 262721 456840 263502
rect 456798 262712 456854 262721
rect 456798 262647 456854 262656
rect 457168 235000 457220 235006
rect 457166 234968 457168 234977
rect 457220 234968 457222 234977
rect 457166 234903 457222 234912
rect 457352 222148 457404 222154
rect 457352 222090 457404 222096
rect 457364 221105 457392 222090
rect 457350 221096 457406 221105
rect 457350 221031 457406 221040
rect 456800 207256 456852 207262
rect 456798 207224 456800 207233
rect 456852 207224 456854 207233
rect 456798 207159 456854 207168
rect 457258 207224 457314 207233
rect 457258 207159 457314 207168
rect 456800 168088 456852 168094
rect 456800 168030 456852 168036
rect 456812 167686 456840 168030
rect 457272 168026 457300 207159
rect 457260 168020 457312 168026
rect 457260 167962 457312 167968
rect 456892 167952 456944 167958
rect 456892 167894 456944 167900
rect 456904 167822 456932 167894
rect 456892 167816 456944 167822
rect 456892 167758 456944 167764
rect 456800 167680 456852 167686
rect 456800 167622 456852 167628
rect 457272 167618 457300 167962
rect 457364 167958 457392 221031
rect 457352 167952 457404 167958
rect 457352 167894 457404 167900
rect 457260 167612 457312 167618
rect 457260 167554 457312 167560
rect 456800 161288 456852 161294
rect 456800 161230 456852 161236
rect 456812 161129 456840 161230
rect 456798 161120 456854 161129
rect 456798 161055 456854 161064
rect 456800 159996 456852 160002
rect 456800 159938 456852 159944
rect 456812 159633 456840 159938
rect 456798 159624 456854 159633
rect 456798 159559 456854 159568
rect 456800 157072 456852 157078
rect 456800 157014 456852 157020
rect 456812 156641 456840 157014
rect 456798 156632 456854 156641
rect 456798 156567 456854 156576
rect 456800 155372 456852 155378
rect 456800 155314 456852 155320
rect 456812 155145 456840 155314
rect 456798 155136 456854 155145
rect 456798 155071 456854 155080
rect 456800 154148 456852 154154
rect 456800 154090 456852 154096
rect 456812 153649 456840 154090
rect 456798 153640 456854 153649
rect 456798 153575 456854 153584
rect 456892 150680 456944 150686
rect 456890 150648 456892 150657
rect 456944 150648 456946 150657
rect 456890 150583 456946 150592
rect 456800 150204 456852 150210
rect 456800 150146 456852 150152
rect 456812 149161 456840 150146
rect 456798 149152 456854 149161
rect 456798 149087 456854 149096
rect 457456 147665 457484 294442
rect 457720 283620 457772 283626
rect 457720 283562 457772 283568
rect 457628 276684 457680 276690
rect 457628 276626 457680 276632
rect 457536 273964 457588 273970
rect 457536 273906 457588 273912
rect 457442 147656 457498 147665
rect 457442 147591 457498 147600
rect 456800 144696 456852 144702
rect 456798 144664 456800 144673
rect 456852 144664 456854 144673
rect 456798 144599 456854 144608
rect 456800 143200 456852 143206
rect 456798 143168 456800 143177
rect 456852 143168 456854 143177
rect 456798 143103 456854 143112
rect 457260 141704 457312 141710
rect 457258 141672 457260 141681
rect 457312 141672 457314 141681
rect 457258 141607 457314 141616
rect 456800 140480 456852 140486
rect 456800 140422 456852 140428
rect 456812 140185 456840 140422
rect 456798 140176 456854 140185
rect 456798 140111 456854 140120
rect 457260 138916 457312 138922
rect 457260 138858 457312 138864
rect 457272 138689 457300 138858
rect 457258 138680 457314 138689
rect 457258 138615 457314 138624
rect 457260 137896 457312 137902
rect 457260 137838 457312 137844
rect 457272 137193 457300 137838
rect 457258 137184 457314 137193
rect 457258 137119 457314 137128
rect 457548 134201 457576 273906
rect 457640 146169 457668 276626
rect 457732 152153 457760 283562
rect 457812 279472 457864 279478
rect 457812 279414 457864 279420
rect 457824 158137 457852 279414
rect 458088 278112 458140 278118
rect 458088 278054 458140 278060
rect 458100 274174 458128 278054
rect 458180 275460 458232 275466
rect 458180 275402 458232 275408
rect 458088 274168 458140 274174
rect 458088 274110 458140 274116
rect 458192 271250 458220 275402
rect 458732 272536 458784 272542
rect 458732 272478 458784 272484
rect 458180 271244 458232 271250
rect 458180 271186 458232 271192
rect 458640 271176 458692 271182
rect 458640 271118 458692 271124
rect 457904 268524 457956 268530
rect 457904 268466 457956 268472
rect 457916 162625 457944 268466
rect 457996 249076 458048 249082
rect 457996 249018 458048 249024
rect 458008 248849 458036 249018
rect 457994 248840 458050 248849
rect 457994 248775 458050 248784
rect 458008 167686 458036 248775
rect 458086 234968 458142 234977
rect 458086 234903 458142 234912
rect 458100 167890 458128 234903
rect 458088 167884 458140 167890
rect 458088 167826 458140 167832
rect 457996 167680 458048 167686
rect 457996 167622 458048 167628
rect 457902 162616 457958 162625
rect 457902 162551 457958 162560
rect 457810 158128 457866 158137
rect 457810 158063 457866 158072
rect 458652 154154 458680 271118
rect 458744 155378 458772 272478
rect 458732 155372 458784 155378
rect 458732 155314 458784 155320
rect 458640 154148 458692 154154
rect 458640 154090 458692 154096
rect 457718 152144 457774 152153
rect 457718 152079 457774 152088
rect 457626 146160 457682 146169
rect 457626 146095 457682 146104
rect 458836 144702 458864 312598
rect 458916 311228 458968 311234
rect 458916 311170 458968 311176
rect 458928 157078 458956 311170
rect 459020 161294 459048 313958
rect 459100 309868 459152 309874
rect 459100 309810 459152 309816
rect 459008 161288 459060 161294
rect 459008 161230 459060 161236
rect 459112 160002 459140 309810
rect 459560 278044 459612 278050
rect 459560 277986 459612 277992
rect 459572 273290 459600 277986
rect 459560 273284 459612 273290
rect 459560 273226 459612 273232
rect 459376 271244 459428 271250
rect 459376 271186 459428 271192
rect 459284 268456 459336 268462
rect 459284 268398 459336 268404
rect 459192 268388 459244 268394
rect 459192 268330 459244 268336
rect 459100 159996 459152 160002
rect 459100 159938 459152 159944
rect 458916 157072 458968 157078
rect 458916 157014 458968 157020
rect 458824 144696 458876 144702
rect 458824 144638 458876 144644
rect 459204 140486 459232 268330
rect 459296 143206 459324 268398
rect 459388 150686 459416 271186
rect 460112 269952 460164 269958
rect 460112 269894 460164 269900
rect 459468 269884 459520 269890
rect 459468 269826 459520 269832
rect 459376 150680 459428 150686
rect 459376 150622 459428 150628
rect 459480 150210 459508 269826
rect 459468 150204 459520 150210
rect 459468 150146 459520 150152
rect 459284 143200 459336 143206
rect 459284 143142 459336 143148
rect 460124 141710 460152 269894
rect 460112 141704 460164 141710
rect 460112 141646 460164 141652
rect 459192 140480 459244 140486
rect 459192 140422 459244 140428
rect 457534 134192 457590 134201
rect 457534 134127 457590 134136
rect 457076 132932 457128 132938
rect 457076 132874 457128 132880
rect 457088 132705 457116 132874
rect 457074 132696 457130 132705
rect 457074 132631 457130 132640
rect 457444 128240 457496 128246
rect 457442 128208 457444 128217
rect 457496 128208 457498 128217
rect 457442 128143 457498 128152
rect 457352 125248 457404 125254
rect 457350 125216 457352 125225
rect 457404 125216 457406 125225
rect 457350 125151 457406 125160
rect 457076 122596 457128 122602
rect 457076 122538 457128 122544
rect 457088 122233 457116 122538
rect 457074 122224 457130 122233
rect 457074 122159 457130 122168
rect 460216 52086 460244 317426
rect 463068 316470 463096 320076
rect 463344 318782 463372 320076
rect 463332 318776 463384 318782
rect 463332 318718 463384 318724
rect 463620 316538 463648 320076
rect 463896 316606 463924 320076
rect 463884 316600 463936 316606
rect 463884 316542 463936 316548
rect 463608 316532 463660 316538
rect 463608 316474 463660 316480
rect 463056 316464 463108 316470
rect 463056 316406 463108 316412
rect 464172 315246 464200 320076
rect 461584 315240 461636 315246
rect 461584 315182 461636 315188
rect 463608 315240 463660 315246
rect 463608 315182 463660 315188
rect 464160 315240 464212 315246
rect 464160 315182 464212 315188
rect 460480 314152 460532 314158
rect 460480 314094 460532 314100
rect 460296 312792 460348 312798
rect 460296 312734 460348 312740
rect 460308 122602 460336 312734
rect 460388 312724 460440 312730
rect 460388 312666 460440 312672
rect 460400 125254 460428 312666
rect 460492 137902 460520 314094
rect 460572 311364 460624 311370
rect 460572 311306 460624 311312
rect 460584 306066 460612 311306
rect 460572 306060 460624 306066
rect 460572 306002 460624 306008
rect 461596 299470 461624 315182
rect 462228 314628 462280 314634
rect 462228 314570 462280 314576
rect 461768 311296 461820 311302
rect 461768 311238 461820 311244
rect 461780 306134 461808 311238
rect 462240 307834 462268 314570
rect 463620 311302 463648 315182
rect 464724 311894 464752 320076
rect 465000 314634 465028 320076
rect 464988 314628 465040 314634
rect 464988 314570 465040 314576
rect 465276 311894 465304 320076
rect 465552 315178 465580 320076
rect 465828 317490 465856 320076
rect 465816 317484 465868 317490
rect 465816 317426 465868 317432
rect 465540 315172 465592 315178
rect 465540 315114 465592 315120
rect 466104 313290 466132 320076
rect 463988 311866 464752 311894
rect 465184 311866 465304 311894
rect 465368 313262 466132 313290
rect 463608 311296 463660 311302
rect 463608 311238 463660 311244
rect 463988 309806 464016 311866
rect 465184 311370 465212 311866
rect 465172 311364 465224 311370
rect 465172 311306 465224 311312
rect 463976 309800 464028 309806
rect 463976 309742 464028 309748
rect 462228 307828 462280 307834
rect 462228 307770 462280 307776
rect 461768 306128 461820 306134
rect 461768 306070 461820 306076
rect 465368 302802 465396 313262
rect 465816 312860 465868 312866
rect 465816 312802 465868 312808
rect 465724 307828 465776 307834
rect 465724 307770 465776 307776
rect 465356 302796 465408 302802
rect 465356 302738 465408 302744
rect 461584 299464 461636 299470
rect 461584 299406 461636 299412
rect 461676 285728 461728 285734
rect 461676 285670 461728 285676
rect 461688 283694 461716 285670
rect 461676 283688 461728 283694
rect 461676 283630 461728 283636
rect 464344 282124 464396 282130
rect 464344 282066 464396 282072
rect 464356 275466 464384 282066
rect 464344 275460 464396 275466
rect 464344 275402 464396 275408
rect 460664 275392 460716 275398
rect 460664 275334 460716 275340
rect 460572 274032 460624 274038
rect 460572 273974 460624 273980
rect 460480 137896 460532 137902
rect 460480 137838 460532 137844
rect 460584 128246 460612 273974
rect 460676 132938 460704 275334
rect 463332 271856 463384 271862
rect 463332 271798 463384 271804
rect 460756 270020 460808 270026
rect 460756 269962 460808 269968
rect 460768 138922 460796 269962
rect 463344 269822 463372 271798
rect 463332 269816 463384 269822
rect 463332 269758 463384 269764
rect 465736 268666 465764 307770
rect 465828 285734 465856 312802
rect 466380 290494 466408 320076
rect 466656 311894 466684 320076
rect 466932 313886 466960 320076
rect 467208 316010 467236 320076
rect 467484 318794 467512 320076
rect 467484 318766 467604 318794
rect 467208 315982 467512 316010
rect 466920 313880 466972 313886
rect 466920 313822 466972 313828
rect 466656 311866 467420 311894
rect 467392 304434 467420 311866
rect 467380 304428 467432 304434
rect 467380 304370 467432 304376
rect 467484 293282 467512 315982
rect 467576 314226 467604 318766
rect 467760 314378 467788 320076
rect 467668 314350 467788 314378
rect 467564 314220 467616 314226
rect 467564 314162 467616 314168
rect 467564 313880 467616 313886
rect 467564 313822 467616 313828
rect 467472 293276 467524 293282
rect 467472 293218 467524 293224
rect 467576 291786 467604 313822
rect 467564 291780 467616 291786
rect 467564 291722 467616 291728
rect 466368 290488 466420 290494
rect 466368 290430 466420 290436
rect 467668 287706 467696 314350
rect 467748 314220 467800 314226
rect 467748 314162 467800 314168
rect 467656 287700 467708 287706
rect 467656 287642 467708 287648
rect 465816 285728 465868 285734
rect 465816 285670 465868 285676
rect 466184 285660 466236 285666
rect 466184 285602 466236 285608
rect 466196 282130 466224 285602
rect 466460 284368 466512 284374
rect 466460 284310 466512 284316
rect 466184 282124 466236 282130
rect 466184 282066 466236 282072
rect 466472 281602 466500 284310
rect 466380 281574 466500 281602
rect 466380 278118 466408 281574
rect 467760 280838 467788 314162
rect 468036 311894 468064 320076
rect 468312 313274 468340 320076
rect 468588 319938 468616 320076
rect 468576 319932 468628 319938
rect 468576 319874 468628 319880
rect 468864 318442 468892 320076
rect 469140 319666 469168 320076
rect 469128 319660 469180 319666
rect 469128 319602 469180 319608
rect 468852 318436 468904 318442
rect 468852 318378 468904 318384
rect 469416 318374 469444 320076
rect 469692 319802 469720 320076
rect 469680 319796 469732 319802
rect 469680 319738 469732 319744
rect 469968 318646 469996 320076
rect 470244 319938 470272 320076
rect 470232 319932 470284 319938
rect 470232 319874 470284 319880
rect 469956 318640 470008 318646
rect 469956 318582 470008 318588
rect 470520 318578 470548 320076
rect 470508 318572 470560 318578
rect 470508 318514 470560 318520
rect 469404 318368 469456 318374
rect 469404 318310 469456 318316
rect 470796 317694 470824 320076
rect 471072 318510 471100 320076
rect 471244 319524 471296 319530
rect 471244 319466 471296 319472
rect 471256 319054 471284 319466
rect 471244 319048 471296 319054
rect 471244 318990 471296 318996
rect 471060 318504 471112 318510
rect 471060 318446 471112 318452
rect 471348 317830 471376 320076
rect 471624 317966 471652 320076
rect 471612 317960 471664 317966
rect 471612 317902 471664 317908
rect 471336 317824 471388 317830
rect 471336 317766 471388 317772
rect 470784 317688 470836 317694
rect 470784 317630 470836 317636
rect 471900 317014 471928 320076
rect 472176 318238 472204 320076
rect 472164 318232 472216 318238
rect 472164 318174 472216 318180
rect 471980 317552 472032 317558
rect 471980 317494 472032 317500
rect 471888 317008 471940 317014
rect 471888 316950 471940 316956
rect 471992 315382 472020 317494
rect 472452 316674 472480 320076
rect 472728 318345 472756 320076
rect 473004 319122 473032 320076
rect 472992 319116 473044 319122
rect 472992 319058 473044 319064
rect 472714 318336 472770 318345
rect 472714 318271 472770 318280
rect 472716 317484 472768 317490
rect 472716 317426 472768 317432
rect 472440 316668 472492 316674
rect 472440 316610 472492 316616
rect 471980 315376 472032 315382
rect 471980 315318 472032 315324
rect 468300 313268 468352 313274
rect 468300 313210 468352 313216
rect 472624 313064 472676 313070
rect 472624 313006 472676 313012
rect 468036 311866 468984 311894
rect 468484 290420 468536 290426
rect 468484 290362 468536 290368
rect 467840 288380 467892 288386
rect 467840 288322 467892 288328
rect 467852 285734 467880 288322
rect 467840 285728 467892 285734
rect 467840 285670 467892 285676
rect 468496 284374 468524 290362
rect 468484 284368 468536 284374
rect 468484 284310 468536 284316
rect 467748 280832 467800 280838
rect 467748 280774 467800 280780
rect 466368 278112 466420 278118
rect 466368 278054 466420 278060
rect 468956 269822 468984 311866
rect 470600 298988 470652 298994
rect 470600 298930 470652 298936
rect 470612 295338 470640 298930
rect 470520 295310 470640 295338
rect 470520 290426 470548 295310
rect 471980 292596 472032 292602
rect 471980 292538 472032 292544
rect 470508 290420 470560 290426
rect 470508 290362 470560 290368
rect 471992 289898 472020 292538
rect 471900 289870 472020 289898
rect 471900 288454 471928 289870
rect 471888 288448 471940 288454
rect 471888 288390 471940 288396
rect 471520 285728 471572 285734
rect 471520 285670 471572 285676
rect 469864 284776 469916 284782
rect 469864 284718 469916 284724
rect 469876 271930 469904 284718
rect 471532 278050 471560 285670
rect 472636 284782 472664 313006
rect 472728 307834 472756 317426
rect 473280 316878 473308 320076
rect 473556 318034 473584 320076
rect 473544 318028 473596 318034
rect 473544 317970 473596 317976
rect 473832 316946 473860 320076
rect 473820 316940 473872 316946
rect 473820 316882 473872 316888
rect 473268 316872 473320 316878
rect 473268 316814 473320 316820
rect 474108 316810 474136 320076
rect 474384 319870 474412 320076
rect 474372 319864 474424 319870
rect 474372 319806 474424 319812
rect 474096 316804 474148 316810
rect 474096 316746 474148 316752
rect 473360 315240 473412 315246
rect 473360 315182 473412 315188
rect 473372 312866 473400 315182
rect 474660 313070 474688 320076
rect 474936 317558 474964 320076
rect 474924 317552 474976 317558
rect 474924 317494 474976 317500
rect 475212 317490 475240 320076
rect 475200 317484 475252 317490
rect 475200 317426 475252 317432
rect 474648 313064 474700 313070
rect 474648 313006 474700 313012
rect 473360 312860 473412 312866
rect 473360 312802 473412 312808
rect 475488 311894 475516 320076
rect 475764 314090 475792 320076
rect 476040 315790 476068 320076
rect 476316 317966 476344 320076
rect 476304 317960 476356 317966
rect 476304 317902 476356 317908
rect 476592 316034 476620 320076
rect 476868 318050 476896 320076
rect 477144 318186 477172 320076
rect 477420 318322 477448 320076
rect 477420 318294 477540 318322
rect 477144 318158 477448 318186
rect 476868 318022 477356 318050
rect 477132 317960 477184 317966
rect 477132 317902 477184 317908
rect 476224 316006 476620 316034
rect 476028 315784 476080 315790
rect 476028 315726 476080 315732
rect 475752 314084 475804 314090
rect 475752 314026 475804 314032
rect 475028 311866 475516 311894
rect 472716 307828 472768 307834
rect 472716 307770 472768 307776
rect 473360 306332 473412 306338
rect 473360 306274 473412 306280
rect 472716 303680 472768 303686
rect 472716 303622 472768 303628
rect 472624 284776 472676 284782
rect 472624 284718 472676 284724
rect 472728 282198 472756 303622
rect 473372 298994 473400 306274
rect 474004 306060 474056 306066
rect 474004 306002 474056 306008
rect 473360 298988 473412 298994
rect 473360 298930 473412 298936
rect 474016 285734 474044 306002
rect 475028 303686 475056 311866
rect 475016 303680 475068 303686
rect 475016 303622 475068 303628
rect 475108 298988 475160 298994
rect 475108 298930 475160 298936
rect 475120 292602 475148 298930
rect 475108 292596 475160 292602
rect 475108 292538 475160 292544
rect 476224 286482 476252 316006
rect 477144 309806 477172 317902
rect 477224 310480 477276 310486
rect 477224 310422 477276 310428
rect 477132 309800 477184 309806
rect 477132 309742 477184 309748
rect 477236 306406 477264 310422
rect 477224 306400 477276 306406
rect 477224 306342 477276 306348
rect 477328 305930 477356 318022
rect 477316 305924 477368 305930
rect 477316 305866 477368 305872
rect 477420 300014 477448 318158
rect 477512 317966 477540 318294
rect 477696 318034 477724 320076
rect 477972 318102 478000 320076
rect 477960 318096 478012 318102
rect 477960 318038 478012 318044
rect 477684 318028 477736 318034
rect 477684 317970 477736 317976
rect 477500 317960 477552 317966
rect 477500 317902 477552 317908
rect 478248 316034 478276 320076
rect 478524 318170 478552 320076
rect 478800 318782 478828 320076
rect 479076 319258 479104 320076
rect 479064 319252 479116 319258
rect 479064 319194 479116 319200
rect 478788 318776 478840 318782
rect 478788 318718 478840 318724
rect 479352 318238 479380 320076
rect 479340 318232 479392 318238
rect 479340 318174 479392 318180
rect 478512 318164 478564 318170
rect 478512 318106 478564 318112
rect 479524 318164 479576 318170
rect 479524 318106 479576 318112
rect 478604 318096 478656 318102
rect 478604 318038 478656 318044
rect 478248 316006 478552 316034
rect 478144 302252 478196 302258
rect 478144 302194 478196 302200
rect 477500 301980 477552 301986
rect 477500 301922 477552 301928
rect 477408 300008 477460 300014
rect 477408 299950 477460 299956
rect 477512 298994 477540 301922
rect 477500 298988 477552 298994
rect 477500 298930 477552 298936
rect 478156 292602 478184 302194
rect 478524 294574 478552 316006
rect 478616 315382 478644 318038
rect 478696 318028 478748 318034
rect 478696 317970 478748 317976
rect 478604 315376 478656 315382
rect 478604 315318 478656 315324
rect 478708 307086 478736 317970
rect 478696 307080 478748 307086
rect 478696 307022 478748 307028
rect 478512 294568 478564 294574
rect 478512 294510 478564 294516
rect 476764 292596 476816 292602
rect 476764 292538 476816 292544
rect 478144 292596 478196 292602
rect 478144 292538 478196 292544
rect 476212 286476 476264 286482
rect 476212 286418 476264 286424
rect 474004 285728 474056 285734
rect 474004 285670 474056 285676
rect 472716 282192 472768 282198
rect 472716 282134 472768 282140
rect 471520 278044 471572 278050
rect 471520 277986 471572 277992
rect 476776 271930 476804 292538
rect 479536 288998 479564 318106
rect 479628 317830 479656 320076
rect 479904 318306 479932 320076
rect 480180 318510 480208 320076
rect 480456 318782 480484 320076
rect 480444 318776 480496 318782
rect 480444 318718 480496 318724
rect 480168 318504 480220 318510
rect 480168 318446 480220 318452
rect 480732 318345 480760 320076
rect 480718 318336 480774 318345
rect 479892 318300 479944 318306
rect 480718 318271 480774 318280
rect 479892 318242 479944 318248
rect 481008 318238 481036 320076
rect 480996 318232 481048 318238
rect 480996 318174 481048 318180
rect 481284 318050 481312 320076
rect 481456 319456 481508 319462
rect 481456 319398 481508 319404
rect 481468 318850 481496 319398
rect 481456 318844 481508 318850
rect 481456 318786 481508 318792
rect 481456 318232 481508 318238
rect 481456 318174 481508 318180
rect 480272 318022 481312 318050
rect 481468 318034 481496 318174
rect 481456 318028 481508 318034
rect 479616 317824 479668 317830
rect 479616 317766 479668 317772
rect 480272 315926 480300 318022
rect 481456 317970 481508 317976
rect 481560 317966 481588 320076
rect 480352 317960 480404 317966
rect 480352 317902 480404 317908
rect 481548 317960 481600 317966
rect 481548 317902 481600 317908
rect 480260 315920 480312 315926
rect 480260 315862 480312 315868
rect 480364 315858 480392 317902
rect 481836 317082 481864 320076
rect 482112 317762 482140 320076
rect 482388 318481 482416 320076
rect 482664 319054 482692 320076
rect 482652 319048 482704 319054
rect 482652 318990 482704 318996
rect 482374 318472 482430 318481
rect 482374 318407 482430 318416
rect 482100 317756 482152 317762
rect 482100 317698 482152 317704
rect 481824 317076 481876 317082
rect 481824 317018 481876 317024
rect 482940 316962 482968 320076
rect 483216 318753 483244 320076
rect 483202 318744 483258 318753
rect 483202 318679 483258 318688
rect 483492 318617 483520 320076
rect 483768 319394 483796 320076
rect 484044 319598 484072 320076
rect 484032 319592 484084 319598
rect 484032 319534 484084 319540
rect 483756 319388 483808 319394
rect 483756 319330 483808 319336
rect 484320 319190 484348 320076
rect 484596 319734 484624 320076
rect 484584 319728 484636 319734
rect 484584 319670 484636 319676
rect 484308 319184 484360 319190
rect 484308 319126 484360 319132
rect 483478 318608 483534 318617
rect 483478 318543 483534 318552
rect 484492 318096 484544 318102
rect 484872 318050 484900 320076
rect 485044 319864 485096 319870
rect 485044 319806 485096 319812
rect 485056 319258 485084 319806
rect 485044 319252 485096 319258
rect 485044 319194 485096 319200
rect 484492 318038 484544 318044
rect 481836 316934 482968 316962
rect 481640 316872 481692 316878
rect 481640 316814 481692 316820
rect 480352 315852 480404 315858
rect 480352 315794 480404 315800
rect 481652 314702 481680 316814
rect 481836 315994 481864 316934
rect 481824 315988 481876 315994
rect 481824 315930 481876 315936
rect 481640 314696 481692 314702
rect 481640 314638 481692 314644
rect 479616 314628 479668 314634
rect 479616 314570 479668 314576
rect 481548 314628 481600 314634
rect 481548 314570 481600 314576
rect 479628 302258 479656 314570
rect 481560 310554 481588 314570
rect 481548 310548 481600 310554
rect 481548 310490 481600 310496
rect 483756 307760 483808 307766
rect 483756 307702 483808 307708
rect 483768 303822 483796 307702
rect 484504 306066 484532 318038
rect 484596 318022 484900 318050
rect 484596 314702 484624 318022
rect 484676 317960 484728 317966
rect 484676 317902 484728 317908
rect 484584 314696 484636 314702
rect 484584 314638 484636 314644
rect 484492 306060 484544 306066
rect 484492 306002 484544 306008
rect 481272 303816 481324 303822
rect 481272 303758 481324 303764
rect 483756 303816 483808 303822
rect 483756 303758 483808 303764
rect 479616 302252 479668 302258
rect 479616 302194 479668 302200
rect 481284 301986 481312 303758
rect 481272 301980 481324 301986
rect 481272 301922 481324 301928
rect 479524 288992 479576 288998
rect 479524 288934 479576 288940
rect 484688 274718 484716 317902
rect 485044 317688 485096 317694
rect 485044 317630 485096 317636
rect 485056 307766 485084 317630
rect 485148 316878 485176 320076
rect 485424 318102 485452 320076
rect 485412 318096 485464 318102
rect 485412 318038 485464 318044
rect 485700 317966 485728 320076
rect 485872 318096 485924 318102
rect 485872 318038 485924 318044
rect 485976 318050 486004 320076
rect 485688 317960 485740 317966
rect 485688 317902 485740 317908
rect 485136 316872 485188 316878
rect 485136 316814 485188 316820
rect 485044 307760 485096 307766
rect 485044 307702 485096 307708
rect 485884 293350 485912 318038
rect 485976 318022 486188 318050
rect 485964 317960 486016 317966
rect 485964 317902 486016 317908
rect 485976 305998 486004 317902
rect 486056 317756 486108 317762
rect 486056 317698 486108 317704
rect 485964 305992 486016 305998
rect 485964 305934 486016 305940
rect 485872 293344 485924 293350
rect 485872 293286 485924 293292
rect 486068 291718 486096 317698
rect 486160 315246 486188 318022
rect 486252 317694 486280 320076
rect 486528 317966 486556 320076
rect 486804 318102 486832 320076
rect 486792 318096 486844 318102
rect 486792 318038 486844 318044
rect 486516 317960 486568 317966
rect 486516 317902 486568 317908
rect 487080 317762 487108 320076
rect 487160 318232 487212 318238
rect 487160 318174 487212 318180
rect 487068 317756 487120 317762
rect 487068 317698 487120 317704
rect 486240 317688 486292 317694
rect 486240 317630 486292 317636
rect 486148 315240 486200 315246
rect 486148 315182 486200 315188
rect 486056 291712 486108 291718
rect 486056 291654 486108 291660
rect 482468 274712 482520 274718
rect 482468 274654 482520 274660
rect 484676 274712 484728 274718
rect 484676 274654 484728 274660
rect 469864 271924 469916 271930
rect 469864 271866 469916 271872
rect 476764 271924 476816 271930
rect 476764 271866 476816 271872
rect 472716 271856 472768 271862
rect 472716 271798 472768 271804
rect 468944 269816 468996 269822
rect 468944 269758 468996 269764
rect 472728 268734 472756 271798
rect 482480 270094 482508 274654
rect 473268 270088 473320 270094
rect 473268 270030 473320 270036
rect 482468 270088 482520 270094
rect 482468 270030 482520 270036
rect 472716 268728 472768 268734
rect 472716 268670 472768 268676
rect 465724 268660 465776 268666
rect 465724 268602 465776 268608
rect 473280 268598 473308 270030
rect 473268 268592 473320 268598
rect 473268 268534 473320 268540
rect 487172 268530 487200 318174
rect 487356 316034 487384 320076
rect 487632 318102 487660 320076
rect 487620 318096 487672 318102
rect 487620 318038 487672 318044
rect 487908 318034 487936 320076
rect 488184 318050 488212 320076
rect 488460 318238 488488 320076
rect 488736 318288 488764 320076
rect 488552 318260 488764 318288
rect 488448 318232 488500 318238
rect 488448 318174 488500 318180
rect 488356 318096 488408 318102
rect 487896 318028 487948 318034
rect 488184 318022 488304 318050
rect 488356 318038 488408 318044
rect 487896 317970 487948 317976
rect 487356 316006 488212 316034
rect 488184 307222 488212 316006
rect 488172 307216 488224 307222
rect 488172 307158 488224 307164
rect 488276 304570 488304 318022
rect 488264 304564 488316 304570
rect 488264 304506 488316 304512
rect 488368 293350 488396 318038
rect 488448 318028 488500 318034
rect 488448 317970 488500 317976
rect 488356 293344 488408 293350
rect 488356 293286 488408 293292
rect 488460 278118 488488 317970
rect 488552 312798 488580 318260
rect 489012 318152 489040 320076
rect 488736 318124 489040 318152
rect 488632 317960 488684 317966
rect 488632 317902 488684 317908
rect 488540 312792 488592 312798
rect 488540 312734 488592 312740
rect 488448 278112 488500 278118
rect 488644 278089 488672 317902
rect 488736 301481 488764 318124
rect 489288 318050 489316 320076
rect 488828 318022 489316 318050
rect 488828 312730 488856 318022
rect 489564 317966 489592 320076
rect 489644 318776 489696 318782
rect 489644 318718 489696 318724
rect 489656 317966 489684 318718
rect 489552 317960 489604 317966
rect 489552 317902 489604 317908
rect 489644 317960 489696 317966
rect 489644 317902 489696 317908
rect 489840 316034 489868 320076
rect 489920 318232 489972 318238
rect 489920 318174 489972 318180
rect 488920 316006 489868 316034
rect 488816 312724 488868 312730
rect 488816 312666 488868 312672
rect 488722 301472 488778 301481
rect 488722 301407 488778 301416
rect 488448 278054 488500 278060
rect 488630 278080 488686 278089
rect 488630 278015 488686 278024
rect 488920 274038 488948 316006
rect 488908 274032 488960 274038
rect 488908 273974 488960 273980
rect 487160 268524 487212 268530
rect 487160 268466 487212 268472
rect 489932 268433 489960 318174
rect 490012 318096 490064 318102
rect 490012 318038 490064 318044
rect 490116 318050 490144 320076
rect 490392 318102 490420 320076
rect 490380 318096 490432 318102
rect 490024 272513 490052 318038
rect 490116 318022 490328 318050
rect 490380 318038 490432 318044
rect 490196 317756 490248 317762
rect 490196 317698 490248 317704
rect 490104 317688 490156 317694
rect 490104 317630 490156 317636
rect 490116 273970 490144 317630
rect 490208 275398 490236 317698
rect 490300 307057 490328 318022
rect 490668 317762 490696 320076
rect 490656 317756 490708 317762
rect 490656 317698 490708 317704
rect 490944 317694 490972 320076
rect 491220 318238 491248 320076
rect 491208 318232 491260 318238
rect 491208 318174 491260 318180
rect 491496 318050 491524 320076
rect 491772 318050 491800 320076
rect 491312 318022 491524 318050
rect 491588 318022 491800 318050
rect 490932 317688 490984 317694
rect 490932 317630 490984 317636
rect 491312 314158 491340 318022
rect 491392 317756 491444 317762
rect 491392 317698 491444 317704
rect 491300 314152 491352 314158
rect 491300 314094 491352 314100
rect 490286 307048 490342 307057
rect 490286 306983 490342 306992
rect 490196 275392 490248 275398
rect 490196 275334 490248 275340
rect 490104 273964 490156 273970
rect 490104 273906 490156 273912
rect 490010 272504 490066 272513
rect 490010 272439 490066 272448
rect 489918 268424 489974 268433
rect 491404 268394 491432 317698
rect 491484 317688 491536 317694
rect 491484 317630 491536 317636
rect 491496 269958 491524 317630
rect 491588 270026 491616 318022
rect 492048 317762 492076 320076
rect 492036 317756 492088 317762
rect 492036 317698 492088 317704
rect 492324 317694 492352 320076
rect 492312 317688 492364 317694
rect 492312 317630 492364 317636
rect 492600 316034 492628 320076
rect 492876 318050 492904 320076
rect 493152 318186 493180 320076
rect 491680 316006 492628 316034
rect 492692 318022 492904 318050
rect 492968 318158 493180 318186
rect 491576 270020 491628 270026
rect 491576 269962 491628 269968
rect 491484 269952 491536 269958
rect 491484 269894 491536 269900
rect 491680 268462 491708 316006
rect 492692 312662 492720 318022
rect 492968 317948 492996 318158
rect 492876 317920 492996 317948
rect 492772 317756 492824 317762
rect 492772 317698 492824 317704
rect 492680 312656 492732 312662
rect 492680 312598 492732 312604
rect 492784 271250 492812 317698
rect 492876 276690 492904 317920
rect 493428 317778 493456 320076
rect 492968 317750 493456 317778
rect 492968 294506 492996 317750
rect 493704 316034 493732 320076
rect 493980 317762 494008 320076
rect 494152 318232 494204 318238
rect 494152 318174 494204 318180
rect 494060 318096 494112 318102
rect 494060 318038 494112 318044
rect 493968 317756 494020 317762
rect 493968 317698 494020 317704
rect 493060 316006 493732 316034
rect 492956 294500 493008 294506
rect 492956 294442 493008 294448
rect 492864 276684 492916 276690
rect 492864 276626 492916 276632
rect 492772 271244 492824 271250
rect 492772 271186 492824 271192
rect 493060 269890 493088 316006
rect 494072 271182 494100 318038
rect 494164 272542 494192 318174
rect 494256 318050 494284 320076
rect 494532 318102 494560 320076
rect 494808 318238 494836 320076
rect 494796 318232 494848 318238
rect 494796 318174 494848 318180
rect 494520 318096 494572 318102
rect 494256 318022 494376 318050
rect 494520 318038 494572 318044
rect 494244 316804 494296 316810
rect 494244 316746 494296 316752
rect 494256 279478 494284 316746
rect 494348 283626 494376 318022
rect 495084 316034 495112 320076
rect 495360 316810 495388 320076
rect 495348 316804 495400 316810
rect 495348 316746 495400 316752
rect 494440 316006 495112 316034
rect 494440 311234 494468 316006
rect 495636 311894 495664 320076
rect 495912 314022 495940 320076
rect 496188 314022 496216 320076
rect 495900 314016 495952 314022
rect 495900 313958 495952 313964
rect 496176 314016 496228 314022
rect 496176 313958 496228 313964
rect 495452 311866 495664 311894
rect 496464 311894 496492 320076
rect 496464 311866 496676 311894
rect 494428 311228 494480 311234
rect 494428 311170 494480 311176
rect 495452 309874 495480 311866
rect 495440 309868 495492 309874
rect 495440 309810 495492 309816
rect 496648 307154 496676 311866
rect 496636 307148 496688 307154
rect 496636 307090 496688 307096
rect 494336 283620 494388 283626
rect 494336 283562 494388 283568
rect 494244 279472 494296 279478
rect 494244 279414 494296 279420
rect 494152 272536 494204 272542
rect 494152 272478 494204 272484
rect 496740 271182 496768 320076
rect 497016 311894 497044 320076
rect 497292 318102 497320 320076
rect 497280 318096 497332 318102
rect 497280 318038 497332 318044
rect 497568 315926 497596 320076
rect 497556 315920 497608 315926
rect 497556 315862 497608 315868
rect 497016 311866 497780 311894
rect 497752 271250 497780 311866
rect 497844 308514 497872 320076
rect 498120 316010 498148 320076
rect 498396 318238 498424 320076
rect 498384 318232 498436 318238
rect 498384 318174 498436 318180
rect 497936 315982 498148 316010
rect 498672 315994 498700 320076
rect 498660 315988 498712 315994
rect 497832 308508 497884 308514
rect 497832 308450 497884 308456
rect 497936 273970 497964 315982
rect 498660 315930 498712 315936
rect 498016 315920 498068 315926
rect 498016 315862 498068 315868
rect 497924 273964 497976 273970
rect 497924 273906 497976 273912
rect 498028 272542 498056 315862
rect 498948 312662 498976 320076
rect 498936 312656 498988 312662
rect 498936 312598 498988 312604
rect 499224 311894 499252 320076
rect 499396 315988 499448 315994
rect 499396 315930 499448 315936
rect 499132 311866 499252 311894
rect 498016 272536 498068 272542
rect 498016 272478 498068 272484
rect 497740 271244 497792 271250
rect 497740 271186 497792 271192
rect 494060 271176 494112 271182
rect 494060 271118 494112 271124
rect 496728 271176 496780 271182
rect 496728 271118 496780 271124
rect 493048 269884 493100 269890
rect 493048 269826 493100 269832
rect 491668 268456 491720 268462
rect 491668 268398 491720 268404
rect 499132 268394 499160 311866
rect 499408 272610 499436 315930
rect 499500 312798 499528 320076
rect 499776 314090 499804 320076
rect 500052 315790 500080 320076
rect 500224 319524 500276 319530
rect 500224 319466 500276 319472
rect 500236 318170 500264 319466
rect 500224 318164 500276 318170
rect 500224 318106 500276 318112
rect 500040 315784 500092 315790
rect 500040 315726 500092 315732
rect 499764 314084 499816 314090
rect 499764 314026 499816 314032
rect 499488 312792 499540 312798
rect 499488 312734 499540 312740
rect 500328 311894 500356 320076
rect 500604 315926 500632 320076
rect 500880 316010 500908 320076
rect 500696 315982 500908 316010
rect 500592 315920 500644 315926
rect 500592 315862 500644 315868
rect 500592 315784 500644 315790
rect 500592 315726 500644 315732
rect 500328 311866 500540 311894
rect 499396 272604 499448 272610
rect 499396 272546 499448 272552
rect 500512 268462 500540 311866
rect 500604 311302 500632 315726
rect 500592 311296 500644 311302
rect 500592 311238 500644 311244
rect 500696 278050 500724 315982
rect 500776 315920 500828 315926
rect 500776 315862 500828 315868
rect 500684 278044 500736 278050
rect 500684 277986 500736 277992
rect 500788 269890 500816 315862
rect 501156 312730 501184 320076
rect 501432 315994 501460 320076
rect 501420 315988 501472 315994
rect 501420 315930 501472 315936
rect 501708 315926 501736 320076
rect 501984 316010 502012 320076
rect 502260 316010 502288 320076
rect 501892 315982 502012 316010
rect 502064 315988 502116 315994
rect 501696 315920 501748 315926
rect 501696 315862 501748 315868
rect 501144 312724 501196 312730
rect 501144 312666 501196 312672
rect 501892 311234 501920 315982
rect 502064 315930 502116 315936
rect 502168 315982 502288 316010
rect 501972 312724 502024 312730
rect 501972 312666 502024 312672
rect 501880 311228 501932 311234
rect 501880 311170 501932 311176
rect 501984 309874 502012 312666
rect 501972 309868 502024 309874
rect 501972 309810 502024 309816
rect 502076 308582 502104 315930
rect 502064 308576 502116 308582
rect 502064 308518 502116 308524
rect 502168 271318 502196 315982
rect 502248 315920 502300 315926
rect 502248 315862 502300 315868
rect 502156 271312 502208 271318
rect 502156 271254 502208 271260
rect 502260 270026 502288 315862
rect 502536 312798 502564 320076
rect 502524 312792 502576 312798
rect 502524 312734 502576 312740
rect 502812 311894 502840 320076
rect 503088 318170 503116 320076
rect 503076 318164 503128 318170
rect 503076 318106 503128 318112
rect 503364 311894 503392 320076
rect 503640 311894 503668 320076
rect 502812 311866 503300 311894
rect 503364 311866 503484 311894
rect 502248 270020 502300 270026
rect 502248 269962 502300 269968
rect 500776 269884 500828 269890
rect 500776 269826 500828 269832
rect 503272 268530 503300 311866
rect 503456 309777 503484 311866
rect 503548 311866 503668 311894
rect 503916 311894 503944 320076
rect 508502 319968 508558 319977
rect 508502 319903 508558 319912
rect 503916 311866 505048 311894
rect 503442 309768 503498 309777
rect 503442 309703 503498 309712
rect 503548 300393 503576 311866
rect 503534 300384 503590 300393
rect 503534 300319 503590 300328
rect 505020 269958 505048 311866
rect 508516 295118 508544 319903
rect 509896 300762 509924 354646
rect 510710 348120 510766 348129
rect 510710 348055 510766 348064
rect 510618 342408 510674 342417
rect 510618 342343 510674 342352
rect 510158 327720 510214 327729
rect 510158 327655 510214 327664
rect 510066 324864 510122 324873
rect 510066 324799 510122 324808
rect 509976 320884 510028 320890
rect 509976 320826 510028 320832
rect 509988 318442 510016 320826
rect 510080 320249 510108 324799
rect 510066 320240 510122 320249
rect 510066 320175 510122 320184
rect 509976 318436 510028 318442
rect 509976 318378 510028 318384
rect 509884 300756 509936 300762
rect 509884 300698 509936 300704
rect 508504 295112 508556 295118
rect 508504 295054 508556 295060
rect 510172 292466 510200 327655
rect 510342 327312 510398 327321
rect 510342 327247 510398 327256
rect 510250 326088 510306 326097
rect 510250 326023 510306 326032
rect 510264 300830 510292 326023
rect 510252 300824 510304 300830
rect 510252 300766 510304 300772
rect 510356 300626 510384 327247
rect 510434 326904 510490 326913
rect 510434 326839 510490 326848
rect 510448 320657 510476 326839
rect 510434 320648 510490 320657
rect 510434 320583 510490 320592
rect 510344 300620 510396 300626
rect 510344 300562 510396 300568
rect 510632 298110 510660 342343
rect 510724 303210 510752 348055
rect 510816 315722 510844 360295
rect 510894 345672 510950 345681
rect 510894 345607 510950 345616
rect 510804 315716 510856 315722
rect 510804 315658 510856 315664
rect 510908 303618 510936 345607
rect 511000 320385 511028 361111
rect 511078 355872 511134 355881
rect 511078 355807 511134 355816
rect 511092 320521 511120 355807
rect 511170 337104 511226 337113
rect 511170 337039 511226 337048
rect 511078 320512 511134 320521
rect 511078 320447 511134 320456
rect 510986 320376 511042 320385
rect 510986 320311 511042 320320
rect 511184 305794 511212 337039
rect 511276 318345 511304 465666
rect 512644 423088 512696 423094
rect 512644 423030 512696 423036
rect 512276 378140 512328 378146
rect 512276 378082 512328 378088
rect 512288 377097 512316 378082
rect 512656 377505 512684 423030
rect 512828 423020 512880 423026
rect 512828 422962 512880 422968
rect 512736 422952 512788 422958
rect 512736 422894 512788 422900
rect 512748 378321 512776 422894
rect 512840 383654 512868 422962
rect 512840 383626 512960 383654
rect 512828 379500 512880 379506
rect 512828 379442 512880 379448
rect 512840 378729 512868 379442
rect 512826 378720 512882 378729
rect 512826 378655 512882 378664
rect 512734 378312 512790 378321
rect 512734 378247 512790 378256
rect 512932 377913 512960 383626
rect 512918 377904 512974 377913
rect 512918 377839 512974 377848
rect 512642 377496 512698 377505
rect 512642 377431 512698 377440
rect 512736 377460 512788 377466
rect 512736 377402 512788 377408
rect 512274 377088 512330 377097
rect 512274 377023 512330 377032
rect 512276 375964 512328 375970
rect 512276 375906 512328 375912
rect 512288 375465 512316 375906
rect 512274 375456 512330 375465
rect 512274 375391 512330 375400
rect 512092 375352 512144 375358
rect 512092 375294 512144 375300
rect 512104 375057 512132 375294
rect 512090 375048 512146 375057
rect 512090 374983 512146 374992
rect 512000 373380 512052 373386
rect 512000 373322 512052 373328
rect 512012 373017 512040 373322
rect 511998 373008 512054 373017
rect 511998 372943 512054 372952
rect 512748 372201 512776 377402
rect 513286 376680 513342 376689
rect 513196 376644 513248 376650
rect 513286 376615 513342 376624
rect 513196 376586 513248 376592
rect 513104 376576 513156 376582
rect 513104 376518 513156 376524
rect 513116 375873 513144 376518
rect 513208 376281 513236 376586
rect 513300 376514 513328 376615
rect 513288 376508 513340 376514
rect 513288 376450 513340 376456
rect 513194 376272 513250 376281
rect 513194 376207 513250 376216
rect 513102 375864 513158 375873
rect 513102 375799 513158 375808
rect 513288 375284 513340 375290
rect 513288 375226 513340 375232
rect 512828 375216 512880 375222
rect 512828 375158 512880 375164
rect 512840 374241 512868 375158
rect 513300 374649 513328 375226
rect 513286 374640 513342 374649
rect 513286 374575 513342 374584
rect 512826 374232 512882 374241
rect 512826 374167 512882 374176
rect 513288 373992 513340 373998
rect 513288 373934 513340 373940
rect 513300 373833 513328 373934
rect 513286 373824 513342 373833
rect 513286 373759 513342 373768
rect 513288 373516 513340 373522
rect 513288 373458 513340 373464
rect 513300 373425 513328 373458
rect 513286 373416 513342 373425
rect 513286 373351 513342 373360
rect 513286 372600 513342 372609
rect 513286 372535 513288 372544
rect 513340 372535 513342 372544
rect 513288 372506 513340 372512
rect 513196 372496 513248 372502
rect 513196 372438 513248 372444
rect 512734 372192 512790 372201
rect 512734 372127 512790 372136
rect 512460 371816 512512 371822
rect 512458 371784 512460 371793
rect 512512 371784 512514 371793
rect 512458 371719 512514 371728
rect 513208 371385 513236 372438
rect 513194 371376 513250 371385
rect 513194 371311 513250 371320
rect 513196 371204 513248 371210
rect 513196 371146 513248 371152
rect 513104 371068 513156 371074
rect 513104 371010 513156 371016
rect 513116 370161 513144 371010
rect 513208 370569 513236 371146
rect 513288 371136 513340 371142
rect 513288 371078 513340 371084
rect 513300 370977 513328 371078
rect 513286 370968 513342 370977
rect 513286 370903 513342 370912
rect 513194 370560 513250 370569
rect 513194 370495 513250 370504
rect 513102 370152 513158 370161
rect 513102 370087 513158 370096
rect 513288 369844 513340 369850
rect 513288 369786 513340 369792
rect 513196 369776 513248 369782
rect 513102 369744 513158 369753
rect 513196 369718 513248 369724
rect 513102 369679 513104 369688
rect 513156 369679 513158 369688
rect 513104 369650 513156 369656
rect 513208 368529 513236 369718
rect 513300 369345 513328 369786
rect 513286 369336 513342 369345
rect 513286 369271 513342 369280
rect 513288 369096 513340 369102
rect 513288 369038 513340 369044
rect 513300 368937 513328 369038
rect 513286 368928 513342 368937
rect 513286 368863 513342 368872
rect 513194 368520 513250 368529
rect 512184 368484 512236 368490
rect 513194 368455 513250 368464
rect 512184 368426 512236 368432
rect 512196 368121 512224 368426
rect 512182 368112 512238 368121
rect 512182 368047 512238 368056
rect 512276 367804 512328 367810
rect 512276 367746 512328 367752
rect 512288 367713 512316 367746
rect 512274 367704 512330 367713
rect 512274 367639 512330 367648
rect 513286 367296 513342 367305
rect 513286 367231 513342 367240
rect 513300 367130 513328 367231
rect 513288 367124 513340 367130
rect 513288 367066 513340 367072
rect 513010 366888 513066 366897
rect 513010 366823 513066 366832
rect 512826 366072 512882 366081
rect 512826 366007 512882 366016
rect 512090 364032 512146 364041
rect 512090 363967 512146 363976
rect 512104 363866 512132 363967
rect 512092 363860 512144 363866
rect 512092 363802 512144 363808
rect 512642 362808 512698 362817
rect 512642 362743 512698 362752
rect 512090 361992 512146 362001
rect 512090 361927 512092 361936
rect 512144 361927 512146 361936
rect 512092 361898 512144 361904
rect 512656 361690 512684 362743
rect 512644 361684 512696 361690
rect 512644 361626 512696 361632
rect 512840 360942 512868 366007
rect 513024 365770 513052 366823
rect 513194 366480 513250 366489
rect 513194 366415 513250 366424
rect 513208 366314 513236 366415
rect 513196 366308 513248 366314
rect 513196 366250 513248 366256
rect 513012 365764 513064 365770
rect 513012 365706 513064 365712
rect 512918 365664 512974 365673
rect 512918 365599 512974 365608
rect 512932 364478 512960 365599
rect 513194 365256 513250 365265
rect 513194 365191 513250 365200
rect 513102 364848 513158 364857
rect 513102 364783 513158 364792
rect 512920 364472 512972 364478
rect 512920 364414 512972 364420
rect 513010 363216 513066 363225
rect 513010 363151 513012 363160
rect 513064 363151 513066 363160
rect 513012 363122 513064 363128
rect 512828 360936 512880 360942
rect 512828 360878 512880 360884
rect 513116 360874 513144 364783
rect 513208 362234 513236 365191
rect 513286 364440 513342 364449
rect 513286 364375 513288 364384
rect 513340 364375 513342 364384
rect 513288 364346 513340 364352
rect 513286 363624 513342 363633
rect 513286 363559 513342 363568
rect 513300 362982 513328 363559
rect 513288 362976 513340 362982
rect 513288 362918 513340 362924
rect 513286 362400 513342 362409
rect 513286 362335 513342 362344
rect 513196 362228 513248 362234
rect 513196 362170 513248 362176
rect 513300 361758 513328 362335
rect 513288 361752 513340 361758
rect 513288 361694 513340 361700
rect 513286 361584 513342 361593
rect 513286 361519 513342 361528
rect 513300 361434 513328 361519
rect 513300 361406 513512 361434
rect 513104 360868 513156 360874
rect 513104 360810 513156 360816
rect 513102 360768 513158 360777
rect 513102 360703 513158 360712
rect 513116 360262 513144 360703
rect 513104 360256 513156 360262
rect 513104 360198 513156 360204
rect 513010 359952 513066 359961
rect 513010 359887 513066 359896
rect 513024 358834 513052 359887
rect 513286 359544 513342 359553
rect 513342 359502 513420 359530
rect 513286 359479 513342 359488
rect 513012 358828 513064 358834
rect 513012 358770 513064 358776
rect 511998 358728 512054 358737
rect 511998 358663 512054 358672
rect 511538 335880 511594 335889
rect 511538 335815 511594 335824
rect 511356 320952 511408 320958
rect 511356 320894 511408 320900
rect 511262 318336 511318 318345
rect 511262 318271 511318 318280
rect 511368 317830 511396 320894
rect 511356 317824 511408 317830
rect 511356 317766 511408 317772
rect 511552 305862 511580 335815
rect 511906 326496 511962 326505
rect 511906 326431 511962 326440
rect 511920 322538 511948 326431
rect 511736 322510 511948 322538
rect 511736 319977 511764 322510
rect 511908 322244 511960 322250
rect 511908 322186 511960 322192
rect 511722 319968 511778 319977
rect 511722 319903 511778 319912
rect 511920 318374 511948 322186
rect 511908 318368 511960 318374
rect 511908 318310 511960 318316
rect 511540 305856 511592 305862
rect 511540 305798 511592 305804
rect 511172 305788 511224 305794
rect 511172 305730 511224 305736
rect 510896 303612 510948 303618
rect 510896 303554 510948 303560
rect 510712 303204 510764 303210
rect 510712 303146 510764 303152
rect 512012 302938 512040 358663
rect 513010 358320 513066 358329
rect 513010 358255 513066 358264
rect 513024 358018 513052 358255
rect 513012 358012 513064 358018
rect 513012 357954 513064 357960
rect 512090 357912 512146 357921
rect 512090 357847 512146 357856
rect 512104 357746 512132 357847
rect 512092 357740 512144 357746
rect 512092 357682 512144 357688
rect 513286 357504 513342 357513
rect 513286 357439 513288 357448
rect 513340 357439 513342 357448
rect 513288 357410 513340 357416
rect 512182 357096 512238 357105
rect 512182 357031 512238 357040
rect 512090 356280 512146 356289
rect 512196 356250 512224 357031
rect 512642 356688 512698 356697
rect 512642 356623 512698 356632
rect 512090 356215 512146 356224
rect 512184 356244 512236 356250
rect 512104 303006 512132 356215
rect 512184 356186 512236 356192
rect 512656 356114 512684 356623
rect 512644 356108 512696 356114
rect 512644 356050 512696 356056
rect 512734 355464 512790 355473
rect 512734 355399 512790 355408
rect 512748 355026 512776 355399
rect 513286 355056 513342 355065
rect 512736 355020 512788 355026
rect 513286 354991 513342 355000
rect 512736 354962 512788 354968
rect 513300 354754 513328 354991
rect 513288 354748 513340 354754
rect 513288 354690 513340 354696
rect 513102 354648 513158 354657
rect 513102 354583 513158 354592
rect 512550 354240 512606 354249
rect 512550 354175 512606 354184
rect 512564 354142 512592 354175
rect 512552 354136 512604 354142
rect 512552 354078 512604 354084
rect 512182 353832 512238 353841
rect 512182 353767 512238 353776
rect 512196 352050 512224 353767
rect 513116 353326 513144 354583
rect 513104 353320 513156 353326
rect 513104 353262 513156 353268
rect 513286 352608 513342 352617
rect 513286 352543 513342 352552
rect 512276 352300 512328 352306
rect 512276 352242 512328 352248
rect 512288 352209 512316 352242
rect 512274 352200 512330 352209
rect 512274 352135 512330 352144
rect 512196 352022 512316 352050
rect 512182 349344 512238 349353
rect 512182 349279 512238 349288
rect 512196 349246 512224 349279
rect 512184 349240 512236 349246
rect 512184 349182 512236 349188
rect 512182 346896 512238 346905
rect 512182 346831 512238 346840
rect 512196 346458 512224 346831
rect 512184 346452 512236 346458
rect 512184 346394 512236 346400
rect 512288 345014 512316 352022
rect 513300 351966 513328 352543
rect 513288 351960 513340 351966
rect 513288 351902 513340 351908
rect 512642 351792 512698 351801
rect 512642 351727 512644 351736
rect 512696 351727 512698 351736
rect 512644 351698 512696 351704
rect 513286 351384 513342 351393
rect 513286 351319 513342 351328
rect 513300 351082 513328 351319
rect 513288 351076 513340 351082
rect 513288 351018 513340 351024
rect 512642 350976 512698 350985
rect 512642 350911 512644 350920
rect 512696 350911 512698 350920
rect 512644 350882 512696 350888
rect 513288 350600 513340 350606
rect 513286 350568 513288 350577
rect 513340 350568 513342 350577
rect 513286 350503 513342 350512
rect 512826 350160 512882 350169
rect 512826 350095 512882 350104
rect 512840 349314 512868 350095
rect 513286 349752 513342 349761
rect 513286 349687 513342 349696
rect 513300 349586 513328 349687
rect 513288 349580 513340 349586
rect 513288 349522 513340 349528
rect 512828 349308 512880 349314
rect 512828 349250 512880 349256
rect 513194 348936 513250 348945
rect 513194 348871 513250 348880
rect 513208 347818 513236 348871
rect 513286 348528 513342 348537
rect 513286 348463 513342 348472
rect 513300 348226 513328 348463
rect 513288 348220 513340 348226
rect 513288 348162 513340 348168
rect 513196 347812 513248 347818
rect 513196 347754 513248 347760
rect 513010 347712 513066 347721
rect 513010 347647 513066 347656
rect 512826 347304 512882 347313
rect 512826 347239 512882 347248
rect 512840 346730 512868 347239
rect 512828 346724 512880 346730
rect 512828 346666 512880 346672
rect 513024 346594 513052 347647
rect 513012 346588 513064 346594
rect 513012 346530 513064 346536
rect 512458 346488 512514 346497
rect 512458 346423 512514 346432
rect 512196 344986 512316 345014
rect 512196 315518 512224 344986
rect 512274 344448 512330 344457
rect 512274 344383 512330 344392
rect 512288 344010 512316 344383
rect 512276 344004 512328 344010
rect 512276 343946 512328 343952
rect 512366 343224 512422 343233
rect 512366 343159 512422 343168
rect 512380 342922 512408 343159
rect 512368 342916 512420 342922
rect 512368 342858 512420 342864
rect 512366 342816 512422 342825
rect 512366 342751 512422 342760
rect 512274 342000 512330 342009
rect 512274 341935 512330 341944
rect 512288 341426 512316 341935
rect 512276 341420 512328 341426
rect 512276 341362 512328 341368
rect 512276 341284 512328 341290
rect 512276 341226 512328 341232
rect 512288 341193 512316 341226
rect 512274 341184 512330 341193
rect 512274 341119 512330 341128
rect 512380 341034 512408 342751
rect 512288 341006 512408 341034
rect 512184 315512 512236 315518
rect 512184 315454 512236 315460
rect 512092 303000 512144 303006
rect 512092 302942 512144 302948
rect 512000 302932 512052 302938
rect 512000 302874 512052 302880
rect 510620 298104 510672 298110
rect 510620 298046 510672 298052
rect 512288 296002 512316 341006
rect 512366 340776 512422 340785
rect 512366 340711 512422 340720
rect 512380 339726 512408 340711
rect 512368 339720 512420 339726
rect 512368 339662 512420 339668
rect 512366 339552 512422 339561
rect 512366 339487 512368 339496
rect 512420 339487 512422 339496
rect 512368 339458 512420 339464
rect 512472 335354 512500 346423
rect 513194 346080 513250 346089
rect 513194 346015 513250 346024
rect 513208 345234 513236 346015
rect 513286 345264 513342 345273
rect 513196 345228 513248 345234
rect 513286 345199 513342 345208
rect 513196 345170 513248 345176
rect 513300 345098 513328 345199
rect 513288 345092 513340 345098
rect 513288 345034 513340 345040
rect 513286 344856 513342 344865
rect 513286 344791 513342 344800
rect 513300 344418 513328 344791
rect 513288 344412 513340 344418
rect 513288 344354 513340 344360
rect 512826 344040 512882 344049
rect 512826 343975 512882 343984
rect 512840 343806 512868 343975
rect 512828 343800 512880 343806
rect 512828 343742 512880 343748
rect 513286 343632 513342 343641
rect 513286 343567 513342 343576
rect 513300 342378 513328 343567
rect 513288 342372 513340 342378
rect 513288 342314 513340 342320
rect 513286 341592 513342 341601
rect 513286 341527 513342 341536
rect 513300 340950 513328 341527
rect 513288 340944 513340 340950
rect 513288 340886 513340 340892
rect 513010 340368 513066 340377
rect 513010 340303 513066 340312
rect 513024 339794 513052 340303
rect 513286 339960 513342 339969
rect 513286 339895 513288 339904
rect 513340 339895 513342 339904
rect 513288 339866 513340 339872
rect 513012 339788 513064 339794
rect 513012 339730 513064 339736
rect 513286 339144 513342 339153
rect 513286 339079 513342 339088
rect 513194 338736 513250 338745
rect 513194 338671 513250 338680
rect 513208 338434 513236 338671
rect 513196 338428 513248 338434
rect 513196 338370 513248 338376
rect 512550 338328 512606 338337
rect 512550 338263 512552 338272
rect 512604 338263 512606 338272
rect 512552 338234 512604 338240
rect 513300 338162 513328 339079
rect 513288 338156 513340 338162
rect 513288 338098 513340 338104
rect 513010 337920 513066 337929
rect 513010 337855 513066 337864
rect 512918 337512 512974 337521
rect 512918 337447 512974 337456
rect 512932 337074 512960 337447
rect 512920 337068 512972 337074
rect 512920 337010 512972 337016
rect 513024 336802 513052 337855
rect 513012 336796 513064 336802
rect 513012 336738 513064 336744
rect 513286 336696 513342 336705
rect 513286 336631 513342 336640
rect 513194 336288 513250 336297
rect 513194 336223 513250 336232
rect 513208 335986 513236 336223
rect 513196 335980 513248 335986
rect 513196 335922 513248 335928
rect 513300 335714 513328 336631
rect 513288 335708 513340 335714
rect 513288 335650 513340 335656
rect 512734 335472 512790 335481
rect 512734 335407 512736 335416
rect 512788 335407 512790 335416
rect 512736 335378 512788 335384
rect 512380 335326 512500 335354
rect 512380 305658 512408 335326
rect 512826 335064 512882 335073
rect 512826 334999 512882 335008
rect 512642 334248 512698 334257
rect 512642 334183 512698 334192
rect 512458 330576 512514 330585
rect 512458 330511 512514 330520
rect 512368 305652 512420 305658
rect 512368 305594 512420 305600
rect 512472 304298 512500 330511
rect 512550 329760 512606 329769
rect 512550 329695 512606 329704
rect 512564 329050 512592 329695
rect 512552 329044 512604 329050
rect 512552 328986 512604 328992
rect 512550 328944 512606 328953
rect 512550 328879 512606 328888
rect 512564 328778 512592 328879
rect 512552 328772 512604 328778
rect 512552 328714 512604 328720
rect 512656 325694 512684 334183
rect 512840 334082 512868 334999
rect 513010 334656 513066 334665
rect 513010 334591 513066 334600
rect 513024 334218 513052 334591
rect 513012 334212 513064 334218
rect 513012 334154 513064 334160
rect 512828 334076 512880 334082
rect 512828 334018 512880 334024
rect 512918 333840 512974 333849
rect 512918 333775 512974 333784
rect 512826 333024 512882 333033
rect 512826 332959 512882 332968
rect 512840 332654 512868 332959
rect 512932 332858 512960 333775
rect 512920 332852 512972 332858
rect 512920 332794 512972 332800
rect 513288 332784 513340 332790
rect 513288 332726 513340 332732
rect 512828 332648 512880 332654
rect 513300 332625 513328 332726
rect 512828 332590 512880 332596
rect 513286 332616 513342 332625
rect 513286 332551 513342 332560
rect 512826 332208 512882 332217
rect 512826 332143 512882 332152
rect 512734 331800 512790 331809
rect 512734 331735 512790 331744
rect 512564 325666 512684 325694
rect 512564 315586 512592 325666
rect 512642 325544 512698 325553
rect 512642 325479 512698 325488
rect 512552 315580 512604 315586
rect 512552 315522 512604 315528
rect 512656 305726 512684 325479
rect 512748 315654 512776 331735
rect 512840 331294 512868 332143
rect 513288 331492 513340 331498
rect 513288 331434 513340 331440
rect 513300 331401 513328 331434
rect 513286 331392 513342 331401
rect 513286 331327 513342 331336
rect 512828 331288 512880 331294
rect 512828 331230 512880 331236
rect 513286 329352 513342 329361
rect 513286 329287 513342 329296
rect 513300 328506 513328 329287
rect 513288 328500 513340 328506
rect 513288 328442 513340 328448
rect 513286 328128 513342 328137
rect 513286 328063 513342 328072
rect 513300 327418 513328 328063
rect 513288 327412 513340 327418
rect 513288 327354 513340 327360
rect 512826 322824 512882 322833
rect 512826 322759 512882 322768
rect 512736 315648 512788 315654
rect 512736 315590 512788 315596
rect 512644 305720 512696 305726
rect 512644 305662 512696 305668
rect 512460 304292 512512 304298
rect 512460 304234 512512 304240
rect 512276 295996 512328 296002
rect 512276 295938 512328 295944
rect 510160 292460 510212 292466
rect 510160 292402 510212 292408
rect 512840 275330 512868 322759
rect 513392 295254 513420 359502
rect 513484 354674 513512 361406
rect 513484 354646 513696 354674
rect 513470 353424 513526 353433
rect 513470 353359 513526 353368
rect 513484 295322 513512 353359
rect 513562 353016 513618 353025
rect 513562 352951 513618 352960
rect 513576 300558 513604 352951
rect 513668 315450 513696 354646
rect 513748 346452 513800 346458
rect 513748 346394 513800 346400
rect 513656 315444 513708 315450
rect 513656 315386 513708 315392
rect 513760 303278 513788 346394
rect 513840 341420 513892 341426
rect 513840 341362 513892 341368
rect 513852 303346 513880 341362
rect 513932 328772 513984 328778
rect 513932 328714 513984 328720
rect 513840 303340 513892 303346
rect 513840 303282 513892 303288
rect 513748 303272 513800 303278
rect 513748 303214 513800 303220
rect 513564 300552 513616 300558
rect 513564 300494 513616 300500
rect 513472 295316 513524 295322
rect 513472 295258 513524 295264
rect 513380 295248 513432 295254
rect 513380 295190 513432 295196
rect 513944 292126 513972 328714
rect 514036 319666 514064 470562
rect 514116 381540 514168 381546
rect 514116 381482 514168 381488
rect 514128 373386 514156 381482
rect 514116 373380 514168 373386
rect 514116 373322 514168 373328
rect 514760 363860 514812 363866
rect 514760 363802 514812 363808
rect 514772 359922 514800 363802
rect 514852 363180 514904 363186
rect 514852 363122 514904 363128
rect 514760 359916 514812 359922
rect 514760 359858 514812 359864
rect 514864 358698 514892 363122
rect 514944 361956 514996 361962
rect 514944 361898 514996 361904
rect 514852 358692 514904 358698
rect 514852 358634 514904 358640
rect 514956 358578 514984 361898
rect 514772 358550 514984 358578
rect 514116 339516 514168 339522
rect 514116 339458 514168 339464
rect 514024 319660 514076 319666
rect 514024 319602 514076 319608
rect 514128 303550 514156 339458
rect 514208 329044 514260 329050
rect 514208 328986 514260 328992
rect 514116 303544 514168 303550
rect 514116 303486 514168 303492
rect 514220 300354 514248 328986
rect 514208 300348 514260 300354
rect 514208 300290 514260 300296
rect 514772 292534 514800 358550
rect 514944 357740 514996 357746
rect 514944 357682 514996 357688
rect 514852 356244 514904 356250
rect 514852 356186 514904 356192
rect 514864 294982 514892 356186
rect 514956 304502 514984 357682
rect 515036 349240 515088 349246
rect 515036 349182 515088 349188
rect 514944 304496 514996 304502
rect 514944 304438 514996 304444
rect 515048 300694 515076 349182
rect 515128 344004 515180 344010
rect 515128 343946 515180 343952
rect 515140 303142 515168 343946
rect 515220 342916 515272 342922
rect 515220 342858 515272 342864
rect 515128 303136 515180 303142
rect 515128 303078 515180 303084
rect 515232 303074 515260 342858
rect 515312 339720 515364 339726
rect 515312 339662 515364 339668
rect 515324 303482 515352 339662
rect 515416 317966 515444 599558
rect 515496 563100 515548 563106
rect 515496 563042 515548 563048
rect 515404 317960 515456 317966
rect 515404 317902 515456 317908
rect 515508 317150 515536 563042
rect 516782 467256 516838 467265
rect 516782 467191 516838 467200
rect 515588 421932 515640 421938
rect 515588 421874 515640 421880
rect 515600 367810 515628 421874
rect 515680 385688 515732 385694
rect 515680 385630 515732 385636
rect 515692 375970 515720 385630
rect 515772 380180 515824 380186
rect 515772 380122 515824 380128
rect 515680 375964 515732 375970
rect 515680 375906 515732 375912
rect 515784 371822 515812 380122
rect 515772 371816 515824 371822
rect 515772 371758 515824 371764
rect 515588 367804 515640 367810
rect 515588 367746 515640 367752
rect 516232 356108 516284 356114
rect 516232 356050 516284 356056
rect 515588 338292 515640 338298
rect 515588 338234 515640 338240
rect 515496 317144 515548 317150
rect 515496 317086 515548 317092
rect 515312 303476 515364 303482
rect 515312 303418 515364 303424
rect 515600 303414 515628 338234
rect 516140 335436 516192 335442
rect 516140 335378 516192 335384
rect 516152 315314 516180 335378
rect 516140 315308 516192 315314
rect 516140 315250 516192 315256
rect 516244 304366 516272 356050
rect 516324 351756 516376 351762
rect 516324 351698 516376 351704
rect 516232 304360 516284 304366
rect 516232 304302 516284 304308
rect 515588 303408 515640 303414
rect 515588 303350 515640 303356
rect 515220 303068 515272 303074
rect 515220 303010 515272 303016
rect 515036 300688 515088 300694
rect 515036 300630 515088 300636
rect 516336 300422 516364 351698
rect 516600 337068 516652 337074
rect 516600 337010 516652 337016
rect 516416 334076 516468 334082
rect 516416 334018 516468 334024
rect 516324 300416 516376 300422
rect 516324 300358 516376 300364
rect 514852 294976 514904 294982
rect 514852 294918 514904 294924
rect 514760 292528 514812 292534
rect 514760 292470 514812 292476
rect 516428 292398 516456 334018
rect 516508 332852 516560 332858
rect 516508 332794 516560 332800
rect 516416 292392 516468 292398
rect 516416 292334 516468 292340
rect 516520 292330 516548 332794
rect 516612 298042 516640 337010
rect 516692 334212 516744 334218
rect 516692 334154 516744 334160
rect 516600 298036 516652 298042
rect 516600 297978 516652 297984
rect 516704 297974 516732 334154
rect 516796 318578 516824 467191
rect 517520 373312 517572 373318
rect 517520 373254 517572 373260
rect 517532 372570 517560 373254
rect 517520 372564 517572 372570
rect 517520 372506 517572 372512
rect 517520 361684 517572 361690
rect 517520 361626 517572 361632
rect 517532 360126 517560 361626
rect 517520 360120 517572 360126
rect 517520 360062 517572 360068
rect 517520 355020 517572 355026
rect 517520 354962 517572 354968
rect 516968 350940 517020 350946
rect 516968 350882 517020 350888
rect 516876 331288 516928 331294
rect 516876 331230 516928 331236
rect 516784 318572 516836 318578
rect 516784 318514 516836 318520
rect 516888 300150 516916 331230
rect 516876 300144 516928 300150
rect 516876 300086 516928 300092
rect 516692 297968 516744 297974
rect 516692 297910 516744 297916
rect 516980 295050 517008 350882
rect 517532 300218 517560 354962
rect 517612 354136 517664 354142
rect 517612 354078 517664 354084
rect 517624 300286 517652 354078
rect 517704 350600 517756 350606
rect 517704 350542 517756 350548
rect 517716 300490 517744 350542
rect 517796 339924 517848 339930
rect 517796 339866 517848 339872
rect 517704 300484 517756 300490
rect 517704 300426 517756 300432
rect 517612 300280 517664 300286
rect 517612 300222 517664 300228
rect 517520 300212 517572 300218
rect 517520 300154 517572 300160
rect 517808 297770 517836 339866
rect 518072 339788 518124 339794
rect 518072 339730 518124 339736
rect 517888 338428 517940 338434
rect 517888 338370 517940 338376
rect 517900 297838 517928 338370
rect 517980 335980 518032 335986
rect 517980 335922 518032 335928
rect 517992 297906 518020 335922
rect 518084 312594 518112 339730
rect 518176 318034 518204 599626
rect 518256 576904 518308 576910
rect 518256 576846 518308 576852
rect 518268 319802 518296 576846
rect 518348 536852 518400 536858
rect 518348 536794 518400 536800
rect 518256 319796 518308 319802
rect 518256 319738 518308 319744
rect 518360 318306 518388 536794
rect 523696 516769 523724 600086
rect 531332 600086 532082 600114
rect 531332 520946 531360 600086
rect 540532 598262 540560 600100
rect 543752 599690 543780 700266
rect 559668 699825 559696 703520
rect 559654 699816 559710 699825
rect 559654 699751 559710 699760
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 579632 683194 579660 683839
rect 570604 683188 570656 683194
rect 570604 683130 570656 683136
rect 579620 683188 579672 683194
rect 579620 683130 579672 683136
rect 543740 599684 543792 599690
rect 543740 599626 543792 599632
rect 540520 598256 540572 598262
rect 540520 598198 540572 598204
rect 531320 520940 531372 520946
rect 531320 520882 531372 520888
rect 523682 516760 523738 516769
rect 523682 516695 523738 516704
rect 550638 516760 550694 516769
rect 550638 516695 550694 516704
rect 547880 514072 547932 514078
rect 547880 514014 547932 514020
rect 543740 512712 543792 512718
rect 543740 512654 543792 512660
rect 538220 512644 538272 512650
rect 538220 512586 538272 512592
rect 519544 510672 519596 510678
rect 519544 510614 519596 510620
rect 518440 423156 518492 423162
rect 518440 423098 518492 423104
rect 518452 369714 518480 423098
rect 518532 420232 518584 420238
rect 518532 420174 518584 420180
rect 518544 373522 518572 420174
rect 518532 373516 518584 373522
rect 518532 373458 518584 373464
rect 518440 369708 518492 369714
rect 518440 369650 518492 369656
rect 518900 366308 518952 366314
rect 518900 366250 518952 366256
rect 518912 358494 518940 366250
rect 518900 358488 518952 358494
rect 518900 358430 518952 358436
rect 518900 353320 518952 353326
rect 518900 353262 518952 353268
rect 518348 318300 518400 318306
rect 518348 318242 518400 318248
rect 518164 318028 518216 318034
rect 518164 317970 518216 317976
rect 518072 312588 518124 312594
rect 518072 312530 518124 312536
rect 517980 297900 518032 297906
rect 517980 297842 518032 297848
rect 517888 297832 517940 297838
rect 517888 297774 517940 297780
rect 517796 297764 517848 297770
rect 517796 297706 517848 297712
rect 516968 295044 517020 295050
rect 516968 294986 517020 294992
rect 518912 294778 518940 353262
rect 518992 349580 519044 349586
rect 518992 349522 519044 349528
rect 519004 294914 519032 349522
rect 519084 346724 519136 346730
rect 519084 346666 519136 346672
rect 519096 297634 519124 346666
rect 519176 345228 519228 345234
rect 519176 345170 519228 345176
rect 519084 297628 519136 297634
rect 519084 297570 519136 297576
rect 519188 297566 519216 345170
rect 519268 342372 519320 342378
rect 519268 342314 519320 342320
rect 519280 297702 519308 342314
rect 519452 341284 519504 341290
rect 519452 341226 519504 341232
rect 519360 335708 519412 335714
rect 519360 335650 519412 335656
rect 519268 297696 519320 297702
rect 519268 297638 519320 297644
rect 519176 297560 519228 297566
rect 519176 297502 519228 297508
rect 518992 294908 519044 294914
rect 518992 294850 519044 294856
rect 518900 294772 518952 294778
rect 518900 294714 518952 294720
rect 516508 292324 516560 292330
rect 516508 292266 516560 292272
rect 519372 292194 519400 335650
rect 519464 297498 519492 341226
rect 519556 317218 519584 510614
rect 534080 508564 534132 508570
rect 534080 508506 534132 508512
rect 531320 505164 531372 505170
rect 531320 505106 531372 505112
rect 521750 467120 521806 467129
rect 521750 467055 521806 467064
rect 521764 464916 521792 467055
rect 528376 466540 528428 466546
rect 528376 466482 528428 466488
rect 525064 466472 525116 466478
rect 525064 466414 525116 466420
rect 525076 464916 525104 466414
rect 528388 464916 528416 466482
rect 531332 464930 531360 505106
rect 534092 480254 534120 508506
rect 534092 480226 534672 480254
rect 534644 464930 534672 480226
rect 538232 464930 538260 512586
rect 540980 509924 541032 509930
rect 540980 509866 541032 509872
rect 540992 480254 541020 509866
rect 543752 480254 543780 512654
rect 540992 480226 541296 480254
rect 543752 480226 544608 480254
rect 541268 464930 541296 480226
rect 544580 464930 544608 480226
rect 547892 464930 547920 514014
rect 550652 480254 550680 516695
rect 550652 480226 551232 480254
rect 551204 464930 551232 480226
rect 554872 465180 554924 465186
rect 554872 465122 554924 465128
rect 531332 464902 531714 464930
rect 534644 464902 535026 464930
rect 538232 464902 538338 464930
rect 541268 464902 541650 464930
rect 544580 464902 544962 464930
rect 547892 464902 548274 464930
rect 551204 464902 551586 464930
rect 554884 464916 554912 465122
rect 558184 465112 558236 465118
rect 558184 465054 558236 465060
rect 558196 464916 558224 465054
rect 561678 444952 561734 444961
rect 561678 444887 561734 444896
rect 519636 422408 519688 422414
rect 519636 422350 519688 422356
rect 519648 369102 519676 422350
rect 520844 421938 520872 425068
rect 521948 425054 522330 425082
rect 523420 425054 523802 425082
rect 520832 421932 520884 421938
rect 520832 421874 520884 421880
rect 521948 412634 521976 425054
rect 522396 422816 522448 422822
rect 522396 422758 522448 422764
rect 521672 412606 521976 412634
rect 519728 384328 519780 384334
rect 519728 384270 519780 384276
rect 519740 373998 519768 384270
rect 519728 373992 519780 373998
rect 519728 373934 519780 373940
rect 519636 369096 519688 369102
rect 519636 369038 519688 369044
rect 521672 368490 521700 412606
rect 522304 411936 522356 411942
rect 522304 411878 522356 411884
rect 521660 368484 521712 368490
rect 521660 368426 521712 368432
rect 520280 360256 520332 360262
rect 520280 360198 520332 360204
rect 519636 332784 519688 332790
rect 519636 332726 519688 332732
rect 519544 317212 519596 317218
rect 519544 317154 519596 317160
rect 519452 297492 519504 297498
rect 519452 297434 519504 297440
rect 519360 292188 519412 292194
rect 519360 292130 519412 292136
rect 513932 292120 513984 292126
rect 513932 292062 513984 292068
rect 519648 291922 519676 332726
rect 519728 331492 519780 331498
rect 519728 331434 519780 331440
rect 519636 291916 519688 291922
rect 519636 291858 519688 291864
rect 519740 291854 519768 331434
rect 520292 295186 520320 360198
rect 520372 358012 520424 358018
rect 520372 357954 520424 357960
rect 520280 295180 520332 295186
rect 520280 295122 520332 295128
rect 520384 294710 520412 357954
rect 520648 352300 520700 352306
rect 520648 352242 520700 352248
rect 520464 351076 520516 351082
rect 520464 351018 520516 351024
rect 520372 294704 520424 294710
rect 520372 294646 520424 294652
rect 519728 291848 519780 291854
rect 519728 291790 519780 291796
rect 520476 289610 520504 351018
rect 520556 349308 520608 349314
rect 520556 349250 520608 349256
rect 520464 289604 520516 289610
rect 520464 289546 520516 289552
rect 520568 289542 520596 349250
rect 520660 294642 520688 352242
rect 520740 348220 520792 348226
rect 520740 348162 520792 348168
rect 520752 294846 520780 348162
rect 521660 347812 521712 347818
rect 521660 347754 521712 347760
rect 520832 344412 520884 344418
rect 520832 344354 520884 344360
rect 520844 297430 520872 344354
rect 520924 327412 520976 327418
rect 520924 327354 520976 327360
rect 520832 297424 520884 297430
rect 520832 297366 520884 297372
rect 520740 294840 520792 294846
rect 520740 294782 520792 294788
rect 520648 294636 520700 294642
rect 520648 294578 520700 294584
rect 520556 289536 520608 289542
rect 520556 289478 520608 289484
rect 520936 289066 520964 327354
rect 521672 289338 521700 347754
rect 521752 346588 521804 346594
rect 521752 346530 521804 346536
rect 521660 289332 521712 289338
rect 521660 289274 521712 289280
rect 521764 289202 521792 346530
rect 521844 345092 521896 345098
rect 521844 345034 521896 345040
rect 521856 289270 521884 345034
rect 521936 343800 521988 343806
rect 521936 343742 521988 343748
rect 521844 289264 521896 289270
rect 521844 289206 521896 289212
rect 521752 289196 521804 289202
rect 521752 289138 521804 289144
rect 521948 289134 521976 343742
rect 522028 340944 522080 340950
rect 522028 340886 522080 340892
rect 522040 292262 522068 340886
rect 522120 338156 522172 338162
rect 522120 338098 522172 338104
rect 522028 292256 522080 292262
rect 522028 292198 522080 292204
rect 522132 291990 522160 338098
rect 522212 336796 522264 336802
rect 522212 336738 522264 336744
rect 522224 292058 522252 336738
rect 522316 318510 522344 411878
rect 522408 371074 522436 422758
rect 523420 412634 523448 425054
rect 523684 423224 523736 423230
rect 523684 423166 523736 423172
rect 523052 412606 523448 412634
rect 522396 371068 522448 371074
rect 522396 371010 522448 371016
rect 523052 369782 523080 412606
rect 523696 371142 523724 423166
rect 525260 422414 525288 425068
rect 526364 425054 526746 425082
rect 525248 422408 525300 422414
rect 525248 422350 525300 422356
rect 526364 412634 526392 425054
rect 528204 423162 528232 425068
rect 528192 423156 528244 423162
rect 528192 423098 528244 423104
rect 529676 422822 529704 425068
rect 530780 425054 531162 425082
rect 529664 422816 529716 422822
rect 529664 422758 529716 422764
rect 530780 412634 530808 425054
rect 532620 423230 532648 425068
rect 533344 423292 533396 423298
rect 533344 423234 533396 423240
rect 532608 423224 532660 423230
rect 532608 423166 532660 423172
rect 525812 412606 526392 412634
rect 529952 412606 530808 412634
rect 523684 371136 523736 371142
rect 523684 371078 523736 371084
rect 525812 369850 525840 412606
rect 529952 371210 529980 412606
rect 533356 375222 533384 423234
rect 533344 375216 533396 375222
rect 533344 375158 533396 375164
rect 534092 372570 534120 425068
rect 535472 425054 535578 425082
rect 536852 425054 537050 425082
rect 538232 425054 538522 425082
rect 539612 425054 539994 425082
rect 535472 380186 535500 425054
rect 536104 423428 536156 423434
rect 536104 423370 536156 423376
rect 535460 380180 535512 380186
rect 535460 380122 535512 380128
rect 536116 375290 536144 423370
rect 536852 377466 536880 425054
rect 537484 423360 537536 423366
rect 537484 423302 537536 423308
rect 536840 377460 536892 377466
rect 536840 377402 536892 377408
rect 537496 375358 537524 423302
rect 537484 375352 537536 375358
rect 537484 375294 537536 375300
rect 536104 375284 536156 375290
rect 536104 375226 536156 375232
rect 538232 373318 538260 425054
rect 538864 423156 538916 423162
rect 538864 423098 538916 423104
rect 538876 376582 538904 423098
rect 539612 381546 539640 425054
rect 540244 423224 540296 423230
rect 540244 423166 540296 423172
rect 539600 381540 539652 381546
rect 539600 381482 539652 381488
rect 540256 376650 540284 423166
rect 541452 420238 541480 425068
rect 542556 425054 542938 425082
rect 541440 420232 541492 420238
rect 541440 420174 541492 420180
rect 542556 412634 542584 425054
rect 544396 423298 544424 425068
rect 545868 423434 545896 425068
rect 545856 423428 545908 423434
rect 545856 423370 545908 423376
rect 547340 423366 547368 425068
rect 548444 425054 548826 425082
rect 547328 423360 547380 423366
rect 547328 423302 547380 423308
rect 544384 423292 544436 423298
rect 544384 423234 544436 423240
rect 544476 423292 544528 423298
rect 544476 423234 544528 423240
rect 544488 412634 544516 423234
rect 547144 421592 547196 421598
rect 547144 421534 547196 421540
rect 542372 412606 542584 412634
rect 544396 412606 544516 412634
rect 542372 384334 542400 412606
rect 542360 384328 542412 384334
rect 542360 384270 542412 384276
rect 543004 380180 543056 380186
rect 543004 380122 543056 380128
rect 543016 379506 543044 380122
rect 543004 379500 543056 379506
rect 543004 379442 543056 379448
rect 540244 376644 540296 376650
rect 540244 376586 540296 376592
rect 538864 376576 538916 376582
rect 538864 376518 538916 376524
rect 544396 376514 544424 412606
rect 547156 378146 547184 421534
rect 548444 412634 548472 425054
rect 550284 423162 550312 425068
rect 551756 423230 551784 425068
rect 553228 423298 553256 425068
rect 553216 423292 553268 423298
rect 553216 423234 553268 423240
rect 551744 423224 551796 423230
rect 551744 423166 551796 423172
rect 550272 423156 550324 423162
rect 550272 423098 550324 423104
rect 554700 421598 554728 425068
rect 556172 423094 556200 425068
rect 556160 423088 556212 423094
rect 556160 423030 556212 423036
rect 557644 423026 557672 425068
rect 557632 423020 557684 423026
rect 557632 422962 557684 422968
rect 559116 422958 559144 425068
rect 559104 422952 559156 422958
rect 559104 422894 559156 422900
rect 554688 421592 554740 421598
rect 554688 421534 554740 421540
rect 547892 412606 548472 412634
rect 547892 385694 547920 412606
rect 547880 385688 547932 385694
rect 547880 385630 547932 385636
rect 554964 382968 555016 382974
rect 554964 382910 555016 382916
rect 554976 379916 555004 382910
rect 561692 380186 561720 444887
rect 561680 380180 561732 380186
rect 561680 380122 561732 380128
rect 564532 379568 564584 379574
rect 564584 379516 564926 379522
rect 564532 379510 564926 379516
rect 564544 379494 564926 379510
rect 547144 378140 547196 378146
rect 547144 378082 547196 378088
rect 544384 376508 544436 376514
rect 544384 376450 544436 376456
rect 538220 373312 538272 373318
rect 538220 373254 538272 373260
rect 534080 372564 534132 372570
rect 534080 372506 534132 372512
rect 529940 371204 529992 371210
rect 529940 371146 529992 371152
rect 525800 369844 525852 369850
rect 525800 369786 525852 369792
rect 523040 369776 523092 369782
rect 523040 369718 523092 369724
rect 547144 367124 547196 367130
rect 547144 367066 547196 367072
rect 523040 361752 523092 361758
rect 523040 361694 523092 361700
rect 522304 318504 522356 318510
rect 522304 318446 522356 318452
rect 522212 292052 522264 292058
rect 522212 291994 522264 292000
rect 522120 291984 522172 291990
rect 522120 291926 522172 291932
rect 523052 289814 523080 361694
rect 547156 360058 547184 367066
rect 547972 365764 548024 365770
rect 547972 365706 548024 365712
rect 547144 360052 547196 360058
rect 547144 359994 547196 360000
rect 547984 359854 548012 365706
rect 548064 364472 548116 364478
rect 548064 364414 548116 364420
rect 547972 359848 548024 359854
rect 547972 359790 548024 359796
rect 523132 358828 523184 358834
rect 523132 358770 523184 358776
rect 523040 289808 523092 289814
rect 523040 289750 523092 289756
rect 523144 289746 523172 358770
rect 548076 358630 548104 364414
rect 549352 364404 549404 364410
rect 549352 364346 549404 364352
rect 549168 362228 549220 362234
rect 549168 362170 549220 362176
rect 548064 358624 548116 358630
rect 548064 358566 548116 358572
rect 549180 358562 549208 362170
rect 549364 360194 549392 364346
rect 550548 362976 550600 362982
rect 550548 362918 550600 362924
rect 549352 360188 549404 360194
rect 549352 360130 549404 360136
rect 550560 359990 550588 362918
rect 550732 360936 550784 360942
rect 550732 360878 550784 360884
rect 550744 360670 550772 360878
rect 551928 360732 551980 360738
rect 551928 360674 551980 360680
rect 550732 360664 550784 360670
rect 550732 360606 550784 360612
rect 551468 360664 551520 360670
rect 551468 360606 551520 360612
rect 550640 360120 550692 360126
rect 550692 360068 550850 360074
rect 550640 360062 550850 360068
rect 550652 360046 550850 360062
rect 550548 359984 550600 359990
rect 550548 359926 550600 359932
rect 549168 358556 549220 358562
rect 549168 358498 549220 358504
rect 551480 358426 551508 360606
rect 551940 358766 551968 360674
rect 557184 360194 557474 360210
rect 557172 360188 557474 360194
rect 557224 360182 557474 360188
rect 557172 360130 557224 360136
rect 551928 358760 551980 358766
rect 551928 358702 551980 358708
rect 552492 358698 552520 360060
rect 553872 360046 554162 360074
rect 553872 359990 553900 360046
rect 553860 359984 553912 359990
rect 553860 359926 553912 359932
rect 555804 359922 555832 360060
rect 555792 359916 555844 359922
rect 555792 359858 555844 359864
rect 559116 358766 559144 360060
rect 559104 358760 559156 358766
rect 559104 358702 559156 358708
rect 552480 358692 552532 358698
rect 552480 358634 552532 358640
rect 560772 358562 560800 360060
rect 562428 358630 562456 360060
rect 562416 358624 562468 358630
rect 562416 358566 562468 358572
rect 560760 358556 560812 358562
rect 560760 358498 560812 358504
rect 564084 358426 564112 360060
rect 565740 358494 565768 360060
rect 567396 359854 567424 360060
rect 568776 360058 569066 360074
rect 568764 360052 569066 360058
rect 568816 360046 569066 360052
rect 568764 359994 568816 360000
rect 567384 359848 567436 359854
rect 567384 359790 567436 359796
rect 565728 358488 565780 358494
rect 565728 358430 565780 358436
rect 551468 358420 551520 358426
rect 551468 358362 551520 358368
rect 564072 358420 564124 358426
rect 564072 358362 564124 358368
rect 523224 357468 523276 357474
rect 523224 357410 523276 357416
rect 523132 289740 523184 289746
rect 523132 289682 523184 289688
rect 523236 289678 523264 357410
rect 523316 354748 523368 354754
rect 523316 354690 523368 354696
rect 523224 289672 523276 289678
rect 523224 289614 523276 289620
rect 523328 289406 523356 354690
rect 523408 351960 523460 351966
rect 523408 351902 523460 351908
rect 523420 289474 523448 351902
rect 523500 332648 523552 332654
rect 523500 332590 523552 332596
rect 523408 289468 523460 289474
rect 523408 289410 523460 289416
rect 523316 289400 523368 289406
rect 523316 289342 523368 289348
rect 521936 289128 521988 289134
rect 521936 289070 521988 289076
rect 520924 289060 520976 289066
rect 520924 289002 520976 289008
rect 523512 286346 523540 332590
rect 523592 328500 523644 328506
rect 523592 328442 523644 328448
rect 523604 286414 523632 328442
rect 570616 319938 570644 683130
rect 573364 670744 573416 670750
rect 580172 670744 580224 670750
rect 573364 670686 573416 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 571984 616888 572036 616894
rect 571984 616830 572036 616836
rect 570696 456816 570748 456822
rect 570696 456758 570748 456764
rect 570604 319932 570656 319938
rect 570604 319874 570656 319880
rect 543004 318232 543056 318238
rect 543004 318174 543056 318180
rect 538864 315376 538916 315382
rect 538864 315318 538916 315324
rect 529940 307216 529992 307222
rect 529940 307158 529992 307164
rect 523592 286408 523644 286414
rect 523592 286350 523644 286356
rect 523500 286340 523552 286346
rect 523500 286282 523552 286288
rect 512828 275324 512880 275330
rect 512828 275266 512880 275272
rect 505008 269952 505060 269958
rect 505008 269894 505060 269900
rect 503260 268524 503312 268530
rect 503260 268466 503312 268472
rect 500500 268456 500552 268462
rect 500500 268398 500552 268404
rect 489918 268359 489974 268368
rect 491392 268388 491444 268394
rect 491392 268330 491444 268336
rect 499120 268388 499172 268394
rect 499120 268330 499172 268336
rect 529952 209273 529980 307158
rect 531412 304564 531464 304570
rect 531412 304506 531464 304512
rect 531320 293344 531372 293350
rect 531320 293286 531372 293292
rect 530032 278112 530084 278118
rect 530032 278054 530084 278060
rect 530044 244225 530072 278054
rect 530030 244216 530086 244225
rect 530030 244151 530086 244160
rect 531332 226273 531360 293286
rect 531424 261089 531452 304506
rect 536104 301504 536156 301510
rect 536104 301446 536156 301452
rect 533344 297356 533396 297362
rect 533344 297298 533396 297304
rect 531410 261080 531466 261089
rect 531410 261015 531466 261024
rect 531318 226264 531374 226273
rect 531318 226199 531374 226208
rect 529938 209264 529994 209273
rect 529938 209199 529994 209208
rect 533356 206990 533384 297298
rect 533344 206984 533396 206990
rect 533344 206926 533396 206932
rect 532700 174548 532752 174554
rect 532700 174490 532752 174496
rect 532712 171134 532740 174490
rect 532712 171106 533016 171134
rect 482376 168020 482428 168026
rect 482376 167962 482428 167968
rect 469864 164960 469916 164966
rect 469864 164902 469916 164908
rect 460756 138916 460808 138922
rect 460756 138858 460808 138864
rect 460664 132932 460716 132938
rect 460664 132874 460716 132880
rect 460572 128240 460624 128246
rect 460572 128182 460624 128188
rect 460388 125248 460440 125254
rect 460388 125190 460440 125196
rect 460296 122596 460348 122602
rect 460296 122538 460348 122544
rect 460204 52080 460256 52086
rect 456338 52048 456394 52057
rect 460204 52022 460256 52028
rect 456338 51983 456394 51992
rect 469876 42770 469904 164902
rect 482388 149954 482416 167962
rect 487160 167952 487212 167958
rect 487160 167894 487212 167900
rect 486422 163432 486478 163441
rect 486422 163367 486478 163376
rect 486436 153882 486464 163367
rect 486424 153876 486476 153882
rect 486424 153818 486476 153824
rect 487172 149954 487200 167894
rect 491576 167816 491628 167822
rect 491576 167758 491628 167764
rect 491588 149954 491616 167758
rect 500960 167748 501012 167754
rect 500960 167690 501012 167696
rect 496174 164384 496230 164393
rect 496174 164319 496230 164328
rect 496188 149954 496216 164319
rect 500972 149954 501000 167690
rect 504364 166388 504416 166394
rect 504364 166330 504416 166336
rect 504376 153202 504404 166330
rect 508504 166320 508556 166326
rect 508504 166262 508556 166268
rect 504364 153196 504416 153202
rect 504364 153138 504416 153144
rect 505468 153196 505520 153202
rect 505468 153138 505520 153144
rect 505480 149954 505508 153138
rect 508516 151910 508544 166262
rect 514760 165708 514812 165714
rect 514760 165650 514812 165656
rect 508504 151904 508556 151910
rect 508504 151846 508556 151852
rect 510068 151904 510120 151910
rect 510068 151846 510120 151852
rect 510080 149954 510108 151846
rect 514772 149954 514800 165650
rect 519176 165640 519228 165646
rect 519176 165582 519228 165588
rect 519188 149954 519216 165582
rect 523776 164892 523828 164898
rect 523776 164834 523828 164840
rect 523788 149954 523816 164834
rect 528560 153876 528612 153882
rect 528560 153818 528612 153824
rect 528572 149954 528600 153818
rect 532988 149954 533016 171106
rect 536116 167006 536144 301446
rect 537484 296064 537536 296070
rect 537484 296006 537536 296012
rect 537496 245614 537524 296006
rect 537484 245608 537536 245614
rect 537484 245550 537536 245556
rect 538876 193186 538904 315318
rect 540244 294568 540296 294574
rect 540244 294510 540296 294516
rect 540256 233238 540284 294510
rect 540244 233232 540296 233238
rect 540244 233174 540296 233180
rect 538864 193180 538916 193186
rect 538864 193122 538916 193128
rect 536840 185632 536892 185638
rect 536840 185574 536892 185580
rect 536852 171134 536880 185574
rect 536852 171106 537432 171134
rect 536104 167000 536156 167006
rect 536104 166942 536156 166948
rect 537404 151814 537432 171106
rect 537484 167680 537536 167686
rect 537484 167622 537536 167628
rect 537496 152522 537524 167622
rect 537484 152516 537536 152522
rect 537484 152458 537536 152464
rect 542912 152516 542964 152522
rect 542912 152458 542964 152464
rect 542924 151842 542952 152458
rect 542912 151836 542964 151842
rect 537404 151786 537616 151814
rect 537588 149954 537616 151786
rect 542912 151778 542964 151784
rect 542924 149954 542952 151778
rect 482388 149926 482816 149954
rect 487172 149926 487416 149954
rect 491588 149926 492016 149954
rect 496188 149926 496616 149954
rect 500972 149926 501216 149954
rect 505480 149926 505816 149954
rect 510080 149926 510416 149954
rect 514772 149926 515016 149954
rect 519188 149926 519616 149954
rect 523788 149926 524216 149954
rect 528572 149926 528816 149954
rect 532988 149926 533416 149954
rect 537588 149926 538016 149954
rect 542616 149926 542952 149954
rect 543016 149734 543044 318174
rect 548524 318164 548576 318170
rect 548524 318106 548576 318112
rect 544384 307080 544436 307086
rect 544384 307022 544436 307028
rect 543096 280832 543148 280838
rect 543096 280774 543148 280780
rect 543108 179382 543136 280774
rect 543096 179376 543148 179382
rect 543096 179318 543148 179324
rect 544396 153202 544424 307022
rect 546500 300076 546552 300082
rect 546500 300018 546552 300024
rect 546512 171134 546540 300018
rect 546512 171106 546816 171134
rect 544384 153196 544436 153202
rect 544384 153138 544436 153144
rect 546788 149954 546816 171106
rect 546788 149926 547216 149954
rect 543004 149728 543056 149734
rect 543004 149670 543056 149676
rect 548536 149462 548564 318106
rect 548616 318096 548668 318102
rect 548616 318038 548668 318044
rect 548628 149530 548656 318038
rect 570708 317286 570736 456758
rect 570788 378208 570840 378214
rect 570788 378150 570840 378156
rect 570800 319870 570828 378150
rect 570788 319864 570840 319870
rect 570788 319806 570840 319812
rect 571996 317422 572024 616830
rect 572076 364404 572128 364410
rect 572076 364346 572128 364352
rect 572088 320006 572116 364346
rect 572076 320000 572128 320006
rect 572076 319942 572128 319948
rect 571984 317416 572036 317422
rect 571984 317358 572036 317364
rect 573376 317354 573404 670686
rect 580170 670647 580226 670656
rect 577504 630692 577556 630698
rect 577504 630634 577556 630640
rect 577516 318646 577544 630634
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 579632 576910 579660 577623
rect 579620 576904 579672 576910
rect 579620 576846 579672 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580276 465730 580304 697167
rect 580354 644056 580410 644065
rect 580354 643991 580410 644000
rect 580368 599622 580396 643991
rect 580446 630864 580502 630873
rect 580446 630799 580502 630808
rect 580460 630698 580488 630799
rect 580448 630692 580500 630698
rect 580448 630634 580500 630640
rect 580356 599616 580408 599622
rect 580356 599558 580408 599564
rect 580446 591016 580502 591025
rect 580446 590951 580502 590960
rect 580354 524512 580410 524521
rect 580354 524447 580410 524456
rect 580264 465724 580316 465730
rect 580264 465666 580316 465672
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580262 431624 580318 431633
rect 580262 431559 580318 431568
rect 579618 378448 579674 378457
rect 579618 378383 579674 378392
rect 579632 378214 579660 378383
rect 579620 378208 579672 378214
rect 579620 378150 579672 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 579986 325272 580042 325281
rect 579986 325207 580042 325216
rect 580000 319462 580028 325207
rect 580276 319530 580304 431559
rect 580368 322250 580396 524447
rect 580460 411942 580488 590951
rect 580538 484664 580594 484673
rect 580538 484599 580594 484608
rect 580448 411936 580500 411942
rect 580448 411878 580500 411884
rect 580446 404968 580502 404977
rect 580446 404903 580502 404912
rect 580356 322244 580408 322250
rect 580356 322186 580408 322192
rect 580264 319524 580316 319530
rect 580264 319466 580316 319472
rect 579988 319456 580040 319462
rect 579988 319398 580040 319404
rect 580460 318714 580488 404903
rect 580552 320958 580580 484599
rect 580630 418296 580686 418305
rect 580630 418231 580686 418240
rect 580540 320952 580592 320958
rect 580540 320894 580592 320900
rect 580644 320890 580672 418231
rect 580722 351928 580778 351937
rect 580722 351863 580778 351872
rect 580632 320884 580684 320890
rect 580632 320826 580684 320832
rect 580448 318708 580500 318714
rect 580448 318650 580500 318656
rect 577504 318640 577556 318646
rect 577504 318582 577556 318588
rect 580736 317898 580764 351863
rect 580724 317892 580776 317898
rect 580724 317834 580776 317840
rect 573364 317348 573416 317354
rect 573364 317290 573416 317296
rect 570696 317280 570748 317286
rect 570696 317222 570748 317228
rect 550916 314084 550968 314090
rect 550916 314026 550968 314032
rect 550640 314016 550692 314022
rect 550640 313958 550692 313964
rect 549536 312792 549588 312798
rect 549536 312734 549588 312740
rect 549352 308508 549404 308514
rect 549352 308450 549404 308456
rect 549260 307148 549312 307154
rect 549260 307090 549312 307096
rect 548616 149524 548668 149530
rect 548616 149466 548668 149472
rect 548524 149456 548576 149462
rect 548524 149398 548576 149404
rect 549166 148200 549222 148209
rect 549166 148135 549222 148144
rect 549180 146062 549208 148135
rect 549168 146056 549220 146062
rect 549168 145998 549220 146004
rect 549272 93854 549300 307090
rect 549364 96801 549392 308450
rect 549444 273964 549496 273970
rect 549444 273906 549496 273912
rect 549456 99385 549484 273906
rect 549548 138689 549576 312734
rect 549628 272604 549680 272610
rect 549628 272546 549680 272552
rect 549534 138680 549590 138689
rect 549534 138615 549590 138624
rect 549640 104417 549668 272546
rect 549812 271312 549864 271318
rect 549812 271254 549864 271260
rect 549720 270020 549772 270026
rect 549720 269962 549772 269968
rect 549732 131073 549760 269962
rect 549824 136241 549852 271254
rect 549904 146056 549956 146062
rect 549902 146024 549904 146033
rect 549956 146024 549958 146033
rect 549902 145959 549958 145968
rect 549810 136232 549866 136241
rect 549810 136167 549866 136176
rect 549718 131064 549774 131073
rect 549718 130999 549774 131008
rect 549626 104408 549682 104417
rect 549626 104343 549682 104352
rect 549442 99376 549498 99385
rect 549442 99311 549498 99320
rect 549350 96792 549406 96801
rect 549350 96727 549406 96736
rect 549272 93826 549392 93854
rect 549364 84833 549392 93826
rect 549350 84824 549406 84833
rect 549350 84759 549406 84768
rect 550652 81841 550680 313958
rect 550824 312724 550876 312730
rect 550824 312666 550876 312672
rect 550732 312656 550784 312662
rect 550732 312598 550784 312604
rect 550744 106321 550772 312598
rect 550836 111217 550864 312666
rect 550928 113665 550956 314026
rect 566464 313948 566516 313954
rect 566464 313890 566516 313896
rect 551008 311296 551060 311302
rect 551008 311238 551060 311244
rect 551020 116113 551048 311238
rect 552480 311228 552532 311234
rect 552480 311170 552532 311176
rect 552296 308576 552348 308582
rect 552296 308518 552348 308524
rect 551192 278044 551244 278050
rect 551192 277986 551244 277992
rect 551100 268388 551152 268394
rect 551100 268330 551152 268336
rect 551006 116104 551062 116113
rect 551006 116039 551062 116048
rect 550914 113656 550970 113665
rect 550914 113591 550970 113600
rect 550822 111208 550878 111217
rect 550822 111143 550878 111152
rect 551112 108769 551140 268330
rect 551204 123457 551232 277986
rect 552204 271244 552256 271250
rect 552204 271186 552256 271192
rect 552020 271176 552072 271182
rect 552020 271118 552072 271124
rect 551376 269884 551428 269890
rect 551376 269826 551428 269832
rect 551284 268456 551336 268462
rect 551284 268398 551336 268404
rect 551190 123448 551246 123457
rect 551190 123383 551246 123392
rect 551296 118561 551324 268398
rect 551388 121009 551416 269826
rect 551468 151836 551520 151842
rect 551468 151778 551520 151784
rect 551374 121000 551430 121009
rect 551374 120935 551430 120944
rect 551282 118552 551338 118561
rect 551282 118487 551338 118496
rect 551098 108760 551154 108769
rect 551098 108695 551154 108704
rect 550730 106312 550786 106321
rect 550730 106247 550786 106256
rect 550638 81832 550694 81841
rect 550638 81767 550694 81776
rect 551480 53242 551508 151778
rect 552032 86737 552060 271118
rect 552112 149456 552164 149462
rect 552112 149398 552164 149404
rect 552124 143041 552152 149398
rect 552110 143032 552166 143041
rect 552110 142967 552166 142976
rect 552112 142928 552164 142934
rect 552112 142870 552164 142876
rect 552124 101425 552152 142870
rect 552110 101416 552166 101425
rect 552110 101351 552166 101360
rect 552216 89185 552244 271186
rect 552308 128353 552336 308518
rect 552388 272536 552440 272542
rect 552388 272478 552440 272484
rect 552294 128344 552350 128353
rect 552294 128279 552350 128288
rect 552400 94081 552428 272478
rect 552492 133249 552520 311170
rect 558184 311160 558236 311166
rect 558184 311102 558236 311108
rect 552756 309868 552808 309874
rect 552756 309810 552808 309816
rect 552572 268524 552624 268530
rect 552572 268466 552624 268472
rect 552584 140593 552612 268466
rect 552664 149728 552716 149734
rect 552664 149670 552716 149676
rect 552676 142934 552704 149670
rect 552664 142928 552716 142934
rect 552664 142870 552716 142876
rect 552664 142792 552716 142798
rect 552664 142734 552716 142740
rect 552570 140584 552626 140593
rect 552570 140519 552626 140528
rect 552478 133240 552534 133249
rect 552478 133175 552534 133184
rect 552386 94072 552442 94081
rect 552386 94007 552442 94016
rect 552676 91633 552704 142734
rect 552768 125905 552796 309810
rect 555424 302864 555476 302870
rect 555424 302806 555476 302812
rect 554780 269952 554832 269958
rect 554780 269894 554832 269900
rect 552848 149524 552900 149530
rect 552848 149466 552900 149472
rect 552860 142798 552888 149466
rect 552848 142792 552900 142798
rect 552848 142734 552900 142740
rect 552754 125896 552810 125905
rect 552754 125831 552810 125840
rect 552662 91624 552718 91633
rect 552662 91559 552718 91568
rect 552202 89176 552258 89185
rect 552202 89111 552258 89120
rect 552018 86728 552074 86737
rect 552018 86663 552074 86672
rect 538128 53236 538180 53242
rect 538128 53178 538180 53184
rect 551468 53236 551520 53242
rect 551468 53178 551520 53184
rect 469864 42764 469916 42770
rect 469864 42706 469916 42712
rect 536840 42764 536892 42770
rect 536840 42706 536892 42712
rect 536852 41993 536880 42706
rect 536838 41984 536894 41993
rect 536838 41919 536894 41928
rect 456248 36576 456300 36582
rect 456248 36518 456300 36524
rect 538140 34105 538168 53178
rect 554792 53106 554820 269894
rect 555436 86970 555464 302806
rect 558196 126954 558224 311102
rect 562324 309800 562376 309806
rect 562324 309742 562376 309748
rect 559564 300008 559616 300014
rect 559564 299950 559616 299956
rect 558184 126948 558236 126954
rect 558184 126890 558236 126896
rect 555424 86964 555476 86970
rect 555424 86906 555476 86912
rect 559576 73166 559604 299950
rect 562336 113150 562364 309742
rect 562324 113144 562376 113150
rect 562324 113086 562376 113092
rect 559564 73160 559616 73166
rect 559564 73102 559616 73108
rect 540612 53100 540664 53106
rect 540612 53042 540664 53048
rect 554780 53100 554832 53106
rect 554780 53042 554832 53048
rect 540624 50425 540652 53042
rect 540610 50416 540666 50425
rect 540610 50351 540666 50360
rect 538126 34096 538182 34105
rect 538126 34031 538182 34040
rect 566476 6866 566504 313890
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 569224 308440 569276 308446
rect 569224 308382 569276 308388
rect 569236 46918 569264 308382
rect 570604 305924 570656 305930
rect 570604 305866 570656 305872
rect 569224 46912 569276 46918
rect 569224 46854 569276 46860
rect 570616 33114 570644 305866
rect 573364 304428 573416 304434
rect 573364 304370 573416 304376
rect 571984 290488 572036 290494
rect 571984 290430 572036 290436
rect 570604 33108 570656 33114
rect 570604 33050 570656 33056
rect 571996 20670 572024 290430
rect 573376 60722 573404 304370
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 576124 293276 576176 293282
rect 576124 293218 576176 293224
rect 574744 291780 574796 291786
rect 574744 291722 574796 291728
rect 574756 100706 574784 291722
rect 576136 139398 576164 293218
rect 580356 288992 580408 288998
rect 580356 288934 580408 288940
rect 580264 287700 580316 287706
rect 580264 287642 580316 287648
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580276 219065 580304 287642
rect 580368 272241 580396 288934
rect 580354 272232 580410 272241
rect 580354 272167 580410 272176
rect 580356 269816 580408 269822
rect 580356 269758 580408 269764
rect 580368 258913 580396 269758
rect 580354 258904 580410 258913
rect 580354 258839 580410 258848
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 576124 139392 576176 139398
rect 580172 139392 580224 139398
rect 576124 139334 576176 139340
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 574744 100700 574796 100706
rect 574744 100642 574796 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 573364 60716 573416 60722
rect 573364 60658 573416 60664
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 571984 20664 572036 20670
rect 571984 20606 572036 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 566464 6860 566516 6866
rect 566464 6802 566516 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 456156 3528 456208 3534
rect 456156 3470 456208 3476
rect 454774 3431 454830 3440
rect 456064 3460 456116 3466
rect 456064 3402 456116 3408
rect 392584 2100 392636 2106
rect 392584 2042 392636 2048
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 8114 668480 8170 668536
rect 3422 658144 3478 658200
rect 3146 619112 3202 619168
rect 3698 632032 3754 632088
rect 3606 579944 3662 580000
rect 3514 527856 3570 527912
rect 3422 501744 3478 501800
rect 3790 606056 3846 606112
rect 3790 566888 3846 566944
rect 3698 514800 3754 514856
rect 3606 462576 3662 462632
rect 3514 423544 3570 423600
rect 3974 553832 4030 553888
rect 40498 700304 40554 700360
rect 105450 700440 105506 700496
rect 202786 671336 202842 671392
rect 300122 700576 300178 700632
rect 24306 668616 24362 668672
rect 3882 475632 3938 475688
rect 3790 449520 3846 449576
rect 3698 410488 3754 410544
rect 382278 662360 382334 662416
rect 382278 651752 382334 651808
rect 382922 641144 382978 641200
rect 382278 630536 382334 630592
rect 382278 619928 382334 619984
rect 382278 609320 382334 609376
rect 382278 598712 382334 598768
rect 382278 588104 382334 588160
rect 382278 577496 382334 577552
rect 382278 566888 382334 566944
rect 382278 556280 382334 556336
rect 382278 545672 382334 545728
rect 382278 535064 382334 535120
rect 382278 524476 382334 524512
rect 382278 524456 382280 524476
rect 382280 524456 382332 524476
rect 382332 524456 382334 524476
rect 382278 513848 382334 513904
rect 382278 503240 382334 503296
rect 382278 492668 382280 492688
rect 382280 492668 382332 492688
rect 382332 492668 382334 492688
rect 382278 492632 382334 492668
rect 382278 482024 382334 482080
rect 382370 471416 382426 471472
rect 382278 460808 382334 460864
rect 382278 450200 382334 450256
rect 383014 439592 383070 439648
rect 382278 407768 382334 407824
rect 3514 397432 3570 397488
rect 3422 371320 3478 371376
rect 382278 397160 382334 397216
rect 382278 386552 382334 386608
rect 382278 375944 382334 376000
rect 383106 428984 383162 429040
rect 382646 365336 382702 365392
rect 383198 418376 383254 418432
rect 3606 358400 3662 358456
rect 382922 354728 382978 354784
rect 3698 345344 3754 345400
rect 3606 293120 3662 293176
rect 3514 241032 3570 241088
rect 3422 214920 3478 214976
rect 382278 344120 382334 344176
rect 3974 319232 4030 319288
rect 3882 306176 3938 306232
rect 3790 267144 3846 267200
rect 3698 254088 3754 254144
rect 422206 336776 422262 336832
rect 383106 333512 383162 333568
rect 383014 322904 383070 322960
rect 382922 312296 382978 312352
rect 3882 201864 3938 201920
rect 3790 162832 3846 162888
rect 3606 149776 3662 149832
rect 3514 110608 3570 110664
rect 3422 97552 3478 97608
rect 3330 84632 3386 84688
rect 3422 71576 3478 71632
rect 3698 136720 3754 136776
rect 3974 188808 4030 188864
rect 3606 58520 3662 58576
rect 3606 51992 3662 52048
rect 7654 50496 7710 50552
rect 2870 50360 2926 50416
rect 1674 3576 1730 3632
rect 570 3304 626 3360
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 5262 3984 5318 4040
rect 4066 3440 4122 3496
rect 6458 3712 6514 3768
rect 18602 51856 18658 51912
rect 51354 50768 51410 50824
rect 47858 50632 47914 50688
rect 46662 50224 46718 50280
rect 9954 3848 10010 3904
rect 380438 3984 380494 4040
rect 382278 301688 382334 301744
rect 382278 280472 382334 280528
rect 382278 269864 382334 269920
rect 382278 259256 382334 259312
rect 382278 248648 382334 248704
rect 382278 238040 382334 238096
rect 382278 227432 382334 227488
rect 382278 206216 382334 206272
rect 382278 195608 382334 195664
rect 382278 185000 382334 185056
rect 382278 174392 382334 174448
rect 382278 153176 382334 153232
rect 382278 142568 382334 142624
rect 382278 131960 382334 132016
rect 382278 110744 382334 110800
rect 382278 100136 382334 100192
rect 382278 89528 382334 89584
rect 382278 78920 382334 78976
rect 382278 68312 382334 68368
rect 382278 57704 382334 57760
rect 384302 294480 384358 294536
rect 383290 291080 383346 291136
rect 383382 216824 383438 216880
rect 383474 121352 383530 121408
rect 385866 291760 385922 291816
rect 389822 297472 389878 297528
rect 388442 291896 388498 291952
rect 388442 3848 388498 3904
rect 391478 294616 391534 294672
rect 393042 300192 393098 300248
rect 392858 300056 392914 300112
rect 392950 297336 393006 297392
rect 398194 302776 398250 302832
rect 402334 289176 402390 289232
rect 402518 289040 402574 289096
rect 403714 50768 403770 50824
rect 406382 305768 406438 305824
rect 403898 50632 403954 50688
rect 406750 305904 406806 305960
rect 406566 305632 406622 305688
rect 406474 51856 406530 51912
rect 407762 286320 407818 286376
rect 406750 50496 406806 50552
rect 406566 50360 406622 50416
rect 407762 3712 407818 3768
rect 409142 163376 409198 163432
rect 433982 334736 434038 334792
rect 433430 330792 433486 330848
rect 434442 326848 434498 326904
rect 434074 322904 434130 322960
rect 433522 318960 433578 319016
rect 434258 315052 434260 315072
rect 434260 315052 434312 315072
rect 434312 315052 434314 315072
rect 434258 315016 434314 315052
rect 433982 311072 434038 311128
rect 433890 307128 433946 307184
rect 445390 668480 445446 668536
rect 445390 318688 445446 318744
rect 447138 375808 447194 375864
rect 447138 375284 447194 375320
rect 447138 375264 447140 375284
rect 447140 375264 447192 375284
rect 447192 375264 447194 375284
rect 447230 374720 447286 374776
rect 447322 374176 447378 374232
rect 447138 373632 447194 373688
rect 447230 373088 447286 373144
rect 447138 372544 447194 372600
rect 447322 372000 447378 372056
rect 447230 371456 447286 371512
rect 447138 370912 447194 370968
rect 447230 370368 447286 370424
rect 447322 369824 447378 369880
rect 447138 369280 447194 369336
rect 447230 368736 447286 368792
rect 447138 368192 447194 368248
rect 447230 367648 447286 367704
rect 447322 367104 447378 367160
rect 447138 366560 447194 366616
rect 447230 366016 447286 366072
rect 447138 365508 447140 365528
rect 447140 365508 447192 365528
rect 447192 365508 447194 365528
rect 447138 365472 447194 365508
rect 447230 364928 447286 364984
rect 447322 364384 447378 364440
rect 447138 363840 447194 363896
rect 447230 363296 447286 363352
rect 447138 362752 447194 362808
rect 447230 362208 447286 362264
rect 447322 361664 447378 361720
rect 447138 361120 447194 361176
rect 447230 360576 447286 360632
rect 447230 360032 447286 360088
rect 447138 359488 447194 359544
rect 447322 358964 447378 359000
rect 447322 358944 447324 358964
rect 447324 358944 447376 358964
rect 447376 358944 447378 358964
rect 447230 358400 447286 358456
rect 447138 357856 447194 357912
rect 447230 357312 447286 357368
rect 447138 356224 447194 356280
rect 447322 356768 447378 356824
rect 447414 353504 447470 353560
rect 447138 350240 447194 350296
rect 447230 349696 447286 349752
rect 447322 349152 447378 349208
rect 447230 348608 447286 348664
rect 447138 348064 447194 348120
rect 447138 347556 447140 347576
rect 447140 347556 447192 347576
rect 447192 347556 447194 347576
rect 447138 347520 447194 347556
rect 447230 346976 447286 347032
rect 447322 346432 447378 346488
rect 447138 345344 447194 345400
rect 447138 342624 447194 342680
rect 447598 342080 447654 342136
rect 447138 338272 447194 338328
rect 447690 338000 447746 338056
rect 447230 337728 447286 337784
rect 447138 337184 447194 337240
rect 447690 336776 447746 336832
rect 447230 336640 447286 336696
rect 447138 336096 447194 336152
rect 447322 335552 447378 335608
rect 447230 335008 447286 335064
rect 447138 334464 447194 334520
rect 447230 333920 447286 333976
rect 447138 333376 447194 333432
rect 447322 332832 447378 332888
rect 447138 331744 447194 331800
rect 447230 331200 447286 331256
rect 447414 332288 447470 332344
rect 447506 330112 447562 330168
rect 446954 318552 447010 318608
rect 446494 276664 446550 276720
rect 447874 352960 447930 353016
rect 447966 344256 448022 344312
rect 448058 343712 448114 343768
rect 448150 341536 448206 341592
rect 448058 340992 448114 341048
rect 447874 340448 447930 340504
rect 447966 329704 448022 329760
rect 447966 329024 448022 329080
rect 448150 330656 448206 330712
rect 448334 355136 448390 355192
rect 448334 345888 448390 345944
rect 448242 329704 448298 329760
rect 448242 329604 448244 329624
rect 448244 329604 448296 329624
rect 448296 329604 448298 329624
rect 448242 329568 448298 329604
rect 448242 328500 448298 328536
rect 448242 328480 448244 328500
rect 448244 328480 448296 328500
rect 448296 328480 448298 328500
rect 449070 354048 449126 354104
rect 448518 327936 448574 327992
rect 543462 699760 543518 699816
rect 458730 678544 458786 678600
rect 457902 632848 457958 632904
rect 457810 629992 457866 630048
rect 457718 627136 457774 627192
rect 457626 621424 457682 621480
rect 457534 615712 457590 615768
rect 457442 612856 457498 612912
rect 457350 610000 457406 610056
rect 458086 624280 458142 624336
rect 457994 618568 458050 618624
rect 457902 607144 457958 607200
rect 459282 669976 459338 670032
rect 459098 664264 459154 664320
rect 459006 652840 459062 652896
rect 458914 647128 458970 647184
rect 458822 641416 458878 641472
rect 458730 599528 458786 599584
rect 458822 596808 458878 596864
rect 459190 658552 459246 658608
rect 460570 666576 460626 666632
rect 460386 661000 460442 661056
rect 460478 655852 460534 655888
rect 460478 655832 460480 655852
rect 460480 655832 460532 655852
rect 460532 655832 460534 655852
rect 460386 650120 460442 650176
rect 460294 643748 460350 643784
rect 460294 643728 460296 643748
rect 460296 643728 460348 643748
rect 460348 643728 460350 643748
rect 459466 638560 459522 638616
rect 459374 604288 459430 604344
rect 459374 593952 459430 594008
rect 460570 600888 460626 600944
rect 459466 518064 459522 518120
rect 449990 512352 450046 512408
rect 449254 355680 449310 355736
rect 449346 352416 449402 352472
rect 449622 354592 449678 354648
rect 449530 351872 449586 351928
rect 449714 351328 449770 351384
rect 449438 350784 449494 350840
rect 449714 344800 449770 344856
rect 449622 324128 449678 324184
rect 449806 343168 449862 343224
rect 449806 339904 449862 339960
rect 450082 510176 450138 510232
rect 450450 516976 450506 517032
rect 450542 514664 450598 514720
rect 450450 512352 450506 512408
rect 450358 510176 450414 510232
rect 450266 507592 450322 507648
rect 450174 505416 450230 505472
rect 450082 339108 450138 339144
rect 450082 339088 450084 339108
rect 450084 339088 450136 339108
rect 450136 339088 450138 339108
rect 449990 327120 450046 327176
rect 449898 326576 449954 326632
rect 450542 503240 450598 503296
rect 450266 338000 450322 338056
rect 464434 501064 464490 501120
rect 482742 517520 482798 517576
rect 480442 516860 480498 516896
rect 480442 516840 480444 516860
rect 480444 516840 480496 516860
rect 480496 516840 480498 516860
rect 492126 516840 492182 516896
rect 491850 516568 491906 516624
rect 492126 508884 492182 508940
rect 478142 467064 478198 467120
rect 472806 382336 472862 382392
rect 489182 391176 489238 391232
rect 475382 382336 475438 382392
rect 490838 382336 490894 382392
rect 492126 382336 492182 382392
rect 494702 520920 494758 520976
rect 494150 512488 494206 512544
rect 494150 505164 494206 505200
rect 494150 505144 494152 505164
rect 494152 505144 494204 505164
rect 494204 505144 494206 505164
rect 494794 515924 494796 515944
rect 494796 515924 494848 515944
rect 494848 515924 494850 515944
rect 494794 515888 494850 515924
rect 494794 501200 494850 501256
rect 506478 537376 506534 537432
rect 506570 516976 506626 517032
rect 510986 361120 511042 361176
rect 510802 360304 510858 360360
rect 510066 359080 510122 359136
rect 450358 326576 450414 326632
rect 450266 326032 450322 326088
rect 450542 326032 450598 326088
rect 450174 325488 450230 325544
rect 450082 324944 450138 325000
rect 450450 323856 450506 323912
rect 450634 325488 450690 325544
rect 450634 324944 450690 325000
rect 464434 320320 464490 320376
rect 423264 164328 423320 164384
rect 454774 315288 454830 315344
rect 406382 3576 406438 3632
rect 455050 50224 455106 50280
rect 454774 3440 454830 3496
rect 460018 320048 460074 320104
rect 461122 319776 461178 319832
rect 462134 319912 462190 319968
rect 461950 319504 462006 319560
rect 456798 262656 456854 262712
rect 457166 234948 457168 234968
rect 457168 234948 457220 234968
rect 457220 234948 457222 234968
rect 457166 234912 457222 234948
rect 457350 221040 457406 221096
rect 456798 207204 456800 207224
rect 456800 207204 456852 207224
rect 456852 207204 456854 207224
rect 456798 207168 456854 207204
rect 457258 207168 457314 207224
rect 456798 161064 456854 161120
rect 456798 159568 456854 159624
rect 456798 156576 456854 156632
rect 456798 155080 456854 155136
rect 456798 153584 456854 153640
rect 456890 150628 456892 150648
rect 456892 150628 456944 150648
rect 456944 150628 456946 150648
rect 456890 150592 456946 150628
rect 456798 149096 456854 149152
rect 457442 147600 457498 147656
rect 456798 144644 456800 144664
rect 456800 144644 456852 144664
rect 456852 144644 456854 144664
rect 456798 144608 456854 144644
rect 456798 143148 456800 143168
rect 456800 143148 456852 143168
rect 456852 143148 456854 143168
rect 456798 143112 456854 143148
rect 457258 141652 457260 141672
rect 457260 141652 457312 141672
rect 457312 141652 457314 141672
rect 457258 141616 457314 141652
rect 456798 140120 456854 140176
rect 457258 138624 457314 138680
rect 457258 137128 457314 137184
rect 457994 248784 458050 248840
rect 458086 234912 458142 234968
rect 457902 162560 457958 162616
rect 457810 158072 457866 158128
rect 457718 152088 457774 152144
rect 457626 146104 457682 146160
rect 457534 134136 457590 134192
rect 457074 132640 457130 132696
rect 457442 128188 457444 128208
rect 457444 128188 457496 128208
rect 457496 128188 457498 128208
rect 457442 128152 457498 128188
rect 457350 125196 457352 125216
rect 457352 125196 457404 125216
rect 457404 125196 457406 125216
rect 457350 125160 457406 125196
rect 457074 122168 457130 122224
rect 472714 318280 472770 318336
rect 480718 318280 480774 318336
rect 482374 318416 482430 318472
rect 483202 318688 483258 318744
rect 483478 318552 483534 318608
rect 488722 301416 488778 301472
rect 488630 278024 488686 278080
rect 490286 306992 490342 307048
rect 490010 272448 490066 272504
rect 489918 268368 489974 268424
rect 508502 319912 508558 319968
rect 503442 309712 503498 309768
rect 503534 300328 503590 300384
rect 510710 348064 510766 348120
rect 510618 342352 510674 342408
rect 510158 327664 510214 327720
rect 510066 324808 510122 324864
rect 510066 320184 510122 320240
rect 510342 327256 510398 327312
rect 510250 326032 510306 326088
rect 510434 326848 510490 326904
rect 510434 320592 510490 320648
rect 510894 345616 510950 345672
rect 511078 355816 511134 355872
rect 511170 337048 511226 337104
rect 511078 320456 511134 320512
rect 510986 320320 511042 320376
rect 512826 378664 512882 378720
rect 512734 378256 512790 378312
rect 512918 377848 512974 377904
rect 512642 377440 512698 377496
rect 512274 377032 512330 377088
rect 512274 375400 512330 375456
rect 512090 374992 512146 375048
rect 511998 372952 512054 373008
rect 513286 376624 513342 376680
rect 513194 376216 513250 376272
rect 513102 375808 513158 375864
rect 513286 374584 513342 374640
rect 512826 374176 512882 374232
rect 513286 373768 513342 373824
rect 513286 373360 513342 373416
rect 513286 372564 513342 372600
rect 513286 372544 513288 372564
rect 513288 372544 513340 372564
rect 513340 372544 513342 372564
rect 512734 372136 512790 372192
rect 512458 371764 512460 371784
rect 512460 371764 512512 371784
rect 512512 371764 512514 371784
rect 512458 371728 512514 371764
rect 513194 371320 513250 371376
rect 513286 370912 513342 370968
rect 513194 370504 513250 370560
rect 513102 370096 513158 370152
rect 513102 369708 513158 369744
rect 513102 369688 513104 369708
rect 513104 369688 513156 369708
rect 513156 369688 513158 369708
rect 513286 369280 513342 369336
rect 513286 368872 513342 368928
rect 513194 368464 513250 368520
rect 512182 368056 512238 368112
rect 512274 367648 512330 367704
rect 513286 367240 513342 367296
rect 513010 366832 513066 366888
rect 512826 366016 512882 366072
rect 512090 363976 512146 364032
rect 512642 362752 512698 362808
rect 512090 361956 512146 361992
rect 512090 361936 512092 361956
rect 512092 361936 512144 361956
rect 512144 361936 512146 361956
rect 513194 366424 513250 366480
rect 512918 365608 512974 365664
rect 513194 365200 513250 365256
rect 513102 364792 513158 364848
rect 513010 363180 513066 363216
rect 513010 363160 513012 363180
rect 513012 363160 513064 363180
rect 513064 363160 513066 363180
rect 513286 364404 513342 364440
rect 513286 364384 513288 364404
rect 513288 364384 513340 364404
rect 513340 364384 513342 364404
rect 513286 363568 513342 363624
rect 513286 362344 513342 362400
rect 513286 361528 513342 361584
rect 513102 360712 513158 360768
rect 513010 359896 513066 359952
rect 513286 359488 513342 359544
rect 511998 358672 512054 358728
rect 511538 335824 511594 335880
rect 511262 318280 511318 318336
rect 511906 326440 511962 326496
rect 511722 319912 511778 319968
rect 513010 358264 513066 358320
rect 512090 357856 512146 357912
rect 513286 357468 513342 357504
rect 513286 357448 513288 357468
rect 513288 357448 513340 357468
rect 513340 357448 513342 357468
rect 512182 357040 512238 357096
rect 512090 356224 512146 356280
rect 512642 356632 512698 356688
rect 512734 355408 512790 355464
rect 513286 355000 513342 355056
rect 513102 354592 513158 354648
rect 512550 354184 512606 354240
rect 512182 353776 512238 353832
rect 513286 352552 513342 352608
rect 512274 352144 512330 352200
rect 512182 349288 512238 349344
rect 512182 346840 512238 346896
rect 512642 351756 512698 351792
rect 512642 351736 512644 351756
rect 512644 351736 512696 351756
rect 512696 351736 512698 351756
rect 513286 351328 513342 351384
rect 512642 350940 512698 350976
rect 512642 350920 512644 350940
rect 512644 350920 512696 350940
rect 512696 350920 512698 350940
rect 513286 350548 513288 350568
rect 513288 350548 513340 350568
rect 513340 350548 513342 350568
rect 513286 350512 513342 350548
rect 512826 350104 512882 350160
rect 513286 349696 513342 349752
rect 513194 348880 513250 348936
rect 513286 348472 513342 348528
rect 513010 347656 513066 347712
rect 512826 347248 512882 347304
rect 512458 346432 512514 346488
rect 512274 344392 512330 344448
rect 512366 343168 512422 343224
rect 512366 342760 512422 342816
rect 512274 341944 512330 342000
rect 512274 341128 512330 341184
rect 512366 340720 512422 340776
rect 512366 339516 512422 339552
rect 512366 339496 512368 339516
rect 512368 339496 512420 339516
rect 512420 339496 512422 339516
rect 513194 346024 513250 346080
rect 513286 345208 513342 345264
rect 513286 344800 513342 344856
rect 512826 343984 512882 344040
rect 513286 343576 513342 343632
rect 513286 341536 513342 341592
rect 513010 340312 513066 340368
rect 513286 339924 513342 339960
rect 513286 339904 513288 339924
rect 513288 339904 513340 339924
rect 513340 339904 513342 339924
rect 513286 339088 513342 339144
rect 513194 338680 513250 338736
rect 512550 338292 512606 338328
rect 512550 338272 512552 338292
rect 512552 338272 512604 338292
rect 512604 338272 512606 338292
rect 513010 337864 513066 337920
rect 512918 337456 512974 337512
rect 513286 336640 513342 336696
rect 513194 336232 513250 336288
rect 512734 335436 512790 335472
rect 512734 335416 512736 335436
rect 512736 335416 512788 335436
rect 512788 335416 512790 335436
rect 512826 335008 512882 335064
rect 512642 334192 512698 334248
rect 512458 330520 512514 330576
rect 512550 329704 512606 329760
rect 512550 328888 512606 328944
rect 513010 334600 513066 334656
rect 512918 333784 512974 333840
rect 512826 332968 512882 333024
rect 513286 332560 513342 332616
rect 512826 332152 512882 332208
rect 512734 331744 512790 331800
rect 512642 325488 512698 325544
rect 513286 331336 513342 331392
rect 513286 329296 513342 329352
rect 513286 328072 513342 328128
rect 512826 322768 512882 322824
rect 513470 353368 513526 353424
rect 513562 352960 513618 353016
rect 516782 467200 516838 467256
rect 559654 699760 559710 699816
rect 580262 697176 580318 697232
rect 579618 683848 579674 683904
rect 523682 516704 523738 516760
rect 550638 516704 550694 516760
rect 521750 467064 521806 467120
rect 561678 444896 561734 444952
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 530030 244160 530086 244216
rect 531410 261024 531466 261080
rect 531318 226208 531374 226264
rect 529938 209208 529994 209264
rect 456338 51992 456394 52048
rect 486422 163376 486478 163432
rect 496174 164328 496230 164384
rect 580170 670656 580226 670692
rect 580170 617480 580226 617536
rect 579618 577632 579674 577688
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 580170 511264 580226 511320
rect 579986 471416 580042 471472
rect 580354 644000 580410 644056
rect 580446 630808 580502 630864
rect 580446 590960 580502 591016
rect 580354 524456 580410 524512
rect 580170 458088 580226 458144
rect 580262 431568 580318 431624
rect 579618 378392 579674 378448
rect 580170 365064 580226 365120
rect 579986 325216 580042 325272
rect 580538 484608 580594 484664
rect 580446 404912 580502 404968
rect 580630 418240 580686 418296
rect 580722 351872 580778 351928
rect 549166 148144 549222 148200
rect 549534 138624 549590 138680
rect 549902 146004 549904 146024
rect 549904 146004 549956 146024
rect 549956 146004 549958 146024
rect 549902 145968 549958 146004
rect 549810 136176 549866 136232
rect 549718 131008 549774 131064
rect 549626 104352 549682 104408
rect 549442 99320 549498 99376
rect 549350 96736 549406 96792
rect 549350 84768 549406 84824
rect 551006 116048 551062 116104
rect 550914 113600 550970 113656
rect 550822 111152 550878 111208
rect 551190 123392 551246 123448
rect 551374 120944 551430 121000
rect 551282 118496 551338 118552
rect 551098 108704 551154 108760
rect 550730 106256 550786 106312
rect 550638 81776 550694 81832
rect 552110 142976 552166 143032
rect 552110 101360 552166 101416
rect 552294 128288 552350 128344
rect 552570 140528 552626 140584
rect 552478 133184 552534 133240
rect 552386 94016 552442 94072
rect 552754 125840 552810 125896
rect 552662 91568 552718 91624
rect 552202 89120 552258 89176
rect 552018 86672 552074 86728
rect 536838 41928 536894 41984
rect 540610 50360 540666 50416
rect 538126 34040 538182 34096
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 580354 272176 580410 272232
rect 580354 258848 580410 258904
rect 580262 219000 580318 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect 300117 700634 300183 700637
rect 447910 700634 447916 700636
rect 300117 700632 447916 700634
rect 300117 700576 300122 700632
rect 300178 700576 447916 700632
rect 300117 700574 447916 700576
rect 300117 700571 300183 700574
rect 447910 700572 447916 700574
rect 447980 700572 447986 700636
rect 105445 700498 105511 700501
rect 444230 700498 444236 700500
rect 105445 700496 444236 700498
rect 105445 700440 105450 700496
rect 105506 700440 444236 700496
rect 105445 700438 444236 700440
rect 105445 700435 105511 700438
rect 444230 700436 444236 700438
rect 444300 700436 444306 700500
rect 40493 700362 40559 700365
rect 447726 700362 447732 700364
rect 40493 700360 447732 700362
rect 40493 700304 40498 700360
rect 40554 700304 447732 700360
rect 40493 700302 447732 700304
rect 40493 700299 40559 700302
rect 447726 700300 447732 700302
rect 447796 700300 447802 700364
rect 542670 699756 542676 699820
rect 542740 699818 542746 699820
rect 543457 699818 543523 699821
rect 542740 699816 543523 699818
rect 542740 699760 543462 699816
rect 543518 699760 543523 699816
rect 542740 699758 543523 699760
rect 542740 699756 542746 699758
rect 543457 699755 543523 699758
rect 558862 699756 558868 699820
rect 558932 699818 558938 699820
rect 559649 699818 559715 699821
rect 558932 699816 559715 699818
rect 558932 699760 559654 699816
rect 559710 699760 559715 699816
rect 558932 699758 559715 699760
rect 558932 699756 558938 699758
rect 559649 699755 559715 699758
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect 458725 678602 458791 678605
rect 458725 678600 460092 678602
rect 458725 678544 458730 678600
rect 458786 678544 460092 678600
rect 458725 678542 460092 678544
rect 458725 678539 458791 678542
rect 457846 675684 457852 675748
rect 457916 675746 457922 675748
rect 457916 675686 460092 675746
rect 457916 675684 457922 675686
rect 458030 672828 458036 672892
rect 458100 672890 458106 672892
rect 458100 672830 460092 672890
rect 458100 672828 458106 672830
rect 202781 671394 202847 671397
rect 448094 671394 448100 671396
rect 202781 671392 448100 671394
rect -960 671258 480 671348
rect 202781 671336 202786 671392
rect 202842 671336 448100 671392
rect 202781 671334 448100 671336
rect 202781 671331 202847 671334
rect 448094 671332 448100 671334
rect 448164 671332 448170 671396
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect 459277 670034 459343 670037
rect 459277 670032 460092 670034
rect 459277 669976 459282 670032
rect 459338 669976 460092 670032
rect 459277 669974 460092 669976
rect 459277 669971 459343 669974
rect 24301 668674 24367 668677
rect 446254 668674 446260 668676
rect 24301 668672 446260 668674
rect 24301 668616 24306 668672
rect 24362 668616 446260 668672
rect 24301 668614 446260 668616
rect 24301 668611 24367 668614
rect 446254 668612 446260 668614
rect 446324 668612 446330 668676
rect 8109 668538 8175 668541
rect 445385 668538 445451 668541
rect 8109 668536 445451 668538
rect 8109 668480 8114 668536
rect 8170 668480 445390 668536
rect 445446 668480 445451 668536
rect 8109 668478 445451 668480
rect 8109 668475 8175 668478
rect 445385 668475 445451 668478
rect 460614 666637 460674 667148
rect 460565 666632 460674 666637
rect 460565 666576 460570 666632
rect 460626 666576 460674 666632
rect 460565 666574 460674 666576
rect 460565 666571 460631 666574
rect 459093 664322 459159 664325
rect 459093 664320 460092 664322
rect 459093 664264 459098 664320
rect 459154 664264 460092 664320
rect 459093 664262 460092 664264
rect 459093 664259 459159 664262
rect 382273 662418 382339 662421
rect 379868 662416 382339 662418
rect 379868 662360 382278 662416
rect 382334 662360 382339 662416
rect 379868 662358 382339 662360
rect 382273 662355 382339 662358
rect 460430 661061 460490 661436
rect 460381 661056 460490 661061
rect 460381 661000 460386 661056
rect 460442 661000 460490 661056
rect 460381 660998 460490 661000
rect 460381 660995 460447 660998
rect 459185 658610 459251 658613
rect 459185 658608 460092 658610
rect 459185 658552 459190 658608
rect 459246 658552 460092 658608
rect 459185 658550 460092 658552
rect 459185 658547 459251 658550
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect 460473 655890 460539 655893
rect 460430 655888 460539 655890
rect 460430 655832 460478 655888
rect 460534 655832 460539 655888
rect 460430 655827 460539 655832
rect 460430 655724 460490 655827
rect 459001 652898 459067 652901
rect 459001 652896 460092 652898
rect 459001 652840 459006 652896
rect 459062 652840 460092 652896
rect 459001 652838 460092 652840
rect 459001 652835 459067 652838
rect 382273 651810 382339 651813
rect 379868 651808 382339 651810
rect 379868 651752 382278 651808
rect 382334 651752 382339 651808
rect 379868 651750 382339 651752
rect 382273 651747 382339 651750
rect 460381 650178 460447 650181
rect 460381 650176 460490 650178
rect 460381 650120 460386 650176
rect 460442 650120 460490 650176
rect 460381 650115 460490 650120
rect 460430 650012 460490 650115
rect 458909 647186 458975 647189
rect 458909 647184 460092 647186
rect 458909 647128 458914 647184
rect 458970 647128 460092 647184
rect 458909 647126 460092 647128
rect 458909 647123 458975 647126
rect -960 644996 480 645236
rect 460246 643789 460306 644300
rect 580349 644058 580415 644061
rect 583520 644058 584960 644148
rect 580349 644056 584960 644058
rect 580349 644000 580354 644056
rect 580410 644000 584960 644056
rect 580349 643998 584960 644000
rect 580349 643995 580415 643998
rect 583520 643908 584960 643998
rect 460246 643784 460355 643789
rect 460246 643728 460294 643784
rect 460350 643728 460355 643784
rect 460246 643726 460355 643728
rect 460289 643723 460355 643726
rect 458817 641474 458883 641477
rect 458817 641472 460092 641474
rect 458817 641416 458822 641472
rect 458878 641416 460092 641472
rect 458817 641414 460092 641416
rect 458817 641411 458883 641414
rect 382917 641202 382983 641205
rect 379868 641200 382983 641202
rect 379868 641144 382922 641200
rect 382978 641144 382983 641200
rect 379868 641142 382983 641144
rect 382917 641139 382983 641142
rect 459461 638618 459527 638621
rect 459461 638616 460092 638618
rect 459461 638560 459466 638616
rect 459522 638560 460092 638616
rect 459461 638558 460092 638560
rect 459461 638555 459527 638558
rect 459134 635700 459140 635764
rect 459204 635762 459210 635764
rect 459204 635702 460092 635762
rect 459204 635700 459210 635702
rect 457897 632906 457963 632909
rect 457897 632904 460092 632906
rect 457897 632848 457902 632904
rect 457958 632848 460092 632904
rect 457897 632846 460092 632848
rect 457897 632843 457963 632846
rect -960 632090 480 632180
rect 3693 632090 3759 632093
rect -960 632088 3759 632090
rect -960 632032 3698 632088
rect 3754 632032 3759 632088
rect -960 632030 3759 632032
rect -960 631940 480 632030
rect 3693 632027 3759 632030
rect 580441 630866 580507 630869
rect 583520 630866 584960 630956
rect 580441 630864 584960 630866
rect 580441 630808 580446 630864
rect 580502 630808 584960 630864
rect 580441 630806 584960 630808
rect 580441 630803 580507 630806
rect 583520 630716 584960 630806
rect 382273 630594 382339 630597
rect 379868 630592 382339 630594
rect 379868 630536 382278 630592
rect 382334 630536 382339 630592
rect 379868 630534 382339 630536
rect 382273 630531 382339 630534
rect 457805 630050 457871 630053
rect 457805 630048 460092 630050
rect 457805 629992 457810 630048
rect 457866 629992 460092 630048
rect 457805 629990 460092 629992
rect 457805 629987 457871 629990
rect 457713 627194 457779 627197
rect 457713 627192 460092 627194
rect 457713 627136 457718 627192
rect 457774 627136 460092 627192
rect 457713 627134 460092 627136
rect 457713 627131 457779 627134
rect 458081 624338 458147 624341
rect 458081 624336 460092 624338
rect 458081 624280 458086 624336
rect 458142 624280 460092 624336
rect 458081 624278 460092 624280
rect 458081 624275 458147 624278
rect 457621 621482 457687 621485
rect 457621 621480 460092 621482
rect 457621 621424 457626 621480
rect 457682 621424 460092 621480
rect 457621 621422 460092 621424
rect 457621 621419 457687 621422
rect 382273 619986 382339 619989
rect 379868 619984 382339 619986
rect 379868 619928 382278 619984
rect 382334 619928 382339 619984
rect 379868 619926 382339 619928
rect 382273 619923 382339 619926
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 457989 618626 458055 618629
rect 457989 618624 460092 618626
rect 457989 618568 457994 618624
rect 458050 618568 460092 618624
rect 457989 618566 460092 618568
rect 457989 618563 458055 618566
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 457529 615770 457595 615773
rect 457529 615768 460092 615770
rect 457529 615712 457534 615768
rect 457590 615712 460092 615768
rect 457529 615710 460092 615712
rect 457529 615707 457595 615710
rect 457437 612914 457503 612917
rect 457437 612912 460092 612914
rect 457437 612856 457442 612912
rect 457498 612856 460092 612912
rect 457437 612854 460092 612856
rect 457437 612851 457503 612854
rect 457345 610058 457411 610061
rect 457345 610056 460092 610058
rect 457345 610000 457350 610056
rect 457406 610000 460092 610056
rect 457345 609998 460092 610000
rect 457345 609995 457411 609998
rect 382273 609378 382339 609381
rect 379868 609376 382339 609378
rect 379868 609320 382278 609376
rect 382334 609320 382339 609376
rect 379868 609318 382339 609320
rect 382273 609315 382339 609318
rect 457897 607202 457963 607205
rect 457897 607200 460092 607202
rect 457897 607144 457902 607200
rect 457958 607144 460092 607200
rect 457897 607142 460092 607144
rect 457897 607139 457963 607142
rect -960 606114 480 606204
rect 3785 606114 3851 606117
rect -960 606112 3851 606114
rect -960 606056 3790 606112
rect 3846 606056 3851 606112
rect -960 606054 3851 606056
rect -960 605964 480 606054
rect 3785 606051 3851 606054
rect 459369 604346 459435 604349
rect 459369 604344 460092 604346
rect 459369 604288 459374 604344
rect 459430 604288 460092 604344
rect 459369 604286 460092 604288
rect 459369 604283 459435 604286
rect 583520 604060 584960 604300
rect 460614 600949 460674 601460
rect 460565 600944 460674 600949
rect 460565 600888 460570 600944
rect 460626 600888 460674 600944
rect 460565 600886 460674 600888
rect 460565 600883 460631 600886
rect 458725 599586 458791 599589
rect 472014 599586 472020 599588
rect 458725 599584 472020 599586
rect 458725 599528 458730 599584
rect 458786 599528 472020 599584
rect 458725 599526 472020 599528
rect 458725 599523 458791 599526
rect 472014 599524 472020 599526
rect 472084 599524 472090 599588
rect 382273 598770 382339 598773
rect 379868 598768 382339 598770
rect 379868 598712 382278 598768
rect 382334 598712 382339 598768
rect 379868 598710 382339 598712
rect 382273 598707 382339 598710
rect 458817 596866 458883 596869
rect 491334 596866 491340 596868
rect 458817 596864 491340 596866
rect 458817 596808 458822 596864
rect 458878 596808 491340 596864
rect 458817 596806 491340 596808
rect 458817 596803 458883 596806
rect 491334 596804 491340 596806
rect 491404 596804 491410 596868
rect 459369 594010 459435 594013
rect 474774 594010 474780 594012
rect 459369 594008 474780 594010
rect 459369 593952 459374 594008
rect 459430 593952 474780 594008
rect 459369 593950 474780 593952
rect 459369 593947 459435 593950
rect 474774 593948 474780 593950
rect 474844 593948 474850 594012
rect -960 592908 480 593148
rect 580441 591018 580507 591021
rect 583520 591018 584960 591108
rect 580441 591016 584960 591018
rect 580441 590960 580446 591016
rect 580502 590960 584960 591016
rect 580441 590958 584960 590960
rect 580441 590955 580507 590958
rect 583520 590868 584960 590958
rect 382273 588162 382339 588165
rect 379868 588160 382339 588162
rect 379868 588104 382278 588160
rect 382334 588104 382339 588160
rect 379868 588102 382339 588104
rect 382273 588099 382339 588102
rect -960 580002 480 580092
rect 3601 580002 3667 580005
rect -960 580000 3667 580002
rect -960 579944 3606 580000
rect 3662 579944 3667 580000
rect -960 579942 3667 579944
rect -960 579852 480 579942
rect 3601 579939 3667 579942
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 382273 577554 382339 577557
rect 379868 577552 382339 577554
rect 379868 577496 382278 577552
rect 382334 577496 382339 577552
rect 583520 577540 584960 577630
rect 379868 577494 382339 577496
rect 382273 577491 382339 577494
rect -960 566946 480 567036
rect 3785 566946 3851 566949
rect 382273 566946 382339 566949
rect -960 566944 3851 566946
rect -960 566888 3790 566944
rect 3846 566888 3851 566944
rect -960 566886 3851 566888
rect 379868 566944 382339 566946
rect 379868 566888 382278 566944
rect 382334 566888 382339 566944
rect 379868 566886 382339 566888
rect -960 566796 480 566886
rect 3785 566883 3851 566886
rect 382273 566883 382339 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect 382273 556338 382339 556341
rect 379868 556336 382339 556338
rect 379868 556280 382278 556336
rect 382334 556280 382339 556336
rect 379868 556278 382339 556280
rect 382273 556275 382339 556278
rect -960 553890 480 553980
rect 3969 553890 4035 553893
rect -960 553888 4035 553890
rect -960 553832 3974 553888
rect 4030 553832 4035 553888
rect -960 553830 4035 553832
rect -960 553740 480 553830
rect 3969 553827 4035 553830
rect 583520 551020 584960 551260
rect 382273 545730 382339 545733
rect 379868 545728 382339 545730
rect 379868 545672 382278 545728
rect 382334 545672 382339 545728
rect 379868 545670 382339 545672
rect 382273 545667 382339 545670
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 457846 537372 457852 537436
rect 457916 537434 457922 537436
rect 506473 537434 506539 537437
rect 457916 537432 506539 537434
rect 457916 537376 506478 537432
rect 506534 537376 506539 537432
rect 457916 537374 506539 537376
rect 457916 537372 457922 537374
rect 506473 537371 506539 537374
rect 382273 535122 382339 535125
rect 379868 535120 382339 535122
rect 379868 535064 382278 535120
rect 382334 535064 382339 535120
rect 379868 535062 382339 535064
rect 382273 535059 382339 535062
rect -960 527914 480 528004
rect 3509 527914 3575 527917
rect -960 527912 3575 527914
rect -960 527856 3514 527912
rect 3570 527856 3575 527912
rect -960 527854 3575 527856
rect -960 527764 480 527854
rect 3509 527851 3575 527854
rect 382273 524514 382339 524517
rect 379868 524512 382339 524514
rect 379868 524456 382278 524512
rect 382334 524456 382339 524512
rect 379868 524454 382339 524456
rect 382273 524451 382339 524454
rect 580349 524514 580415 524517
rect 583520 524514 584960 524604
rect 580349 524512 584960 524514
rect 580349 524456 580354 524512
rect 580410 524456 584960 524512
rect 580349 524454 584960 524456
rect 580349 524451 580415 524454
rect 583520 524364 584960 524454
rect 458030 520916 458036 520980
rect 458100 520978 458106 520980
rect 494697 520978 494763 520981
rect 458100 520976 494763 520978
rect 458100 520920 494702 520976
rect 494758 520920 494763 520976
rect 458100 520918 494763 520920
rect 458100 520916 458106 520918
rect 494697 520915 494763 520918
rect 459461 518122 459527 518125
rect 490414 518122 490420 518124
rect 459461 518120 490420 518122
rect 459461 518064 459466 518120
rect 459522 518064 490420 518120
rect 459461 518062 490420 518064
rect 459461 518059 459527 518062
rect 490414 518060 490420 518062
rect 490484 518060 490490 518124
rect 482737 517580 482803 517581
rect 482686 517516 482692 517580
rect 482756 517578 482803 517580
rect 482756 517576 482848 517578
rect 482798 517520 482848 517576
rect 482756 517518 482848 517520
rect 482756 517516 482803 517518
rect 482737 517515 482803 517516
rect 450445 517034 450511 517037
rect 506565 517034 506631 517037
rect 450445 517032 506631 517034
rect 450445 516976 450450 517032
rect 450506 516976 506570 517032
rect 506626 516976 506631 517032
rect 450445 516974 506631 516976
rect 450445 516971 450511 516974
rect 506565 516971 506631 516974
rect 480437 516898 480503 516901
rect 492121 516898 492187 516901
rect 480437 516896 492187 516898
rect 480437 516840 480442 516896
rect 480498 516840 492126 516896
rect 492182 516840 492187 516896
rect 480437 516838 492187 516840
rect 480437 516835 480503 516838
rect 492121 516835 492187 516838
rect 451038 516762 451044 516764
rect 450678 516702 451044 516762
rect 450678 516528 450738 516702
rect 451038 516700 451044 516702
rect 451108 516762 451114 516764
rect 523677 516762 523743 516765
rect 550633 516762 550699 516765
rect 451108 516760 550699 516762
rect 451108 516704 523682 516760
rect 523738 516704 550638 516760
rect 550694 516704 550699 516760
rect 451108 516702 550699 516704
rect 451108 516700 451114 516702
rect 523677 516699 523743 516702
rect 550633 516699 550699 516702
rect 491845 516626 491911 516629
rect 491845 516624 491954 516626
rect 491845 516568 491850 516624
rect 491906 516568 491954 516624
rect 491845 516563 491954 516568
rect 491894 515946 491954 516563
rect 494789 515946 494855 515949
rect 491894 515944 494855 515946
rect 491894 515888 494794 515944
rect 494850 515888 494855 515944
rect 491894 515886 494855 515888
rect 494789 515883 494855 515886
rect -960 514858 480 514948
rect 3693 514858 3759 514861
rect -960 514856 3759 514858
rect -960 514800 3698 514856
rect 3754 514800 3759 514856
rect -960 514798 3759 514800
rect -960 514708 480 514798
rect 3693 514795 3759 514798
rect 450537 514722 450603 514725
rect 450494 514720 450603 514722
rect 450494 514664 450542 514720
rect 450598 514664 450603 514720
rect 450494 514659 450603 514664
rect 450494 514384 450554 514659
rect 450486 514320 450492 514384
rect 450556 514320 450562 514384
rect 382273 513906 382339 513909
rect 379868 513904 382339 513906
rect 379868 513848 382278 513904
rect 382334 513848 382339 513904
rect 379868 513846 382339 513848
rect 382273 513843 382339 513846
rect 494145 512546 494211 512549
rect 491894 512544 494211 512546
rect 491894 512488 494150 512544
rect 494206 512488 494211 512544
rect 491894 512486 494211 512488
rect 491894 512448 491954 512486
rect 494145 512483 494211 512486
rect 449985 512410 450051 512413
rect 450445 512410 450511 512413
rect 449985 512408 450554 512410
rect 449985 512352 449990 512408
rect 450046 512352 450450 512408
rect 450506 512352 450554 512408
rect 449985 512350 450554 512352
rect 449985 512347 450051 512350
rect 450445 512347 450554 512350
rect 450494 512176 450554 512347
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 450077 510234 450143 510237
rect 450353 510234 450419 510237
rect 450077 510232 450419 510234
rect 450077 510176 450082 510232
rect 450138 510176 450358 510232
rect 450414 510176 450419 510232
rect 450077 510174 450419 510176
rect 450077 510171 450143 510174
rect 450310 510171 450419 510174
rect 450310 510000 450370 510171
rect 492121 508942 492187 508945
rect 491924 508940 492187 508942
rect 491924 508884 492126 508940
rect 492182 508884 492187 508940
rect 491924 508882 492187 508884
rect 492121 508879 492187 508882
rect 450310 507653 450370 507824
rect 450261 507648 450370 507653
rect 450261 507592 450266 507648
rect 450322 507592 450370 507648
rect 450261 507590 450370 507592
rect 450261 507587 450327 507590
rect 450126 505477 450186 505648
rect 450126 505472 450235 505477
rect 450126 505416 450174 505472
rect 450230 505416 450235 505472
rect 450126 505414 450235 505416
rect 450169 505411 450235 505414
rect 491894 505202 491954 505376
rect 494145 505202 494211 505205
rect 491894 505200 494211 505202
rect 491894 505144 494150 505200
rect 494206 505144 494211 505200
rect 491894 505142 494211 505144
rect 494145 505139 494211 505142
rect 450494 503301 450554 503472
rect 382273 503298 382339 503301
rect 379868 503296 382339 503298
rect 379868 503240 382278 503296
rect 382334 503240 382339 503296
rect 379868 503238 382339 503240
rect 450494 503296 450603 503301
rect 450494 503240 450542 503296
rect 450598 503240 450603 503296
rect 450494 503238 450603 503240
rect 382273 503235 382339 503238
rect 450537 503235 450603 503238
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 491894 501666 491954 501840
rect 470550 501606 491954 501666
rect 450678 501122 450738 501296
rect 464429 501122 464495 501125
rect 470550 501122 470610 501606
rect 491894 501258 491954 501606
rect 494789 501258 494855 501261
rect 491894 501256 494855 501258
rect 491894 501200 494794 501256
rect 494850 501200 494855 501256
rect 491894 501198 494855 501200
rect 494789 501195 494855 501198
rect 450678 501120 470610 501122
rect 450678 501064 464434 501120
rect 464490 501064 470610 501120
rect 450678 501062 470610 501064
rect 464429 501059 464495 501062
rect 583520 497844 584960 498084
rect 382273 492690 382339 492693
rect 379868 492688 382339 492690
rect 379868 492632 382278 492688
rect 382334 492632 382339 492688
rect 379868 492630 382339 492632
rect 382273 492627 382339 492630
rect -960 488596 480 488836
rect 580533 484666 580599 484669
rect 583520 484666 584960 484756
rect 580533 484664 584960 484666
rect 580533 484608 580538 484664
rect 580594 484608 584960 484664
rect 580533 484606 584960 484608
rect 580533 484603 580599 484606
rect 583520 484516 584960 484606
rect 382273 482082 382339 482085
rect 379868 482080 382339 482082
rect 379868 482024 382278 482080
rect 382334 482024 382339 482080
rect 379868 482022 382339 482024
rect 382273 482019 382339 482022
rect -960 475690 480 475780
rect 3877 475690 3943 475693
rect -960 475688 3943 475690
rect -960 475632 3882 475688
rect 3938 475632 3943 475688
rect -960 475630 3943 475632
rect -960 475540 480 475630
rect 3877 475627 3943 475630
rect 382365 471474 382431 471477
rect 379868 471472 382431 471474
rect 379868 471416 382370 471472
rect 382426 471416 382431 471472
rect 379868 471414 382431 471416
rect 382365 471411 382431 471414
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 516777 467258 516843 467261
rect 542670 467258 542676 467260
rect 516777 467256 542676 467258
rect 516777 467200 516782 467256
rect 516838 467200 542676 467256
rect 516777 467198 542676 467200
rect 516777 467195 516843 467198
rect 542670 467196 542676 467198
rect 542740 467196 542746 467260
rect 478137 467122 478203 467125
rect 482686 467122 482692 467124
rect 478137 467120 482692 467122
rect 478137 467064 478142 467120
rect 478198 467064 482692 467120
rect 478137 467062 482692 467064
rect 478137 467059 478203 467062
rect 482686 467060 482692 467062
rect 482756 467122 482762 467124
rect 521745 467122 521811 467125
rect 482756 467120 521811 467122
rect 482756 467064 521750 467120
rect 521806 467064 521811 467120
rect 482756 467062 521811 467064
rect 482756 467060 482762 467062
rect 521745 467059 521811 467062
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 382273 460866 382339 460869
rect 379868 460864 382339 460866
rect 379868 460808 382278 460864
rect 382334 460808 382339 460864
rect 379868 460806 382339 460808
rect 382273 460803 382339 460806
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 382273 450258 382339 450261
rect 379868 450256 382339 450258
rect 379868 450200 382278 450256
rect 382334 450200 382339 450256
rect 379868 450198 382339 450200
rect 382273 450195 382339 450198
rect -960 449578 480 449668
rect 3785 449578 3851 449581
rect -960 449576 3851 449578
rect -960 449520 3790 449576
rect 3846 449520 3851 449576
rect -960 449518 3851 449520
rect -960 449428 480 449518
rect 3785 449515 3851 449518
rect 561673 444954 561739 444957
rect 559820 444952 561739 444954
rect 559820 444896 561678 444952
rect 561734 444896 561739 444952
rect 559820 444894 561739 444896
rect 561673 444891 561739 444894
rect 583520 444668 584960 444908
rect 383009 439650 383075 439653
rect 379868 439648 383075 439650
rect 379868 439592 383014 439648
rect 383070 439592 383075 439648
rect 379868 439590 383075 439592
rect 383009 439587 383075 439590
rect -960 436508 480 436748
rect 580257 431626 580323 431629
rect 583520 431626 584960 431716
rect 580257 431624 584960 431626
rect 580257 431568 580262 431624
rect 580318 431568 584960 431624
rect 580257 431566 584960 431568
rect 580257 431563 580323 431566
rect 583520 431476 584960 431566
rect 383101 429042 383167 429045
rect 379868 429040 383167 429042
rect 379868 428984 383106 429040
rect 383162 428984 383167 429040
rect 379868 428982 383167 428984
rect 383101 428979 383167 428982
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 383193 418434 383259 418437
rect 379868 418432 383259 418434
rect 379868 418376 383198 418432
rect 383254 418376 383259 418432
rect 379868 418374 383259 418376
rect 383193 418371 383259 418374
rect 580625 418298 580691 418301
rect 583520 418298 584960 418388
rect 580625 418296 584960 418298
rect 580625 418240 580630 418296
rect 580686 418240 584960 418296
rect 580625 418238 584960 418240
rect 580625 418235 580691 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3693 410546 3759 410549
rect -960 410544 3759 410546
rect -960 410488 3698 410544
rect 3754 410488 3759 410544
rect -960 410486 3759 410488
rect -960 410396 480 410486
rect 3693 410483 3759 410486
rect 382273 407826 382339 407829
rect 379868 407824 382339 407826
rect 379868 407768 382278 407824
rect 382334 407768 382339 407824
rect 379868 407766 382339 407768
rect 382273 407763 382339 407766
rect 580441 404970 580507 404973
rect 583520 404970 584960 405060
rect 580441 404968 584960 404970
rect 580441 404912 580446 404968
rect 580502 404912 584960 404968
rect 580441 404910 584960 404912
rect 580441 404907 580507 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 382273 397218 382339 397221
rect 379868 397216 382339 397218
rect 379868 397160 382278 397216
rect 382334 397160 382339 397216
rect 379868 397158 382339 397160
rect 382273 397155 382339 397158
rect 583520 391628 584960 391868
rect 459134 391172 459140 391236
rect 459204 391234 459210 391236
rect 489177 391234 489243 391237
rect 459204 391232 489243 391234
rect 459204 391176 489182 391232
rect 489238 391176 489243 391232
rect 459204 391174 489243 391176
rect 459204 391172 459210 391174
rect 489177 391171 489243 391174
rect 382273 386610 382339 386613
rect 379868 386608 382339 386610
rect 379868 386552 382278 386608
rect 382334 386552 382339 386608
rect 379868 386550 382339 386552
rect 382273 386547 382339 386550
rect -960 384284 480 384524
rect 472014 382332 472020 382396
rect 472084 382394 472090 382396
rect 472801 382394 472867 382397
rect 472084 382392 472867 382394
rect 472084 382336 472806 382392
rect 472862 382336 472867 382392
rect 472084 382334 472867 382336
rect 472084 382332 472090 382334
rect 472801 382331 472867 382334
rect 474774 382332 474780 382396
rect 474844 382394 474850 382396
rect 475377 382394 475443 382397
rect 474844 382392 475443 382394
rect 474844 382336 475382 382392
rect 475438 382336 475443 382392
rect 474844 382334 475443 382336
rect 474844 382332 474850 382334
rect 475377 382331 475443 382334
rect 490414 382332 490420 382396
rect 490484 382394 490490 382396
rect 490833 382394 490899 382397
rect 490484 382392 490899 382394
rect 490484 382336 490838 382392
rect 490894 382336 490899 382392
rect 490484 382334 490899 382336
rect 490484 382332 490490 382334
rect 490833 382331 490899 382334
rect 491334 382332 491340 382396
rect 491404 382394 491410 382396
rect 492121 382394 492187 382397
rect 491404 382392 492187 382394
rect 491404 382336 492126 382392
rect 492182 382336 492187 382392
rect 491404 382334 492187 382336
rect 491404 382332 491410 382334
rect 492121 382331 492187 382334
rect 512821 378722 512887 378725
rect 509956 378720 512887 378722
rect 509956 378664 512826 378720
rect 512882 378664 512887 378720
rect 509956 378662 512887 378664
rect 512821 378659 512887 378662
rect 579613 378450 579679 378453
rect 583520 378450 584960 378540
rect 579613 378448 584960 378450
rect 579613 378392 579618 378448
rect 579674 378392 584960 378448
rect 579613 378390 584960 378392
rect 579613 378387 579679 378390
rect 512729 378314 512795 378317
rect 509956 378312 512795 378314
rect 509956 378256 512734 378312
rect 512790 378256 512795 378312
rect 583520 378300 584960 378390
rect 509956 378254 512795 378256
rect 512729 378251 512795 378254
rect 512913 377906 512979 377909
rect 509956 377904 512979 377906
rect 509956 377848 512918 377904
rect 512974 377848 512979 377904
rect 509956 377846 512979 377848
rect 512913 377843 512979 377846
rect 512637 377498 512703 377501
rect 509956 377496 512703 377498
rect 509956 377440 512642 377496
rect 512698 377440 512703 377496
rect 509956 377438 512703 377440
rect 512637 377435 512703 377438
rect 512269 377090 512335 377093
rect 509956 377088 512335 377090
rect 509956 377032 512274 377088
rect 512330 377032 512335 377088
rect 509956 377030 512335 377032
rect 512269 377027 512335 377030
rect 513281 376682 513347 376685
rect 509956 376680 513347 376682
rect 509956 376624 513286 376680
rect 513342 376624 513347 376680
rect 509956 376622 513347 376624
rect 513281 376619 513347 376622
rect 513189 376274 513255 376277
rect 509956 376272 513255 376274
rect 509956 376216 513194 376272
rect 513250 376216 513255 376272
rect 509956 376214 513255 376216
rect 513189 376211 513255 376214
rect 382273 376002 382339 376005
rect 379868 376000 382339 376002
rect 379868 375944 382278 376000
rect 382334 375944 382339 376000
rect 379868 375942 382339 375944
rect 382273 375939 382339 375942
rect 447133 375866 447199 375869
rect 513097 375866 513163 375869
rect 447133 375864 450156 375866
rect 447133 375808 447138 375864
rect 447194 375808 450156 375864
rect 447133 375806 450156 375808
rect 509956 375864 513163 375866
rect 509956 375808 513102 375864
rect 513158 375808 513163 375864
rect 509956 375806 513163 375808
rect 447133 375803 447199 375806
rect 513097 375803 513163 375806
rect 512269 375458 512335 375461
rect 509956 375456 512335 375458
rect 509956 375400 512274 375456
rect 512330 375400 512335 375456
rect 509956 375398 512335 375400
rect 512269 375395 512335 375398
rect 447133 375322 447199 375325
rect 447133 375320 450156 375322
rect 447133 375264 447138 375320
rect 447194 375264 450156 375320
rect 447133 375262 450156 375264
rect 447133 375259 447199 375262
rect 512085 375050 512151 375053
rect 509956 375048 512151 375050
rect 509956 374992 512090 375048
rect 512146 374992 512151 375048
rect 509956 374990 512151 374992
rect 512085 374987 512151 374990
rect 447225 374778 447291 374781
rect 447225 374776 450156 374778
rect 447225 374720 447230 374776
rect 447286 374720 450156 374776
rect 447225 374718 450156 374720
rect 447225 374715 447291 374718
rect 513281 374642 513347 374645
rect 509956 374640 513347 374642
rect 509956 374584 513286 374640
rect 513342 374584 513347 374640
rect 509956 374582 513347 374584
rect 513281 374579 513347 374582
rect 447317 374234 447383 374237
rect 512821 374234 512887 374237
rect 447317 374232 450156 374234
rect 447317 374176 447322 374232
rect 447378 374176 450156 374232
rect 447317 374174 450156 374176
rect 509956 374232 512887 374234
rect 509956 374176 512826 374232
rect 512882 374176 512887 374232
rect 509956 374174 512887 374176
rect 447317 374171 447383 374174
rect 512821 374171 512887 374174
rect 513281 373826 513347 373829
rect 509956 373824 513347 373826
rect 509956 373768 513286 373824
rect 513342 373768 513347 373824
rect 509956 373766 513347 373768
rect 513281 373763 513347 373766
rect 447133 373690 447199 373693
rect 447133 373688 450156 373690
rect 447133 373632 447138 373688
rect 447194 373632 450156 373688
rect 447133 373630 450156 373632
rect 447133 373627 447199 373630
rect 513281 373418 513347 373421
rect 509956 373416 513347 373418
rect 509956 373360 513286 373416
rect 513342 373360 513347 373416
rect 509956 373358 513347 373360
rect 513281 373355 513347 373358
rect 447225 373146 447291 373149
rect 447225 373144 450156 373146
rect 447225 373088 447230 373144
rect 447286 373088 450156 373144
rect 447225 373086 450156 373088
rect 447225 373083 447291 373086
rect 511993 373010 512059 373013
rect 509956 373008 512059 373010
rect 509956 372952 511998 373008
rect 512054 372952 512059 373008
rect 509956 372950 512059 372952
rect 511993 372947 512059 372950
rect 447133 372602 447199 372605
rect 513281 372602 513347 372605
rect 447133 372600 450156 372602
rect 447133 372544 447138 372600
rect 447194 372544 450156 372600
rect 447133 372542 450156 372544
rect 509956 372600 513347 372602
rect 509956 372544 513286 372600
rect 513342 372544 513347 372600
rect 509956 372542 513347 372544
rect 447133 372539 447199 372542
rect 513281 372539 513347 372542
rect 512729 372194 512795 372197
rect 509956 372192 512795 372194
rect 509956 372136 512734 372192
rect 512790 372136 512795 372192
rect 509956 372134 512795 372136
rect 512729 372131 512795 372134
rect 447317 372058 447383 372061
rect 447317 372056 450156 372058
rect 447317 372000 447322 372056
rect 447378 372000 450156 372056
rect 447317 371998 450156 372000
rect 447317 371995 447383 371998
rect 512453 371786 512519 371789
rect 509956 371784 512519 371786
rect 509956 371728 512458 371784
rect 512514 371728 512519 371784
rect 509956 371726 512519 371728
rect 512453 371723 512519 371726
rect 447225 371514 447291 371517
rect 447225 371512 450156 371514
rect -960 371378 480 371468
rect 447225 371456 447230 371512
rect 447286 371456 450156 371512
rect 447225 371454 450156 371456
rect 447225 371451 447291 371454
rect 3417 371378 3483 371381
rect 513189 371378 513255 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect 509956 371376 513255 371378
rect 509956 371320 513194 371376
rect 513250 371320 513255 371376
rect 509956 371318 513255 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 513189 371315 513255 371318
rect 447133 370970 447199 370973
rect 513281 370970 513347 370973
rect 447133 370968 450156 370970
rect 447133 370912 447138 370968
rect 447194 370912 450156 370968
rect 447133 370910 450156 370912
rect 509956 370968 513347 370970
rect 509956 370912 513286 370968
rect 513342 370912 513347 370968
rect 509956 370910 513347 370912
rect 447133 370907 447199 370910
rect 513281 370907 513347 370910
rect 513189 370562 513255 370565
rect 509956 370560 513255 370562
rect 509956 370504 513194 370560
rect 513250 370504 513255 370560
rect 509956 370502 513255 370504
rect 513189 370499 513255 370502
rect 447225 370426 447291 370429
rect 447225 370424 450156 370426
rect 447225 370368 447230 370424
rect 447286 370368 450156 370424
rect 447225 370366 450156 370368
rect 447225 370363 447291 370366
rect 513097 370154 513163 370157
rect 509956 370152 513163 370154
rect 509956 370096 513102 370152
rect 513158 370096 513163 370152
rect 509956 370094 513163 370096
rect 513097 370091 513163 370094
rect 447317 369882 447383 369885
rect 447317 369880 450156 369882
rect 447317 369824 447322 369880
rect 447378 369824 450156 369880
rect 447317 369822 450156 369824
rect 447317 369819 447383 369822
rect 513097 369746 513163 369749
rect 509956 369744 513163 369746
rect 509956 369688 513102 369744
rect 513158 369688 513163 369744
rect 509956 369686 513163 369688
rect 513097 369683 513163 369686
rect 447133 369338 447199 369341
rect 513281 369338 513347 369341
rect 447133 369336 450156 369338
rect 447133 369280 447138 369336
rect 447194 369280 450156 369336
rect 447133 369278 450156 369280
rect 509956 369336 513347 369338
rect 509956 369280 513286 369336
rect 513342 369280 513347 369336
rect 509956 369278 513347 369280
rect 447133 369275 447199 369278
rect 513281 369275 513347 369278
rect 513281 368930 513347 368933
rect 509956 368928 513347 368930
rect 509956 368872 513286 368928
rect 513342 368872 513347 368928
rect 509956 368870 513347 368872
rect 513281 368867 513347 368870
rect 447225 368794 447291 368797
rect 447225 368792 450156 368794
rect 447225 368736 447230 368792
rect 447286 368736 450156 368792
rect 447225 368734 450156 368736
rect 447225 368731 447291 368734
rect 513189 368522 513255 368525
rect 509956 368520 513255 368522
rect 509956 368464 513194 368520
rect 513250 368464 513255 368520
rect 509956 368462 513255 368464
rect 513189 368459 513255 368462
rect 447133 368250 447199 368253
rect 447133 368248 450156 368250
rect 447133 368192 447138 368248
rect 447194 368192 450156 368248
rect 447133 368190 450156 368192
rect 447133 368187 447199 368190
rect 512177 368114 512243 368117
rect 509956 368112 512243 368114
rect 509956 368056 512182 368112
rect 512238 368056 512243 368112
rect 509956 368054 512243 368056
rect 512177 368051 512243 368054
rect 447225 367706 447291 367709
rect 512269 367706 512335 367709
rect 447225 367704 450156 367706
rect 447225 367648 447230 367704
rect 447286 367648 450156 367704
rect 447225 367646 450156 367648
rect 509956 367704 512335 367706
rect 509956 367648 512274 367704
rect 512330 367648 512335 367704
rect 509956 367646 512335 367648
rect 447225 367643 447291 367646
rect 512269 367643 512335 367646
rect 513281 367298 513347 367301
rect 509956 367296 513347 367298
rect 509956 367240 513286 367296
rect 513342 367240 513347 367296
rect 509956 367238 513347 367240
rect 513281 367235 513347 367238
rect 447317 367162 447383 367165
rect 447317 367160 450156 367162
rect 447317 367104 447322 367160
rect 447378 367104 450156 367160
rect 447317 367102 450156 367104
rect 447317 367099 447383 367102
rect 513005 366890 513071 366893
rect 509956 366888 513071 366890
rect 509956 366832 513010 366888
rect 513066 366832 513071 366888
rect 509956 366830 513071 366832
rect 513005 366827 513071 366830
rect 447133 366618 447199 366621
rect 447133 366616 450156 366618
rect 447133 366560 447138 366616
rect 447194 366560 450156 366616
rect 447133 366558 450156 366560
rect 447133 366555 447199 366558
rect 513189 366482 513255 366485
rect 509956 366480 513255 366482
rect 509956 366424 513194 366480
rect 513250 366424 513255 366480
rect 509956 366422 513255 366424
rect 513189 366419 513255 366422
rect 447225 366074 447291 366077
rect 512821 366074 512887 366077
rect 447225 366072 450156 366074
rect 447225 366016 447230 366072
rect 447286 366016 450156 366072
rect 447225 366014 450156 366016
rect 509956 366072 512887 366074
rect 509956 366016 512826 366072
rect 512882 366016 512887 366072
rect 509956 366014 512887 366016
rect 447225 366011 447291 366014
rect 512821 366011 512887 366014
rect 512913 365666 512979 365669
rect 509956 365664 512979 365666
rect 509956 365608 512918 365664
rect 512974 365608 512979 365664
rect 509956 365606 512979 365608
rect 512913 365603 512979 365606
rect 447133 365530 447199 365533
rect 447133 365528 450156 365530
rect 447133 365472 447138 365528
rect 447194 365472 450156 365528
rect 447133 365470 450156 365472
rect 447133 365467 447199 365470
rect 382641 365394 382707 365397
rect 379868 365392 382707 365394
rect 379868 365336 382646 365392
rect 382702 365336 382707 365392
rect 379868 365334 382707 365336
rect 382641 365331 382707 365334
rect 513189 365258 513255 365261
rect 509956 365256 513255 365258
rect 509956 365200 513194 365256
rect 513250 365200 513255 365256
rect 509956 365198 513255 365200
rect 513189 365195 513255 365198
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 447225 364986 447291 364989
rect 447225 364984 450156 364986
rect 447225 364928 447230 364984
rect 447286 364928 450156 364984
rect 583520 364972 584960 365062
rect 447225 364926 450156 364928
rect 447225 364923 447291 364926
rect 513097 364850 513163 364853
rect 509956 364848 513163 364850
rect 509956 364792 513102 364848
rect 513158 364792 513163 364848
rect 509956 364790 513163 364792
rect 513097 364787 513163 364790
rect 447317 364442 447383 364445
rect 513281 364442 513347 364445
rect 447317 364440 450156 364442
rect 447317 364384 447322 364440
rect 447378 364384 450156 364440
rect 447317 364382 450156 364384
rect 509956 364440 513347 364442
rect 509956 364384 513286 364440
rect 513342 364384 513347 364440
rect 509956 364382 513347 364384
rect 447317 364379 447383 364382
rect 513281 364379 513347 364382
rect 512085 364034 512151 364037
rect 509956 364032 512151 364034
rect 509956 363976 512090 364032
rect 512146 363976 512151 364032
rect 509956 363974 512151 363976
rect 512085 363971 512151 363974
rect 447133 363898 447199 363901
rect 447133 363896 450156 363898
rect 447133 363840 447138 363896
rect 447194 363840 450156 363896
rect 447133 363838 450156 363840
rect 447133 363835 447199 363838
rect 513281 363626 513347 363629
rect 509956 363624 513347 363626
rect 509956 363568 513286 363624
rect 513342 363568 513347 363624
rect 509956 363566 513347 363568
rect 513281 363563 513347 363566
rect 447225 363354 447291 363357
rect 447225 363352 450156 363354
rect 447225 363296 447230 363352
rect 447286 363296 450156 363352
rect 447225 363294 450156 363296
rect 447225 363291 447291 363294
rect 513005 363218 513071 363221
rect 509956 363216 513071 363218
rect 509956 363160 513010 363216
rect 513066 363160 513071 363216
rect 509956 363158 513071 363160
rect 513005 363155 513071 363158
rect 447133 362810 447199 362813
rect 512637 362810 512703 362813
rect 447133 362808 450156 362810
rect 447133 362752 447138 362808
rect 447194 362752 450156 362808
rect 447133 362750 450156 362752
rect 509956 362808 512703 362810
rect 509956 362752 512642 362808
rect 512698 362752 512703 362808
rect 509956 362750 512703 362752
rect 447133 362747 447199 362750
rect 512637 362747 512703 362750
rect 513281 362402 513347 362405
rect 509956 362400 513347 362402
rect 509956 362344 513286 362400
rect 513342 362344 513347 362400
rect 509956 362342 513347 362344
rect 513281 362339 513347 362342
rect 447225 362266 447291 362269
rect 447225 362264 450156 362266
rect 447225 362208 447230 362264
rect 447286 362208 450156 362264
rect 447225 362206 450156 362208
rect 447225 362203 447291 362206
rect 512085 361994 512151 361997
rect 509956 361992 512151 361994
rect 509956 361936 512090 361992
rect 512146 361936 512151 361992
rect 509956 361934 512151 361936
rect 512085 361931 512151 361934
rect 447317 361722 447383 361725
rect 447317 361720 450156 361722
rect 447317 361664 447322 361720
rect 447378 361664 450156 361720
rect 447317 361662 450156 361664
rect 447317 361659 447383 361662
rect 513281 361586 513347 361589
rect 509956 361584 513347 361586
rect 509956 361528 513286 361584
rect 513342 361528 513347 361584
rect 509956 361526 513347 361528
rect 513281 361523 513347 361526
rect 447133 361178 447199 361181
rect 510981 361178 511047 361181
rect 447133 361176 450156 361178
rect 447133 361120 447138 361176
rect 447194 361120 450156 361176
rect 447133 361118 450156 361120
rect 509956 361176 511047 361178
rect 509956 361120 510986 361176
rect 511042 361120 511047 361176
rect 509956 361118 511047 361120
rect 447133 361115 447199 361118
rect 510981 361115 511047 361118
rect 513097 360770 513163 360773
rect 509956 360768 513163 360770
rect 509956 360712 513102 360768
rect 513158 360712 513163 360768
rect 509956 360710 513163 360712
rect 513097 360707 513163 360710
rect 447225 360634 447291 360637
rect 447225 360632 450156 360634
rect 447225 360576 447230 360632
rect 447286 360576 450156 360632
rect 447225 360574 450156 360576
rect 447225 360571 447291 360574
rect 510797 360362 510863 360365
rect 509956 360360 510863 360362
rect 509956 360304 510802 360360
rect 510858 360304 510863 360360
rect 509956 360302 510863 360304
rect 510797 360299 510863 360302
rect 447225 360090 447291 360093
rect 447225 360088 450156 360090
rect 447225 360032 447230 360088
rect 447286 360032 450156 360088
rect 447225 360030 450156 360032
rect 447225 360027 447291 360030
rect 513005 359954 513071 359957
rect 509956 359952 513071 359954
rect 509956 359896 513010 359952
rect 513066 359896 513071 359952
rect 509956 359894 513071 359896
rect 513005 359891 513071 359894
rect 447133 359546 447199 359549
rect 513281 359546 513347 359549
rect 447133 359544 450156 359546
rect 447133 359488 447138 359544
rect 447194 359488 450156 359544
rect 447133 359486 450156 359488
rect 509956 359544 513347 359546
rect 509956 359488 513286 359544
rect 513342 359488 513347 359544
rect 509956 359486 513347 359488
rect 447133 359483 447199 359486
rect 513281 359483 513347 359486
rect 510061 359138 510127 359141
rect 509956 359136 510127 359138
rect 509956 359080 510066 359136
rect 510122 359080 510127 359136
rect 509956 359078 510127 359080
rect 510061 359075 510127 359078
rect 447317 359002 447383 359005
rect 447317 359000 450156 359002
rect 447317 358944 447322 359000
rect 447378 358944 450156 359000
rect 447317 358942 450156 358944
rect 447317 358939 447383 358942
rect 511993 358730 512059 358733
rect 509956 358728 512059 358730
rect 509956 358672 511998 358728
rect 512054 358672 512059 358728
rect 509956 358670 512059 358672
rect 511993 358667 512059 358670
rect -960 358458 480 358548
rect 3601 358458 3667 358461
rect -960 358456 3667 358458
rect -960 358400 3606 358456
rect 3662 358400 3667 358456
rect -960 358398 3667 358400
rect -960 358308 480 358398
rect 3601 358395 3667 358398
rect 447225 358458 447291 358461
rect 447225 358456 450156 358458
rect 447225 358400 447230 358456
rect 447286 358400 450156 358456
rect 447225 358398 450156 358400
rect 447225 358395 447291 358398
rect 513005 358322 513071 358325
rect 509956 358320 513071 358322
rect 509956 358264 513010 358320
rect 513066 358264 513071 358320
rect 509956 358262 513071 358264
rect 513005 358259 513071 358262
rect 447133 357914 447199 357917
rect 512085 357914 512151 357917
rect 447133 357912 450156 357914
rect 447133 357856 447138 357912
rect 447194 357856 450156 357912
rect 447133 357854 450156 357856
rect 509956 357912 512151 357914
rect 509956 357856 512090 357912
rect 512146 357856 512151 357912
rect 509956 357854 512151 357856
rect 447133 357851 447199 357854
rect 512085 357851 512151 357854
rect 513281 357506 513347 357509
rect 509956 357504 513347 357506
rect 509956 357448 513286 357504
rect 513342 357448 513347 357504
rect 509956 357446 513347 357448
rect 513281 357443 513347 357446
rect 447225 357370 447291 357373
rect 447225 357368 450156 357370
rect 447225 357312 447230 357368
rect 447286 357312 450156 357368
rect 447225 357310 450156 357312
rect 447225 357307 447291 357310
rect 512177 357098 512243 357101
rect 509956 357096 512243 357098
rect 509956 357040 512182 357096
rect 512238 357040 512243 357096
rect 509956 357038 512243 357040
rect 512177 357035 512243 357038
rect 447317 356826 447383 356829
rect 447317 356824 450156 356826
rect 447317 356768 447322 356824
rect 447378 356768 450156 356824
rect 447317 356766 450156 356768
rect 447317 356763 447383 356766
rect 512637 356690 512703 356693
rect 509956 356688 512703 356690
rect 509956 356632 512642 356688
rect 512698 356632 512703 356688
rect 509956 356630 512703 356632
rect 512637 356627 512703 356630
rect 447133 356282 447199 356285
rect 512085 356282 512151 356285
rect 447133 356280 450156 356282
rect 447133 356224 447138 356280
rect 447194 356224 450156 356280
rect 447133 356222 450156 356224
rect 509956 356280 512151 356282
rect 509956 356224 512090 356280
rect 512146 356224 512151 356280
rect 509956 356222 512151 356224
rect 447133 356219 447199 356222
rect 512085 356219 512151 356222
rect 511073 355874 511139 355877
rect 509956 355872 511139 355874
rect 509956 355816 511078 355872
rect 511134 355816 511139 355872
rect 509956 355814 511139 355816
rect 511073 355811 511139 355814
rect 449249 355738 449315 355741
rect 449249 355736 450156 355738
rect 449249 355680 449254 355736
rect 449310 355680 450156 355736
rect 449249 355678 450156 355680
rect 449249 355675 449315 355678
rect 512729 355466 512795 355469
rect 509956 355464 512795 355466
rect 509956 355408 512734 355464
rect 512790 355408 512795 355464
rect 509956 355406 512795 355408
rect 512729 355403 512795 355406
rect 448329 355194 448395 355197
rect 448329 355192 450156 355194
rect 448329 355136 448334 355192
rect 448390 355136 450156 355192
rect 448329 355134 450156 355136
rect 448329 355131 448395 355134
rect 513281 355058 513347 355061
rect 509956 355056 513347 355058
rect 509956 355000 513286 355056
rect 513342 355000 513347 355056
rect 509956 354998 513347 355000
rect 513281 354995 513347 354998
rect 382917 354786 382983 354789
rect 379868 354784 382983 354786
rect 379868 354728 382922 354784
rect 382978 354728 382983 354784
rect 379868 354726 382983 354728
rect 382917 354723 382983 354726
rect 449617 354650 449683 354653
rect 513097 354650 513163 354653
rect 449617 354648 450156 354650
rect 449617 354592 449622 354648
rect 449678 354592 450156 354648
rect 449617 354590 450156 354592
rect 509956 354648 513163 354650
rect 509956 354592 513102 354648
rect 513158 354592 513163 354648
rect 509956 354590 513163 354592
rect 449617 354587 449683 354590
rect 513097 354587 513163 354590
rect 512545 354242 512611 354245
rect 509956 354240 512611 354242
rect 509956 354184 512550 354240
rect 512606 354184 512611 354240
rect 509956 354182 512611 354184
rect 512545 354179 512611 354182
rect 449065 354106 449131 354109
rect 449065 354104 450156 354106
rect 449065 354048 449070 354104
rect 449126 354048 450156 354104
rect 449065 354046 450156 354048
rect 449065 354043 449131 354046
rect 512177 353834 512243 353837
rect 509956 353832 512243 353834
rect 509956 353776 512182 353832
rect 512238 353776 512243 353832
rect 509956 353774 512243 353776
rect 512177 353771 512243 353774
rect 447409 353562 447475 353565
rect 447409 353560 450156 353562
rect 447409 353504 447414 353560
rect 447470 353504 450156 353560
rect 447409 353502 450156 353504
rect 447409 353499 447475 353502
rect 513465 353426 513531 353429
rect 509956 353424 513531 353426
rect 509956 353368 513470 353424
rect 513526 353368 513531 353424
rect 509956 353366 513531 353368
rect 513465 353363 513531 353366
rect 447869 353018 447935 353021
rect 513557 353018 513623 353021
rect 447869 353016 450156 353018
rect 447869 352960 447874 353016
rect 447930 352960 450156 353016
rect 447869 352958 450156 352960
rect 509956 353016 513623 353018
rect 509956 352960 513562 353016
rect 513618 352960 513623 353016
rect 509956 352958 513623 352960
rect 447869 352955 447935 352958
rect 513557 352955 513623 352958
rect 513281 352610 513347 352613
rect 509956 352608 513347 352610
rect 509956 352552 513286 352608
rect 513342 352552 513347 352608
rect 509956 352550 513347 352552
rect 513281 352547 513347 352550
rect 449341 352474 449407 352477
rect 449341 352472 450156 352474
rect 449341 352416 449346 352472
rect 449402 352416 450156 352472
rect 449341 352414 450156 352416
rect 449341 352411 449407 352414
rect 512269 352202 512335 352205
rect 509956 352200 512335 352202
rect 509956 352144 512274 352200
rect 512330 352144 512335 352200
rect 509956 352142 512335 352144
rect 512269 352139 512335 352142
rect 449525 351930 449591 351933
rect 580717 351930 580783 351933
rect 583520 351930 584960 352020
rect 449525 351928 450156 351930
rect 449525 351872 449530 351928
rect 449586 351872 450156 351928
rect 449525 351870 450156 351872
rect 580717 351928 584960 351930
rect 580717 351872 580722 351928
rect 580778 351872 584960 351928
rect 580717 351870 584960 351872
rect 449525 351867 449591 351870
rect 580717 351867 580783 351870
rect 512637 351794 512703 351797
rect 509956 351792 512703 351794
rect 509956 351736 512642 351792
rect 512698 351736 512703 351792
rect 583520 351780 584960 351870
rect 509956 351734 512703 351736
rect 512637 351731 512703 351734
rect 449709 351386 449775 351389
rect 513281 351386 513347 351389
rect 449709 351384 450156 351386
rect 449709 351328 449714 351384
rect 449770 351328 450156 351384
rect 449709 351326 450156 351328
rect 509956 351384 513347 351386
rect 509956 351328 513286 351384
rect 513342 351328 513347 351384
rect 509956 351326 513347 351328
rect 449709 351323 449775 351326
rect 513281 351323 513347 351326
rect 512637 350978 512703 350981
rect 509956 350976 512703 350978
rect 509956 350920 512642 350976
rect 512698 350920 512703 350976
rect 509956 350918 512703 350920
rect 512637 350915 512703 350918
rect 449433 350842 449499 350845
rect 449433 350840 450156 350842
rect 449433 350784 449438 350840
rect 449494 350784 450156 350840
rect 449433 350782 450156 350784
rect 449433 350779 449499 350782
rect 513281 350570 513347 350573
rect 509956 350568 513347 350570
rect 509956 350512 513286 350568
rect 513342 350512 513347 350568
rect 509956 350510 513347 350512
rect 513281 350507 513347 350510
rect 447133 350298 447199 350301
rect 447133 350296 450156 350298
rect 447133 350240 447138 350296
rect 447194 350240 450156 350296
rect 447133 350238 450156 350240
rect 447133 350235 447199 350238
rect 512821 350162 512887 350165
rect 509956 350160 512887 350162
rect 509956 350104 512826 350160
rect 512882 350104 512887 350160
rect 509956 350102 512887 350104
rect 512821 350099 512887 350102
rect 447225 349754 447291 349757
rect 513281 349754 513347 349757
rect 447225 349752 450156 349754
rect 447225 349696 447230 349752
rect 447286 349696 450156 349752
rect 447225 349694 450156 349696
rect 509956 349752 513347 349754
rect 509956 349696 513286 349752
rect 513342 349696 513347 349752
rect 509956 349694 513347 349696
rect 447225 349691 447291 349694
rect 513281 349691 513347 349694
rect 512177 349346 512243 349349
rect 509956 349344 512243 349346
rect 509956 349288 512182 349344
rect 512238 349288 512243 349344
rect 509956 349286 512243 349288
rect 512177 349283 512243 349286
rect 447317 349210 447383 349213
rect 447317 349208 450156 349210
rect 447317 349152 447322 349208
rect 447378 349152 450156 349208
rect 447317 349150 450156 349152
rect 447317 349147 447383 349150
rect 513189 348938 513255 348941
rect 509956 348936 513255 348938
rect 509956 348880 513194 348936
rect 513250 348880 513255 348936
rect 509956 348878 513255 348880
rect 513189 348875 513255 348878
rect 447225 348666 447291 348669
rect 447225 348664 450156 348666
rect 447225 348608 447230 348664
rect 447286 348608 450156 348664
rect 447225 348606 450156 348608
rect 447225 348603 447291 348606
rect 513281 348530 513347 348533
rect 509956 348528 513347 348530
rect 509956 348472 513286 348528
rect 513342 348472 513347 348528
rect 509956 348470 513347 348472
rect 513281 348467 513347 348470
rect 447133 348122 447199 348125
rect 510705 348122 510771 348125
rect 447133 348120 450156 348122
rect 447133 348064 447138 348120
rect 447194 348064 450156 348120
rect 447133 348062 450156 348064
rect 509956 348120 510771 348122
rect 509956 348064 510710 348120
rect 510766 348064 510771 348120
rect 509956 348062 510771 348064
rect 447133 348059 447199 348062
rect 510705 348059 510771 348062
rect 513005 347714 513071 347717
rect 509956 347712 513071 347714
rect 509956 347656 513010 347712
rect 513066 347656 513071 347712
rect 509956 347654 513071 347656
rect 513005 347651 513071 347654
rect 447133 347578 447199 347581
rect 447133 347576 450156 347578
rect 447133 347520 447138 347576
rect 447194 347520 450156 347576
rect 447133 347518 450156 347520
rect 447133 347515 447199 347518
rect 512821 347306 512887 347309
rect 509956 347304 512887 347306
rect 509956 347248 512826 347304
rect 512882 347248 512887 347304
rect 509956 347246 512887 347248
rect 512821 347243 512887 347246
rect 447225 347034 447291 347037
rect 447225 347032 450156 347034
rect 447225 346976 447230 347032
rect 447286 346976 450156 347032
rect 447225 346974 450156 346976
rect 447225 346971 447291 346974
rect 512177 346898 512243 346901
rect 509956 346896 512243 346898
rect 509956 346840 512182 346896
rect 512238 346840 512243 346896
rect 509956 346838 512243 346840
rect 512177 346835 512243 346838
rect 447317 346490 447383 346493
rect 512453 346490 512519 346493
rect 447317 346488 450156 346490
rect 447317 346432 447322 346488
rect 447378 346432 450156 346488
rect 447317 346430 450156 346432
rect 509956 346488 512519 346490
rect 509956 346432 512458 346488
rect 512514 346432 512519 346488
rect 509956 346430 512519 346432
rect 447317 346427 447383 346430
rect 512453 346427 512519 346430
rect 513189 346082 513255 346085
rect 509956 346080 513255 346082
rect 509956 346024 513194 346080
rect 513250 346024 513255 346080
rect 509956 346022 513255 346024
rect 513189 346019 513255 346022
rect 448329 345946 448395 345949
rect 448329 345944 450156 345946
rect 448329 345888 448334 345944
rect 448390 345888 450156 345944
rect 448329 345886 450156 345888
rect 448329 345883 448395 345886
rect 510889 345674 510955 345677
rect 509956 345672 510955 345674
rect 509956 345616 510894 345672
rect 510950 345616 510955 345672
rect 509956 345614 510955 345616
rect 510889 345611 510955 345614
rect -960 345402 480 345492
rect 3693 345402 3759 345405
rect -960 345400 3759 345402
rect -960 345344 3698 345400
rect 3754 345344 3759 345400
rect -960 345342 3759 345344
rect -960 345252 480 345342
rect 3693 345339 3759 345342
rect 447133 345402 447199 345405
rect 447133 345400 450156 345402
rect 447133 345344 447138 345400
rect 447194 345344 450156 345400
rect 447133 345342 450156 345344
rect 447133 345339 447199 345342
rect 513281 345266 513347 345269
rect 509956 345264 513347 345266
rect 509956 345208 513286 345264
rect 513342 345208 513347 345264
rect 509956 345206 513347 345208
rect 513281 345203 513347 345206
rect 449709 344858 449775 344861
rect 513281 344858 513347 344861
rect 449709 344856 450156 344858
rect 449709 344800 449714 344856
rect 449770 344800 450156 344856
rect 449709 344798 450156 344800
rect 509956 344856 513347 344858
rect 509956 344800 513286 344856
rect 513342 344800 513347 344856
rect 509956 344798 513347 344800
rect 449709 344795 449775 344798
rect 513281 344795 513347 344798
rect 512269 344450 512335 344453
rect 509956 344448 512335 344450
rect 509956 344392 512274 344448
rect 512330 344392 512335 344448
rect 509956 344390 512335 344392
rect 512269 344387 512335 344390
rect 447961 344314 448027 344317
rect 447961 344312 450156 344314
rect 447961 344256 447966 344312
rect 448022 344256 450156 344312
rect 447961 344254 450156 344256
rect 447961 344251 448027 344254
rect 382273 344178 382339 344181
rect 379868 344176 382339 344178
rect 379868 344120 382278 344176
rect 382334 344120 382339 344176
rect 379868 344118 382339 344120
rect 382273 344115 382339 344118
rect 512821 344042 512887 344045
rect 509956 344040 512887 344042
rect 509956 343984 512826 344040
rect 512882 343984 512887 344040
rect 509956 343982 512887 343984
rect 512821 343979 512887 343982
rect 448053 343770 448119 343773
rect 448053 343768 450156 343770
rect 448053 343712 448058 343768
rect 448114 343712 450156 343768
rect 448053 343710 450156 343712
rect 448053 343707 448119 343710
rect 513281 343634 513347 343637
rect 509956 343632 513347 343634
rect 509956 343576 513286 343632
rect 513342 343576 513347 343632
rect 509956 343574 513347 343576
rect 513281 343571 513347 343574
rect 449801 343226 449867 343229
rect 512361 343226 512427 343229
rect 449801 343224 450156 343226
rect 449801 343168 449806 343224
rect 449862 343168 450156 343224
rect 449801 343166 450156 343168
rect 509956 343224 512427 343226
rect 509956 343168 512366 343224
rect 512422 343168 512427 343224
rect 509956 343166 512427 343168
rect 449801 343163 449867 343166
rect 512361 343163 512427 343166
rect 512361 342818 512427 342821
rect 509956 342816 512427 342818
rect 509956 342760 512366 342816
rect 512422 342760 512427 342816
rect 509956 342758 512427 342760
rect 512361 342755 512427 342758
rect 447133 342682 447199 342685
rect 447133 342680 450156 342682
rect 447133 342624 447138 342680
rect 447194 342624 450156 342680
rect 447133 342622 450156 342624
rect 447133 342619 447199 342622
rect 510613 342410 510679 342413
rect 509956 342408 510679 342410
rect 509956 342352 510618 342408
rect 510674 342352 510679 342408
rect 509956 342350 510679 342352
rect 510613 342347 510679 342350
rect 447593 342138 447659 342141
rect 447593 342136 450156 342138
rect 447593 342080 447598 342136
rect 447654 342080 450156 342136
rect 447593 342078 450156 342080
rect 447593 342075 447659 342078
rect 512269 342002 512335 342005
rect 509956 342000 512335 342002
rect 509956 341944 512274 342000
rect 512330 341944 512335 342000
rect 509956 341942 512335 341944
rect 512269 341939 512335 341942
rect 448145 341594 448211 341597
rect 513281 341594 513347 341597
rect 448145 341592 450156 341594
rect 448145 341536 448150 341592
rect 448206 341536 450156 341592
rect 448145 341534 450156 341536
rect 509956 341592 513347 341594
rect 509956 341536 513286 341592
rect 513342 341536 513347 341592
rect 509956 341534 513347 341536
rect 448145 341531 448211 341534
rect 513281 341531 513347 341534
rect 512269 341186 512335 341189
rect 509956 341184 512335 341186
rect 509956 341128 512274 341184
rect 512330 341128 512335 341184
rect 509956 341126 512335 341128
rect 512269 341123 512335 341126
rect 448053 341050 448119 341053
rect 448053 341048 450156 341050
rect 448053 340992 448058 341048
rect 448114 340992 450156 341048
rect 448053 340990 450156 340992
rect 448053 340987 448119 340990
rect 512361 340778 512427 340781
rect 509956 340776 512427 340778
rect 509956 340720 512366 340776
rect 512422 340720 512427 340776
rect 509956 340718 512427 340720
rect 512361 340715 512427 340718
rect 447869 340506 447935 340509
rect 447869 340504 450156 340506
rect 447869 340448 447874 340504
rect 447930 340448 450156 340504
rect 447869 340446 450156 340448
rect 447869 340443 447935 340446
rect 513005 340370 513071 340373
rect 509956 340368 513071 340370
rect 509956 340312 513010 340368
rect 513066 340312 513071 340368
rect 509956 340310 513071 340312
rect 513005 340307 513071 340310
rect 449801 339962 449867 339965
rect 513281 339962 513347 339965
rect 449801 339960 450156 339962
rect 449801 339904 449806 339960
rect 449862 339904 450156 339960
rect 449801 339902 450156 339904
rect 509956 339960 513347 339962
rect 509956 339904 513286 339960
rect 513342 339904 513347 339960
rect 509956 339902 513347 339904
rect 449801 339899 449867 339902
rect 513281 339899 513347 339902
rect 512361 339554 512427 339557
rect 509956 339552 512427 339554
rect 509956 339496 512366 339552
rect 512422 339496 512427 339552
rect 509956 339494 512427 339496
rect 512361 339491 512427 339494
rect 450126 339149 450186 339388
rect 450077 339144 450186 339149
rect 513281 339146 513347 339149
rect 450077 339088 450082 339144
rect 450138 339088 450186 339144
rect 450077 339086 450186 339088
rect 509956 339144 513347 339146
rect 509956 339088 513286 339144
rect 513342 339088 513347 339144
rect 509956 339086 513347 339088
rect 450077 339083 450143 339086
rect 513281 339083 513347 339086
rect 513189 338738 513255 338741
rect 509956 338736 513255 338738
rect 509956 338680 513194 338736
rect 513250 338680 513255 338736
rect 509956 338678 513255 338680
rect 513189 338675 513255 338678
rect 583520 338452 584960 338692
rect 447133 338330 447199 338333
rect 512545 338330 512611 338333
rect 447133 338328 450156 338330
rect 447133 338272 447138 338328
rect 447194 338272 450156 338328
rect 447133 338270 450156 338272
rect 509956 338328 512611 338330
rect 509956 338272 512550 338328
rect 512606 338272 512611 338328
rect 509956 338270 512611 338272
rect 447133 338267 447199 338270
rect 512545 338267 512611 338270
rect 447685 338058 447751 338061
rect 450261 338058 450327 338061
rect 447685 338056 450327 338058
rect 447685 338000 447690 338056
rect 447746 338000 450266 338056
rect 450322 338000 450327 338056
rect 447685 337998 450327 338000
rect 447685 337995 447751 337998
rect 450261 337995 450327 337998
rect 513005 337922 513071 337925
rect 509956 337920 513071 337922
rect 509956 337864 513010 337920
rect 513066 337864 513071 337920
rect 509956 337862 513071 337864
rect 513005 337859 513071 337862
rect 447225 337786 447291 337789
rect 447225 337784 450156 337786
rect 447225 337728 447230 337784
rect 447286 337728 450156 337784
rect 447225 337726 450156 337728
rect 447225 337723 447291 337726
rect 512913 337514 512979 337517
rect 509956 337512 512979 337514
rect 509956 337456 512918 337512
rect 512974 337456 512979 337512
rect 509956 337454 512979 337456
rect 512913 337451 512979 337454
rect 447133 337242 447199 337245
rect 447133 337240 450156 337242
rect 447133 337184 447138 337240
rect 447194 337184 450156 337240
rect 447133 337182 450156 337184
rect 447133 337179 447199 337182
rect 511165 337106 511231 337109
rect 509956 337104 511231 337106
rect 509956 337048 511170 337104
rect 511226 337048 511231 337104
rect 509956 337046 511231 337048
rect 511165 337043 511231 337046
rect 422201 336834 422267 336837
rect 422886 336834 422892 336836
rect 422201 336832 422892 336834
rect 422201 336776 422206 336832
rect 422262 336776 422892 336832
rect 422201 336774 422892 336776
rect 422201 336771 422267 336774
rect 422886 336772 422892 336774
rect 422956 336834 422962 336836
rect 447685 336834 447751 336837
rect 422956 336832 447751 336834
rect 422956 336776 447690 336832
rect 447746 336776 447751 336832
rect 422956 336774 447751 336776
rect 422956 336772 422962 336774
rect 447685 336771 447751 336774
rect 447225 336698 447291 336701
rect 513281 336698 513347 336701
rect 447225 336696 450156 336698
rect 447225 336640 447230 336696
rect 447286 336640 450156 336696
rect 447225 336638 450156 336640
rect 509956 336696 513347 336698
rect 509956 336640 513286 336696
rect 513342 336640 513347 336696
rect 509956 336638 513347 336640
rect 447225 336635 447291 336638
rect 513281 336635 513347 336638
rect 513189 336290 513255 336293
rect 509956 336288 513255 336290
rect 509956 336232 513194 336288
rect 513250 336232 513255 336288
rect 509956 336230 513255 336232
rect 513189 336227 513255 336230
rect 447133 336154 447199 336157
rect 447133 336152 450156 336154
rect 447133 336096 447138 336152
rect 447194 336096 450156 336152
rect 447133 336094 450156 336096
rect 447133 336091 447199 336094
rect 511533 335882 511599 335885
rect 509956 335880 511599 335882
rect 509956 335824 511538 335880
rect 511594 335824 511599 335880
rect 509956 335822 511599 335824
rect 511533 335819 511599 335822
rect 447317 335610 447383 335613
rect 447317 335608 450156 335610
rect 447317 335552 447322 335608
rect 447378 335552 450156 335608
rect 447317 335550 450156 335552
rect 447317 335547 447383 335550
rect 512729 335474 512795 335477
rect 509956 335472 512795 335474
rect 509956 335416 512734 335472
rect 512790 335416 512795 335472
rect 509956 335414 512795 335416
rect 512729 335411 512795 335414
rect 447225 335066 447291 335069
rect 512821 335066 512887 335069
rect 447225 335064 450156 335066
rect 447225 335008 447230 335064
rect 447286 335008 450156 335064
rect 447225 335006 450156 335008
rect 509956 335064 512887 335066
rect 509956 335008 512826 335064
rect 512882 335008 512887 335064
rect 509956 335006 512887 335008
rect 447225 335003 447291 335006
rect 512821 335003 512887 335006
rect 433977 334794 434043 334797
rect 431940 334792 434043 334794
rect 431940 334736 433982 334792
rect 434038 334736 434043 334792
rect 431940 334734 434043 334736
rect 433977 334731 434043 334734
rect 513005 334658 513071 334661
rect 509956 334656 513071 334658
rect 509956 334600 513010 334656
rect 513066 334600 513071 334656
rect 509956 334598 513071 334600
rect 513005 334595 513071 334598
rect 447133 334522 447199 334525
rect 447133 334520 450156 334522
rect 447133 334464 447138 334520
rect 447194 334464 450156 334520
rect 447133 334462 450156 334464
rect 447133 334459 447199 334462
rect 512637 334250 512703 334253
rect 509956 334248 512703 334250
rect 509956 334192 512642 334248
rect 512698 334192 512703 334248
rect 509956 334190 512703 334192
rect 512637 334187 512703 334190
rect 447225 333978 447291 333981
rect 447225 333976 450156 333978
rect 447225 333920 447230 333976
rect 447286 333920 450156 333976
rect 447225 333918 450156 333920
rect 447225 333915 447291 333918
rect 512913 333842 512979 333845
rect 509956 333840 512979 333842
rect 509956 333784 512918 333840
rect 512974 333784 512979 333840
rect 509956 333782 512979 333784
rect 512913 333779 512979 333782
rect 383101 333570 383167 333573
rect 379868 333568 383167 333570
rect 379868 333512 383106 333568
rect 383162 333512 383167 333568
rect 379868 333510 383167 333512
rect 383101 333507 383167 333510
rect 447133 333434 447199 333437
rect 518198 333434 518204 333436
rect 447133 333432 450156 333434
rect 447133 333376 447138 333432
rect 447194 333376 450156 333432
rect 447133 333374 450156 333376
rect 509956 333374 518204 333434
rect 447133 333371 447199 333374
rect 518198 333372 518204 333374
rect 518268 333372 518274 333436
rect 512821 333026 512887 333029
rect 509956 333024 512887 333026
rect 509956 332968 512826 333024
rect 512882 332968 512887 333024
rect 509956 332966 512887 332968
rect 512821 332963 512887 332966
rect 447317 332890 447383 332893
rect 447317 332888 450156 332890
rect 447317 332832 447322 332888
rect 447378 332832 450156 332888
rect 447317 332830 450156 332832
rect 447317 332827 447383 332830
rect 513281 332618 513347 332621
rect 509956 332616 513347 332618
rect 509956 332560 513286 332616
rect 513342 332560 513347 332616
rect 509956 332558 513347 332560
rect 513281 332555 513347 332558
rect -960 332196 480 332436
rect 447409 332346 447475 332349
rect 447409 332344 450156 332346
rect 447409 332288 447414 332344
rect 447470 332288 450156 332344
rect 447409 332286 450156 332288
rect 447409 332283 447475 332286
rect 512821 332210 512887 332213
rect 509956 332208 512887 332210
rect 509956 332152 512826 332208
rect 512882 332152 512887 332208
rect 509956 332150 512887 332152
rect 512821 332147 512887 332150
rect 447133 331802 447199 331805
rect 512729 331802 512795 331805
rect 447133 331800 450156 331802
rect 447133 331744 447138 331800
rect 447194 331744 450156 331800
rect 447133 331742 450156 331744
rect 509956 331800 512795 331802
rect 509956 331744 512734 331800
rect 512790 331744 512795 331800
rect 509956 331742 512795 331744
rect 447133 331739 447199 331742
rect 512729 331739 512795 331742
rect 513281 331394 513347 331397
rect 509956 331392 513347 331394
rect 509956 331336 513286 331392
rect 513342 331336 513347 331392
rect 509956 331334 513347 331336
rect 513281 331331 513347 331334
rect 447225 331258 447291 331261
rect 447225 331256 450156 331258
rect 447225 331200 447230 331256
rect 447286 331200 450156 331256
rect 447225 331198 450156 331200
rect 447225 331195 447291 331198
rect 510654 330986 510660 330988
rect 509956 330926 510660 330986
rect 510654 330924 510660 330926
rect 510724 330924 510730 330988
rect 433425 330850 433491 330853
rect 431940 330848 433491 330850
rect 431940 330792 433430 330848
rect 433486 330792 433491 330848
rect 431940 330790 433491 330792
rect 433425 330787 433491 330790
rect 448145 330714 448211 330717
rect 448145 330712 450156 330714
rect 448145 330656 448150 330712
rect 448206 330656 450156 330712
rect 448145 330654 450156 330656
rect 448145 330651 448211 330654
rect 512453 330578 512519 330581
rect 509956 330576 512519 330578
rect 509956 330520 512458 330576
rect 512514 330520 512519 330576
rect 509956 330518 512519 330520
rect 512453 330515 512519 330518
rect 447501 330170 447567 330173
rect 517830 330170 517836 330172
rect 447501 330168 450156 330170
rect 447501 330112 447506 330168
rect 447562 330112 450156 330168
rect 447501 330110 450156 330112
rect 509956 330110 517836 330170
rect 447501 330107 447567 330110
rect 517830 330108 517836 330110
rect 517900 330108 517906 330172
rect 447961 329762 448027 329765
rect 448237 329762 448303 329765
rect 512545 329762 512611 329765
rect 447961 329760 448303 329762
rect 447961 329704 447966 329760
rect 448022 329704 448242 329760
rect 448298 329704 448303 329760
rect 447961 329702 448303 329704
rect 509956 329760 512611 329762
rect 509956 329704 512550 329760
rect 512606 329704 512611 329760
rect 509956 329702 512611 329704
rect 447961 329699 448027 329702
rect 448237 329699 448303 329702
rect 512545 329699 512611 329702
rect 448237 329628 448303 329629
rect 448237 329626 448284 329628
rect 448156 329624 448284 329626
rect 448348 329626 448354 329628
rect 448156 329568 448242 329624
rect 448156 329566 448284 329568
rect 448237 329564 448284 329566
rect 448348 329566 450156 329626
rect 448348 329564 448354 329566
rect 448237 329563 448303 329564
rect 513281 329354 513347 329357
rect 509956 329352 513347 329354
rect 509956 329296 513286 329352
rect 513342 329296 513347 329352
rect 509956 329294 513347 329296
rect 513281 329291 513347 329294
rect 447961 329082 448027 329085
rect 447961 329080 450156 329082
rect 447961 329024 447966 329080
rect 448022 329024 450156 329080
rect 447961 329022 450156 329024
rect 447961 329019 448027 329022
rect 512545 328946 512611 328949
rect 509956 328944 512611 328946
rect 509956 328888 512550 328944
rect 512606 328888 512611 328944
rect 509956 328886 512611 328888
rect 512545 328883 512611 328886
rect 448237 328538 448303 328541
rect 514886 328538 514892 328540
rect 448237 328536 450156 328538
rect 448237 328480 448242 328536
rect 448298 328480 450156 328536
rect 448237 328478 450156 328480
rect 509956 328478 514892 328538
rect 448237 328475 448303 328478
rect 514886 328476 514892 328478
rect 514956 328476 514962 328540
rect 450624 328266 450630 328268
rect 450126 328206 450630 328266
rect 448513 327994 448579 327997
rect 450126 327994 450186 328206
rect 450624 328204 450630 328206
rect 450694 328204 450700 328268
rect 513281 328130 513347 328133
rect 509956 328128 513347 328130
rect 509956 328072 513286 328128
rect 513342 328072 513347 328128
rect 509956 328070 513347 328072
rect 513281 328067 513347 328070
rect 448513 327992 450186 327994
rect 448513 327936 448518 327992
rect 448574 327964 450186 327992
rect 448574 327936 450156 327964
rect 448513 327934 450156 327936
rect 448513 327931 448579 327934
rect 450486 327722 450492 327724
rect 450310 327662 450492 327722
rect 450310 327450 450370 327662
rect 450486 327660 450492 327662
rect 450556 327660 450562 327724
rect 510153 327722 510219 327725
rect 509956 327720 510219 327722
rect 509956 327664 510158 327720
rect 510214 327664 510219 327720
rect 509956 327662 510219 327664
rect 510153 327659 510219 327662
rect 450156 327420 450370 327450
rect 450126 327390 450340 327420
rect 449985 327178 450051 327181
rect 450126 327178 450186 327390
rect 510337 327314 510403 327317
rect 509956 327312 510403 327314
rect 509956 327256 510342 327312
rect 510398 327256 510403 327312
rect 509956 327254 510403 327256
rect 510337 327251 510403 327254
rect 449985 327176 450186 327178
rect 449985 327120 449990 327176
rect 450046 327120 450186 327176
rect 449985 327118 450186 327120
rect 449985 327115 450051 327118
rect 434437 326906 434503 326909
rect 510429 326906 510495 326909
rect 431940 326904 434503 326906
rect 431940 326848 434442 326904
rect 434498 326848 434503 326904
rect 509956 326904 510495 326906
rect 431940 326846 434503 326848
rect 434437 326843 434503 326846
rect 449893 326634 449959 326637
rect 450126 326634 450186 326876
rect 509956 326848 510434 326904
rect 510490 326848 510495 326904
rect 509956 326846 510495 326848
rect 510429 326843 510495 326846
rect 450353 326634 450419 326637
rect 449893 326632 450419 326634
rect 449893 326576 449898 326632
rect 449954 326576 450358 326632
rect 450414 326576 450419 326632
rect 449893 326574 450419 326576
rect 449893 326571 449959 326574
rect 450353 326571 450419 326574
rect 511901 326498 511967 326501
rect 509956 326496 511967 326498
rect 509956 326440 511906 326496
rect 511962 326440 511967 326496
rect 509956 326438 511967 326440
rect 511901 326435 511967 326438
rect 450494 326093 450554 326332
rect 450261 326090 450327 326093
rect 450261 326088 450370 326090
rect 450261 326032 450266 326088
rect 450322 326032 450370 326088
rect 450261 326027 450370 326032
rect 450494 326088 450603 326093
rect 510245 326090 510311 326093
rect 450494 326032 450542 326088
rect 450598 326032 450603 326088
rect 450494 326030 450603 326032
rect 509956 326088 510311 326090
rect 509956 326032 510250 326088
rect 510306 326032 510311 326088
rect 509956 326030 510311 326032
rect 450537 326027 450603 326030
rect 510245 326027 510311 326030
rect 450310 325788 450370 326027
rect 509956 325622 511090 325682
rect 450169 325546 450235 325549
rect 450629 325546 450695 325549
rect 450126 325544 450695 325546
rect 450126 325488 450174 325544
rect 450230 325488 450634 325544
rect 450690 325488 450695 325544
rect 450126 325486 450695 325488
rect 511030 325546 511090 325622
rect 512637 325546 512703 325549
rect 511030 325544 512703 325546
rect 511030 325488 512642 325544
rect 512698 325488 512703 325544
rect 511030 325486 512703 325488
rect 450126 325483 450235 325486
rect 450629 325483 450695 325486
rect 512637 325483 512703 325486
rect 450126 325244 450186 325483
rect 510286 325274 510292 325276
rect 509956 325214 510292 325274
rect 510286 325212 510292 325214
rect 510356 325212 510362 325276
rect 579981 325274 580047 325277
rect 583520 325274 584960 325364
rect 579981 325272 584960 325274
rect 579981 325216 579986 325272
rect 580042 325216 584960 325272
rect 579981 325214 584960 325216
rect 579981 325211 580047 325214
rect 583520 325124 584960 325214
rect 450077 325002 450143 325005
rect 450629 325002 450695 325005
rect 450077 325000 450695 325002
rect 450077 324944 450082 325000
rect 450138 324944 450634 325000
rect 450690 324944 450695 325000
rect 450077 324942 450695 324944
rect 450077 324939 450186 324942
rect 450629 324939 450695 324942
rect 450126 324700 450186 324939
rect 510061 324866 510127 324869
rect 509956 324864 510127 324866
rect 509956 324808 510066 324864
rect 510122 324808 510127 324864
rect 509956 324806 510127 324808
rect 510061 324803 510127 324806
rect 515070 324458 515076 324460
rect 509956 324398 515076 324458
rect 515070 324396 515076 324398
rect 515140 324396 515146 324460
rect 449617 324186 449683 324189
rect 449617 324184 450340 324186
rect 449617 324128 449622 324184
rect 449678 324156 450340 324184
rect 449678 324128 450370 324156
rect 449617 324126 450370 324128
rect 449617 324123 449683 324126
rect 450310 323914 450370 324126
rect 514150 324050 514156 324052
rect 509956 323990 514156 324050
rect 514150 323988 514156 323990
rect 514220 323988 514226 324052
rect 450445 323914 450511 323917
rect 450310 323912 450511 323914
rect 450310 323856 450450 323912
rect 450506 323856 450511 323912
rect 450310 323854 450511 323856
rect 450445 323851 450511 323854
rect 510838 323642 510844 323644
rect 509956 323582 510844 323642
rect 510838 323580 510844 323582
rect 510908 323580 510914 323644
rect 518014 323234 518020 323236
rect 509956 323174 518020 323234
rect 518014 323172 518020 323174
rect 518084 323172 518090 323236
rect 383009 322962 383075 322965
rect 434069 322962 434135 322965
rect 379868 322960 383075 322962
rect 379868 322904 383014 322960
rect 383070 322904 383075 322960
rect 379868 322902 383075 322904
rect 431940 322960 434135 322962
rect 431940 322904 434074 322960
rect 434130 322904 434135 322960
rect 431940 322902 434135 322904
rect 383009 322899 383075 322902
rect 434069 322899 434135 322902
rect 512821 322826 512887 322829
rect 509956 322824 512887 322826
rect 509956 322768 512826 322824
rect 512882 322768 512887 322824
rect 509956 322766 512887 322768
rect 512821 322763 512887 322766
rect 514702 322418 514708 322420
rect 509956 322358 514708 322418
rect 514702 322356 514708 322358
rect 514772 322356 514778 322420
rect 511022 322010 511028 322012
rect 509956 321950 511028 322010
rect 511022 321948 511028 321950
rect 511092 321948 511098 322012
rect 511206 321602 511212 321604
rect 509956 321542 511212 321602
rect 511206 321540 511212 321542
rect 511276 321540 511282 321604
rect 489870 320998 502350 321058
rect 463734 320316 463740 320380
rect 463804 320378 463810 320380
rect 464429 320378 464495 320381
rect 463804 320376 464495 320378
rect 463804 320320 464434 320376
rect 464490 320320 464495 320376
rect 463804 320318 464495 320320
rect 463804 320316 463810 320318
rect 464429 320315 464495 320318
rect 454534 320180 454540 320244
rect 454604 320242 454610 320244
rect 489870 320242 489930 320998
rect 502290 320786 502350 320998
rect 509558 320786 509618 321164
rect 502290 320726 509618 320786
rect 507158 320588 507164 320652
rect 507228 320650 507234 320652
rect 510429 320650 510495 320653
rect 507228 320648 510495 320650
rect 507228 320592 510434 320648
rect 510490 320592 510495 320648
rect 507228 320590 510495 320592
rect 507228 320588 507234 320590
rect 510429 320587 510495 320590
rect 507342 320452 507348 320516
rect 507412 320514 507418 320516
rect 511073 320514 511139 320517
rect 507412 320512 511139 320514
rect 507412 320456 511078 320512
rect 511134 320456 511139 320512
rect 507412 320454 511139 320456
rect 507412 320452 507418 320454
rect 511073 320451 511139 320454
rect 506974 320316 506980 320380
rect 507044 320378 507050 320380
rect 510981 320378 511047 320381
rect 507044 320376 511047 320378
rect 507044 320320 510986 320376
rect 511042 320320 511047 320376
rect 507044 320318 511047 320320
rect 507044 320316 507050 320318
rect 510981 320315 511047 320318
rect 454604 320182 489930 320242
rect 510061 320242 510127 320245
rect 510470 320242 510476 320244
rect 510061 320240 510476 320242
rect 510061 320184 510066 320240
rect 510122 320184 510476 320240
rect 510061 320182 510476 320184
rect 454604 320180 454610 320182
rect 510061 320179 510127 320182
rect 510470 320180 510476 320182
rect 510540 320180 510546 320244
rect 460013 320106 460079 320109
rect 558862 320106 558868 320108
rect 460013 320104 558868 320106
rect 460013 320048 460018 320104
rect 460074 320048 558868 320104
rect 460013 320046 558868 320048
rect 460013 320043 460079 320046
rect 558862 320044 558868 320046
rect 558932 320044 558938 320108
rect 447726 319908 447732 319972
rect 447796 319970 447802 319972
rect 462129 319970 462195 319973
rect 447796 319968 462195 319970
rect 447796 319912 462134 319968
rect 462190 319912 462195 319968
rect 447796 319910 462195 319912
rect 447796 319908 447802 319910
rect 462129 319907 462195 319910
rect 508497 319970 508563 319973
rect 511717 319970 511783 319973
rect 508497 319968 511783 319970
rect 508497 319912 508502 319968
rect 508558 319912 511722 319968
rect 511778 319912 511783 319968
rect 508497 319910 511783 319912
rect 508497 319907 508563 319910
rect 511717 319907 511783 319910
rect 447910 319772 447916 319836
rect 447980 319834 447986 319836
rect 461117 319834 461183 319837
rect 447980 319832 461183 319834
rect 447980 319776 461122 319832
rect 461178 319776 461183 319832
rect 447980 319774 461183 319776
rect 447980 319772 447986 319774
rect 461117 319771 461183 319774
rect 444230 319636 444236 319700
rect 444300 319698 444306 319700
rect 444300 319638 447150 319698
rect 444300 319636 444306 319638
rect 447090 319562 447150 319638
rect 461945 319562 462011 319565
rect 447090 319560 462011 319562
rect 447090 319504 461950 319560
rect 462006 319504 462011 319560
rect 447090 319502 462011 319504
rect 461945 319499 462011 319502
rect -960 319290 480 319380
rect 3969 319290 4035 319293
rect -960 319288 4035 319290
rect -960 319232 3974 319288
rect 4030 319232 4035 319288
rect -960 319230 4035 319232
rect -960 319140 480 319230
rect 3969 319227 4035 319230
rect 433517 319018 433583 319021
rect 431940 319016 433583 319018
rect 431940 318960 433522 319016
rect 433578 318960 433583 319016
rect 431940 318958 433583 318960
rect 433517 318955 433583 318958
rect 445385 318746 445451 318749
rect 483197 318746 483263 318749
rect 445385 318744 483263 318746
rect 445385 318688 445390 318744
rect 445446 318688 483202 318744
rect 483258 318688 483263 318744
rect 445385 318686 483263 318688
rect 445385 318683 445451 318686
rect 483197 318683 483263 318686
rect 446949 318610 447015 318613
rect 483473 318610 483539 318613
rect 446949 318608 483539 318610
rect 446949 318552 446954 318608
rect 447010 318552 483478 318608
rect 483534 318552 483539 318608
rect 446949 318550 483539 318552
rect 446949 318547 447015 318550
rect 483473 318547 483539 318550
rect 448094 318412 448100 318476
rect 448164 318474 448170 318476
rect 482369 318474 482435 318477
rect 448164 318472 482435 318474
rect 448164 318416 482374 318472
rect 482430 318416 482435 318472
rect 448164 318414 482435 318416
rect 448164 318412 448170 318414
rect 482369 318411 482435 318414
rect 446254 318276 446260 318340
rect 446324 318338 446330 318340
rect 472709 318338 472775 318341
rect 446324 318336 472775 318338
rect 446324 318280 472714 318336
rect 472770 318280 472775 318336
rect 446324 318278 472775 318280
rect 446324 318276 446330 318278
rect 472709 318275 472775 318278
rect 480713 318338 480779 318341
rect 511257 318338 511323 318341
rect 480713 318336 511323 318338
rect 480713 318280 480718 318336
rect 480774 318280 511262 318336
rect 511318 318280 511323 318336
rect 480713 318278 511323 318280
rect 480713 318275 480779 318278
rect 511257 318275 511323 318278
rect 509182 316644 509188 316708
rect 509252 316706 509258 316708
rect 510286 316706 510292 316708
rect 509252 316646 510292 316706
rect 509252 316644 509258 316646
rect 510286 316644 510292 316646
rect 510356 316644 510362 316708
rect 454769 315346 454835 315349
rect 514518 315346 514524 315348
rect 454769 315344 514524 315346
rect 454769 315288 454774 315344
rect 454830 315288 514524 315344
rect 454769 315286 514524 315288
rect 454769 315283 454835 315286
rect 514518 315284 514524 315286
rect 514588 315284 514594 315348
rect 434253 315074 434319 315077
rect 431940 315072 434319 315074
rect 431940 315016 434258 315072
rect 434314 315016 434319 315072
rect 431940 315014 434319 315016
rect 434253 315011 434319 315014
rect 382917 312354 382983 312357
rect 379868 312352 382983 312354
rect 379868 312296 382922 312352
rect 382978 312296 382983 312352
rect 379868 312294 382983 312296
rect 382917 312291 382983 312294
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 433977 311130 434043 311133
rect 431940 311128 434043 311130
rect 431940 311072 433982 311128
rect 434038 311072 434043 311128
rect 431940 311070 434043 311072
rect 433977 311067 434043 311070
rect 503437 309770 503503 309773
rect 547638 309770 547644 309772
rect 503437 309768 547644 309770
rect 503437 309712 503442 309768
rect 503498 309712 547644 309768
rect 503437 309710 547644 309712
rect 503437 309707 503503 309710
rect 547638 309708 547644 309710
rect 547708 309708 547714 309772
rect 433885 307186 433951 307189
rect 431940 307184 433951 307186
rect 431940 307128 433890 307184
rect 433946 307128 433951 307184
rect 431940 307126 433951 307128
rect 433885 307123 433951 307126
rect 458766 306988 458772 307052
rect 458836 307050 458842 307052
rect 490281 307050 490347 307053
rect 458836 307048 490347 307050
rect 458836 306992 490286 307048
rect 490342 306992 490347 307048
rect 458836 306990 490347 306992
rect 458836 306988 458842 306990
rect 490281 306987 490347 306990
rect -960 306234 480 306324
rect 3877 306234 3943 306237
rect -960 306232 3943 306234
rect -960 306176 3882 306232
rect 3938 306176 3943 306232
rect -960 306174 3943 306176
rect -960 306084 480 306174
rect 3877 306171 3943 306174
rect 406745 305962 406811 305965
rect 510838 305962 510844 305964
rect 406745 305960 510844 305962
rect 406745 305904 406750 305960
rect 406806 305904 510844 305960
rect 406745 305902 510844 305904
rect 406745 305899 406811 305902
rect 510838 305900 510844 305902
rect 510908 305900 510914 305964
rect 406377 305826 406443 305829
rect 511206 305826 511212 305828
rect 406377 305824 511212 305826
rect 406377 305768 406382 305824
rect 406438 305768 511212 305824
rect 406377 305766 511212 305768
rect 406377 305763 406443 305766
rect 511206 305764 511212 305766
rect 511276 305764 511282 305828
rect 406561 305690 406627 305693
rect 511022 305690 511028 305692
rect 406561 305688 511028 305690
rect 406561 305632 406566 305688
rect 406622 305632 511028 305688
rect 406561 305630 511028 305632
rect 406561 305627 406627 305630
rect 511022 305628 511028 305630
rect 511092 305628 511098 305692
rect 398189 302834 398255 302837
rect 510470 302834 510476 302836
rect 398189 302832 510476 302834
rect 398189 302776 398194 302832
rect 398250 302776 510476 302832
rect 398189 302774 510476 302776
rect 398189 302771 398255 302774
rect 510470 302772 510476 302774
rect 510540 302772 510546 302836
rect 382273 301746 382339 301749
rect 379868 301744 382339 301746
rect 379868 301688 382278 301744
rect 382334 301688 382339 301744
rect 379868 301686 382339 301688
rect 382273 301683 382339 301686
rect 457294 301412 457300 301476
rect 457364 301474 457370 301476
rect 488717 301474 488783 301477
rect 457364 301472 488783 301474
rect 457364 301416 488722 301472
rect 488778 301416 488783 301472
rect 457364 301414 488783 301416
rect 457364 301412 457370 301414
rect 488717 301411 488783 301414
rect 503529 300386 503595 300389
rect 548006 300386 548012 300388
rect 503529 300384 548012 300386
rect 503529 300328 503534 300384
rect 503590 300328 548012 300384
rect 503529 300326 548012 300328
rect 503529 300323 503595 300326
rect 548006 300324 548012 300326
rect 548076 300324 548082 300388
rect 393037 300250 393103 300253
rect 510654 300250 510660 300252
rect 393037 300248 510660 300250
rect 393037 300192 393042 300248
rect 393098 300192 510660 300248
rect 393037 300190 510660 300192
rect 393037 300187 393103 300190
rect 510654 300188 510660 300190
rect 510724 300188 510730 300252
rect 392853 300114 392919 300117
rect 514886 300114 514892 300116
rect 392853 300112 514892 300114
rect 392853 300056 392858 300112
rect 392914 300056 514892 300112
rect 392853 300054 514892 300056
rect 392853 300051 392919 300054
rect 514886 300052 514892 300054
rect 514956 300052 514962 300116
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 389817 297530 389883 297533
rect 514150 297530 514156 297532
rect 389817 297528 514156 297530
rect 389817 297472 389822 297528
rect 389878 297472 514156 297528
rect 389817 297470 514156 297472
rect 389817 297467 389883 297470
rect 514150 297468 514156 297470
rect 514220 297468 514226 297532
rect 392945 297394 393011 297397
rect 518198 297394 518204 297396
rect 392945 297392 518204 297394
rect 392945 297336 392950 297392
rect 393006 297336 518204 297392
rect 392945 297334 518204 297336
rect 392945 297331 393011 297334
rect 518198 297332 518204 297334
rect 518268 297332 518274 297396
rect 391473 294674 391539 294677
rect 507342 294674 507348 294676
rect 391473 294672 507348 294674
rect 391473 294616 391478 294672
rect 391534 294616 507348 294672
rect 391473 294614 507348 294616
rect 391473 294611 391539 294614
rect 507342 294612 507348 294614
rect 507412 294612 507418 294676
rect 384297 294538 384363 294541
rect 508998 294538 509004 294540
rect 384297 294536 509004 294538
rect 384297 294480 384302 294536
rect 384358 294480 509004 294536
rect 384297 294478 509004 294480
rect 384297 294475 384363 294478
rect 508998 294476 509004 294478
rect 509068 294476 509074 294540
rect -960 293178 480 293268
rect 3601 293178 3667 293181
rect -960 293176 3667 293178
rect -960 293120 3606 293176
rect 3662 293120 3667 293176
rect -960 293118 3667 293120
rect -960 293028 480 293118
rect 3601 293115 3667 293118
rect 388437 291954 388503 291957
rect 515070 291954 515076 291956
rect 388437 291952 515076 291954
rect 388437 291896 388442 291952
rect 388498 291896 515076 291952
rect 388437 291894 515076 291896
rect 388437 291891 388503 291894
rect 515070 291892 515076 291894
rect 515140 291892 515146 291956
rect 385861 291818 385927 291821
rect 517830 291818 517836 291820
rect 385861 291816 517836 291818
rect 385861 291760 385866 291816
rect 385922 291760 517836 291816
rect 385861 291758 517836 291760
rect 385861 291755 385927 291758
rect 517830 291756 517836 291758
rect 517900 291756 517906 291820
rect 383285 291138 383351 291141
rect 379868 291136 383351 291138
rect 379868 291080 383290 291136
rect 383346 291080 383351 291136
rect 379868 291078 383351 291080
rect 383285 291075 383351 291078
rect 402329 289234 402395 289237
rect 506974 289234 506980 289236
rect 402329 289232 506980 289234
rect 402329 289176 402334 289232
rect 402390 289176 506980 289232
rect 402329 289174 506980 289176
rect 402329 289171 402395 289174
rect 506974 289172 506980 289174
rect 507044 289172 507050 289236
rect 402513 289098 402579 289101
rect 507158 289098 507164 289100
rect 402513 289096 507164 289098
rect 402513 289040 402518 289096
rect 402574 289040 507164 289096
rect 402513 289038 507164 289040
rect 402513 289035 402579 289038
rect 507158 289036 507164 289038
rect 507228 289036 507234 289100
rect 407757 286378 407823 286381
rect 518014 286378 518020 286380
rect 407757 286376 518020 286378
rect 407757 286320 407762 286376
rect 407818 286320 518020 286376
rect 407757 286318 518020 286320
rect 407757 286315 407823 286318
rect 518014 286316 518020 286318
rect 518084 286316 518090 286380
rect 583520 285276 584960 285516
rect 382273 280530 382339 280533
rect 379868 280528 382339 280530
rect 379868 280472 382278 280528
rect 382334 280472 382339 280528
rect 379868 280470 382339 280472
rect 382273 280467 382339 280470
rect -960 279972 480 280212
rect 457478 278020 457484 278084
rect 457548 278082 457554 278084
rect 488625 278082 488691 278085
rect 457548 278080 488691 278082
rect 457548 278024 488630 278080
rect 488686 278024 488691 278080
rect 457548 278022 488691 278024
rect 457548 278020 457554 278022
rect 488625 278019 488691 278022
rect 446489 276722 446555 276725
rect 463734 276722 463740 276724
rect 446489 276720 463740 276722
rect 446489 276664 446494 276720
rect 446550 276664 463740 276720
rect 446489 276662 463740 276664
rect 446489 276659 446555 276662
rect 463734 276660 463740 276662
rect 463804 276660 463810 276724
rect 457662 272444 457668 272508
rect 457732 272506 457738 272508
rect 490005 272506 490071 272509
rect 457732 272504 490071 272506
rect 457732 272448 490010 272504
rect 490066 272448 490071 272504
rect 457732 272446 490071 272448
rect 457732 272444 457738 272446
rect 490005 272443 490071 272446
rect 580349 272234 580415 272237
rect 583520 272234 584960 272324
rect 580349 272232 584960 272234
rect 580349 272176 580354 272232
rect 580410 272176 584960 272232
rect 580349 272174 584960 272176
rect 580349 272171 580415 272174
rect 583520 272084 584960 272174
rect 382273 269922 382339 269925
rect 379868 269920 382339 269922
rect 379868 269864 382278 269920
rect 382334 269864 382339 269920
rect 379868 269862 382339 269864
rect 382273 269859 382339 269862
rect 458950 268364 458956 268428
rect 459020 268426 459026 268428
rect 489913 268426 489979 268429
rect 459020 268424 489979 268426
rect 459020 268368 489918 268424
rect 489974 268368 489979 268424
rect 459020 268366 489979 268368
rect 459020 268364 459026 268366
rect 489913 268363 489979 268366
rect -960 267202 480 267292
rect 3785 267202 3851 267205
rect -960 267200 3851 267202
rect -960 267144 3790 267200
rect 3846 267144 3851 267200
rect -960 267142 3851 267144
rect -960 267052 480 267142
rect 3785 267139 3851 267142
rect 456793 262714 456859 262717
rect 456793 262712 460092 262714
rect 456793 262656 456798 262712
rect 456854 262656 460092 262712
rect 456793 262654 460092 262656
rect 456793 262651 456859 262654
rect 531405 261082 531471 261085
rect 529828 261080 531471 261082
rect 529828 261024 531410 261080
rect 531466 261024 531471 261080
rect 529828 261022 531471 261024
rect 531405 261019 531471 261022
rect 382273 259314 382339 259317
rect 379868 259312 382339 259314
rect 379868 259256 382278 259312
rect 382334 259256 382339 259312
rect 379868 259254 382339 259256
rect 382273 259251 382339 259254
rect 580349 258906 580415 258909
rect 583520 258906 584960 258996
rect 580349 258904 584960 258906
rect 580349 258848 580354 258904
rect 580410 258848 584960 258904
rect 580349 258846 584960 258848
rect 580349 258843 580415 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3693 254146 3759 254149
rect -960 254144 3759 254146
rect -960 254088 3698 254144
rect 3754 254088 3759 254144
rect -960 254086 3759 254088
rect -960 253996 480 254086
rect 3693 254083 3759 254086
rect 457989 248842 458055 248845
rect 457989 248840 460092 248842
rect 457989 248784 457994 248840
rect 458050 248784 460092 248840
rect 457989 248782 460092 248784
rect 457989 248779 458055 248782
rect 382273 248706 382339 248709
rect 379868 248704 382339 248706
rect 379868 248648 382278 248704
rect 382334 248648 382339 248704
rect 379868 248646 382339 248648
rect 382273 248643 382339 248646
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 530025 244218 530091 244221
rect 529798 244216 530091 244218
rect 529798 244160 530030 244216
rect 530086 244160 530091 244216
rect 529798 244158 530091 244160
rect 529798 243644 529858 244158
rect 530025 244155 530091 244158
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 382273 238098 382339 238101
rect 379868 238096 382339 238098
rect 379868 238040 382278 238096
rect 382334 238040 382339 238096
rect 379868 238038 382339 238040
rect 382273 238035 382339 238038
rect 457161 234970 457227 234973
rect 458081 234970 458147 234973
rect 457161 234968 460092 234970
rect 457161 234912 457166 234968
rect 457222 234912 458086 234968
rect 458142 234912 460092 234968
rect 457161 234910 460092 234912
rect 457161 234907 457227 234910
rect 458081 234907 458147 234910
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 382273 227490 382339 227493
rect 379868 227488 382339 227490
rect 379868 227432 382278 227488
rect 382334 227432 382339 227488
rect 379868 227430 382339 227432
rect 382273 227427 382339 227430
rect 531313 226266 531379 226269
rect 529828 226264 531379 226266
rect 529828 226208 531318 226264
rect 531374 226208 531379 226264
rect 529828 226206 531379 226208
rect 531313 226203 531379 226206
rect 457345 221098 457411 221101
rect 457345 221096 460092 221098
rect 457345 221040 457350 221096
rect 457406 221040 460092 221096
rect 457345 221038 460092 221040
rect 457345 221035 457411 221038
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect 383377 216882 383443 216885
rect 379868 216880 383443 216882
rect 379868 216824 383382 216880
rect 383438 216824 383443 216880
rect 379868 216822 383443 216824
rect 383377 216819 383443 216822
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 529933 209266 529999 209269
rect 529798 209264 529999 209266
rect 529798 209208 529938 209264
rect 529994 209208 529999 209264
rect 529798 209206 529999 209208
rect 529798 208828 529858 209206
rect 529933 209203 529999 209206
rect 456793 207226 456859 207229
rect 457253 207226 457319 207229
rect 456793 207224 460092 207226
rect 456793 207168 456798 207224
rect 456854 207168 457258 207224
rect 457314 207168 460092 207224
rect 456793 207166 460092 207168
rect 456793 207163 456859 207166
rect 457253 207163 457319 207166
rect 382273 206274 382339 206277
rect 379868 206272 382339 206274
rect 379868 206216 382278 206272
rect 382334 206216 382339 206272
rect 379868 206214 382339 206216
rect 382273 206211 382339 206214
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3877 201922 3943 201925
rect -960 201920 3943 201922
rect -960 201864 3882 201920
rect 3938 201864 3943 201920
rect -960 201862 3943 201864
rect -960 201772 480 201862
rect 3877 201859 3943 201862
rect 382273 195666 382339 195669
rect 379868 195664 382339 195666
rect 379868 195608 382278 195664
rect 382334 195608 382339 195664
rect 379868 195606 382339 195608
rect 382273 195603 382339 195606
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3969 188866 4035 188869
rect -960 188864 4035 188866
rect -960 188808 3974 188864
rect 4030 188808 4035 188864
rect -960 188806 4035 188808
rect -960 188716 480 188806
rect 3969 188803 4035 188806
rect 382273 185058 382339 185061
rect 379868 185056 382339 185058
rect 379868 185000 382278 185056
rect 382334 185000 382339 185056
rect 379868 184998 382339 185000
rect 382273 184995 382339 184998
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 382273 174450 382339 174453
rect 379868 174448 382339 174450
rect 379868 174392 382278 174448
rect 382334 174392 382339 174448
rect 379868 174390 382339 174392
rect 382273 174387 382339 174390
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 423259 164388 423325 164389
rect 423254 164386 423260 164388
rect 423172 164326 423260 164386
rect 423324 164386 423330 164388
rect 496169 164386 496235 164389
rect 423324 164384 496235 164386
rect 423324 164328 496174 164384
rect 496230 164328 496235 164384
rect 423254 164324 423260 164326
rect 423324 164326 496235 164328
rect 423324 164324 423330 164326
rect 423259 164323 423325 164324
rect 496169 164323 496235 164326
rect 448278 164114 448284 164116
rect 379838 164054 448284 164114
rect 379838 163812 379898 164054
rect 448278 164052 448284 164054
rect 448348 164114 448354 164116
rect 448348 164054 451290 164114
rect 448348 164052 448354 164054
rect 409137 163434 409203 163437
rect 423254 163434 423260 163436
rect 409137 163432 423260 163434
rect 409137 163376 409142 163432
rect 409198 163376 423260 163432
rect 409137 163374 423260 163376
rect 409137 163371 409203 163374
rect 423254 163372 423260 163374
rect 423324 163372 423330 163436
rect 451230 163434 451290 164054
rect 486417 163434 486483 163437
rect 451230 163432 486483 163434
rect 451230 163376 486422 163432
rect 486478 163376 486483 163432
rect 451230 163374 486483 163376
rect 486417 163371 486483 163374
rect -960 162890 480 162980
rect 3785 162890 3851 162893
rect -960 162888 3851 162890
rect -960 162832 3790 162888
rect 3846 162832 3851 162888
rect -960 162830 3851 162832
rect -960 162740 480 162830
rect 3785 162827 3851 162830
rect 457897 162618 457963 162621
rect 454940 162616 457963 162618
rect 454940 162560 457902 162616
rect 457958 162560 457963 162616
rect 454940 162558 457963 162560
rect 457897 162555 457963 162558
rect 456793 161122 456859 161125
rect 454940 161120 456859 161122
rect 454940 161064 456798 161120
rect 456854 161064 456859 161120
rect 454940 161062 456859 161064
rect 456793 161059 456859 161062
rect 456793 159626 456859 159629
rect 454940 159624 456859 159626
rect 454940 159568 456798 159624
rect 456854 159568 456859 159624
rect 454940 159566 456859 159568
rect 456793 159563 456859 159566
rect 457805 158130 457871 158133
rect 454940 158128 457871 158130
rect 454940 158072 457810 158128
rect 457866 158072 457871 158128
rect 454940 158070 457871 158072
rect 457805 158067 457871 158070
rect 456793 156634 456859 156637
rect 454940 156632 456859 156634
rect 454940 156576 456798 156632
rect 456854 156576 456859 156632
rect 454940 156574 456859 156576
rect 456793 156571 456859 156574
rect 456793 155138 456859 155141
rect 454940 155136 456859 155138
rect 454940 155080 456798 155136
rect 456854 155080 456859 155136
rect 454940 155078 456859 155080
rect 456793 155075 456859 155078
rect 456793 153642 456859 153645
rect 454940 153640 456859 153642
rect 454940 153584 456798 153640
rect 456854 153584 456859 153640
rect 454940 153582 456859 153584
rect 456793 153579 456859 153582
rect 382273 153234 382339 153237
rect 379868 153232 382339 153234
rect 379868 153176 382278 153232
rect 382334 153176 382339 153232
rect 379868 153174 382339 153176
rect 382273 153171 382339 153174
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 457713 152146 457779 152149
rect 454940 152144 457779 152146
rect 454940 152088 457718 152144
rect 457774 152088 457779 152144
rect 454940 152086 457779 152088
rect 457713 152083 457779 152086
rect 456885 150650 456951 150653
rect 454940 150648 456951 150650
rect 454940 150592 456890 150648
rect 456946 150592 456951 150648
rect 454940 150590 456951 150592
rect 456885 150587 456951 150590
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 456793 149154 456859 149157
rect 454940 149152 456859 149154
rect 454940 149096 456798 149152
rect 456854 149096 456859 149152
rect 454940 149094 456859 149096
rect 456793 149091 456859 149094
rect 548006 148548 548012 148612
rect 548076 148610 548082 148612
rect 548076 148550 549362 148610
rect 548076 148548 548082 148550
rect 548006 148140 548012 148204
rect 548076 148202 548082 148204
rect 549161 148202 549227 148205
rect 548076 148200 549227 148202
rect 548076 148144 549166 148200
rect 549222 148144 549227 148200
rect 548076 148142 549227 148144
rect 548076 148140 548082 148142
rect 549161 148139 549227 148142
rect 549302 147900 549362 148550
rect 457437 147658 457503 147661
rect 454940 147656 457503 147658
rect 454940 147600 457442 147656
rect 457498 147600 457503 147656
rect 454940 147598 457503 147600
rect 457437 147595 457503 147598
rect 457621 146162 457687 146165
rect 454940 146160 457687 146162
rect 454940 146104 457626 146160
rect 457682 146104 457687 146160
rect 454940 146102 457687 146104
rect 457621 146099 457687 146102
rect 549897 146026 549963 146029
rect 549854 146024 549963 146026
rect 549854 145968 549902 146024
rect 549958 145968 549963 146024
rect 549854 145963 549963 145968
rect 549854 145452 549914 145963
rect 456793 144666 456859 144669
rect 454940 144664 456859 144666
rect 454940 144608 456798 144664
rect 456854 144608 456859 144664
rect 454940 144606 456859 144608
rect 456793 144603 456859 144606
rect 456793 143170 456859 143173
rect 454940 143168 456859 143170
rect 454940 143112 456798 143168
rect 456854 143112 456859 143168
rect 454940 143110 456859 143112
rect 456793 143107 456859 143110
rect 552105 143034 552171 143037
rect 549884 143032 552171 143034
rect 549884 142976 552110 143032
rect 552166 142976 552171 143032
rect 549884 142974 552171 142976
rect 552105 142971 552171 142974
rect 382273 142626 382339 142629
rect 379868 142624 382339 142626
rect 379868 142568 382278 142624
rect 382334 142568 382339 142624
rect 379868 142566 382339 142568
rect 382273 142563 382339 142566
rect 457253 141674 457319 141677
rect 454940 141672 457319 141674
rect 454940 141616 457258 141672
rect 457314 141616 457319 141672
rect 454940 141614 457319 141616
rect 457253 141611 457319 141614
rect 552565 140586 552631 140589
rect 549884 140584 552631 140586
rect 549884 140528 552570 140584
rect 552626 140528 552631 140584
rect 549884 140526 552631 140528
rect 552565 140523 552631 140526
rect 456793 140178 456859 140181
rect 454940 140176 456859 140178
rect 454940 140120 456798 140176
rect 456854 140120 456859 140176
rect 454940 140118 456859 140120
rect 456793 140115 456859 140118
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 457253 138682 457319 138685
rect 549529 138682 549595 138685
rect 454940 138680 457319 138682
rect 454940 138624 457258 138680
rect 457314 138624 457319 138680
rect 454940 138622 457319 138624
rect 457253 138619 457319 138622
rect 549486 138680 549595 138682
rect 549486 138624 549534 138680
rect 549590 138624 549595 138680
rect 549486 138619 549595 138624
rect 549486 138108 549546 138619
rect 457253 137186 457319 137189
rect 454940 137184 457319 137186
rect 454940 137128 457258 137184
rect 457314 137128 457319 137184
rect 454940 137126 457319 137128
rect 457253 137123 457319 137126
rect -960 136778 480 136868
rect 3693 136778 3759 136781
rect -960 136776 3759 136778
rect -960 136720 3698 136776
rect 3754 136720 3759 136776
rect -960 136718 3759 136720
rect -960 136628 480 136718
rect 3693 136715 3759 136718
rect 549805 136234 549871 136237
rect 549805 136232 549914 136234
rect 549805 136176 549810 136232
rect 549866 136176 549914 136232
rect 549805 136171 549914 136176
rect 458950 135690 458956 135692
rect 454940 135630 458956 135690
rect 458950 135628 458956 135630
rect 459020 135628 459026 135692
rect 549854 135660 549914 136171
rect 457529 134194 457595 134197
rect 454940 134192 457595 134194
rect 454940 134136 457534 134192
rect 457590 134136 457595 134192
rect 454940 134134 457595 134136
rect 457529 134131 457595 134134
rect 552473 133242 552539 133245
rect 549884 133240 552539 133242
rect 549884 133184 552478 133240
rect 552534 133184 552539 133240
rect 549884 133182 552539 133184
rect 552473 133179 552539 133182
rect 457069 132698 457135 132701
rect 454940 132696 457135 132698
rect 454940 132640 457074 132696
rect 457130 132640 457135 132696
rect 454940 132638 457135 132640
rect 457069 132635 457135 132638
rect 382273 132018 382339 132021
rect 379868 132016 382339 132018
rect 379868 131960 382278 132016
rect 382334 131960 382339 132016
rect 379868 131958 382339 131960
rect 382273 131955 382339 131958
rect 457662 131202 457668 131204
rect 454940 131142 457668 131202
rect 457662 131140 457668 131142
rect 457732 131140 457738 131204
rect 549713 131066 549779 131069
rect 549670 131064 549779 131066
rect 549670 131008 549718 131064
rect 549774 131008 549779 131064
rect 549670 131003 549779 131008
rect 549670 130764 549730 131003
rect 458766 129706 458772 129708
rect 454940 129646 458772 129706
rect 458766 129644 458772 129646
rect 458836 129644 458842 129708
rect 552289 128346 552355 128349
rect 549884 128344 552355 128346
rect 549884 128288 552294 128344
rect 552350 128288 552355 128344
rect 549884 128286 552355 128288
rect 552289 128283 552355 128286
rect 457437 128210 457503 128213
rect 454940 128208 457503 128210
rect 454940 128152 457442 128208
rect 457498 128152 457503 128208
rect 454940 128150 457503 128152
rect 457437 128147 457503 128150
rect 457478 126714 457484 126716
rect 454940 126654 457484 126714
rect 457478 126652 457484 126654
rect 457548 126652 457554 126716
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 552749 125898 552815 125901
rect 549884 125896 552815 125898
rect 549884 125840 552754 125896
rect 552810 125840 552815 125896
rect 583520 125884 584960 125974
rect 549884 125838 552815 125840
rect 552749 125835 552815 125838
rect 457345 125218 457411 125221
rect 454940 125216 457411 125218
rect 454940 125160 457350 125216
rect 457406 125160 457411 125216
rect 454940 125158 457411 125160
rect 457345 125155 457411 125158
rect -960 123572 480 123812
rect 457294 123722 457300 123724
rect 454940 123662 457300 123722
rect 457294 123660 457300 123662
rect 457364 123660 457370 123724
rect 551185 123450 551251 123453
rect 549884 123448 551251 123450
rect 549884 123392 551190 123448
rect 551246 123392 551251 123448
rect 549884 123390 551251 123392
rect 551185 123387 551251 123390
rect 457069 122226 457135 122229
rect 454940 122224 457135 122226
rect 454940 122168 457074 122224
rect 457130 122168 457135 122224
rect 454940 122166 457135 122168
rect 457069 122163 457135 122166
rect 383469 121410 383535 121413
rect 379868 121408 383535 121410
rect 379868 121352 383474 121408
rect 383530 121352 383535 121408
rect 379868 121350 383535 121352
rect 383469 121347 383535 121350
rect 551369 121002 551435 121005
rect 549884 121000 551435 121002
rect 549884 120944 551374 121000
rect 551430 120944 551435 121000
rect 549884 120942 551435 120944
rect 551369 120939 551435 120942
rect 551277 118554 551343 118557
rect 549884 118552 551343 118554
rect 549884 118496 551282 118552
rect 551338 118496 551343 118552
rect 549884 118494 551343 118496
rect 551277 118491 551343 118494
rect 551001 116106 551067 116109
rect 549884 116104 551067 116106
rect 549884 116048 551006 116104
rect 551062 116048 551067 116104
rect 549884 116046 551067 116048
rect 551001 116043 551067 116046
rect 550909 113658 550975 113661
rect 549884 113656 550975 113658
rect 549884 113600 550914 113656
rect 550970 113600 550975 113656
rect 549884 113598 550975 113600
rect 550909 113595 550975 113598
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 550817 111210 550883 111213
rect 549884 111208 550883 111210
rect 549884 111152 550822 111208
rect 550878 111152 550883 111208
rect 549884 111150 550883 111152
rect 550817 111147 550883 111150
rect 382273 110802 382339 110805
rect 379868 110800 382339 110802
rect -960 110666 480 110756
rect 379868 110744 382278 110800
rect 382334 110744 382339 110800
rect 379868 110742 382339 110744
rect 382273 110739 382339 110742
rect 3509 110666 3575 110669
rect -960 110664 3575 110666
rect -960 110608 3514 110664
rect 3570 110608 3575 110664
rect -960 110606 3575 110608
rect -960 110516 480 110606
rect 3509 110603 3575 110606
rect 551093 108762 551159 108765
rect 549884 108760 551159 108762
rect 549884 108704 551098 108760
rect 551154 108704 551159 108760
rect 549884 108702 551159 108704
rect 551093 108699 551159 108702
rect 550725 106314 550791 106317
rect 549884 106312 550791 106314
rect 549884 106256 550730 106312
rect 550786 106256 550791 106312
rect 549884 106254 550791 106256
rect 550725 106251 550791 106254
rect 549621 104410 549687 104413
rect 549621 104408 549730 104410
rect 549621 104352 549626 104408
rect 549682 104352 549730 104408
rect 549621 104347 549730 104352
rect 549670 103836 549730 104347
rect 552105 101418 552171 101421
rect 549884 101416 552171 101418
rect 549884 101360 552110 101416
rect 552166 101360 552171 101416
rect 549884 101358 552171 101360
rect 552105 101355 552171 101358
rect 382273 100194 382339 100197
rect 379868 100192 382339 100194
rect 379868 100136 382278 100192
rect 382334 100136 382339 100192
rect 379868 100134 382339 100136
rect 382273 100131 382339 100134
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 549437 99378 549503 99381
rect 549437 99376 549546 99378
rect 549437 99320 549442 99376
rect 549498 99320 549546 99376
rect 583520 99364 584960 99454
rect 549437 99315 549546 99320
rect 549486 98940 549546 99315
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 549345 96794 549411 96797
rect 549302 96792 549411 96794
rect 549302 96736 549350 96792
rect 549406 96736 549411 96792
rect 549302 96731 549411 96736
rect 549302 96492 549362 96731
rect 552381 94074 552447 94077
rect 549884 94072 552447 94074
rect 549884 94016 552386 94072
rect 552442 94016 552447 94072
rect 549884 94014 552447 94016
rect 552381 94011 552447 94014
rect 552657 91626 552723 91629
rect 549884 91624 552723 91626
rect 549884 91568 552662 91624
rect 552718 91568 552723 91624
rect 549884 91566 552723 91568
rect 552657 91563 552723 91566
rect 382273 89586 382339 89589
rect 379868 89584 382339 89586
rect 379868 89528 382278 89584
rect 382334 89528 382339 89584
rect 379868 89526 382339 89528
rect 382273 89523 382339 89526
rect 552197 89178 552263 89181
rect 549884 89176 552263 89178
rect 549884 89120 552202 89176
rect 552258 89120 552263 89176
rect 549884 89118 552263 89120
rect 552197 89115 552263 89118
rect 552013 86730 552079 86733
rect 549884 86728 552079 86730
rect 549884 86672 552018 86728
rect 552074 86672 552079 86728
rect 549884 86670 552079 86672
rect 552013 86667 552079 86670
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 549345 84826 549411 84829
rect 549302 84824 549411 84826
rect -960 84690 480 84780
rect 549302 84768 549350 84824
rect 549406 84768 549411 84824
rect 549302 84763 549411 84768
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 549302 84252 549362 84763
rect 550633 81834 550699 81837
rect 549884 81832 550699 81834
rect 549884 81776 550638 81832
rect 550694 81776 550699 81832
rect 549884 81774 550699 81776
rect 550633 81771 550699 81774
rect 382273 78978 382339 78981
rect 379868 78976 382339 78978
rect 379868 78920 382278 78976
rect 382334 78920 382339 78976
rect 379868 78918 382339 78920
rect 382273 78915 382339 78918
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 382273 68370 382339 68373
rect 379868 68368 382339 68370
rect 379868 68312 382278 68368
rect 382334 68312 382339 68368
rect 379868 68310 382339 68312
rect 382273 68307 382339 68310
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3601 58578 3667 58581
rect -960 58576 3667 58578
rect -960 58520 3606 58576
rect 3662 58520 3667 58576
rect -960 58518 3667 58520
rect -960 58428 480 58518
rect 3601 58515 3667 58518
rect 382273 57762 382339 57765
rect 379868 57760 382339 57762
rect 379868 57704 382278 57760
rect 382334 57704 382339 57760
rect 379868 57702 382339 57704
rect 382273 57699 382339 57702
rect 3601 52050 3667 52053
rect 456333 52050 456399 52053
rect 3601 52048 456399 52050
rect 3601 51992 3606 52048
rect 3662 51992 456338 52048
rect 456394 51992 456399 52048
rect 3601 51990 456399 51992
rect 3601 51987 3667 51990
rect 456333 51987 456399 51990
rect 18597 51914 18663 51917
rect 406469 51914 406535 51917
rect 18597 51912 406535 51914
rect 18597 51856 18602 51912
rect 18658 51856 406474 51912
rect 406530 51856 406535 51912
rect 18597 51854 406535 51856
rect 18597 51851 18663 51854
rect 406469 51851 406535 51854
rect 51349 50826 51415 50829
rect 403709 50826 403775 50829
rect 51349 50824 403775 50826
rect 51349 50768 51354 50824
rect 51410 50768 403714 50824
rect 403770 50768 403775 50824
rect 51349 50766 403775 50768
rect 51349 50763 51415 50766
rect 403709 50763 403775 50766
rect 47853 50690 47919 50693
rect 403893 50690 403959 50693
rect 47853 50688 403959 50690
rect 47853 50632 47858 50688
rect 47914 50632 403898 50688
rect 403954 50632 403959 50688
rect 47853 50630 403959 50632
rect 47853 50627 47919 50630
rect 403893 50627 403959 50630
rect 7649 50554 7715 50557
rect 406745 50554 406811 50557
rect 7649 50552 406811 50554
rect 7649 50496 7654 50552
rect 7710 50496 406750 50552
rect 406806 50496 406811 50552
rect 7649 50494 406811 50496
rect 7649 50491 7715 50494
rect 406745 50491 406811 50494
rect 2865 50418 2931 50421
rect 406561 50418 406627 50421
rect 2865 50416 406627 50418
rect 2865 50360 2870 50416
rect 2926 50360 406566 50416
rect 406622 50360 406627 50416
rect 2865 50358 406627 50360
rect 2865 50355 2931 50358
rect 406561 50355 406627 50358
rect 540605 50418 540671 50421
rect 540605 50416 540714 50418
rect 540605 50360 540610 50416
rect 540666 50360 540714 50416
rect 540605 50355 540714 50360
rect 46657 50282 46723 50285
rect 455045 50282 455111 50285
rect 46657 50280 455111 50282
rect 46657 50224 46662 50280
rect 46718 50224 455050 50280
rect 455106 50224 455111 50280
rect 46657 50222 455111 50224
rect 46657 50219 46723 50222
rect 455045 50219 455111 50222
rect 540654 49844 540714 50355
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 536833 41986 536899 41989
rect 536833 41984 540132 41986
rect 536833 41928 536838 41984
rect 536894 41928 540132 41984
rect 536833 41926 540132 41928
rect 536833 41923 536899 41926
rect 538121 34098 538187 34101
rect 538121 34096 540132 34098
rect 538121 34040 538126 34096
rect 538182 34040 540132 34096
rect 538121 34038 540132 34040
rect 538121 34035 538187 34038
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 5257 4042 5323 4045
rect 380433 4042 380499 4045
rect 5257 4040 380499 4042
rect 5257 3984 5262 4040
rect 5318 3984 380438 4040
rect 380494 3984 380499 4040
rect 5257 3982 380499 3984
rect 5257 3979 5323 3982
rect 380433 3979 380499 3982
rect 9949 3906 10015 3909
rect 388437 3906 388503 3909
rect 9949 3904 388503 3906
rect 9949 3848 9954 3904
rect 10010 3848 388442 3904
rect 388498 3848 388503 3904
rect 9949 3846 388503 3848
rect 9949 3843 10015 3846
rect 388437 3843 388503 3846
rect 6453 3770 6519 3773
rect 407757 3770 407823 3773
rect 6453 3768 407823 3770
rect 6453 3712 6458 3768
rect 6514 3712 407762 3768
rect 407818 3712 407823 3768
rect 6453 3710 407823 3712
rect 6453 3707 6519 3710
rect 407757 3707 407823 3710
rect 1669 3634 1735 3637
rect 406377 3634 406443 3637
rect 1669 3632 406443 3634
rect 1669 3576 1674 3632
rect 1730 3576 406382 3632
rect 406438 3576 406443 3632
rect 1669 3574 406443 3576
rect 1669 3571 1735 3574
rect 406377 3571 406443 3574
rect 4061 3498 4127 3501
rect 454769 3498 454835 3501
rect 4061 3496 454835 3498
rect 4061 3440 4066 3496
rect 4122 3440 454774 3496
rect 454830 3440 454835 3496
rect 4061 3438 454835 3440
rect 4061 3435 4127 3438
rect 454769 3435 454835 3438
rect 565 3362 631 3365
rect 454534 3362 454540 3364
rect 565 3360 454540 3362
rect 565 3304 570 3360
rect 626 3304 454540 3360
rect 565 3302 454540 3304
rect 565 3299 631 3302
rect 454534 3300 454540 3302
rect 454604 3300 454610 3364
<< via3 >>
rect 447916 700572 447980 700636
rect 444236 700436 444300 700500
rect 447732 700300 447796 700364
rect 542676 699756 542740 699820
rect 558868 699756 558932 699820
rect 457852 675684 457916 675748
rect 458036 672828 458100 672892
rect 448100 671332 448164 671396
rect 446260 668612 446324 668676
rect 459140 635700 459204 635764
rect 472020 599524 472084 599588
rect 491340 596804 491404 596868
rect 474780 593948 474844 594012
rect 457852 537372 457916 537436
rect 458036 520916 458100 520980
rect 490420 518060 490484 518124
rect 482692 517576 482756 517580
rect 482692 517520 482742 517576
rect 482742 517520 482756 517576
rect 482692 517516 482756 517520
rect 451044 516700 451108 516764
rect 450492 514320 450556 514384
rect 542676 467196 542740 467260
rect 482692 467060 482756 467124
rect 459140 391172 459204 391236
rect 472020 382332 472084 382396
rect 474780 382332 474844 382396
rect 490420 382332 490484 382396
rect 491340 382332 491404 382396
rect 422892 336772 422956 336836
rect 518204 333372 518268 333436
rect 510660 330924 510724 330988
rect 517836 330108 517900 330172
rect 448284 329624 448348 329628
rect 448284 329568 448298 329624
rect 448298 329568 448348 329624
rect 448284 329564 448348 329568
rect 514892 328476 514956 328540
rect 450630 328204 450694 328268
rect 450492 327660 450556 327724
rect 510292 325212 510356 325276
rect 515076 324396 515140 324460
rect 514156 323988 514220 324052
rect 510844 323580 510908 323644
rect 518020 323172 518084 323236
rect 514708 322356 514772 322420
rect 511028 321948 511092 322012
rect 511212 321540 511276 321604
rect 463740 320316 463804 320380
rect 454540 320180 454604 320244
rect 507164 320588 507228 320652
rect 507348 320452 507412 320516
rect 506980 320316 507044 320380
rect 510476 320180 510540 320244
rect 558868 320044 558932 320108
rect 447732 319908 447796 319972
rect 447916 319772 447980 319836
rect 444236 319636 444300 319700
rect 448100 318412 448164 318476
rect 446260 318276 446324 318340
rect 509188 316644 509252 316708
rect 510292 316644 510356 316708
rect 514524 315284 514588 315348
rect 547644 309708 547708 309772
rect 458772 306988 458836 307052
rect 510844 305900 510908 305964
rect 511212 305764 511276 305828
rect 511028 305628 511092 305692
rect 510476 302772 510540 302836
rect 457300 301412 457364 301476
rect 548012 300324 548076 300388
rect 510660 300188 510724 300252
rect 514892 300052 514956 300116
rect 514156 297468 514220 297532
rect 518204 297332 518268 297396
rect 507348 294612 507412 294676
rect 509004 294476 509068 294540
rect 515076 291892 515140 291956
rect 517836 291756 517900 291820
rect 506980 289172 507044 289236
rect 507164 289036 507228 289100
rect 518020 286316 518084 286380
rect 457484 278020 457548 278084
rect 463740 276660 463804 276724
rect 457668 272444 457732 272508
rect 458956 268364 459020 268428
rect 423260 164384 423324 164388
rect 423260 164328 423264 164384
rect 423264 164328 423320 164384
rect 423320 164328 423324 164384
rect 423260 164324 423324 164328
rect 448284 164052 448348 164116
rect 423260 163372 423324 163436
rect 548012 148548 548076 148612
rect 548012 148140 548076 148204
rect 458956 135628 459020 135692
rect 457668 131140 457732 131204
rect 458772 129644 458836 129708
rect 457484 126652 457548 126716
rect 457300 123660 457364 123724
rect 454540 3300 454604 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 24114 673774 24734 710042
rect 24114 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 24734 673774
rect 24114 673454 24734 673538
rect 24114 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 24734 673454
rect 24114 669548 24734 673218
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 20394 634054 21014 669498
rect 24208 651454 24528 651486
rect 24208 651218 24250 651454
rect 24486 651218 24528 651454
rect 24208 651134 24528 651218
rect 24208 650898 24250 651134
rect 24486 650898 24528 651134
rect 24208 650866 24528 650898
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 27834 641494 28454 676938
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 24208 615454 24528 615486
rect 24208 615218 24250 615454
rect 24486 615218 24528 615454
rect 24208 615134 24528 615218
rect 24208 614898 24250 615134
rect 24486 614898 24528 615134
rect 24208 614866 24528 614898
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 27834 605494 28454 640938
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 24208 579454 24528 579486
rect 24208 579218 24250 579454
rect 24486 579218 24528 579454
rect 24208 579134 24528 579218
rect 24208 578898 24250 579134
rect 24486 578898 24528 579134
rect 24208 578866 24528 578898
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 27834 569494 28454 604938
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 24208 543454 24528 543486
rect 24208 543218 24250 543454
rect 24486 543218 24528 543454
rect 24208 543134 24528 543218
rect 24208 542898 24250 543134
rect 24486 542898 24528 543134
rect 24208 542866 24528 542898
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 27834 533494 28454 568938
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 24208 507454 24528 507486
rect 24208 507218 24250 507454
rect 24486 507218 24528 507454
rect 24208 507134 24528 507218
rect 24208 506898 24250 507134
rect 24486 506898 24528 507134
rect 24208 506866 24528 506898
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 27834 497494 28454 532938
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 24208 471454 24528 471486
rect 24208 471218 24250 471454
rect 24486 471218 24528 471454
rect 24208 471134 24528 471218
rect 24208 470898 24250 471134
rect 24486 470898 24528 471134
rect 24208 470866 24528 470898
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 27834 461494 28454 496938
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 24208 435454 24528 435486
rect 24208 435218 24250 435454
rect 24486 435218 24528 435454
rect 24208 435134 24528 435218
rect 24208 434898 24250 435134
rect 24486 434898 24528 435134
rect 24208 434866 24528 434898
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 27834 425494 28454 460938
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 24208 399454 24528 399486
rect 24208 399218 24250 399454
rect 24486 399218 24528 399454
rect 24208 399134 24528 399218
rect 24208 398898 24250 399134
rect 24486 398898 24528 399134
rect 24208 398866 24528 398898
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 27834 389494 28454 424938
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 24208 363454 24528 363486
rect 24208 363218 24250 363454
rect 24486 363218 24528 363454
rect 24208 363134 24528 363218
rect 24208 362898 24250 363134
rect 24486 362898 24528 363134
rect 24208 362866 24528 362898
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 27834 353494 28454 388938
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 24208 327454 24528 327486
rect 24208 327218 24250 327454
rect 24486 327218 24528 327454
rect 24208 327134 24528 327218
rect 24208 326898 24250 327134
rect 24486 326898 24528 327134
rect 24208 326866 24528 326898
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 27834 317494 28454 352938
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 24208 291454 24528 291486
rect 24208 291218 24250 291454
rect 24486 291218 24528 291454
rect 24208 291134 24528 291218
rect 24208 290898 24250 291134
rect 24486 290898 24528 291134
rect 24208 290866 24528 290898
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 27834 281494 28454 316938
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 24208 255454 24528 255486
rect 24208 255218 24250 255454
rect 24486 255218 24528 255454
rect 24208 255134 24528 255218
rect 24208 254898 24250 255134
rect 24486 254898 24528 255134
rect 24208 254866 24528 254898
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 27834 245494 28454 280938
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 24208 219454 24528 219486
rect 24208 219218 24250 219454
rect 24486 219218 24528 219454
rect 24208 219134 24528 219218
rect 24208 218898 24250 219134
rect 24486 218898 24528 219134
rect 24208 218866 24528 218898
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 27834 209494 28454 244938
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 24208 183454 24528 183486
rect 24208 183218 24250 183454
rect 24486 183218 24528 183454
rect 24208 183134 24528 183218
rect 24208 182898 24250 183134
rect 24486 182898 24528 183134
rect 24208 182866 24528 182898
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 27834 173494 28454 208938
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 24208 147454 24528 147486
rect 24208 147218 24250 147454
rect 24486 147218 24528 147454
rect 24208 147134 24528 147218
rect 24208 146898 24250 147134
rect 24486 146898 24528 147134
rect 24208 146866 24528 146898
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 27834 137494 28454 172938
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 24208 111454 24528 111486
rect 24208 111218 24250 111454
rect 24486 111218 24528 111454
rect 24208 111134 24528 111218
rect 24208 110898 24250 111134
rect 24486 110898 24528 111134
rect 24208 110866 24528 110898
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 27834 101494 28454 136938
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 24208 75454 24528 75486
rect 24208 75218 24250 75454
rect 24486 75218 24528 75454
rect 24208 75134 24528 75218
rect 24208 74898 24250 75134
rect 24486 74898 24528 75134
rect 24208 74866 24528 74898
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 27834 65494 28454 100938
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 25774 24734 50068
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 39568 655174 39888 655206
rect 39568 654938 39610 655174
rect 39846 654938 39888 655174
rect 39568 654854 39888 654938
rect 39568 654618 39610 654854
rect 39846 654618 39888 654854
rect 39568 654586 39888 654618
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 39568 619174 39888 619206
rect 39568 618938 39610 619174
rect 39846 618938 39888 619174
rect 39568 618854 39888 618938
rect 39568 618618 39610 618854
rect 39846 618618 39888 618854
rect 39568 618586 39888 618618
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 39568 583174 39888 583206
rect 39568 582938 39610 583174
rect 39846 582938 39888 583174
rect 39568 582854 39888 582938
rect 39568 582618 39610 582854
rect 39846 582618 39888 582854
rect 39568 582586 39888 582618
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 39568 547174 39888 547206
rect 39568 546938 39610 547174
rect 39846 546938 39888 547174
rect 39568 546854 39888 546938
rect 39568 546618 39610 546854
rect 39846 546618 39888 546854
rect 39568 546586 39888 546618
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 39568 511174 39888 511206
rect 39568 510938 39610 511174
rect 39846 510938 39888 511174
rect 39568 510854 39888 510938
rect 39568 510618 39610 510854
rect 39846 510618 39888 510854
rect 39568 510586 39888 510618
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 39568 475174 39888 475206
rect 39568 474938 39610 475174
rect 39846 474938 39888 475174
rect 39568 474854 39888 474938
rect 39568 474618 39610 474854
rect 39846 474618 39888 474854
rect 39568 474586 39888 474618
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 39568 439174 39888 439206
rect 39568 438938 39610 439174
rect 39846 438938 39888 439174
rect 39568 438854 39888 438938
rect 39568 438618 39610 438854
rect 39846 438618 39888 438854
rect 39568 438586 39888 438618
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 39568 403174 39888 403206
rect 39568 402938 39610 403174
rect 39846 402938 39888 403174
rect 39568 402854 39888 402938
rect 39568 402618 39610 402854
rect 39846 402618 39888 402854
rect 39568 402586 39888 402618
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 39568 367174 39888 367206
rect 39568 366938 39610 367174
rect 39846 366938 39888 367174
rect 39568 366854 39888 366938
rect 39568 366618 39610 366854
rect 39846 366618 39888 366854
rect 39568 366586 39888 366618
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 39568 331174 39888 331206
rect 39568 330938 39610 331174
rect 39846 330938 39888 331174
rect 39568 330854 39888 330938
rect 39568 330618 39610 330854
rect 39846 330618 39888 330854
rect 39568 330586 39888 330618
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 39568 295174 39888 295206
rect 39568 294938 39610 295174
rect 39846 294938 39888 295174
rect 39568 294854 39888 294938
rect 39568 294618 39610 294854
rect 39846 294618 39888 294854
rect 39568 294586 39888 294618
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 39568 259174 39888 259206
rect 39568 258938 39610 259174
rect 39846 258938 39888 259174
rect 39568 258854 39888 258938
rect 39568 258618 39610 258854
rect 39846 258618 39888 258854
rect 39568 258586 39888 258618
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 39568 223174 39888 223206
rect 39568 222938 39610 223174
rect 39846 222938 39888 223174
rect 39568 222854 39888 222938
rect 39568 222618 39610 222854
rect 39846 222618 39888 222854
rect 39568 222586 39888 222618
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 39568 187174 39888 187206
rect 39568 186938 39610 187174
rect 39846 186938 39888 187174
rect 39568 186854 39888 186938
rect 39568 186618 39610 186854
rect 39846 186618 39888 186854
rect 39568 186586 39888 186618
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 39568 151174 39888 151206
rect 39568 150938 39610 151174
rect 39846 150938 39888 151174
rect 39568 150854 39888 150938
rect 39568 150618 39610 150854
rect 39846 150618 39888 150854
rect 39568 150586 39888 150618
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 39568 115174 39888 115206
rect 39568 114938 39610 115174
rect 39846 114938 39888 115174
rect 39568 114854 39888 114938
rect 39568 114618 39610 114854
rect 39846 114618 39888 114854
rect 39568 114586 39888 114618
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 39568 79174 39888 79206
rect 39568 78938 39610 79174
rect 39846 78938 39888 79174
rect 39568 78854 39888 78938
rect 39568 78618 39610 78854
rect 39846 78618 39888 78854
rect 39568 78586 39888 78618
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 708678 53294 711590
rect 52674 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 53294 708678
rect 52674 708358 53294 708442
rect 52674 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 53294 708358
rect 52674 666334 53294 708122
rect 52674 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 53294 666334
rect 52674 666014 53294 666098
rect 52674 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 53294 666014
rect 52674 630334 53294 665778
rect 56394 709638 57014 711590
rect 56394 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 57014 709638
rect 56394 709318 57014 709402
rect 56394 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 57014 709318
rect 56394 670054 57014 709082
rect 56394 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 57014 670054
rect 56394 669734 57014 669818
rect 56394 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 57014 669734
rect 54928 651454 55248 651486
rect 54928 651218 54970 651454
rect 55206 651218 55248 651454
rect 54928 651134 55248 651218
rect 54928 650898 54970 651134
rect 55206 650898 55248 651134
rect 54928 650866 55248 650898
rect 52674 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 53294 630334
rect 52674 630014 53294 630098
rect 52674 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 53294 630014
rect 52674 594334 53294 629778
rect 56394 634054 57014 669498
rect 56394 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 57014 634054
rect 56394 633734 57014 633818
rect 56394 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 57014 633734
rect 54928 615454 55248 615486
rect 54928 615218 54970 615454
rect 55206 615218 55248 615454
rect 54928 615134 55248 615218
rect 54928 614898 54970 615134
rect 55206 614898 55248 615134
rect 54928 614866 55248 614898
rect 52674 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 53294 594334
rect 52674 594014 53294 594098
rect 52674 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 53294 594014
rect 52674 558334 53294 593778
rect 56394 598054 57014 633498
rect 56394 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 57014 598054
rect 56394 597734 57014 597818
rect 56394 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 57014 597734
rect 54928 579454 55248 579486
rect 54928 579218 54970 579454
rect 55206 579218 55248 579454
rect 54928 579134 55248 579218
rect 54928 578898 54970 579134
rect 55206 578898 55248 579134
rect 54928 578866 55248 578898
rect 52674 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 53294 558334
rect 52674 558014 53294 558098
rect 52674 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 53294 558014
rect 52674 522334 53294 557778
rect 56394 562054 57014 597498
rect 56394 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 57014 562054
rect 56394 561734 57014 561818
rect 56394 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 57014 561734
rect 54928 543454 55248 543486
rect 54928 543218 54970 543454
rect 55206 543218 55248 543454
rect 54928 543134 55248 543218
rect 54928 542898 54970 543134
rect 55206 542898 55248 543134
rect 54928 542866 55248 542898
rect 52674 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 53294 522334
rect 52674 522014 53294 522098
rect 52674 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 53294 522014
rect 52674 486334 53294 521778
rect 56394 526054 57014 561498
rect 56394 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 57014 526054
rect 56394 525734 57014 525818
rect 56394 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 57014 525734
rect 54928 507454 55248 507486
rect 54928 507218 54970 507454
rect 55206 507218 55248 507454
rect 54928 507134 55248 507218
rect 54928 506898 54970 507134
rect 55206 506898 55248 507134
rect 54928 506866 55248 506898
rect 52674 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 53294 486334
rect 52674 486014 53294 486098
rect 52674 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 53294 486014
rect 52674 450334 53294 485778
rect 56394 490054 57014 525498
rect 56394 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 57014 490054
rect 56394 489734 57014 489818
rect 56394 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 57014 489734
rect 54928 471454 55248 471486
rect 54928 471218 54970 471454
rect 55206 471218 55248 471454
rect 54928 471134 55248 471218
rect 54928 470898 54970 471134
rect 55206 470898 55248 471134
rect 54928 470866 55248 470898
rect 52674 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 53294 450334
rect 52674 450014 53294 450098
rect 52674 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 53294 450014
rect 52674 414334 53294 449778
rect 56394 454054 57014 489498
rect 56394 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 57014 454054
rect 56394 453734 57014 453818
rect 56394 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 57014 453734
rect 54928 435454 55248 435486
rect 54928 435218 54970 435454
rect 55206 435218 55248 435454
rect 54928 435134 55248 435218
rect 54928 434898 54970 435134
rect 55206 434898 55248 435134
rect 54928 434866 55248 434898
rect 52674 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 53294 414334
rect 52674 414014 53294 414098
rect 52674 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 53294 414014
rect 52674 378334 53294 413778
rect 56394 418054 57014 453498
rect 56394 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 57014 418054
rect 56394 417734 57014 417818
rect 56394 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 57014 417734
rect 54928 399454 55248 399486
rect 54928 399218 54970 399454
rect 55206 399218 55248 399454
rect 54928 399134 55248 399218
rect 54928 398898 54970 399134
rect 55206 398898 55248 399134
rect 54928 398866 55248 398898
rect 52674 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 53294 378334
rect 52674 378014 53294 378098
rect 52674 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 53294 378014
rect 52674 342334 53294 377778
rect 56394 382054 57014 417498
rect 56394 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 57014 382054
rect 56394 381734 57014 381818
rect 56394 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 57014 381734
rect 54928 363454 55248 363486
rect 54928 363218 54970 363454
rect 55206 363218 55248 363454
rect 54928 363134 55248 363218
rect 54928 362898 54970 363134
rect 55206 362898 55248 363134
rect 54928 362866 55248 362898
rect 52674 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 53294 342334
rect 52674 342014 53294 342098
rect 52674 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 53294 342014
rect 52674 306334 53294 341778
rect 56394 346054 57014 381498
rect 56394 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 57014 346054
rect 56394 345734 57014 345818
rect 56394 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 57014 345734
rect 54928 327454 55248 327486
rect 54928 327218 54970 327454
rect 55206 327218 55248 327454
rect 54928 327134 55248 327218
rect 54928 326898 54970 327134
rect 55206 326898 55248 327134
rect 54928 326866 55248 326898
rect 52674 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 53294 306334
rect 52674 306014 53294 306098
rect 52674 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 53294 306014
rect 52674 270334 53294 305778
rect 56394 310054 57014 345498
rect 56394 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 57014 310054
rect 56394 309734 57014 309818
rect 56394 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 57014 309734
rect 54928 291454 55248 291486
rect 54928 291218 54970 291454
rect 55206 291218 55248 291454
rect 54928 291134 55248 291218
rect 54928 290898 54970 291134
rect 55206 290898 55248 291134
rect 54928 290866 55248 290898
rect 52674 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 53294 270334
rect 52674 270014 53294 270098
rect 52674 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 53294 270014
rect 52674 234334 53294 269778
rect 56394 274054 57014 309498
rect 56394 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 57014 274054
rect 56394 273734 57014 273818
rect 56394 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 57014 273734
rect 54928 255454 55248 255486
rect 54928 255218 54970 255454
rect 55206 255218 55248 255454
rect 54928 255134 55248 255218
rect 54928 254898 54970 255134
rect 55206 254898 55248 255134
rect 54928 254866 55248 254898
rect 52674 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 53294 234334
rect 52674 234014 53294 234098
rect 52674 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 53294 234014
rect 52674 198334 53294 233778
rect 56394 238054 57014 273498
rect 56394 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 57014 238054
rect 56394 237734 57014 237818
rect 56394 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 57014 237734
rect 54928 219454 55248 219486
rect 54928 219218 54970 219454
rect 55206 219218 55248 219454
rect 54928 219134 55248 219218
rect 54928 218898 54970 219134
rect 55206 218898 55248 219134
rect 54928 218866 55248 218898
rect 52674 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 53294 198334
rect 52674 198014 53294 198098
rect 52674 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 53294 198014
rect 52674 162334 53294 197778
rect 56394 202054 57014 237498
rect 56394 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 57014 202054
rect 56394 201734 57014 201818
rect 56394 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 57014 201734
rect 54928 183454 55248 183486
rect 54928 183218 54970 183454
rect 55206 183218 55248 183454
rect 54928 183134 55248 183218
rect 54928 182898 54970 183134
rect 55206 182898 55248 183134
rect 54928 182866 55248 182898
rect 52674 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 53294 162334
rect 52674 162014 53294 162098
rect 52674 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 53294 162014
rect 52674 126334 53294 161778
rect 56394 166054 57014 201498
rect 56394 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 57014 166054
rect 56394 165734 57014 165818
rect 56394 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 57014 165734
rect 54928 147454 55248 147486
rect 54928 147218 54970 147454
rect 55206 147218 55248 147454
rect 54928 147134 55248 147218
rect 54928 146898 54970 147134
rect 55206 146898 55248 147134
rect 54928 146866 55248 146898
rect 52674 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 53294 126334
rect 52674 126014 53294 126098
rect 52674 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 53294 126014
rect 52674 90334 53294 125778
rect 56394 130054 57014 165498
rect 56394 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 57014 130054
rect 56394 129734 57014 129818
rect 56394 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 57014 129734
rect 54928 111454 55248 111486
rect 54928 111218 54970 111454
rect 55206 111218 55248 111454
rect 54928 111134 55248 111218
rect 54928 110898 54970 111134
rect 55206 110898 55248 111134
rect 54928 110866 55248 110898
rect 52674 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 53294 90334
rect 52674 90014 53294 90098
rect 52674 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 53294 90014
rect 52674 54334 53294 89778
rect 56394 94054 57014 129498
rect 56394 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 57014 94054
rect 56394 93734 57014 93818
rect 56394 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 57014 93734
rect 54928 75454 55248 75486
rect 54928 75218 54970 75454
rect 55206 75218 55248 75454
rect 54928 75134 55248 75218
rect 54928 74898 54970 75134
rect 55206 74898 55248 75134
rect 54928 74866 55248 74898
rect 52674 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 53294 54334
rect 52674 54014 53294 54098
rect 52674 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 53294 54014
rect 52674 18334 53294 53778
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 58054 57014 93498
rect 56394 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 57014 58054
rect 56394 57734 57014 57818
rect 56394 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 57014 57734
rect 56394 22054 57014 57498
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 710598 60734 711590
rect 60114 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 60734 710598
rect 60114 710278 60734 710362
rect 60114 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 60734 710278
rect 60114 673774 60734 710042
rect 60114 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 60734 673774
rect 60114 673454 60734 673538
rect 60114 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 60734 673454
rect 60114 637774 60734 673218
rect 60114 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 60734 637774
rect 60114 637454 60734 637538
rect 60114 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 60734 637454
rect 60114 601774 60734 637218
rect 60114 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 60734 601774
rect 60114 601454 60734 601538
rect 60114 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 60734 601454
rect 60114 565774 60734 601218
rect 60114 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 60734 565774
rect 60114 565454 60734 565538
rect 60114 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 60734 565454
rect 60114 529774 60734 565218
rect 60114 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 60734 529774
rect 60114 529454 60734 529538
rect 60114 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 60734 529454
rect 60114 493774 60734 529218
rect 60114 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 60734 493774
rect 60114 493454 60734 493538
rect 60114 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 60734 493454
rect 60114 457774 60734 493218
rect 60114 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 60734 457774
rect 60114 457454 60734 457538
rect 60114 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 60734 457454
rect 60114 421774 60734 457218
rect 60114 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 60734 421774
rect 60114 421454 60734 421538
rect 60114 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 60734 421454
rect 60114 385774 60734 421218
rect 60114 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 60734 385774
rect 60114 385454 60734 385538
rect 60114 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 60734 385454
rect 60114 349774 60734 385218
rect 60114 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 60734 349774
rect 60114 349454 60734 349538
rect 60114 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 60734 349454
rect 60114 313774 60734 349218
rect 60114 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 60734 313774
rect 60114 313454 60734 313538
rect 60114 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 60734 313454
rect 60114 277774 60734 313218
rect 60114 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 60734 277774
rect 60114 277454 60734 277538
rect 60114 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 60734 277454
rect 60114 241774 60734 277218
rect 60114 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 60734 241774
rect 60114 241454 60734 241538
rect 60114 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 60734 241454
rect 60114 205774 60734 241218
rect 60114 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 60734 205774
rect 60114 205454 60734 205538
rect 60114 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 60734 205454
rect 60114 169774 60734 205218
rect 60114 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 60734 169774
rect 60114 169454 60734 169538
rect 60114 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 60734 169454
rect 60114 133774 60734 169218
rect 60114 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 60734 133774
rect 60114 133454 60734 133538
rect 60114 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 60734 133454
rect 60114 97774 60734 133218
rect 60114 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 60734 97774
rect 60114 97454 60734 97538
rect 60114 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 60734 97454
rect 60114 61774 60734 97218
rect 60114 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 60734 61774
rect 60114 61454 60734 61538
rect 60114 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 60734 61454
rect 60114 25774 60734 61218
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 641494 64454 676938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 667017 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 667017 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 667017 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 667017 85574 698058
rect 92394 709638 93014 711590
rect 92394 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 93014 709638
rect 92394 709318 93014 709402
rect 92394 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 93014 709318
rect 92394 670054 93014 709082
rect 92394 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 93014 670054
rect 92394 669734 93014 669818
rect 92394 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 93014 669734
rect 92394 667017 93014 669498
rect 96114 710598 96734 711590
rect 96114 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 96734 710598
rect 96114 710278 96734 710362
rect 96114 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 96734 710278
rect 96114 673774 96734 710042
rect 96114 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 96734 673774
rect 96114 673454 96734 673538
rect 96114 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 96734 673454
rect 96114 667017 96734 673218
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 667017 100454 676938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 667017 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 667017 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 667017 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 667017 121574 698058
rect 128394 709638 129014 711590
rect 128394 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 129014 709638
rect 128394 709318 129014 709402
rect 128394 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 129014 709318
rect 128394 670054 129014 709082
rect 128394 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 129014 670054
rect 128394 669734 129014 669818
rect 128394 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 129014 669734
rect 128394 667017 129014 669498
rect 132114 710598 132734 711590
rect 132114 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 132734 710598
rect 132114 710278 132734 710362
rect 132114 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 132734 710278
rect 132114 673774 132734 710042
rect 132114 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 132734 673774
rect 132114 673454 132734 673538
rect 132114 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 132734 673454
rect 132114 667017 132734 673218
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 667017 136454 676938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 667017 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 667017 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 667017 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 667017 157574 698058
rect 164394 709638 165014 711590
rect 164394 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 165014 709638
rect 164394 709318 165014 709402
rect 164394 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 165014 709318
rect 164394 670054 165014 709082
rect 164394 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 165014 670054
rect 164394 669734 165014 669818
rect 164394 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 165014 669734
rect 164394 667017 165014 669498
rect 168114 710598 168734 711590
rect 168114 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 168734 710598
rect 168114 710278 168734 710362
rect 168114 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 168734 710278
rect 168114 673774 168734 710042
rect 168114 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 168734 673774
rect 168114 673454 168734 673538
rect 168114 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 168734 673454
rect 168114 667017 168734 673218
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 667017 172454 676938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 667017 182414 686898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 667017 186134 690618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 667017 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 669548 193574 698058
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 200394 670054 201014 709082
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 667017 201014 669498
rect 204114 710598 204734 711590
rect 204114 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 204734 710598
rect 204114 710278 204734 710362
rect 204114 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 204734 710278
rect 204114 673774 204734 710042
rect 204114 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 204734 673774
rect 204114 673454 204734 673538
rect 204114 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 204734 673454
rect 204114 667017 204734 673218
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 667017 208454 676938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 667017 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 667017 222134 690618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 667017 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 667017 229574 698058
rect 236394 709638 237014 711590
rect 236394 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 237014 709638
rect 236394 709318 237014 709402
rect 236394 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 237014 709318
rect 236394 670054 237014 709082
rect 236394 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 237014 670054
rect 236394 669734 237014 669818
rect 236394 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 237014 669734
rect 236394 667017 237014 669498
rect 240114 710598 240734 711590
rect 240114 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 240734 710598
rect 240114 710278 240734 710362
rect 240114 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 240734 710278
rect 240114 673774 240734 710042
rect 240114 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 240734 673774
rect 240114 673454 240734 673538
rect 240114 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 240734 673454
rect 240114 667017 240734 673218
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 667017 244454 676938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 667017 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 667017 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 667017 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 667017 265574 698058
rect 272394 709638 273014 711590
rect 272394 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 273014 709638
rect 272394 709318 273014 709402
rect 272394 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 273014 709318
rect 272394 670054 273014 709082
rect 272394 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 273014 670054
rect 272394 669734 273014 669818
rect 272394 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 273014 669734
rect 272394 667017 273014 669498
rect 276114 710598 276734 711590
rect 276114 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 276734 710598
rect 276114 710278 276734 710362
rect 276114 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 276734 710278
rect 276114 673774 276734 710042
rect 276114 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 276734 673774
rect 276114 673454 276734 673538
rect 276114 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 276734 673454
rect 276114 667017 276734 673218
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 667017 280454 676938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 667017 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 667017 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 667017 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 669548 301574 698058
rect 308394 709638 309014 711590
rect 308394 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 309014 709638
rect 308394 709318 309014 709402
rect 308394 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 309014 709318
rect 308394 670054 309014 709082
rect 308394 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 309014 670054
rect 308394 669734 309014 669818
rect 308394 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 309014 669734
rect 308394 667017 309014 669498
rect 312114 710598 312734 711590
rect 312114 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 312734 710598
rect 312114 710278 312734 710362
rect 312114 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 312734 710278
rect 312114 673774 312734 710042
rect 312114 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 312734 673774
rect 312114 673454 312734 673538
rect 312114 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 312734 673454
rect 312114 667017 312734 673218
rect 315834 711558 316454 711590
rect 315834 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 316454 711558
rect 315834 711238 316454 711322
rect 315834 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 316454 711238
rect 315834 677494 316454 711002
rect 315834 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 316454 677494
rect 315834 677174 316454 677258
rect 315834 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 316454 677174
rect 315834 669548 316454 676938
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 667017 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 667017 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 667017 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 667017 337574 698058
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 344394 667017 345014 669498
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 348114 667017 348734 673218
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 667017 352454 676938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 669548 362414 686898
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 667017 366134 690618
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 667017 369854 694338
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 667017 373574 698058
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 70288 655174 70608 655206
rect 70288 654938 70330 655174
rect 70566 654938 70608 655174
rect 70288 654854 70608 654938
rect 70288 654618 70330 654854
rect 70566 654618 70608 654854
rect 70288 654586 70608 654618
rect 101008 655174 101328 655206
rect 101008 654938 101050 655174
rect 101286 654938 101328 655174
rect 101008 654854 101328 654938
rect 101008 654618 101050 654854
rect 101286 654618 101328 654854
rect 101008 654586 101328 654618
rect 131728 655174 132048 655206
rect 131728 654938 131770 655174
rect 132006 654938 132048 655174
rect 131728 654854 132048 654938
rect 131728 654618 131770 654854
rect 132006 654618 132048 654854
rect 131728 654586 132048 654618
rect 162448 655174 162768 655206
rect 162448 654938 162490 655174
rect 162726 654938 162768 655174
rect 162448 654854 162768 654938
rect 162448 654618 162490 654854
rect 162726 654618 162768 654854
rect 162448 654586 162768 654618
rect 193168 655174 193488 655206
rect 193168 654938 193210 655174
rect 193446 654938 193488 655174
rect 193168 654854 193488 654938
rect 193168 654618 193210 654854
rect 193446 654618 193488 654854
rect 193168 654586 193488 654618
rect 223888 655174 224208 655206
rect 223888 654938 223930 655174
rect 224166 654938 224208 655174
rect 223888 654854 224208 654938
rect 223888 654618 223930 654854
rect 224166 654618 224208 654854
rect 223888 654586 224208 654618
rect 254608 655174 254928 655206
rect 254608 654938 254650 655174
rect 254886 654938 254928 655174
rect 254608 654854 254928 654938
rect 254608 654618 254650 654854
rect 254886 654618 254928 654854
rect 254608 654586 254928 654618
rect 285328 655174 285648 655206
rect 285328 654938 285370 655174
rect 285606 654938 285648 655174
rect 285328 654854 285648 654938
rect 285328 654618 285370 654854
rect 285606 654618 285648 654854
rect 285328 654586 285648 654618
rect 316048 655174 316368 655206
rect 316048 654938 316090 655174
rect 316326 654938 316368 655174
rect 316048 654854 316368 654938
rect 316048 654618 316090 654854
rect 316326 654618 316368 654854
rect 316048 654586 316368 654618
rect 346768 655174 347088 655206
rect 346768 654938 346810 655174
rect 347046 654938 347088 655174
rect 346768 654854 347088 654938
rect 346768 654618 346810 654854
rect 347046 654618 347088 654854
rect 346768 654586 347088 654618
rect 85648 651454 85968 651486
rect 85648 651218 85690 651454
rect 85926 651218 85968 651454
rect 85648 651134 85968 651218
rect 85648 650898 85690 651134
rect 85926 650898 85968 651134
rect 85648 650866 85968 650898
rect 116368 651454 116688 651486
rect 116368 651218 116410 651454
rect 116646 651218 116688 651454
rect 116368 651134 116688 651218
rect 116368 650898 116410 651134
rect 116646 650898 116688 651134
rect 116368 650866 116688 650898
rect 147088 651454 147408 651486
rect 147088 651218 147130 651454
rect 147366 651218 147408 651454
rect 147088 651134 147408 651218
rect 147088 650898 147130 651134
rect 147366 650898 147408 651134
rect 147088 650866 147408 650898
rect 177808 651454 178128 651486
rect 177808 651218 177850 651454
rect 178086 651218 178128 651454
rect 177808 651134 178128 651218
rect 177808 650898 177850 651134
rect 178086 650898 178128 651134
rect 177808 650866 178128 650898
rect 208528 651454 208848 651486
rect 208528 651218 208570 651454
rect 208806 651218 208848 651454
rect 208528 651134 208848 651218
rect 208528 650898 208570 651134
rect 208806 650898 208848 651134
rect 208528 650866 208848 650898
rect 239248 651454 239568 651486
rect 239248 651218 239290 651454
rect 239526 651218 239568 651454
rect 239248 651134 239568 651218
rect 239248 650898 239290 651134
rect 239526 650898 239568 651134
rect 239248 650866 239568 650898
rect 269968 651454 270288 651486
rect 269968 651218 270010 651454
rect 270246 651218 270288 651454
rect 269968 651134 270288 651218
rect 269968 650898 270010 651134
rect 270246 650898 270288 651134
rect 269968 650866 270288 650898
rect 300688 651454 301008 651486
rect 300688 651218 300730 651454
rect 300966 651218 301008 651454
rect 300688 651134 301008 651218
rect 300688 650898 300730 651134
rect 300966 650898 301008 651134
rect 300688 650866 301008 650898
rect 331408 651454 331728 651486
rect 331408 651218 331450 651454
rect 331686 651218 331728 651454
rect 331408 651134 331728 651218
rect 331408 650898 331450 651134
rect 331686 650898 331728 651134
rect 331408 650866 331728 650898
rect 362128 651454 362448 651486
rect 362128 651218 362170 651454
rect 362406 651218 362448 651454
rect 362128 651134 362448 651218
rect 362128 650898 362170 651134
rect 362406 650898 362448 651134
rect 362128 650866 362448 650898
rect 63834 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 64454 641494
rect 63834 641174 64454 641258
rect 63834 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 64454 641174
rect 63834 605494 64454 640938
rect 376674 630334 377294 665778
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 377488 655174 377808 655206
rect 377488 654938 377530 655174
rect 377766 654938 377808 655174
rect 377488 654854 377808 654938
rect 377488 654618 377530 654854
rect 377766 654618 377808 654854
rect 377488 654586 377808 654618
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 70288 619174 70608 619206
rect 70288 618938 70330 619174
rect 70566 618938 70608 619174
rect 70288 618854 70608 618938
rect 70288 618618 70330 618854
rect 70566 618618 70608 618854
rect 70288 618586 70608 618618
rect 101008 619174 101328 619206
rect 101008 618938 101050 619174
rect 101286 618938 101328 619174
rect 101008 618854 101328 618938
rect 101008 618618 101050 618854
rect 101286 618618 101328 618854
rect 101008 618586 101328 618618
rect 131728 619174 132048 619206
rect 131728 618938 131770 619174
rect 132006 618938 132048 619174
rect 131728 618854 132048 618938
rect 131728 618618 131770 618854
rect 132006 618618 132048 618854
rect 131728 618586 132048 618618
rect 162448 619174 162768 619206
rect 162448 618938 162490 619174
rect 162726 618938 162768 619174
rect 162448 618854 162768 618938
rect 162448 618618 162490 618854
rect 162726 618618 162768 618854
rect 162448 618586 162768 618618
rect 193168 619174 193488 619206
rect 193168 618938 193210 619174
rect 193446 618938 193488 619174
rect 193168 618854 193488 618938
rect 193168 618618 193210 618854
rect 193446 618618 193488 618854
rect 193168 618586 193488 618618
rect 223888 619174 224208 619206
rect 223888 618938 223930 619174
rect 224166 618938 224208 619174
rect 223888 618854 224208 618938
rect 223888 618618 223930 618854
rect 224166 618618 224208 618854
rect 223888 618586 224208 618618
rect 254608 619174 254928 619206
rect 254608 618938 254650 619174
rect 254886 618938 254928 619174
rect 254608 618854 254928 618938
rect 254608 618618 254650 618854
rect 254886 618618 254928 618854
rect 254608 618586 254928 618618
rect 285328 619174 285648 619206
rect 285328 618938 285370 619174
rect 285606 618938 285648 619174
rect 285328 618854 285648 618938
rect 285328 618618 285370 618854
rect 285606 618618 285648 618854
rect 285328 618586 285648 618618
rect 316048 619174 316368 619206
rect 316048 618938 316090 619174
rect 316326 618938 316368 619174
rect 316048 618854 316368 618938
rect 316048 618618 316090 618854
rect 316326 618618 316368 618854
rect 316048 618586 316368 618618
rect 346768 619174 347088 619206
rect 346768 618938 346810 619174
rect 347046 618938 347088 619174
rect 346768 618854 347088 618938
rect 346768 618618 346810 618854
rect 347046 618618 347088 618854
rect 346768 618586 347088 618618
rect 85648 615454 85968 615486
rect 85648 615218 85690 615454
rect 85926 615218 85968 615454
rect 85648 615134 85968 615218
rect 85648 614898 85690 615134
rect 85926 614898 85968 615134
rect 85648 614866 85968 614898
rect 116368 615454 116688 615486
rect 116368 615218 116410 615454
rect 116646 615218 116688 615454
rect 116368 615134 116688 615218
rect 116368 614898 116410 615134
rect 116646 614898 116688 615134
rect 116368 614866 116688 614898
rect 147088 615454 147408 615486
rect 147088 615218 147130 615454
rect 147366 615218 147408 615454
rect 147088 615134 147408 615218
rect 147088 614898 147130 615134
rect 147366 614898 147408 615134
rect 147088 614866 147408 614898
rect 177808 615454 178128 615486
rect 177808 615218 177850 615454
rect 178086 615218 178128 615454
rect 177808 615134 178128 615218
rect 177808 614898 177850 615134
rect 178086 614898 178128 615134
rect 177808 614866 178128 614898
rect 208528 615454 208848 615486
rect 208528 615218 208570 615454
rect 208806 615218 208848 615454
rect 208528 615134 208848 615218
rect 208528 614898 208570 615134
rect 208806 614898 208848 615134
rect 208528 614866 208848 614898
rect 239248 615454 239568 615486
rect 239248 615218 239290 615454
rect 239526 615218 239568 615454
rect 239248 615134 239568 615218
rect 239248 614898 239290 615134
rect 239526 614898 239568 615134
rect 239248 614866 239568 614898
rect 269968 615454 270288 615486
rect 269968 615218 270010 615454
rect 270246 615218 270288 615454
rect 269968 615134 270288 615218
rect 269968 614898 270010 615134
rect 270246 614898 270288 615134
rect 269968 614866 270288 614898
rect 300688 615454 301008 615486
rect 300688 615218 300730 615454
rect 300966 615218 301008 615454
rect 300688 615134 301008 615218
rect 300688 614898 300730 615134
rect 300966 614898 301008 615134
rect 300688 614866 301008 614898
rect 331408 615454 331728 615486
rect 331408 615218 331450 615454
rect 331686 615218 331728 615454
rect 331408 615134 331728 615218
rect 331408 614898 331450 615134
rect 331686 614898 331728 615134
rect 331408 614866 331728 614898
rect 362128 615454 362448 615486
rect 362128 615218 362170 615454
rect 362406 615218 362448 615454
rect 362128 615134 362448 615218
rect 362128 614898 362170 615134
rect 362406 614898 362448 615134
rect 362128 614866 362448 614898
rect 63834 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 64454 605494
rect 63834 605174 64454 605258
rect 63834 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 64454 605174
rect 63834 569494 64454 604938
rect 376674 594334 377294 629778
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 377488 619174 377808 619206
rect 377488 618938 377530 619174
rect 377766 618938 377808 619174
rect 377488 618854 377808 618938
rect 377488 618618 377530 618854
rect 377766 618618 377808 618854
rect 377488 618586 377808 618618
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 70288 583174 70608 583206
rect 70288 582938 70330 583174
rect 70566 582938 70608 583174
rect 70288 582854 70608 582938
rect 70288 582618 70330 582854
rect 70566 582618 70608 582854
rect 70288 582586 70608 582618
rect 101008 583174 101328 583206
rect 101008 582938 101050 583174
rect 101286 582938 101328 583174
rect 101008 582854 101328 582938
rect 101008 582618 101050 582854
rect 101286 582618 101328 582854
rect 101008 582586 101328 582618
rect 131728 583174 132048 583206
rect 131728 582938 131770 583174
rect 132006 582938 132048 583174
rect 131728 582854 132048 582938
rect 131728 582618 131770 582854
rect 132006 582618 132048 582854
rect 131728 582586 132048 582618
rect 162448 583174 162768 583206
rect 162448 582938 162490 583174
rect 162726 582938 162768 583174
rect 162448 582854 162768 582938
rect 162448 582618 162490 582854
rect 162726 582618 162768 582854
rect 162448 582586 162768 582618
rect 193168 583174 193488 583206
rect 193168 582938 193210 583174
rect 193446 582938 193488 583174
rect 193168 582854 193488 582938
rect 193168 582618 193210 582854
rect 193446 582618 193488 582854
rect 193168 582586 193488 582618
rect 223888 583174 224208 583206
rect 223888 582938 223930 583174
rect 224166 582938 224208 583174
rect 223888 582854 224208 582938
rect 223888 582618 223930 582854
rect 224166 582618 224208 582854
rect 223888 582586 224208 582618
rect 254608 583174 254928 583206
rect 254608 582938 254650 583174
rect 254886 582938 254928 583174
rect 254608 582854 254928 582938
rect 254608 582618 254650 582854
rect 254886 582618 254928 582854
rect 254608 582586 254928 582618
rect 285328 583174 285648 583206
rect 285328 582938 285370 583174
rect 285606 582938 285648 583174
rect 285328 582854 285648 582938
rect 285328 582618 285370 582854
rect 285606 582618 285648 582854
rect 285328 582586 285648 582618
rect 316048 583174 316368 583206
rect 316048 582938 316090 583174
rect 316326 582938 316368 583174
rect 316048 582854 316368 582938
rect 316048 582618 316090 582854
rect 316326 582618 316368 582854
rect 316048 582586 316368 582618
rect 346768 583174 347088 583206
rect 346768 582938 346810 583174
rect 347046 582938 347088 583174
rect 346768 582854 347088 582938
rect 346768 582618 346810 582854
rect 347046 582618 347088 582854
rect 346768 582586 347088 582618
rect 85648 579454 85968 579486
rect 85648 579218 85690 579454
rect 85926 579218 85968 579454
rect 85648 579134 85968 579218
rect 85648 578898 85690 579134
rect 85926 578898 85968 579134
rect 85648 578866 85968 578898
rect 116368 579454 116688 579486
rect 116368 579218 116410 579454
rect 116646 579218 116688 579454
rect 116368 579134 116688 579218
rect 116368 578898 116410 579134
rect 116646 578898 116688 579134
rect 116368 578866 116688 578898
rect 147088 579454 147408 579486
rect 147088 579218 147130 579454
rect 147366 579218 147408 579454
rect 147088 579134 147408 579218
rect 147088 578898 147130 579134
rect 147366 578898 147408 579134
rect 147088 578866 147408 578898
rect 177808 579454 178128 579486
rect 177808 579218 177850 579454
rect 178086 579218 178128 579454
rect 177808 579134 178128 579218
rect 177808 578898 177850 579134
rect 178086 578898 178128 579134
rect 177808 578866 178128 578898
rect 208528 579454 208848 579486
rect 208528 579218 208570 579454
rect 208806 579218 208848 579454
rect 208528 579134 208848 579218
rect 208528 578898 208570 579134
rect 208806 578898 208848 579134
rect 208528 578866 208848 578898
rect 239248 579454 239568 579486
rect 239248 579218 239290 579454
rect 239526 579218 239568 579454
rect 239248 579134 239568 579218
rect 239248 578898 239290 579134
rect 239526 578898 239568 579134
rect 239248 578866 239568 578898
rect 269968 579454 270288 579486
rect 269968 579218 270010 579454
rect 270246 579218 270288 579454
rect 269968 579134 270288 579218
rect 269968 578898 270010 579134
rect 270246 578898 270288 579134
rect 269968 578866 270288 578898
rect 300688 579454 301008 579486
rect 300688 579218 300730 579454
rect 300966 579218 301008 579454
rect 300688 579134 301008 579218
rect 300688 578898 300730 579134
rect 300966 578898 301008 579134
rect 300688 578866 301008 578898
rect 331408 579454 331728 579486
rect 331408 579218 331450 579454
rect 331686 579218 331728 579454
rect 331408 579134 331728 579218
rect 331408 578898 331450 579134
rect 331686 578898 331728 579134
rect 331408 578866 331728 578898
rect 362128 579454 362448 579486
rect 362128 579218 362170 579454
rect 362406 579218 362448 579454
rect 362128 579134 362448 579218
rect 362128 578898 362170 579134
rect 362406 578898 362448 579134
rect 362128 578866 362448 578898
rect 63834 569258 63866 569494
rect 64102 569258 64186 569494
rect 64422 569258 64454 569494
rect 63834 569174 64454 569258
rect 63834 568938 63866 569174
rect 64102 568938 64186 569174
rect 64422 568938 64454 569174
rect 63834 533494 64454 568938
rect 376674 558334 377294 593778
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 377488 583174 377808 583206
rect 377488 582938 377530 583174
rect 377766 582938 377808 583174
rect 377488 582854 377808 582938
rect 377488 582618 377530 582854
rect 377766 582618 377808 582854
rect 377488 582586 377808 582618
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 70288 547174 70608 547206
rect 70288 546938 70330 547174
rect 70566 546938 70608 547174
rect 70288 546854 70608 546938
rect 70288 546618 70330 546854
rect 70566 546618 70608 546854
rect 70288 546586 70608 546618
rect 101008 547174 101328 547206
rect 101008 546938 101050 547174
rect 101286 546938 101328 547174
rect 101008 546854 101328 546938
rect 101008 546618 101050 546854
rect 101286 546618 101328 546854
rect 101008 546586 101328 546618
rect 131728 547174 132048 547206
rect 131728 546938 131770 547174
rect 132006 546938 132048 547174
rect 131728 546854 132048 546938
rect 131728 546618 131770 546854
rect 132006 546618 132048 546854
rect 131728 546586 132048 546618
rect 162448 547174 162768 547206
rect 162448 546938 162490 547174
rect 162726 546938 162768 547174
rect 162448 546854 162768 546938
rect 162448 546618 162490 546854
rect 162726 546618 162768 546854
rect 162448 546586 162768 546618
rect 193168 547174 193488 547206
rect 193168 546938 193210 547174
rect 193446 546938 193488 547174
rect 193168 546854 193488 546938
rect 193168 546618 193210 546854
rect 193446 546618 193488 546854
rect 193168 546586 193488 546618
rect 223888 547174 224208 547206
rect 223888 546938 223930 547174
rect 224166 546938 224208 547174
rect 223888 546854 224208 546938
rect 223888 546618 223930 546854
rect 224166 546618 224208 546854
rect 223888 546586 224208 546618
rect 254608 547174 254928 547206
rect 254608 546938 254650 547174
rect 254886 546938 254928 547174
rect 254608 546854 254928 546938
rect 254608 546618 254650 546854
rect 254886 546618 254928 546854
rect 254608 546586 254928 546618
rect 285328 547174 285648 547206
rect 285328 546938 285370 547174
rect 285606 546938 285648 547174
rect 285328 546854 285648 546938
rect 285328 546618 285370 546854
rect 285606 546618 285648 546854
rect 285328 546586 285648 546618
rect 316048 547174 316368 547206
rect 316048 546938 316090 547174
rect 316326 546938 316368 547174
rect 316048 546854 316368 546938
rect 316048 546618 316090 546854
rect 316326 546618 316368 546854
rect 316048 546586 316368 546618
rect 346768 547174 347088 547206
rect 346768 546938 346810 547174
rect 347046 546938 347088 547174
rect 346768 546854 347088 546938
rect 346768 546618 346810 546854
rect 347046 546618 347088 546854
rect 346768 546586 347088 546618
rect 85648 543454 85968 543486
rect 85648 543218 85690 543454
rect 85926 543218 85968 543454
rect 85648 543134 85968 543218
rect 85648 542898 85690 543134
rect 85926 542898 85968 543134
rect 85648 542866 85968 542898
rect 116368 543454 116688 543486
rect 116368 543218 116410 543454
rect 116646 543218 116688 543454
rect 116368 543134 116688 543218
rect 116368 542898 116410 543134
rect 116646 542898 116688 543134
rect 116368 542866 116688 542898
rect 147088 543454 147408 543486
rect 147088 543218 147130 543454
rect 147366 543218 147408 543454
rect 147088 543134 147408 543218
rect 147088 542898 147130 543134
rect 147366 542898 147408 543134
rect 147088 542866 147408 542898
rect 177808 543454 178128 543486
rect 177808 543218 177850 543454
rect 178086 543218 178128 543454
rect 177808 543134 178128 543218
rect 177808 542898 177850 543134
rect 178086 542898 178128 543134
rect 177808 542866 178128 542898
rect 208528 543454 208848 543486
rect 208528 543218 208570 543454
rect 208806 543218 208848 543454
rect 208528 543134 208848 543218
rect 208528 542898 208570 543134
rect 208806 542898 208848 543134
rect 208528 542866 208848 542898
rect 239248 543454 239568 543486
rect 239248 543218 239290 543454
rect 239526 543218 239568 543454
rect 239248 543134 239568 543218
rect 239248 542898 239290 543134
rect 239526 542898 239568 543134
rect 239248 542866 239568 542898
rect 269968 543454 270288 543486
rect 269968 543218 270010 543454
rect 270246 543218 270288 543454
rect 269968 543134 270288 543218
rect 269968 542898 270010 543134
rect 270246 542898 270288 543134
rect 269968 542866 270288 542898
rect 300688 543454 301008 543486
rect 300688 543218 300730 543454
rect 300966 543218 301008 543454
rect 300688 543134 301008 543218
rect 300688 542898 300730 543134
rect 300966 542898 301008 543134
rect 300688 542866 301008 542898
rect 331408 543454 331728 543486
rect 331408 543218 331450 543454
rect 331686 543218 331728 543454
rect 331408 543134 331728 543218
rect 331408 542898 331450 543134
rect 331686 542898 331728 543134
rect 331408 542866 331728 542898
rect 362128 543454 362448 543486
rect 362128 543218 362170 543454
rect 362406 543218 362448 543454
rect 362128 543134 362448 543218
rect 362128 542898 362170 543134
rect 362406 542898 362448 543134
rect 362128 542866 362448 542898
rect 63834 533258 63866 533494
rect 64102 533258 64186 533494
rect 64422 533258 64454 533494
rect 63834 533174 64454 533258
rect 63834 532938 63866 533174
rect 64102 532938 64186 533174
rect 64422 532938 64454 533174
rect 63834 497494 64454 532938
rect 376674 522334 377294 557778
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 377488 547174 377808 547206
rect 377488 546938 377530 547174
rect 377766 546938 377808 547174
rect 377488 546854 377808 546938
rect 377488 546618 377530 546854
rect 377766 546618 377808 546854
rect 377488 546586 377808 546618
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 70288 511174 70608 511206
rect 70288 510938 70330 511174
rect 70566 510938 70608 511174
rect 70288 510854 70608 510938
rect 70288 510618 70330 510854
rect 70566 510618 70608 510854
rect 70288 510586 70608 510618
rect 101008 511174 101328 511206
rect 101008 510938 101050 511174
rect 101286 510938 101328 511174
rect 101008 510854 101328 510938
rect 101008 510618 101050 510854
rect 101286 510618 101328 510854
rect 101008 510586 101328 510618
rect 131728 511174 132048 511206
rect 131728 510938 131770 511174
rect 132006 510938 132048 511174
rect 131728 510854 132048 510938
rect 131728 510618 131770 510854
rect 132006 510618 132048 510854
rect 131728 510586 132048 510618
rect 162448 511174 162768 511206
rect 162448 510938 162490 511174
rect 162726 510938 162768 511174
rect 162448 510854 162768 510938
rect 162448 510618 162490 510854
rect 162726 510618 162768 510854
rect 162448 510586 162768 510618
rect 193168 511174 193488 511206
rect 193168 510938 193210 511174
rect 193446 510938 193488 511174
rect 193168 510854 193488 510938
rect 193168 510618 193210 510854
rect 193446 510618 193488 510854
rect 193168 510586 193488 510618
rect 223888 511174 224208 511206
rect 223888 510938 223930 511174
rect 224166 510938 224208 511174
rect 223888 510854 224208 510938
rect 223888 510618 223930 510854
rect 224166 510618 224208 510854
rect 223888 510586 224208 510618
rect 254608 511174 254928 511206
rect 254608 510938 254650 511174
rect 254886 510938 254928 511174
rect 254608 510854 254928 510938
rect 254608 510618 254650 510854
rect 254886 510618 254928 510854
rect 254608 510586 254928 510618
rect 285328 511174 285648 511206
rect 285328 510938 285370 511174
rect 285606 510938 285648 511174
rect 285328 510854 285648 510938
rect 285328 510618 285370 510854
rect 285606 510618 285648 510854
rect 285328 510586 285648 510618
rect 316048 511174 316368 511206
rect 316048 510938 316090 511174
rect 316326 510938 316368 511174
rect 316048 510854 316368 510938
rect 316048 510618 316090 510854
rect 316326 510618 316368 510854
rect 316048 510586 316368 510618
rect 346768 511174 347088 511206
rect 346768 510938 346810 511174
rect 347046 510938 347088 511174
rect 346768 510854 347088 510938
rect 346768 510618 346810 510854
rect 347046 510618 347088 510854
rect 346768 510586 347088 510618
rect 85648 507454 85968 507486
rect 85648 507218 85690 507454
rect 85926 507218 85968 507454
rect 85648 507134 85968 507218
rect 85648 506898 85690 507134
rect 85926 506898 85968 507134
rect 85648 506866 85968 506898
rect 116368 507454 116688 507486
rect 116368 507218 116410 507454
rect 116646 507218 116688 507454
rect 116368 507134 116688 507218
rect 116368 506898 116410 507134
rect 116646 506898 116688 507134
rect 116368 506866 116688 506898
rect 147088 507454 147408 507486
rect 147088 507218 147130 507454
rect 147366 507218 147408 507454
rect 147088 507134 147408 507218
rect 147088 506898 147130 507134
rect 147366 506898 147408 507134
rect 147088 506866 147408 506898
rect 177808 507454 178128 507486
rect 177808 507218 177850 507454
rect 178086 507218 178128 507454
rect 177808 507134 178128 507218
rect 177808 506898 177850 507134
rect 178086 506898 178128 507134
rect 177808 506866 178128 506898
rect 208528 507454 208848 507486
rect 208528 507218 208570 507454
rect 208806 507218 208848 507454
rect 208528 507134 208848 507218
rect 208528 506898 208570 507134
rect 208806 506898 208848 507134
rect 208528 506866 208848 506898
rect 239248 507454 239568 507486
rect 239248 507218 239290 507454
rect 239526 507218 239568 507454
rect 239248 507134 239568 507218
rect 239248 506898 239290 507134
rect 239526 506898 239568 507134
rect 239248 506866 239568 506898
rect 269968 507454 270288 507486
rect 269968 507218 270010 507454
rect 270246 507218 270288 507454
rect 269968 507134 270288 507218
rect 269968 506898 270010 507134
rect 270246 506898 270288 507134
rect 269968 506866 270288 506898
rect 300688 507454 301008 507486
rect 300688 507218 300730 507454
rect 300966 507218 301008 507454
rect 300688 507134 301008 507218
rect 300688 506898 300730 507134
rect 300966 506898 301008 507134
rect 300688 506866 301008 506898
rect 331408 507454 331728 507486
rect 331408 507218 331450 507454
rect 331686 507218 331728 507454
rect 331408 507134 331728 507218
rect 331408 506898 331450 507134
rect 331686 506898 331728 507134
rect 331408 506866 331728 506898
rect 362128 507454 362448 507486
rect 362128 507218 362170 507454
rect 362406 507218 362448 507454
rect 362128 507134 362448 507218
rect 362128 506898 362170 507134
rect 362406 506898 362448 507134
rect 362128 506866 362448 506898
rect 63834 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 64454 497494
rect 63834 497174 64454 497258
rect 63834 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 64454 497174
rect 63834 461494 64454 496938
rect 376674 486334 377294 521778
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 377488 511174 377808 511206
rect 377488 510938 377530 511174
rect 377766 510938 377808 511174
rect 377488 510854 377808 510938
rect 377488 510618 377530 510854
rect 377766 510618 377808 510854
rect 377488 510586 377808 510618
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 70288 475174 70608 475206
rect 70288 474938 70330 475174
rect 70566 474938 70608 475174
rect 70288 474854 70608 474938
rect 70288 474618 70330 474854
rect 70566 474618 70608 474854
rect 70288 474586 70608 474618
rect 101008 475174 101328 475206
rect 101008 474938 101050 475174
rect 101286 474938 101328 475174
rect 101008 474854 101328 474938
rect 101008 474618 101050 474854
rect 101286 474618 101328 474854
rect 101008 474586 101328 474618
rect 131728 475174 132048 475206
rect 131728 474938 131770 475174
rect 132006 474938 132048 475174
rect 131728 474854 132048 474938
rect 131728 474618 131770 474854
rect 132006 474618 132048 474854
rect 131728 474586 132048 474618
rect 162448 475174 162768 475206
rect 162448 474938 162490 475174
rect 162726 474938 162768 475174
rect 162448 474854 162768 474938
rect 162448 474618 162490 474854
rect 162726 474618 162768 474854
rect 162448 474586 162768 474618
rect 193168 475174 193488 475206
rect 193168 474938 193210 475174
rect 193446 474938 193488 475174
rect 193168 474854 193488 474938
rect 193168 474618 193210 474854
rect 193446 474618 193488 474854
rect 193168 474586 193488 474618
rect 223888 475174 224208 475206
rect 223888 474938 223930 475174
rect 224166 474938 224208 475174
rect 223888 474854 224208 474938
rect 223888 474618 223930 474854
rect 224166 474618 224208 474854
rect 223888 474586 224208 474618
rect 254608 475174 254928 475206
rect 254608 474938 254650 475174
rect 254886 474938 254928 475174
rect 254608 474854 254928 474938
rect 254608 474618 254650 474854
rect 254886 474618 254928 474854
rect 254608 474586 254928 474618
rect 285328 475174 285648 475206
rect 285328 474938 285370 475174
rect 285606 474938 285648 475174
rect 285328 474854 285648 474938
rect 285328 474618 285370 474854
rect 285606 474618 285648 474854
rect 285328 474586 285648 474618
rect 316048 475174 316368 475206
rect 316048 474938 316090 475174
rect 316326 474938 316368 475174
rect 316048 474854 316368 474938
rect 316048 474618 316090 474854
rect 316326 474618 316368 474854
rect 316048 474586 316368 474618
rect 346768 475174 347088 475206
rect 346768 474938 346810 475174
rect 347046 474938 347088 475174
rect 346768 474854 347088 474938
rect 346768 474618 346810 474854
rect 347046 474618 347088 474854
rect 346768 474586 347088 474618
rect 85648 471454 85968 471486
rect 85648 471218 85690 471454
rect 85926 471218 85968 471454
rect 85648 471134 85968 471218
rect 85648 470898 85690 471134
rect 85926 470898 85968 471134
rect 85648 470866 85968 470898
rect 116368 471454 116688 471486
rect 116368 471218 116410 471454
rect 116646 471218 116688 471454
rect 116368 471134 116688 471218
rect 116368 470898 116410 471134
rect 116646 470898 116688 471134
rect 116368 470866 116688 470898
rect 147088 471454 147408 471486
rect 147088 471218 147130 471454
rect 147366 471218 147408 471454
rect 147088 471134 147408 471218
rect 147088 470898 147130 471134
rect 147366 470898 147408 471134
rect 147088 470866 147408 470898
rect 177808 471454 178128 471486
rect 177808 471218 177850 471454
rect 178086 471218 178128 471454
rect 177808 471134 178128 471218
rect 177808 470898 177850 471134
rect 178086 470898 178128 471134
rect 177808 470866 178128 470898
rect 208528 471454 208848 471486
rect 208528 471218 208570 471454
rect 208806 471218 208848 471454
rect 208528 471134 208848 471218
rect 208528 470898 208570 471134
rect 208806 470898 208848 471134
rect 208528 470866 208848 470898
rect 239248 471454 239568 471486
rect 239248 471218 239290 471454
rect 239526 471218 239568 471454
rect 239248 471134 239568 471218
rect 239248 470898 239290 471134
rect 239526 470898 239568 471134
rect 239248 470866 239568 470898
rect 269968 471454 270288 471486
rect 269968 471218 270010 471454
rect 270246 471218 270288 471454
rect 269968 471134 270288 471218
rect 269968 470898 270010 471134
rect 270246 470898 270288 471134
rect 269968 470866 270288 470898
rect 300688 471454 301008 471486
rect 300688 471218 300730 471454
rect 300966 471218 301008 471454
rect 300688 471134 301008 471218
rect 300688 470898 300730 471134
rect 300966 470898 301008 471134
rect 300688 470866 301008 470898
rect 331408 471454 331728 471486
rect 331408 471218 331450 471454
rect 331686 471218 331728 471454
rect 331408 471134 331728 471218
rect 331408 470898 331450 471134
rect 331686 470898 331728 471134
rect 331408 470866 331728 470898
rect 362128 471454 362448 471486
rect 362128 471218 362170 471454
rect 362406 471218 362448 471454
rect 362128 471134 362448 471218
rect 362128 470898 362170 471134
rect 362406 470898 362448 471134
rect 362128 470866 362448 470898
rect 63834 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 64454 461494
rect 63834 461174 64454 461258
rect 63834 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 64454 461174
rect 63834 425494 64454 460938
rect 376674 450334 377294 485778
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 377488 475174 377808 475206
rect 377488 474938 377530 475174
rect 377766 474938 377808 475174
rect 377488 474854 377808 474938
rect 377488 474618 377530 474854
rect 377766 474618 377808 474854
rect 377488 474586 377808 474618
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 70288 439174 70608 439206
rect 70288 438938 70330 439174
rect 70566 438938 70608 439174
rect 70288 438854 70608 438938
rect 70288 438618 70330 438854
rect 70566 438618 70608 438854
rect 70288 438586 70608 438618
rect 101008 439174 101328 439206
rect 101008 438938 101050 439174
rect 101286 438938 101328 439174
rect 101008 438854 101328 438938
rect 101008 438618 101050 438854
rect 101286 438618 101328 438854
rect 101008 438586 101328 438618
rect 131728 439174 132048 439206
rect 131728 438938 131770 439174
rect 132006 438938 132048 439174
rect 131728 438854 132048 438938
rect 131728 438618 131770 438854
rect 132006 438618 132048 438854
rect 131728 438586 132048 438618
rect 162448 439174 162768 439206
rect 162448 438938 162490 439174
rect 162726 438938 162768 439174
rect 162448 438854 162768 438938
rect 162448 438618 162490 438854
rect 162726 438618 162768 438854
rect 162448 438586 162768 438618
rect 193168 439174 193488 439206
rect 193168 438938 193210 439174
rect 193446 438938 193488 439174
rect 193168 438854 193488 438938
rect 193168 438618 193210 438854
rect 193446 438618 193488 438854
rect 193168 438586 193488 438618
rect 223888 439174 224208 439206
rect 223888 438938 223930 439174
rect 224166 438938 224208 439174
rect 223888 438854 224208 438938
rect 223888 438618 223930 438854
rect 224166 438618 224208 438854
rect 223888 438586 224208 438618
rect 254608 439174 254928 439206
rect 254608 438938 254650 439174
rect 254886 438938 254928 439174
rect 254608 438854 254928 438938
rect 254608 438618 254650 438854
rect 254886 438618 254928 438854
rect 254608 438586 254928 438618
rect 285328 439174 285648 439206
rect 285328 438938 285370 439174
rect 285606 438938 285648 439174
rect 285328 438854 285648 438938
rect 285328 438618 285370 438854
rect 285606 438618 285648 438854
rect 285328 438586 285648 438618
rect 316048 439174 316368 439206
rect 316048 438938 316090 439174
rect 316326 438938 316368 439174
rect 316048 438854 316368 438938
rect 316048 438618 316090 438854
rect 316326 438618 316368 438854
rect 316048 438586 316368 438618
rect 346768 439174 347088 439206
rect 346768 438938 346810 439174
rect 347046 438938 347088 439174
rect 346768 438854 347088 438938
rect 346768 438618 346810 438854
rect 347046 438618 347088 438854
rect 346768 438586 347088 438618
rect 85648 435454 85968 435486
rect 85648 435218 85690 435454
rect 85926 435218 85968 435454
rect 85648 435134 85968 435218
rect 85648 434898 85690 435134
rect 85926 434898 85968 435134
rect 85648 434866 85968 434898
rect 116368 435454 116688 435486
rect 116368 435218 116410 435454
rect 116646 435218 116688 435454
rect 116368 435134 116688 435218
rect 116368 434898 116410 435134
rect 116646 434898 116688 435134
rect 116368 434866 116688 434898
rect 147088 435454 147408 435486
rect 147088 435218 147130 435454
rect 147366 435218 147408 435454
rect 147088 435134 147408 435218
rect 147088 434898 147130 435134
rect 147366 434898 147408 435134
rect 147088 434866 147408 434898
rect 177808 435454 178128 435486
rect 177808 435218 177850 435454
rect 178086 435218 178128 435454
rect 177808 435134 178128 435218
rect 177808 434898 177850 435134
rect 178086 434898 178128 435134
rect 177808 434866 178128 434898
rect 208528 435454 208848 435486
rect 208528 435218 208570 435454
rect 208806 435218 208848 435454
rect 208528 435134 208848 435218
rect 208528 434898 208570 435134
rect 208806 434898 208848 435134
rect 208528 434866 208848 434898
rect 239248 435454 239568 435486
rect 239248 435218 239290 435454
rect 239526 435218 239568 435454
rect 239248 435134 239568 435218
rect 239248 434898 239290 435134
rect 239526 434898 239568 435134
rect 239248 434866 239568 434898
rect 269968 435454 270288 435486
rect 269968 435218 270010 435454
rect 270246 435218 270288 435454
rect 269968 435134 270288 435218
rect 269968 434898 270010 435134
rect 270246 434898 270288 435134
rect 269968 434866 270288 434898
rect 300688 435454 301008 435486
rect 300688 435218 300730 435454
rect 300966 435218 301008 435454
rect 300688 435134 301008 435218
rect 300688 434898 300730 435134
rect 300966 434898 301008 435134
rect 300688 434866 301008 434898
rect 331408 435454 331728 435486
rect 331408 435218 331450 435454
rect 331686 435218 331728 435454
rect 331408 435134 331728 435218
rect 331408 434898 331450 435134
rect 331686 434898 331728 435134
rect 331408 434866 331728 434898
rect 362128 435454 362448 435486
rect 362128 435218 362170 435454
rect 362406 435218 362448 435454
rect 362128 435134 362448 435218
rect 362128 434898 362170 435134
rect 362406 434898 362448 435134
rect 362128 434866 362448 434898
rect 63834 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 64454 425494
rect 63834 425174 64454 425258
rect 63834 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 64454 425174
rect 63834 389494 64454 424938
rect 376674 414334 377294 449778
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 377488 439174 377808 439206
rect 377488 438938 377530 439174
rect 377766 438938 377808 439174
rect 377488 438854 377808 438938
rect 377488 438618 377530 438854
rect 377766 438618 377808 438854
rect 377488 438586 377808 438618
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 70288 403174 70608 403206
rect 70288 402938 70330 403174
rect 70566 402938 70608 403174
rect 70288 402854 70608 402938
rect 70288 402618 70330 402854
rect 70566 402618 70608 402854
rect 70288 402586 70608 402618
rect 101008 403174 101328 403206
rect 101008 402938 101050 403174
rect 101286 402938 101328 403174
rect 101008 402854 101328 402938
rect 101008 402618 101050 402854
rect 101286 402618 101328 402854
rect 101008 402586 101328 402618
rect 131728 403174 132048 403206
rect 131728 402938 131770 403174
rect 132006 402938 132048 403174
rect 131728 402854 132048 402938
rect 131728 402618 131770 402854
rect 132006 402618 132048 402854
rect 131728 402586 132048 402618
rect 162448 403174 162768 403206
rect 162448 402938 162490 403174
rect 162726 402938 162768 403174
rect 162448 402854 162768 402938
rect 162448 402618 162490 402854
rect 162726 402618 162768 402854
rect 162448 402586 162768 402618
rect 193168 403174 193488 403206
rect 193168 402938 193210 403174
rect 193446 402938 193488 403174
rect 193168 402854 193488 402938
rect 193168 402618 193210 402854
rect 193446 402618 193488 402854
rect 193168 402586 193488 402618
rect 223888 403174 224208 403206
rect 223888 402938 223930 403174
rect 224166 402938 224208 403174
rect 223888 402854 224208 402938
rect 223888 402618 223930 402854
rect 224166 402618 224208 402854
rect 223888 402586 224208 402618
rect 254608 403174 254928 403206
rect 254608 402938 254650 403174
rect 254886 402938 254928 403174
rect 254608 402854 254928 402938
rect 254608 402618 254650 402854
rect 254886 402618 254928 402854
rect 254608 402586 254928 402618
rect 285328 403174 285648 403206
rect 285328 402938 285370 403174
rect 285606 402938 285648 403174
rect 285328 402854 285648 402938
rect 285328 402618 285370 402854
rect 285606 402618 285648 402854
rect 285328 402586 285648 402618
rect 316048 403174 316368 403206
rect 316048 402938 316090 403174
rect 316326 402938 316368 403174
rect 316048 402854 316368 402938
rect 316048 402618 316090 402854
rect 316326 402618 316368 402854
rect 316048 402586 316368 402618
rect 346768 403174 347088 403206
rect 346768 402938 346810 403174
rect 347046 402938 347088 403174
rect 346768 402854 347088 402938
rect 346768 402618 346810 402854
rect 347046 402618 347088 402854
rect 346768 402586 347088 402618
rect 85648 399454 85968 399486
rect 85648 399218 85690 399454
rect 85926 399218 85968 399454
rect 85648 399134 85968 399218
rect 85648 398898 85690 399134
rect 85926 398898 85968 399134
rect 85648 398866 85968 398898
rect 116368 399454 116688 399486
rect 116368 399218 116410 399454
rect 116646 399218 116688 399454
rect 116368 399134 116688 399218
rect 116368 398898 116410 399134
rect 116646 398898 116688 399134
rect 116368 398866 116688 398898
rect 147088 399454 147408 399486
rect 147088 399218 147130 399454
rect 147366 399218 147408 399454
rect 147088 399134 147408 399218
rect 147088 398898 147130 399134
rect 147366 398898 147408 399134
rect 147088 398866 147408 398898
rect 177808 399454 178128 399486
rect 177808 399218 177850 399454
rect 178086 399218 178128 399454
rect 177808 399134 178128 399218
rect 177808 398898 177850 399134
rect 178086 398898 178128 399134
rect 177808 398866 178128 398898
rect 208528 399454 208848 399486
rect 208528 399218 208570 399454
rect 208806 399218 208848 399454
rect 208528 399134 208848 399218
rect 208528 398898 208570 399134
rect 208806 398898 208848 399134
rect 208528 398866 208848 398898
rect 239248 399454 239568 399486
rect 239248 399218 239290 399454
rect 239526 399218 239568 399454
rect 239248 399134 239568 399218
rect 239248 398898 239290 399134
rect 239526 398898 239568 399134
rect 239248 398866 239568 398898
rect 269968 399454 270288 399486
rect 269968 399218 270010 399454
rect 270246 399218 270288 399454
rect 269968 399134 270288 399218
rect 269968 398898 270010 399134
rect 270246 398898 270288 399134
rect 269968 398866 270288 398898
rect 300688 399454 301008 399486
rect 300688 399218 300730 399454
rect 300966 399218 301008 399454
rect 300688 399134 301008 399218
rect 300688 398898 300730 399134
rect 300966 398898 301008 399134
rect 300688 398866 301008 398898
rect 331408 399454 331728 399486
rect 331408 399218 331450 399454
rect 331686 399218 331728 399454
rect 331408 399134 331728 399218
rect 331408 398898 331450 399134
rect 331686 398898 331728 399134
rect 331408 398866 331728 398898
rect 362128 399454 362448 399486
rect 362128 399218 362170 399454
rect 362406 399218 362448 399454
rect 362128 399134 362448 399218
rect 362128 398898 362170 399134
rect 362406 398898 362448 399134
rect 362128 398866 362448 398898
rect 63834 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 64454 389494
rect 63834 389174 64454 389258
rect 63834 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 64454 389174
rect 63834 353494 64454 388938
rect 376674 378334 377294 413778
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 377488 403174 377808 403206
rect 377488 402938 377530 403174
rect 377766 402938 377808 403174
rect 377488 402854 377808 402938
rect 377488 402618 377530 402854
rect 377766 402618 377808 402854
rect 377488 402586 377808 402618
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 70288 367174 70608 367206
rect 70288 366938 70330 367174
rect 70566 366938 70608 367174
rect 70288 366854 70608 366938
rect 70288 366618 70330 366854
rect 70566 366618 70608 366854
rect 70288 366586 70608 366618
rect 101008 367174 101328 367206
rect 101008 366938 101050 367174
rect 101286 366938 101328 367174
rect 101008 366854 101328 366938
rect 101008 366618 101050 366854
rect 101286 366618 101328 366854
rect 101008 366586 101328 366618
rect 131728 367174 132048 367206
rect 131728 366938 131770 367174
rect 132006 366938 132048 367174
rect 131728 366854 132048 366938
rect 131728 366618 131770 366854
rect 132006 366618 132048 366854
rect 131728 366586 132048 366618
rect 162448 367174 162768 367206
rect 162448 366938 162490 367174
rect 162726 366938 162768 367174
rect 162448 366854 162768 366938
rect 162448 366618 162490 366854
rect 162726 366618 162768 366854
rect 162448 366586 162768 366618
rect 193168 367174 193488 367206
rect 193168 366938 193210 367174
rect 193446 366938 193488 367174
rect 193168 366854 193488 366938
rect 193168 366618 193210 366854
rect 193446 366618 193488 366854
rect 193168 366586 193488 366618
rect 223888 367174 224208 367206
rect 223888 366938 223930 367174
rect 224166 366938 224208 367174
rect 223888 366854 224208 366938
rect 223888 366618 223930 366854
rect 224166 366618 224208 366854
rect 223888 366586 224208 366618
rect 254608 367174 254928 367206
rect 254608 366938 254650 367174
rect 254886 366938 254928 367174
rect 254608 366854 254928 366938
rect 254608 366618 254650 366854
rect 254886 366618 254928 366854
rect 254608 366586 254928 366618
rect 285328 367174 285648 367206
rect 285328 366938 285370 367174
rect 285606 366938 285648 367174
rect 285328 366854 285648 366938
rect 285328 366618 285370 366854
rect 285606 366618 285648 366854
rect 285328 366586 285648 366618
rect 316048 367174 316368 367206
rect 316048 366938 316090 367174
rect 316326 366938 316368 367174
rect 316048 366854 316368 366938
rect 316048 366618 316090 366854
rect 316326 366618 316368 366854
rect 316048 366586 316368 366618
rect 346768 367174 347088 367206
rect 346768 366938 346810 367174
rect 347046 366938 347088 367174
rect 346768 366854 347088 366938
rect 346768 366618 346810 366854
rect 347046 366618 347088 366854
rect 346768 366586 347088 366618
rect 85648 363454 85968 363486
rect 85648 363218 85690 363454
rect 85926 363218 85968 363454
rect 85648 363134 85968 363218
rect 85648 362898 85690 363134
rect 85926 362898 85968 363134
rect 85648 362866 85968 362898
rect 116368 363454 116688 363486
rect 116368 363218 116410 363454
rect 116646 363218 116688 363454
rect 116368 363134 116688 363218
rect 116368 362898 116410 363134
rect 116646 362898 116688 363134
rect 116368 362866 116688 362898
rect 147088 363454 147408 363486
rect 147088 363218 147130 363454
rect 147366 363218 147408 363454
rect 147088 363134 147408 363218
rect 147088 362898 147130 363134
rect 147366 362898 147408 363134
rect 147088 362866 147408 362898
rect 177808 363454 178128 363486
rect 177808 363218 177850 363454
rect 178086 363218 178128 363454
rect 177808 363134 178128 363218
rect 177808 362898 177850 363134
rect 178086 362898 178128 363134
rect 177808 362866 178128 362898
rect 208528 363454 208848 363486
rect 208528 363218 208570 363454
rect 208806 363218 208848 363454
rect 208528 363134 208848 363218
rect 208528 362898 208570 363134
rect 208806 362898 208848 363134
rect 208528 362866 208848 362898
rect 239248 363454 239568 363486
rect 239248 363218 239290 363454
rect 239526 363218 239568 363454
rect 239248 363134 239568 363218
rect 239248 362898 239290 363134
rect 239526 362898 239568 363134
rect 239248 362866 239568 362898
rect 269968 363454 270288 363486
rect 269968 363218 270010 363454
rect 270246 363218 270288 363454
rect 269968 363134 270288 363218
rect 269968 362898 270010 363134
rect 270246 362898 270288 363134
rect 269968 362866 270288 362898
rect 300688 363454 301008 363486
rect 300688 363218 300730 363454
rect 300966 363218 301008 363454
rect 300688 363134 301008 363218
rect 300688 362898 300730 363134
rect 300966 362898 301008 363134
rect 300688 362866 301008 362898
rect 331408 363454 331728 363486
rect 331408 363218 331450 363454
rect 331686 363218 331728 363454
rect 331408 363134 331728 363218
rect 331408 362898 331450 363134
rect 331686 362898 331728 363134
rect 331408 362866 331728 362898
rect 362128 363454 362448 363486
rect 362128 363218 362170 363454
rect 362406 363218 362448 363454
rect 362128 363134 362448 363218
rect 362128 362898 362170 363134
rect 362406 362898 362448 363134
rect 362128 362866 362448 362898
rect 63834 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 64454 353494
rect 63834 353174 64454 353258
rect 63834 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 64454 353174
rect 63834 317494 64454 352938
rect 376674 342334 377294 377778
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 377488 367174 377808 367206
rect 377488 366938 377530 367174
rect 377766 366938 377808 367174
rect 377488 366854 377808 366938
rect 377488 366618 377530 366854
rect 377766 366618 377808 366854
rect 377488 366586 377808 366618
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 70288 331174 70608 331206
rect 70288 330938 70330 331174
rect 70566 330938 70608 331174
rect 70288 330854 70608 330938
rect 70288 330618 70330 330854
rect 70566 330618 70608 330854
rect 70288 330586 70608 330618
rect 101008 331174 101328 331206
rect 101008 330938 101050 331174
rect 101286 330938 101328 331174
rect 101008 330854 101328 330938
rect 101008 330618 101050 330854
rect 101286 330618 101328 330854
rect 101008 330586 101328 330618
rect 131728 331174 132048 331206
rect 131728 330938 131770 331174
rect 132006 330938 132048 331174
rect 131728 330854 132048 330938
rect 131728 330618 131770 330854
rect 132006 330618 132048 330854
rect 131728 330586 132048 330618
rect 162448 331174 162768 331206
rect 162448 330938 162490 331174
rect 162726 330938 162768 331174
rect 162448 330854 162768 330938
rect 162448 330618 162490 330854
rect 162726 330618 162768 330854
rect 162448 330586 162768 330618
rect 193168 331174 193488 331206
rect 193168 330938 193210 331174
rect 193446 330938 193488 331174
rect 193168 330854 193488 330938
rect 193168 330618 193210 330854
rect 193446 330618 193488 330854
rect 193168 330586 193488 330618
rect 223888 331174 224208 331206
rect 223888 330938 223930 331174
rect 224166 330938 224208 331174
rect 223888 330854 224208 330938
rect 223888 330618 223930 330854
rect 224166 330618 224208 330854
rect 223888 330586 224208 330618
rect 254608 331174 254928 331206
rect 254608 330938 254650 331174
rect 254886 330938 254928 331174
rect 254608 330854 254928 330938
rect 254608 330618 254650 330854
rect 254886 330618 254928 330854
rect 254608 330586 254928 330618
rect 285328 331174 285648 331206
rect 285328 330938 285370 331174
rect 285606 330938 285648 331174
rect 285328 330854 285648 330938
rect 285328 330618 285370 330854
rect 285606 330618 285648 330854
rect 285328 330586 285648 330618
rect 316048 331174 316368 331206
rect 316048 330938 316090 331174
rect 316326 330938 316368 331174
rect 316048 330854 316368 330938
rect 316048 330618 316090 330854
rect 316326 330618 316368 330854
rect 316048 330586 316368 330618
rect 346768 331174 347088 331206
rect 346768 330938 346810 331174
rect 347046 330938 347088 331174
rect 346768 330854 347088 330938
rect 346768 330618 346810 330854
rect 347046 330618 347088 330854
rect 346768 330586 347088 330618
rect 85648 327454 85968 327486
rect 85648 327218 85690 327454
rect 85926 327218 85968 327454
rect 85648 327134 85968 327218
rect 85648 326898 85690 327134
rect 85926 326898 85968 327134
rect 85648 326866 85968 326898
rect 116368 327454 116688 327486
rect 116368 327218 116410 327454
rect 116646 327218 116688 327454
rect 116368 327134 116688 327218
rect 116368 326898 116410 327134
rect 116646 326898 116688 327134
rect 116368 326866 116688 326898
rect 147088 327454 147408 327486
rect 147088 327218 147130 327454
rect 147366 327218 147408 327454
rect 147088 327134 147408 327218
rect 147088 326898 147130 327134
rect 147366 326898 147408 327134
rect 147088 326866 147408 326898
rect 177808 327454 178128 327486
rect 177808 327218 177850 327454
rect 178086 327218 178128 327454
rect 177808 327134 178128 327218
rect 177808 326898 177850 327134
rect 178086 326898 178128 327134
rect 177808 326866 178128 326898
rect 208528 327454 208848 327486
rect 208528 327218 208570 327454
rect 208806 327218 208848 327454
rect 208528 327134 208848 327218
rect 208528 326898 208570 327134
rect 208806 326898 208848 327134
rect 208528 326866 208848 326898
rect 239248 327454 239568 327486
rect 239248 327218 239290 327454
rect 239526 327218 239568 327454
rect 239248 327134 239568 327218
rect 239248 326898 239290 327134
rect 239526 326898 239568 327134
rect 239248 326866 239568 326898
rect 269968 327454 270288 327486
rect 269968 327218 270010 327454
rect 270246 327218 270288 327454
rect 269968 327134 270288 327218
rect 269968 326898 270010 327134
rect 270246 326898 270288 327134
rect 269968 326866 270288 326898
rect 300688 327454 301008 327486
rect 300688 327218 300730 327454
rect 300966 327218 301008 327454
rect 300688 327134 301008 327218
rect 300688 326898 300730 327134
rect 300966 326898 301008 327134
rect 300688 326866 301008 326898
rect 331408 327454 331728 327486
rect 331408 327218 331450 327454
rect 331686 327218 331728 327454
rect 331408 327134 331728 327218
rect 331408 326898 331450 327134
rect 331686 326898 331728 327134
rect 331408 326866 331728 326898
rect 362128 327454 362448 327486
rect 362128 327218 362170 327454
rect 362406 327218 362448 327454
rect 362128 327134 362448 327218
rect 362128 326898 362170 327134
rect 362406 326898 362448 327134
rect 362128 326866 362448 326898
rect 63834 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 64454 317494
rect 63834 317174 64454 317258
rect 63834 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 64454 317174
rect 63834 281494 64454 316938
rect 376674 306334 377294 341778
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 377488 331174 377808 331206
rect 377488 330938 377530 331174
rect 377766 330938 377808 331174
rect 377488 330854 377808 330938
rect 377488 330618 377530 330854
rect 377766 330618 377808 330854
rect 377488 330586 377808 330618
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 70288 295174 70608 295206
rect 70288 294938 70330 295174
rect 70566 294938 70608 295174
rect 70288 294854 70608 294938
rect 70288 294618 70330 294854
rect 70566 294618 70608 294854
rect 70288 294586 70608 294618
rect 101008 295174 101328 295206
rect 101008 294938 101050 295174
rect 101286 294938 101328 295174
rect 101008 294854 101328 294938
rect 101008 294618 101050 294854
rect 101286 294618 101328 294854
rect 101008 294586 101328 294618
rect 131728 295174 132048 295206
rect 131728 294938 131770 295174
rect 132006 294938 132048 295174
rect 131728 294854 132048 294938
rect 131728 294618 131770 294854
rect 132006 294618 132048 294854
rect 131728 294586 132048 294618
rect 162448 295174 162768 295206
rect 162448 294938 162490 295174
rect 162726 294938 162768 295174
rect 162448 294854 162768 294938
rect 162448 294618 162490 294854
rect 162726 294618 162768 294854
rect 162448 294586 162768 294618
rect 193168 295174 193488 295206
rect 193168 294938 193210 295174
rect 193446 294938 193488 295174
rect 193168 294854 193488 294938
rect 193168 294618 193210 294854
rect 193446 294618 193488 294854
rect 193168 294586 193488 294618
rect 223888 295174 224208 295206
rect 223888 294938 223930 295174
rect 224166 294938 224208 295174
rect 223888 294854 224208 294938
rect 223888 294618 223930 294854
rect 224166 294618 224208 294854
rect 223888 294586 224208 294618
rect 254608 295174 254928 295206
rect 254608 294938 254650 295174
rect 254886 294938 254928 295174
rect 254608 294854 254928 294938
rect 254608 294618 254650 294854
rect 254886 294618 254928 294854
rect 254608 294586 254928 294618
rect 285328 295174 285648 295206
rect 285328 294938 285370 295174
rect 285606 294938 285648 295174
rect 285328 294854 285648 294938
rect 285328 294618 285370 294854
rect 285606 294618 285648 294854
rect 285328 294586 285648 294618
rect 316048 295174 316368 295206
rect 316048 294938 316090 295174
rect 316326 294938 316368 295174
rect 316048 294854 316368 294938
rect 316048 294618 316090 294854
rect 316326 294618 316368 294854
rect 316048 294586 316368 294618
rect 346768 295174 347088 295206
rect 346768 294938 346810 295174
rect 347046 294938 347088 295174
rect 346768 294854 347088 294938
rect 346768 294618 346810 294854
rect 347046 294618 347088 294854
rect 346768 294586 347088 294618
rect 85648 291454 85968 291486
rect 85648 291218 85690 291454
rect 85926 291218 85968 291454
rect 85648 291134 85968 291218
rect 85648 290898 85690 291134
rect 85926 290898 85968 291134
rect 85648 290866 85968 290898
rect 116368 291454 116688 291486
rect 116368 291218 116410 291454
rect 116646 291218 116688 291454
rect 116368 291134 116688 291218
rect 116368 290898 116410 291134
rect 116646 290898 116688 291134
rect 116368 290866 116688 290898
rect 147088 291454 147408 291486
rect 147088 291218 147130 291454
rect 147366 291218 147408 291454
rect 147088 291134 147408 291218
rect 147088 290898 147130 291134
rect 147366 290898 147408 291134
rect 147088 290866 147408 290898
rect 177808 291454 178128 291486
rect 177808 291218 177850 291454
rect 178086 291218 178128 291454
rect 177808 291134 178128 291218
rect 177808 290898 177850 291134
rect 178086 290898 178128 291134
rect 177808 290866 178128 290898
rect 208528 291454 208848 291486
rect 208528 291218 208570 291454
rect 208806 291218 208848 291454
rect 208528 291134 208848 291218
rect 208528 290898 208570 291134
rect 208806 290898 208848 291134
rect 208528 290866 208848 290898
rect 239248 291454 239568 291486
rect 239248 291218 239290 291454
rect 239526 291218 239568 291454
rect 239248 291134 239568 291218
rect 239248 290898 239290 291134
rect 239526 290898 239568 291134
rect 239248 290866 239568 290898
rect 269968 291454 270288 291486
rect 269968 291218 270010 291454
rect 270246 291218 270288 291454
rect 269968 291134 270288 291218
rect 269968 290898 270010 291134
rect 270246 290898 270288 291134
rect 269968 290866 270288 290898
rect 300688 291454 301008 291486
rect 300688 291218 300730 291454
rect 300966 291218 301008 291454
rect 300688 291134 301008 291218
rect 300688 290898 300730 291134
rect 300966 290898 301008 291134
rect 300688 290866 301008 290898
rect 331408 291454 331728 291486
rect 331408 291218 331450 291454
rect 331686 291218 331728 291454
rect 331408 291134 331728 291218
rect 331408 290898 331450 291134
rect 331686 290898 331728 291134
rect 331408 290866 331728 290898
rect 362128 291454 362448 291486
rect 362128 291218 362170 291454
rect 362406 291218 362448 291454
rect 362128 291134 362448 291218
rect 362128 290898 362170 291134
rect 362406 290898 362448 291134
rect 362128 290866 362448 290898
rect 63834 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 64454 281494
rect 63834 281174 64454 281258
rect 63834 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 64454 281174
rect 63834 245494 64454 280938
rect 376674 270334 377294 305778
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 377488 295174 377808 295206
rect 377488 294938 377530 295174
rect 377766 294938 377808 295174
rect 377488 294854 377808 294938
rect 377488 294618 377530 294854
rect 377766 294618 377808 294854
rect 377488 294586 377808 294618
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 70288 259174 70608 259206
rect 70288 258938 70330 259174
rect 70566 258938 70608 259174
rect 70288 258854 70608 258938
rect 70288 258618 70330 258854
rect 70566 258618 70608 258854
rect 70288 258586 70608 258618
rect 101008 259174 101328 259206
rect 101008 258938 101050 259174
rect 101286 258938 101328 259174
rect 101008 258854 101328 258938
rect 101008 258618 101050 258854
rect 101286 258618 101328 258854
rect 101008 258586 101328 258618
rect 131728 259174 132048 259206
rect 131728 258938 131770 259174
rect 132006 258938 132048 259174
rect 131728 258854 132048 258938
rect 131728 258618 131770 258854
rect 132006 258618 132048 258854
rect 131728 258586 132048 258618
rect 162448 259174 162768 259206
rect 162448 258938 162490 259174
rect 162726 258938 162768 259174
rect 162448 258854 162768 258938
rect 162448 258618 162490 258854
rect 162726 258618 162768 258854
rect 162448 258586 162768 258618
rect 193168 259174 193488 259206
rect 193168 258938 193210 259174
rect 193446 258938 193488 259174
rect 193168 258854 193488 258938
rect 193168 258618 193210 258854
rect 193446 258618 193488 258854
rect 193168 258586 193488 258618
rect 223888 259174 224208 259206
rect 223888 258938 223930 259174
rect 224166 258938 224208 259174
rect 223888 258854 224208 258938
rect 223888 258618 223930 258854
rect 224166 258618 224208 258854
rect 223888 258586 224208 258618
rect 254608 259174 254928 259206
rect 254608 258938 254650 259174
rect 254886 258938 254928 259174
rect 254608 258854 254928 258938
rect 254608 258618 254650 258854
rect 254886 258618 254928 258854
rect 254608 258586 254928 258618
rect 285328 259174 285648 259206
rect 285328 258938 285370 259174
rect 285606 258938 285648 259174
rect 285328 258854 285648 258938
rect 285328 258618 285370 258854
rect 285606 258618 285648 258854
rect 285328 258586 285648 258618
rect 316048 259174 316368 259206
rect 316048 258938 316090 259174
rect 316326 258938 316368 259174
rect 316048 258854 316368 258938
rect 316048 258618 316090 258854
rect 316326 258618 316368 258854
rect 316048 258586 316368 258618
rect 346768 259174 347088 259206
rect 346768 258938 346810 259174
rect 347046 258938 347088 259174
rect 346768 258854 347088 258938
rect 346768 258618 346810 258854
rect 347046 258618 347088 258854
rect 346768 258586 347088 258618
rect 85648 255454 85968 255486
rect 85648 255218 85690 255454
rect 85926 255218 85968 255454
rect 85648 255134 85968 255218
rect 85648 254898 85690 255134
rect 85926 254898 85968 255134
rect 85648 254866 85968 254898
rect 116368 255454 116688 255486
rect 116368 255218 116410 255454
rect 116646 255218 116688 255454
rect 116368 255134 116688 255218
rect 116368 254898 116410 255134
rect 116646 254898 116688 255134
rect 116368 254866 116688 254898
rect 147088 255454 147408 255486
rect 147088 255218 147130 255454
rect 147366 255218 147408 255454
rect 147088 255134 147408 255218
rect 147088 254898 147130 255134
rect 147366 254898 147408 255134
rect 147088 254866 147408 254898
rect 177808 255454 178128 255486
rect 177808 255218 177850 255454
rect 178086 255218 178128 255454
rect 177808 255134 178128 255218
rect 177808 254898 177850 255134
rect 178086 254898 178128 255134
rect 177808 254866 178128 254898
rect 208528 255454 208848 255486
rect 208528 255218 208570 255454
rect 208806 255218 208848 255454
rect 208528 255134 208848 255218
rect 208528 254898 208570 255134
rect 208806 254898 208848 255134
rect 208528 254866 208848 254898
rect 239248 255454 239568 255486
rect 239248 255218 239290 255454
rect 239526 255218 239568 255454
rect 239248 255134 239568 255218
rect 239248 254898 239290 255134
rect 239526 254898 239568 255134
rect 239248 254866 239568 254898
rect 269968 255454 270288 255486
rect 269968 255218 270010 255454
rect 270246 255218 270288 255454
rect 269968 255134 270288 255218
rect 269968 254898 270010 255134
rect 270246 254898 270288 255134
rect 269968 254866 270288 254898
rect 300688 255454 301008 255486
rect 300688 255218 300730 255454
rect 300966 255218 301008 255454
rect 300688 255134 301008 255218
rect 300688 254898 300730 255134
rect 300966 254898 301008 255134
rect 300688 254866 301008 254898
rect 331408 255454 331728 255486
rect 331408 255218 331450 255454
rect 331686 255218 331728 255454
rect 331408 255134 331728 255218
rect 331408 254898 331450 255134
rect 331686 254898 331728 255134
rect 331408 254866 331728 254898
rect 362128 255454 362448 255486
rect 362128 255218 362170 255454
rect 362406 255218 362448 255454
rect 362128 255134 362448 255218
rect 362128 254898 362170 255134
rect 362406 254898 362448 255134
rect 362128 254866 362448 254898
rect 63834 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 64454 245494
rect 63834 245174 64454 245258
rect 63834 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 64454 245174
rect 63834 209494 64454 244938
rect 376674 234334 377294 269778
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 377488 259174 377808 259206
rect 377488 258938 377530 259174
rect 377766 258938 377808 259174
rect 377488 258854 377808 258938
rect 377488 258618 377530 258854
rect 377766 258618 377808 258854
rect 377488 258586 377808 258618
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 70288 223174 70608 223206
rect 70288 222938 70330 223174
rect 70566 222938 70608 223174
rect 70288 222854 70608 222938
rect 70288 222618 70330 222854
rect 70566 222618 70608 222854
rect 70288 222586 70608 222618
rect 101008 223174 101328 223206
rect 101008 222938 101050 223174
rect 101286 222938 101328 223174
rect 101008 222854 101328 222938
rect 101008 222618 101050 222854
rect 101286 222618 101328 222854
rect 101008 222586 101328 222618
rect 131728 223174 132048 223206
rect 131728 222938 131770 223174
rect 132006 222938 132048 223174
rect 131728 222854 132048 222938
rect 131728 222618 131770 222854
rect 132006 222618 132048 222854
rect 131728 222586 132048 222618
rect 162448 223174 162768 223206
rect 162448 222938 162490 223174
rect 162726 222938 162768 223174
rect 162448 222854 162768 222938
rect 162448 222618 162490 222854
rect 162726 222618 162768 222854
rect 162448 222586 162768 222618
rect 193168 223174 193488 223206
rect 193168 222938 193210 223174
rect 193446 222938 193488 223174
rect 193168 222854 193488 222938
rect 193168 222618 193210 222854
rect 193446 222618 193488 222854
rect 193168 222586 193488 222618
rect 223888 223174 224208 223206
rect 223888 222938 223930 223174
rect 224166 222938 224208 223174
rect 223888 222854 224208 222938
rect 223888 222618 223930 222854
rect 224166 222618 224208 222854
rect 223888 222586 224208 222618
rect 254608 223174 254928 223206
rect 254608 222938 254650 223174
rect 254886 222938 254928 223174
rect 254608 222854 254928 222938
rect 254608 222618 254650 222854
rect 254886 222618 254928 222854
rect 254608 222586 254928 222618
rect 285328 223174 285648 223206
rect 285328 222938 285370 223174
rect 285606 222938 285648 223174
rect 285328 222854 285648 222938
rect 285328 222618 285370 222854
rect 285606 222618 285648 222854
rect 285328 222586 285648 222618
rect 316048 223174 316368 223206
rect 316048 222938 316090 223174
rect 316326 222938 316368 223174
rect 316048 222854 316368 222938
rect 316048 222618 316090 222854
rect 316326 222618 316368 222854
rect 316048 222586 316368 222618
rect 346768 223174 347088 223206
rect 346768 222938 346810 223174
rect 347046 222938 347088 223174
rect 346768 222854 347088 222938
rect 346768 222618 346810 222854
rect 347046 222618 347088 222854
rect 346768 222586 347088 222618
rect 85648 219454 85968 219486
rect 85648 219218 85690 219454
rect 85926 219218 85968 219454
rect 85648 219134 85968 219218
rect 85648 218898 85690 219134
rect 85926 218898 85968 219134
rect 85648 218866 85968 218898
rect 116368 219454 116688 219486
rect 116368 219218 116410 219454
rect 116646 219218 116688 219454
rect 116368 219134 116688 219218
rect 116368 218898 116410 219134
rect 116646 218898 116688 219134
rect 116368 218866 116688 218898
rect 147088 219454 147408 219486
rect 147088 219218 147130 219454
rect 147366 219218 147408 219454
rect 147088 219134 147408 219218
rect 147088 218898 147130 219134
rect 147366 218898 147408 219134
rect 147088 218866 147408 218898
rect 177808 219454 178128 219486
rect 177808 219218 177850 219454
rect 178086 219218 178128 219454
rect 177808 219134 178128 219218
rect 177808 218898 177850 219134
rect 178086 218898 178128 219134
rect 177808 218866 178128 218898
rect 208528 219454 208848 219486
rect 208528 219218 208570 219454
rect 208806 219218 208848 219454
rect 208528 219134 208848 219218
rect 208528 218898 208570 219134
rect 208806 218898 208848 219134
rect 208528 218866 208848 218898
rect 239248 219454 239568 219486
rect 239248 219218 239290 219454
rect 239526 219218 239568 219454
rect 239248 219134 239568 219218
rect 239248 218898 239290 219134
rect 239526 218898 239568 219134
rect 239248 218866 239568 218898
rect 269968 219454 270288 219486
rect 269968 219218 270010 219454
rect 270246 219218 270288 219454
rect 269968 219134 270288 219218
rect 269968 218898 270010 219134
rect 270246 218898 270288 219134
rect 269968 218866 270288 218898
rect 300688 219454 301008 219486
rect 300688 219218 300730 219454
rect 300966 219218 301008 219454
rect 300688 219134 301008 219218
rect 300688 218898 300730 219134
rect 300966 218898 301008 219134
rect 300688 218866 301008 218898
rect 331408 219454 331728 219486
rect 331408 219218 331450 219454
rect 331686 219218 331728 219454
rect 331408 219134 331728 219218
rect 331408 218898 331450 219134
rect 331686 218898 331728 219134
rect 331408 218866 331728 218898
rect 362128 219454 362448 219486
rect 362128 219218 362170 219454
rect 362406 219218 362448 219454
rect 362128 219134 362448 219218
rect 362128 218898 362170 219134
rect 362406 218898 362448 219134
rect 362128 218866 362448 218898
rect 63834 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 64454 209494
rect 63834 209174 64454 209258
rect 63834 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 64454 209174
rect 63834 173494 64454 208938
rect 376674 198334 377294 233778
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 377488 223174 377808 223206
rect 377488 222938 377530 223174
rect 377766 222938 377808 223174
rect 377488 222854 377808 222938
rect 377488 222618 377530 222854
rect 377766 222618 377808 222854
rect 377488 222586 377808 222618
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 70288 187174 70608 187206
rect 70288 186938 70330 187174
rect 70566 186938 70608 187174
rect 70288 186854 70608 186938
rect 70288 186618 70330 186854
rect 70566 186618 70608 186854
rect 70288 186586 70608 186618
rect 101008 187174 101328 187206
rect 101008 186938 101050 187174
rect 101286 186938 101328 187174
rect 101008 186854 101328 186938
rect 101008 186618 101050 186854
rect 101286 186618 101328 186854
rect 101008 186586 101328 186618
rect 131728 187174 132048 187206
rect 131728 186938 131770 187174
rect 132006 186938 132048 187174
rect 131728 186854 132048 186938
rect 131728 186618 131770 186854
rect 132006 186618 132048 186854
rect 131728 186586 132048 186618
rect 162448 187174 162768 187206
rect 162448 186938 162490 187174
rect 162726 186938 162768 187174
rect 162448 186854 162768 186938
rect 162448 186618 162490 186854
rect 162726 186618 162768 186854
rect 162448 186586 162768 186618
rect 193168 187174 193488 187206
rect 193168 186938 193210 187174
rect 193446 186938 193488 187174
rect 193168 186854 193488 186938
rect 193168 186618 193210 186854
rect 193446 186618 193488 186854
rect 193168 186586 193488 186618
rect 223888 187174 224208 187206
rect 223888 186938 223930 187174
rect 224166 186938 224208 187174
rect 223888 186854 224208 186938
rect 223888 186618 223930 186854
rect 224166 186618 224208 186854
rect 223888 186586 224208 186618
rect 254608 187174 254928 187206
rect 254608 186938 254650 187174
rect 254886 186938 254928 187174
rect 254608 186854 254928 186938
rect 254608 186618 254650 186854
rect 254886 186618 254928 186854
rect 254608 186586 254928 186618
rect 285328 187174 285648 187206
rect 285328 186938 285370 187174
rect 285606 186938 285648 187174
rect 285328 186854 285648 186938
rect 285328 186618 285370 186854
rect 285606 186618 285648 186854
rect 285328 186586 285648 186618
rect 316048 187174 316368 187206
rect 316048 186938 316090 187174
rect 316326 186938 316368 187174
rect 316048 186854 316368 186938
rect 316048 186618 316090 186854
rect 316326 186618 316368 186854
rect 316048 186586 316368 186618
rect 346768 187174 347088 187206
rect 346768 186938 346810 187174
rect 347046 186938 347088 187174
rect 346768 186854 347088 186938
rect 346768 186618 346810 186854
rect 347046 186618 347088 186854
rect 346768 186586 347088 186618
rect 85648 183454 85968 183486
rect 85648 183218 85690 183454
rect 85926 183218 85968 183454
rect 85648 183134 85968 183218
rect 85648 182898 85690 183134
rect 85926 182898 85968 183134
rect 85648 182866 85968 182898
rect 116368 183454 116688 183486
rect 116368 183218 116410 183454
rect 116646 183218 116688 183454
rect 116368 183134 116688 183218
rect 116368 182898 116410 183134
rect 116646 182898 116688 183134
rect 116368 182866 116688 182898
rect 147088 183454 147408 183486
rect 147088 183218 147130 183454
rect 147366 183218 147408 183454
rect 147088 183134 147408 183218
rect 147088 182898 147130 183134
rect 147366 182898 147408 183134
rect 147088 182866 147408 182898
rect 177808 183454 178128 183486
rect 177808 183218 177850 183454
rect 178086 183218 178128 183454
rect 177808 183134 178128 183218
rect 177808 182898 177850 183134
rect 178086 182898 178128 183134
rect 177808 182866 178128 182898
rect 208528 183454 208848 183486
rect 208528 183218 208570 183454
rect 208806 183218 208848 183454
rect 208528 183134 208848 183218
rect 208528 182898 208570 183134
rect 208806 182898 208848 183134
rect 208528 182866 208848 182898
rect 239248 183454 239568 183486
rect 239248 183218 239290 183454
rect 239526 183218 239568 183454
rect 239248 183134 239568 183218
rect 239248 182898 239290 183134
rect 239526 182898 239568 183134
rect 239248 182866 239568 182898
rect 269968 183454 270288 183486
rect 269968 183218 270010 183454
rect 270246 183218 270288 183454
rect 269968 183134 270288 183218
rect 269968 182898 270010 183134
rect 270246 182898 270288 183134
rect 269968 182866 270288 182898
rect 300688 183454 301008 183486
rect 300688 183218 300730 183454
rect 300966 183218 301008 183454
rect 300688 183134 301008 183218
rect 300688 182898 300730 183134
rect 300966 182898 301008 183134
rect 300688 182866 301008 182898
rect 331408 183454 331728 183486
rect 331408 183218 331450 183454
rect 331686 183218 331728 183454
rect 331408 183134 331728 183218
rect 331408 182898 331450 183134
rect 331686 182898 331728 183134
rect 331408 182866 331728 182898
rect 362128 183454 362448 183486
rect 362128 183218 362170 183454
rect 362406 183218 362448 183454
rect 362128 183134 362448 183218
rect 362128 182898 362170 183134
rect 362406 182898 362448 183134
rect 362128 182866 362448 182898
rect 63834 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 64454 173494
rect 63834 173174 64454 173258
rect 63834 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 64454 173174
rect 63834 137494 64454 172938
rect 376674 162334 377294 197778
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 377488 187174 377808 187206
rect 377488 186938 377530 187174
rect 377766 186938 377808 187174
rect 377488 186854 377808 186938
rect 377488 186618 377530 186854
rect 377766 186618 377808 186854
rect 377488 186586 377808 186618
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 70288 151174 70608 151206
rect 70288 150938 70330 151174
rect 70566 150938 70608 151174
rect 70288 150854 70608 150938
rect 70288 150618 70330 150854
rect 70566 150618 70608 150854
rect 70288 150586 70608 150618
rect 101008 151174 101328 151206
rect 101008 150938 101050 151174
rect 101286 150938 101328 151174
rect 101008 150854 101328 150938
rect 101008 150618 101050 150854
rect 101286 150618 101328 150854
rect 101008 150586 101328 150618
rect 131728 151174 132048 151206
rect 131728 150938 131770 151174
rect 132006 150938 132048 151174
rect 131728 150854 132048 150938
rect 131728 150618 131770 150854
rect 132006 150618 132048 150854
rect 131728 150586 132048 150618
rect 162448 151174 162768 151206
rect 162448 150938 162490 151174
rect 162726 150938 162768 151174
rect 162448 150854 162768 150938
rect 162448 150618 162490 150854
rect 162726 150618 162768 150854
rect 162448 150586 162768 150618
rect 193168 151174 193488 151206
rect 193168 150938 193210 151174
rect 193446 150938 193488 151174
rect 193168 150854 193488 150938
rect 193168 150618 193210 150854
rect 193446 150618 193488 150854
rect 193168 150586 193488 150618
rect 223888 151174 224208 151206
rect 223888 150938 223930 151174
rect 224166 150938 224208 151174
rect 223888 150854 224208 150938
rect 223888 150618 223930 150854
rect 224166 150618 224208 150854
rect 223888 150586 224208 150618
rect 254608 151174 254928 151206
rect 254608 150938 254650 151174
rect 254886 150938 254928 151174
rect 254608 150854 254928 150938
rect 254608 150618 254650 150854
rect 254886 150618 254928 150854
rect 254608 150586 254928 150618
rect 285328 151174 285648 151206
rect 285328 150938 285370 151174
rect 285606 150938 285648 151174
rect 285328 150854 285648 150938
rect 285328 150618 285370 150854
rect 285606 150618 285648 150854
rect 285328 150586 285648 150618
rect 316048 151174 316368 151206
rect 316048 150938 316090 151174
rect 316326 150938 316368 151174
rect 316048 150854 316368 150938
rect 316048 150618 316090 150854
rect 316326 150618 316368 150854
rect 316048 150586 316368 150618
rect 346768 151174 347088 151206
rect 346768 150938 346810 151174
rect 347046 150938 347088 151174
rect 346768 150854 347088 150938
rect 346768 150618 346810 150854
rect 347046 150618 347088 150854
rect 346768 150586 347088 150618
rect 85648 147454 85968 147486
rect 85648 147218 85690 147454
rect 85926 147218 85968 147454
rect 85648 147134 85968 147218
rect 85648 146898 85690 147134
rect 85926 146898 85968 147134
rect 85648 146866 85968 146898
rect 116368 147454 116688 147486
rect 116368 147218 116410 147454
rect 116646 147218 116688 147454
rect 116368 147134 116688 147218
rect 116368 146898 116410 147134
rect 116646 146898 116688 147134
rect 116368 146866 116688 146898
rect 147088 147454 147408 147486
rect 147088 147218 147130 147454
rect 147366 147218 147408 147454
rect 147088 147134 147408 147218
rect 147088 146898 147130 147134
rect 147366 146898 147408 147134
rect 147088 146866 147408 146898
rect 177808 147454 178128 147486
rect 177808 147218 177850 147454
rect 178086 147218 178128 147454
rect 177808 147134 178128 147218
rect 177808 146898 177850 147134
rect 178086 146898 178128 147134
rect 177808 146866 178128 146898
rect 208528 147454 208848 147486
rect 208528 147218 208570 147454
rect 208806 147218 208848 147454
rect 208528 147134 208848 147218
rect 208528 146898 208570 147134
rect 208806 146898 208848 147134
rect 208528 146866 208848 146898
rect 239248 147454 239568 147486
rect 239248 147218 239290 147454
rect 239526 147218 239568 147454
rect 239248 147134 239568 147218
rect 239248 146898 239290 147134
rect 239526 146898 239568 147134
rect 239248 146866 239568 146898
rect 269968 147454 270288 147486
rect 269968 147218 270010 147454
rect 270246 147218 270288 147454
rect 269968 147134 270288 147218
rect 269968 146898 270010 147134
rect 270246 146898 270288 147134
rect 269968 146866 270288 146898
rect 300688 147454 301008 147486
rect 300688 147218 300730 147454
rect 300966 147218 301008 147454
rect 300688 147134 301008 147218
rect 300688 146898 300730 147134
rect 300966 146898 301008 147134
rect 300688 146866 301008 146898
rect 331408 147454 331728 147486
rect 331408 147218 331450 147454
rect 331686 147218 331728 147454
rect 331408 147134 331728 147218
rect 331408 146898 331450 147134
rect 331686 146898 331728 147134
rect 331408 146866 331728 146898
rect 362128 147454 362448 147486
rect 362128 147218 362170 147454
rect 362406 147218 362448 147454
rect 362128 147134 362448 147218
rect 362128 146898 362170 147134
rect 362406 146898 362448 147134
rect 362128 146866 362448 146898
rect 63834 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 64454 137494
rect 63834 137174 64454 137258
rect 63834 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 64454 137174
rect 63834 101494 64454 136938
rect 376674 126334 377294 161778
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 377488 151174 377808 151206
rect 377488 150938 377530 151174
rect 377766 150938 377808 151174
rect 377488 150854 377808 150938
rect 377488 150618 377530 150854
rect 377766 150618 377808 150854
rect 377488 150586 377808 150618
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 70288 115174 70608 115206
rect 70288 114938 70330 115174
rect 70566 114938 70608 115174
rect 70288 114854 70608 114938
rect 70288 114618 70330 114854
rect 70566 114618 70608 114854
rect 70288 114586 70608 114618
rect 101008 115174 101328 115206
rect 101008 114938 101050 115174
rect 101286 114938 101328 115174
rect 101008 114854 101328 114938
rect 101008 114618 101050 114854
rect 101286 114618 101328 114854
rect 101008 114586 101328 114618
rect 131728 115174 132048 115206
rect 131728 114938 131770 115174
rect 132006 114938 132048 115174
rect 131728 114854 132048 114938
rect 131728 114618 131770 114854
rect 132006 114618 132048 114854
rect 131728 114586 132048 114618
rect 162448 115174 162768 115206
rect 162448 114938 162490 115174
rect 162726 114938 162768 115174
rect 162448 114854 162768 114938
rect 162448 114618 162490 114854
rect 162726 114618 162768 114854
rect 162448 114586 162768 114618
rect 193168 115174 193488 115206
rect 193168 114938 193210 115174
rect 193446 114938 193488 115174
rect 193168 114854 193488 114938
rect 193168 114618 193210 114854
rect 193446 114618 193488 114854
rect 193168 114586 193488 114618
rect 223888 115174 224208 115206
rect 223888 114938 223930 115174
rect 224166 114938 224208 115174
rect 223888 114854 224208 114938
rect 223888 114618 223930 114854
rect 224166 114618 224208 114854
rect 223888 114586 224208 114618
rect 254608 115174 254928 115206
rect 254608 114938 254650 115174
rect 254886 114938 254928 115174
rect 254608 114854 254928 114938
rect 254608 114618 254650 114854
rect 254886 114618 254928 114854
rect 254608 114586 254928 114618
rect 285328 115174 285648 115206
rect 285328 114938 285370 115174
rect 285606 114938 285648 115174
rect 285328 114854 285648 114938
rect 285328 114618 285370 114854
rect 285606 114618 285648 114854
rect 285328 114586 285648 114618
rect 316048 115174 316368 115206
rect 316048 114938 316090 115174
rect 316326 114938 316368 115174
rect 316048 114854 316368 114938
rect 316048 114618 316090 114854
rect 316326 114618 316368 114854
rect 316048 114586 316368 114618
rect 346768 115174 347088 115206
rect 346768 114938 346810 115174
rect 347046 114938 347088 115174
rect 346768 114854 347088 114938
rect 346768 114618 346810 114854
rect 347046 114618 347088 114854
rect 346768 114586 347088 114618
rect 85648 111454 85968 111486
rect 85648 111218 85690 111454
rect 85926 111218 85968 111454
rect 85648 111134 85968 111218
rect 85648 110898 85690 111134
rect 85926 110898 85968 111134
rect 85648 110866 85968 110898
rect 116368 111454 116688 111486
rect 116368 111218 116410 111454
rect 116646 111218 116688 111454
rect 116368 111134 116688 111218
rect 116368 110898 116410 111134
rect 116646 110898 116688 111134
rect 116368 110866 116688 110898
rect 147088 111454 147408 111486
rect 147088 111218 147130 111454
rect 147366 111218 147408 111454
rect 147088 111134 147408 111218
rect 147088 110898 147130 111134
rect 147366 110898 147408 111134
rect 147088 110866 147408 110898
rect 177808 111454 178128 111486
rect 177808 111218 177850 111454
rect 178086 111218 178128 111454
rect 177808 111134 178128 111218
rect 177808 110898 177850 111134
rect 178086 110898 178128 111134
rect 177808 110866 178128 110898
rect 208528 111454 208848 111486
rect 208528 111218 208570 111454
rect 208806 111218 208848 111454
rect 208528 111134 208848 111218
rect 208528 110898 208570 111134
rect 208806 110898 208848 111134
rect 208528 110866 208848 110898
rect 239248 111454 239568 111486
rect 239248 111218 239290 111454
rect 239526 111218 239568 111454
rect 239248 111134 239568 111218
rect 239248 110898 239290 111134
rect 239526 110898 239568 111134
rect 239248 110866 239568 110898
rect 269968 111454 270288 111486
rect 269968 111218 270010 111454
rect 270246 111218 270288 111454
rect 269968 111134 270288 111218
rect 269968 110898 270010 111134
rect 270246 110898 270288 111134
rect 269968 110866 270288 110898
rect 300688 111454 301008 111486
rect 300688 111218 300730 111454
rect 300966 111218 301008 111454
rect 300688 111134 301008 111218
rect 300688 110898 300730 111134
rect 300966 110898 301008 111134
rect 300688 110866 301008 110898
rect 331408 111454 331728 111486
rect 331408 111218 331450 111454
rect 331686 111218 331728 111454
rect 331408 111134 331728 111218
rect 331408 110898 331450 111134
rect 331686 110898 331728 111134
rect 331408 110866 331728 110898
rect 362128 111454 362448 111486
rect 362128 111218 362170 111454
rect 362406 111218 362448 111454
rect 362128 111134 362448 111218
rect 362128 110898 362170 111134
rect 362406 110898 362448 111134
rect 362128 110866 362448 110898
rect 63834 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 64454 101494
rect 63834 101174 64454 101258
rect 63834 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 64454 101174
rect 63834 65494 64454 100938
rect 376674 90334 377294 125778
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 377488 115174 377808 115206
rect 377488 114938 377530 115174
rect 377766 114938 377808 115174
rect 377488 114854 377808 114938
rect 377488 114618 377530 114854
rect 377766 114618 377808 114854
rect 377488 114586 377808 114618
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 70288 79174 70608 79206
rect 70288 78938 70330 79174
rect 70566 78938 70608 79174
rect 70288 78854 70608 78938
rect 70288 78618 70330 78854
rect 70566 78618 70608 78854
rect 70288 78586 70608 78618
rect 101008 79174 101328 79206
rect 101008 78938 101050 79174
rect 101286 78938 101328 79174
rect 101008 78854 101328 78938
rect 101008 78618 101050 78854
rect 101286 78618 101328 78854
rect 101008 78586 101328 78618
rect 131728 79174 132048 79206
rect 131728 78938 131770 79174
rect 132006 78938 132048 79174
rect 131728 78854 132048 78938
rect 131728 78618 131770 78854
rect 132006 78618 132048 78854
rect 131728 78586 132048 78618
rect 162448 79174 162768 79206
rect 162448 78938 162490 79174
rect 162726 78938 162768 79174
rect 162448 78854 162768 78938
rect 162448 78618 162490 78854
rect 162726 78618 162768 78854
rect 162448 78586 162768 78618
rect 193168 79174 193488 79206
rect 193168 78938 193210 79174
rect 193446 78938 193488 79174
rect 193168 78854 193488 78938
rect 193168 78618 193210 78854
rect 193446 78618 193488 78854
rect 193168 78586 193488 78618
rect 223888 79174 224208 79206
rect 223888 78938 223930 79174
rect 224166 78938 224208 79174
rect 223888 78854 224208 78938
rect 223888 78618 223930 78854
rect 224166 78618 224208 78854
rect 223888 78586 224208 78618
rect 254608 79174 254928 79206
rect 254608 78938 254650 79174
rect 254886 78938 254928 79174
rect 254608 78854 254928 78938
rect 254608 78618 254650 78854
rect 254886 78618 254928 78854
rect 254608 78586 254928 78618
rect 285328 79174 285648 79206
rect 285328 78938 285370 79174
rect 285606 78938 285648 79174
rect 285328 78854 285648 78938
rect 285328 78618 285370 78854
rect 285606 78618 285648 78854
rect 285328 78586 285648 78618
rect 316048 79174 316368 79206
rect 316048 78938 316090 79174
rect 316326 78938 316368 79174
rect 316048 78854 316368 78938
rect 316048 78618 316090 78854
rect 316326 78618 316368 78854
rect 316048 78586 316368 78618
rect 346768 79174 347088 79206
rect 346768 78938 346810 79174
rect 347046 78938 347088 79174
rect 346768 78854 347088 78938
rect 346768 78618 346810 78854
rect 347046 78618 347088 78854
rect 346768 78586 347088 78618
rect 85648 75454 85968 75486
rect 85648 75218 85690 75454
rect 85926 75218 85968 75454
rect 85648 75134 85968 75218
rect 85648 74898 85690 75134
rect 85926 74898 85968 75134
rect 85648 74866 85968 74898
rect 116368 75454 116688 75486
rect 116368 75218 116410 75454
rect 116646 75218 116688 75454
rect 116368 75134 116688 75218
rect 116368 74898 116410 75134
rect 116646 74898 116688 75134
rect 116368 74866 116688 74898
rect 147088 75454 147408 75486
rect 147088 75218 147130 75454
rect 147366 75218 147408 75454
rect 147088 75134 147408 75218
rect 147088 74898 147130 75134
rect 147366 74898 147408 75134
rect 147088 74866 147408 74898
rect 177808 75454 178128 75486
rect 177808 75218 177850 75454
rect 178086 75218 178128 75454
rect 177808 75134 178128 75218
rect 177808 74898 177850 75134
rect 178086 74898 178128 75134
rect 177808 74866 178128 74898
rect 208528 75454 208848 75486
rect 208528 75218 208570 75454
rect 208806 75218 208848 75454
rect 208528 75134 208848 75218
rect 208528 74898 208570 75134
rect 208806 74898 208848 75134
rect 208528 74866 208848 74898
rect 239248 75454 239568 75486
rect 239248 75218 239290 75454
rect 239526 75218 239568 75454
rect 239248 75134 239568 75218
rect 239248 74898 239290 75134
rect 239526 74898 239568 75134
rect 239248 74866 239568 74898
rect 269968 75454 270288 75486
rect 269968 75218 270010 75454
rect 270246 75218 270288 75454
rect 269968 75134 270288 75218
rect 269968 74898 270010 75134
rect 270246 74898 270288 75134
rect 269968 74866 270288 74898
rect 300688 75454 301008 75486
rect 300688 75218 300730 75454
rect 300966 75218 301008 75454
rect 300688 75134 301008 75218
rect 300688 74898 300730 75134
rect 300966 74898 301008 75134
rect 300688 74866 301008 74898
rect 331408 75454 331728 75486
rect 331408 75218 331450 75454
rect 331686 75218 331728 75454
rect 331408 75134 331728 75218
rect 331408 74898 331450 75134
rect 331686 74898 331728 75134
rect 331408 74866 331728 74898
rect 362128 75454 362448 75486
rect 362128 75218 362170 75454
rect 362406 75218 362448 75454
rect 362128 75134 362448 75218
rect 362128 74898 362170 75134
rect 362406 74898 362448 75134
rect 362128 74866 362448 74898
rect 63834 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 64454 65494
rect 63834 65174 64454 65258
rect 63834 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 64454 65174
rect 63834 29494 64454 64938
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 58855
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 58855
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 58855
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 50614 85574 58855
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 54334 89294 58855
rect 88674 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 89294 54334
rect 88674 54014 89294 54098
rect 88674 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 89294 54014
rect 88674 18334 89294 53778
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 58054 93014 58855
rect 92394 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 93014 58054
rect 92394 57734 93014 57818
rect 92394 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 93014 57734
rect 92394 22054 93014 57498
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 25774 96734 58855
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 29494 100454 58855
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 39454 110414 58855
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 43174 114134 58855
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 46894 117854 58855
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 50614 121574 58855
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 54334 125294 58855
rect 124674 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 125294 54334
rect 124674 54014 125294 54098
rect 124674 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 125294 54014
rect 124674 18334 125294 53778
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 58054 129014 58855
rect 128394 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 129014 58054
rect 128394 57734 129014 57818
rect 128394 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 129014 57734
rect 128394 22054 129014 57498
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 25774 132734 58855
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 29494 136454 58855
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 39454 146414 58855
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 43174 150134 58855
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 46894 153854 58855
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 50614 157574 58855
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 54334 161294 58855
rect 160674 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 161294 54334
rect 160674 54014 161294 54098
rect 160674 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 161294 54014
rect 160674 18334 161294 53778
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 58054 165014 58855
rect 164394 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 165014 58054
rect 164394 57734 165014 57818
rect 164394 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 165014 57734
rect 164394 22054 165014 57498
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 25774 168734 58855
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 29494 172454 58855
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 39454 182414 58855
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 43174 186134 58855
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 46894 189854 58855
rect 196674 54334 197294 58855
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 14614 193574 50068
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 18334 197294 53778
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 58054 201014 58855
rect 200394 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 201014 58054
rect 200394 57734 201014 57818
rect 200394 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 201014 57734
rect 200394 22054 201014 57498
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 25774 204734 58855
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 29494 208454 58855
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 39454 218414 58855
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 43174 222134 58855
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 46894 225854 58855
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 50614 229574 58855
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 54334 233294 58855
rect 232674 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 233294 54334
rect 232674 54014 233294 54098
rect 232674 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 233294 54014
rect 232674 18334 233294 53778
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 58054 237014 58855
rect 236394 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 237014 58054
rect 236394 57734 237014 57818
rect 236394 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 237014 57734
rect 236394 22054 237014 57498
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 25774 240734 58855
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 29494 244454 58855
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 39454 254414 58855
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 43174 258134 58855
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 46894 261854 58855
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 50614 265574 58855
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 54334 269294 58855
rect 268674 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 269294 54334
rect 268674 54014 269294 54098
rect 268674 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 269294 54014
rect 268674 18334 269294 53778
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 58054 273014 58855
rect 272394 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 273014 58054
rect 272394 57734 273014 57818
rect 272394 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 273014 57734
rect 272394 22054 273014 57498
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 25774 276734 58855
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 29494 280454 58855
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 39454 290414 58855
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 43174 294134 58855
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 46894 297854 58855
rect 304674 54334 305294 58855
rect 304674 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 305294 54334
rect 304674 54014 305294 54098
rect 304674 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 305294 54014
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 14614 301574 50068
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 18334 305294 53778
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 58054 309014 58855
rect 308394 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 309014 58054
rect 308394 57734 309014 57818
rect 308394 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 309014 57734
rect 308394 22054 309014 57498
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 25774 312734 58855
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 29494 316454 50068
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 39454 326414 58855
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 43174 330134 58855
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 46894 333854 58855
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 50614 337574 58855
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 54334 341294 58855
rect 340674 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 341294 54334
rect 340674 54014 341294 54098
rect 340674 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 341294 54014
rect 340674 18334 341294 53778
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 58054 345014 58855
rect 344394 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 345014 58054
rect 344394 57734 345014 57818
rect 344394 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 345014 57734
rect 344394 22054 345014 57498
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 25774 348734 58855
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 29494 352454 58855
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 39454 362414 50068
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 43174 366134 58855
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 46894 369854 58855
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 50614 373574 58855
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 54334 377294 89778
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 377488 79174 377808 79206
rect 377488 78938 377530 79174
rect 377766 78938 377808 79174
rect 377488 78854 377808 78938
rect 377488 78618 377530 78854
rect 377766 78618 377808 78854
rect 377488 78586 377808 78618
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 65494 388454 100938
rect 387834 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 388454 65494
rect 387834 65174 388454 65258
rect 387834 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 388454 65174
rect 387834 29494 388454 64938
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 404658 327454 404978 327486
rect 404658 327218 404700 327454
rect 404936 327218 404978 327454
rect 404658 327134 404978 327218
rect 404658 326898 404700 327134
rect 404936 326898 404978 327134
rect 404658 326866 404978 326898
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 298894 405854 334338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408372 331174 408692 331206
rect 408372 330938 408414 331174
rect 408650 330938 408692 331174
rect 408372 330854 408692 330938
rect 408372 330618 408414 330854
rect 408650 330618 408692 330854
rect 408372 330586 408692 330618
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 302614 409574 338058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 412086 327454 412406 327486
rect 412086 327218 412128 327454
rect 412364 327218 412406 327454
rect 412086 327134 412406 327218
rect 412086 326898 412128 327134
rect 412364 326898 412406 327134
rect 412086 326866 412406 326898
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 306334 413294 341778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 416394 454054 417014 489498
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 415800 331174 416120 331206
rect 415800 330938 415842 331174
rect 416078 330938 416120 331174
rect 415800 330854 416120 330938
rect 415800 330618 415842 330854
rect 416078 330618 416120 330854
rect 415800 330586 416120 330618
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 416394 310054 417014 345498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 493774 420734 529218
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 420114 421774 420734 457218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 497494 424454 532938
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 444412 424454 460938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 442833 434414 470898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 444412 438134 474618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444235 700500 444301 700501
rect 444235 700436 444236 700500
rect 444300 700436 444301 700500
rect 444235 700435 444301 700436
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442833 441854 478338
rect 426624 439174 426944 439206
rect 426624 438938 426666 439174
rect 426902 438938 426944 439174
rect 426624 438854 426944 438938
rect 426624 438618 426666 438854
rect 426902 438618 426944 438854
rect 426624 438586 426944 438618
rect 432305 439174 432625 439206
rect 432305 438938 432347 439174
rect 432583 438938 432625 439174
rect 432305 438854 432625 438938
rect 432305 438618 432347 438854
rect 432583 438618 432625 438854
rect 432305 438586 432625 438618
rect 437986 439174 438306 439206
rect 437986 438938 438028 439174
rect 438264 438938 438306 439174
rect 437986 438854 438306 438938
rect 437986 438618 438028 438854
rect 438264 438618 438306 438854
rect 437986 438586 438306 438618
rect 443667 439174 443987 439206
rect 443667 438938 443709 439174
rect 443945 438938 443987 439174
rect 443667 438854 443987 438938
rect 443667 438618 443709 438854
rect 443945 438618 443987 438854
rect 443667 438586 443987 438618
rect 423784 435454 424104 435486
rect 423784 435218 423826 435454
rect 424062 435218 424104 435454
rect 423784 435134 424104 435218
rect 423784 434898 423826 435134
rect 424062 434898 424104 435134
rect 423784 434866 424104 434898
rect 429465 435454 429785 435486
rect 429465 435218 429507 435454
rect 429743 435218 429785 435454
rect 429465 435134 429785 435218
rect 429465 434898 429507 435134
rect 429743 434898 429785 435134
rect 429465 434866 429785 434898
rect 435146 435454 435466 435486
rect 435146 435218 435188 435454
rect 435424 435218 435466 435454
rect 435146 435134 435466 435218
rect 435146 434898 435188 435134
rect 435424 434898 435466 435134
rect 435146 434866 435466 434898
rect 440827 435454 441147 435486
rect 440827 435218 440869 435454
rect 441105 435218 441147 435454
rect 440827 435134 441147 435218
rect 440827 434898 440869 435134
rect 441105 434898 441147 435134
rect 440827 434866 441147 434898
rect 420114 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 420734 421774
rect 420114 421454 420734 421538
rect 420114 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 420734 421454
rect 420114 385774 420734 421218
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 419514 327454 419834 327486
rect 419514 327218 419556 327454
rect 419792 327218 419834 327454
rect 419514 327134 419834 327218
rect 419514 326898 419556 327134
rect 419792 326898 419834 327134
rect 419514 326866 419834 326898
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 163505 417014 165498
rect 420114 313774 420734 349218
rect 423834 389494 424454 420068
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 423834 353494 424454 388938
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 422891 336836 422957 336837
rect 422891 336772 422892 336836
rect 422956 336772 422957 336836
rect 422891 336771 422957 336772
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 169774 420734 205218
rect 422894 171150 422954 336771
rect 423228 331174 423548 331206
rect 423228 330938 423270 331174
rect 423506 330938 423548 331174
rect 423228 330854 423548 330938
rect 423228 330618 423270 330854
rect 423506 330618 423548 330854
rect 423228 330586 423548 330618
rect 423834 317494 424454 352938
rect 433794 399454 434414 422599
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 430656 331174 430976 331206
rect 430656 330938 430698 331174
rect 430934 330938 430976 331174
rect 430656 330854 430976 330938
rect 430656 330618 430698 330854
rect 430934 330618 430976 330854
rect 430656 330586 430976 330618
rect 426942 327454 427262 327486
rect 426942 327218 426984 327454
rect 427220 327218 427262 327454
rect 426942 327134 427262 327218
rect 426942 326898 426984 327134
rect 427220 326898 427262 327134
rect 426942 326866 427262 326898
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 173494 424454 208938
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 422894 171090 423322 171150
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 163505 420734 169218
rect 423262 164389 423322 171090
rect 423259 164388 423325 164389
rect 423259 164324 423260 164388
rect 423324 164324 423325 164388
rect 423259 164323 423325 164324
rect 423262 163437 423322 164323
rect 423834 163505 424454 172938
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 163505 434414 182898
rect 437514 403174 438134 420068
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 163505 438134 186618
rect 441234 406894 441854 422599
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 444238 319701 444298 700435
rect 444954 698614 445574 707162
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 447915 700636 447981 700637
rect 447915 700572 447916 700636
rect 447980 700572 447981 700636
rect 447915 700571 447981 700572
rect 447731 700364 447797 700365
rect 447731 700300 447732 700364
rect 447796 700300 447797 700364
rect 447731 700299 447797 700300
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 446259 668676 446325 668677
rect 446259 668612 446260 668676
rect 446324 668612 446325 668676
rect 446259 668611 446325 668612
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444235 319700 444301 319701
rect 444235 319636 444236 319700
rect 444300 319636 444301 319700
rect 444235 319635 444301 319636
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 163505 441854 190338
rect 444954 302614 445574 338058
rect 446262 318341 446322 668611
rect 447734 319973 447794 700299
rect 447731 319972 447797 319973
rect 447731 319908 447732 319972
rect 447796 319908 447797 319972
rect 447731 319907 447797 319908
rect 447918 319837 447978 700571
rect 448099 671396 448165 671397
rect 448099 671332 448100 671396
rect 448164 671332 448165 671396
rect 448099 671331 448165 671332
rect 447915 319836 447981 319837
rect 447915 319772 447916 319836
rect 447980 319772 447981 319836
rect 447915 319771 447981 319772
rect 448102 318477 448162 671331
rect 448674 666334 449294 708122
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522334 449294 557778
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 448674 486334 449294 521778
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 517884 453014 525498
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 457851 675748 457917 675749
rect 457851 675684 457852 675748
rect 457916 675684 457917 675748
rect 457851 675683 457917 675684
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 457854 537437 457914 675683
rect 458035 672892 458101 672893
rect 458035 672828 458036 672892
rect 458100 672828 458101 672892
rect 458035 672827 458101 672828
rect 457851 537436 457917 537437
rect 457851 537372 457852 537436
rect 457916 537372 457917 537436
rect 457851 537371 457917 537372
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 517884 456734 529218
rect 458038 520981 458098 672827
rect 459834 665809 460454 676938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 665809 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 665809 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 665809 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 665809 481574 698058
rect 484674 708678 485294 711590
rect 484674 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 485294 708678
rect 484674 708358 485294 708442
rect 484674 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 485294 708358
rect 484674 665809 485294 708122
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 665809 489014 669498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 665809 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 665809 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 665809 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 665809 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 665809 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 665809 517574 698058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 665809 521294 708122
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 665809 525014 669498
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 479568 655174 479888 655206
rect 479568 654938 479610 655174
rect 479846 654938 479888 655174
rect 479568 654854 479888 654938
rect 479568 654618 479610 654854
rect 479846 654618 479888 654854
rect 479568 654586 479888 654618
rect 510288 655174 510608 655206
rect 510288 654938 510330 655174
rect 510566 654938 510608 655174
rect 510288 654854 510608 654938
rect 510288 654618 510330 654854
rect 510566 654618 510608 654854
rect 510288 654586 510608 654618
rect 464208 651454 464528 651486
rect 464208 651218 464250 651454
rect 464486 651218 464528 651454
rect 464208 651134 464528 651218
rect 464208 650898 464250 651134
rect 464486 650898 464528 651134
rect 464208 650866 464528 650898
rect 494928 651454 495248 651486
rect 494928 651218 494970 651454
rect 495206 651218 495248 651454
rect 494928 651134 495248 651218
rect 494928 650898 494970 651134
rect 495206 650898 495248 651134
rect 494928 650866 495248 650898
rect 525648 651454 525968 651486
rect 525648 651218 525690 651454
rect 525926 651218 525968 651454
rect 525648 651134 525968 651218
rect 525648 650898 525690 651134
rect 525926 650898 525968 651134
rect 525648 650866 525968 650898
rect 528114 637774 528734 673218
rect 528114 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 528734 637774
rect 528114 637454 528734 637538
rect 528114 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 528734 637454
rect 459139 635764 459205 635765
rect 459139 635700 459140 635764
rect 459204 635700 459205 635764
rect 459139 635699 459205 635700
rect 458035 520980 458101 520981
rect 458035 520916 458036 520980
rect 458100 520916 458101 520980
rect 458035 520915 458101 520916
rect 451043 516764 451109 516765
rect 451043 516700 451044 516764
rect 451108 516700 451109 516764
rect 451043 516699 451109 516700
rect 450491 514384 450557 514385
rect 450491 514320 450492 514384
rect 450556 514320 450557 514384
rect 450491 514319 450557 514320
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448674 414334 449294 449778
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 448674 378334 449294 413778
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 448283 329628 448349 329629
rect 448283 329564 448284 329628
rect 448348 329564 448349 329628
rect 448283 329563 448349 329564
rect 448099 318476 448165 318477
rect 448099 318412 448100 318476
rect 448164 318412 448165 318476
rect 448099 318411 448165 318412
rect 446259 318340 446325 318341
rect 446259 318276 446260 318340
rect 446324 318276 446325 318340
rect 446259 318275 446325 318276
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 164540 445574 194058
rect 448286 164117 448346 329563
rect 448674 306334 449294 341778
rect 450494 327725 450554 514319
rect 451046 335370 451106 516699
rect 453382 511174 453702 511206
rect 453382 510938 453424 511174
rect 453660 510938 453702 511174
rect 453382 510854 453702 510938
rect 453382 510618 453424 510854
rect 453660 510618 453702 510854
rect 453382 510586 453702 510618
rect 455820 511174 456140 511206
rect 455820 510938 455862 511174
rect 456098 510938 456140 511174
rect 455820 510854 456140 510938
rect 455820 510618 455862 510854
rect 456098 510618 456140 510854
rect 455820 510586 456140 510618
rect 458258 511174 458578 511206
rect 458258 510938 458300 511174
rect 458536 510938 458578 511174
rect 458258 510854 458578 510938
rect 458258 510618 458300 510854
rect 458536 510618 458578 510854
rect 458258 510586 458578 510618
rect 452163 507454 452483 507486
rect 452163 507218 452205 507454
rect 452441 507218 452483 507454
rect 452163 507134 452483 507218
rect 452163 506898 452205 507134
rect 452441 506898 452483 507134
rect 452163 506866 452483 506898
rect 454601 507454 454921 507486
rect 454601 507218 454643 507454
rect 454879 507218 454921 507454
rect 454601 507134 454921 507218
rect 454601 506898 454643 507134
rect 454879 506898 454921 507134
rect 454601 506866 454921 506898
rect 457039 507454 457359 507486
rect 457039 507218 457081 507454
rect 457317 507218 457359 507454
rect 457039 507134 457359 507218
rect 457039 506898 457081 507134
rect 457317 506898 457359 507134
rect 457039 506866 457359 506898
rect 450678 335310 451106 335370
rect 452394 490054 453014 500068
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 452394 418054 453014 453498
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 452394 382054 453014 417498
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 456114 493774 456734 500068
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 456114 421774 456734 457218
rect 456114 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 456734 421774
rect 456114 421454 456734 421538
rect 456114 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 456734 421454
rect 456114 385774 456734 421218
rect 459142 391237 459202 635699
rect 479568 619174 479888 619206
rect 479568 618938 479610 619174
rect 479846 618938 479888 619174
rect 479568 618854 479888 618938
rect 479568 618618 479610 618854
rect 479846 618618 479888 618854
rect 479568 618586 479888 618618
rect 510288 619174 510608 619206
rect 510288 618938 510330 619174
rect 510566 618938 510608 619174
rect 510288 618854 510608 618938
rect 510288 618618 510330 618854
rect 510566 618618 510608 618854
rect 510288 618586 510608 618618
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 525648 615454 525968 615486
rect 525648 615218 525690 615454
rect 525926 615218 525968 615454
rect 525648 615134 525968 615218
rect 525648 614898 525690 615134
rect 525926 614898 525968 615134
rect 525648 614866 525968 614898
rect 459834 605494 460454 608991
rect 459834 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 460454 605494
rect 459834 605174 460454 605258
rect 459834 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 460454 605174
rect 459834 569494 460454 604938
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 459834 517884 460454 532938
rect 469794 579454 470414 608991
rect 472019 599588 472085 599589
rect 472019 599524 472020 599588
rect 472084 599524 472085 599588
rect 472019 599523 472085 599524
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 460696 511174 461016 511206
rect 460696 510938 460738 511174
rect 460974 510938 461016 511174
rect 460696 510854 461016 510938
rect 460696 510618 460738 510854
rect 460974 510618 461016 510854
rect 460696 510586 461016 510618
rect 459477 507454 459797 507486
rect 459477 507218 459519 507454
rect 459755 507218 459797 507454
rect 459477 507134 459797 507218
rect 459477 506898 459519 507134
rect 459755 506898 459797 507134
rect 459477 506866 459797 506898
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 459834 497494 460454 500068
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 459834 461494 460454 496938
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 459834 425494 460454 460938
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 459139 391236 459205 391237
rect 459139 391172 459140 391236
rect 459204 391172 459205 391236
rect 459139 391171 459205 391172
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 454208 363454 454528 363486
rect 454208 363218 454250 363454
rect 454486 363218 454528 363454
rect 454208 363134 454528 363218
rect 454208 362898 454250 363134
rect 454486 362898 454528 363134
rect 454208 362866 454528 362898
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 450678 328470 450738 335310
rect 450632 328410 450738 328470
rect 450632 328269 450692 328410
rect 450629 328268 450695 328269
rect 450629 328204 450630 328268
rect 450694 328204 450695 328268
rect 450629 328203 450695 328204
rect 450491 327724 450557 327725
rect 450491 327660 450492 327724
rect 450556 327660 450557 327724
rect 450491 327659 450557 327660
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448283 164116 448349 164117
rect 448283 164052 448284 164116
rect 448348 164052 448349 164116
rect 448283 164051 448349 164052
rect 448674 163505 449294 197778
rect 452394 310054 453014 345498
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 454208 327454 454528 327486
rect 454208 327218 454250 327454
rect 454486 327218 454528 327454
rect 454208 327134 454528 327218
rect 454208 326898 454250 327134
rect 454486 326898 454528 327134
rect 454208 326866 454528 326898
rect 454539 320244 454605 320245
rect 454539 320180 454540 320244
rect 454604 320180 454605 320244
rect 454539 320179 454605 320180
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 166054 453014 201498
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 423259 163436 423325 163437
rect 423259 163372 423260 163436
rect 423324 163372 423325 163436
rect 423259 163371 423325 163372
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 429568 151174 429888 151206
rect 429568 150938 429610 151174
rect 429846 150938 429888 151174
rect 429568 150854 429888 150938
rect 429568 150618 429610 150854
rect 429846 150618 429888 150854
rect 429568 150586 429888 150618
rect 414208 147454 414528 147486
rect 414208 147218 414250 147454
rect 414486 147218 414528 147454
rect 414208 147134 414528 147218
rect 414208 146898 414250 147134
rect 414486 146898 414528 147134
rect 414208 146866 414528 146898
rect 444928 147454 445248 147486
rect 444928 147218 444970 147454
rect 445206 147218 445248 147454
rect 444928 147134 445248 147218
rect 444928 146898 444970 147134
rect 445206 146898 445248 147134
rect 444928 146866 445248 146898
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 90334 413294 125778
rect 412674 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 413294 90334
rect 412674 90014 413294 90098
rect 412674 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 413294 90014
rect 412674 54334 413294 89778
rect 412674 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 413294 54334
rect 412674 54014 413294 54098
rect 412674 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 413294 54014
rect 412674 18334 413294 53778
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 130054 417014 135791
rect 416394 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 417014 130054
rect 416394 129734 417014 129818
rect 416394 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 417014 129734
rect 416394 94054 417014 129498
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 58054 417014 93498
rect 416394 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 417014 58054
rect 416394 57734 417014 57818
rect 416394 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 417014 57734
rect 416394 22054 417014 57498
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 133774 420734 135791
rect 420114 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 420734 133774
rect 420114 133454 420734 133538
rect 420114 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 420734 133454
rect 420114 97774 420734 133218
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 61774 420734 97218
rect 420114 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 420734 61774
rect 420114 61454 420734 61538
rect 420114 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 420734 61454
rect 420114 25774 420734 61218
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 101494 424454 135791
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 65494 424454 100938
rect 423834 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 424454 65494
rect 423834 65174 424454 65258
rect 423834 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 424454 65174
rect 423834 29494 424454 64938
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 111454 434414 135791
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 115174 438134 135791
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 118894 441854 135791
rect 448674 126334 449294 135791
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 86614 445574 120068
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 90334 449294 125778
rect 448674 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 449294 90334
rect 448674 90014 449294 90098
rect 448674 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 449294 90014
rect 448674 54334 449294 89778
rect 448674 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 449294 54334
rect 448674 54014 449294 54098
rect 448674 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 449294 54014
rect 448674 18334 449294 53778
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 58054 453014 93498
rect 452394 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 453014 58054
rect 452394 57734 453014 57818
rect 452394 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 453014 57734
rect 452394 22054 453014 57498
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 454542 3365 454602 320179
rect 456114 313774 456734 349218
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 459834 389494 460454 424938
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 459834 353494 460454 388938
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 379772 470414 398898
rect 472022 382397 472082 599523
rect 473514 583174 474134 608991
rect 474779 594012 474845 594013
rect 474779 593948 474780 594012
rect 474844 593948 474845 594012
rect 474779 593947 474845 593948
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 455868 474134 474618
rect 473658 435454 473978 435486
rect 473658 435218 473700 435454
rect 473936 435218 473978 435454
rect 473658 435134 473978 435218
rect 473658 434898 473700 435134
rect 473936 434898 473978 435134
rect 473658 434866 473978 434898
rect 473514 403174 474134 432068
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 472019 382396 472085 382397
rect 472019 382332 472020 382396
rect 472084 382332 472085 382396
rect 472019 382331 472085 382332
rect 469568 367174 469888 367206
rect 469568 366938 469610 367174
rect 469846 366938 469888 367174
rect 469568 366854 469888 366938
rect 469568 366618 469610 366854
rect 469846 366618 469888 366854
rect 469568 366586 469888 366618
rect 473514 367174 474134 402618
rect 474782 382397 474842 593947
rect 477234 586894 477854 608991
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 476372 439174 476692 439206
rect 476372 438938 476414 439174
rect 476650 438938 476692 439174
rect 476372 438854 476692 438938
rect 476372 438618 476414 438854
rect 476650 438618 476692 438854
rect 476372 438586 476692 438618
rect 477234 406894 477854 442338
rect 480954 590614 481574 608991
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 484674 594334 485294 608991
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 484674 522334 485294 557778
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 484674 517884 485294 521778
rect 488394 598054 489014 608991
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 492114 601774 492734 608991
rect 492114 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 492734 601774
rect 492114 601454 492734 601538
rect 492114 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 492734 601454
rect 491339 596868 491405 596869
rect 491339 596804 491340 596868
rect 491404 596804 491405 596868
rect 491339 596803 491405 596804
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 488394 517884 489014 525498
rect 490419 518124 490485 518125
rect 490419 518060 490420 518124
rect 490484 518060 490485 518124
rect 490419 518059 490485 518060
rect 482691 517580 482757 517581
rect 482691 517516 482692 517580
rect 482756 517516 482757 517580
rect 482691 517515 482757 517516
rect 482163 507454 482483 507486
rect 482163 507218 482205 507454
rect 482441 507218 482483 507454
rect 482163 507134 482483 507218
rect 482163 506898 482205 507134
rect 482441 506898 482483 507134
rect 482163 506866 482483 506898
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 482694 467125 482754 517515
rect 483382 511174 483702 511206
rect 483382 510938 483424 511174
rect 483660 510938 483702 511174
rect 483382 510854 483702 510938
rect 483382 510618 483424 510854
rect 483660 510618 483702 510854
rect 483382 510586 483702 510618
rect 485820 511174 486140 511206
rect 485820 510938 485862 511174
rect 486098 510938 486140 511174
rect 485820 510854 486140 510938
rect 485820 510618 485862 510854
rect 486098 510618 486140 510854
rect 485820 510586 486140 510618
rect 488258 511174 488578 511206
rect 488258 510938 488300 511174
rect 488536 510938 488578 511174
rect 488258 510854 488578 510938
rect 488258 510618 488300 510854
rect 488536 510618 488578 510854
rect 488258 510586 488578 510618
rect 484601 507454 484921 507486
rect 484601 507218 484643 507454
rect 484879 507218 484921 507454
rect 484601 507134 484921 507218
rect 484601 506898 484643 507134
rect 484879 506898 484921 507134
rect 484601 506866 484921 506898
rect 487039 507454 487359 507486
rect 487039 507218 487081 507454
rect 487317 507218 487359 507454
rect 487039 507134 487359 507218
rect 487039 506898 487081 507134
rect 487317 506898 487359 507134
rect 487039 506866 487359 506898
rect 489477 507454 489797 507486
rect 489477 507218 489519 507454
rect 489755 507218 489797 507454
rect 489477 507134 489797 507218
rect 489477 506898 489519 507134
rect 489755 506898 489797 507134
rect 489477 506866 489797 506898
rect 488394 490054 489014 500068
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 482691 467124 482757 467125
rect 482691 467060 482692 467124
rect 482756 467060 482757 467124
rect 482691 467059 482757 467060
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 479086 435454 479406 435486
rect 479086 435218 479128 435454
rect 479364 435218 479406 435454
rect 479086 435134 479406 435218
rect 479086 434898 479128 435134
rect 479364 434898 479406 435134
rect 479086 434866 479406 434898
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 474779 382396 474845 382397
rect 474779 382332 474780 382396
rect 474844 382332 474845 382396
rect 474779 382331 474845 382332
rect 477234 378737 477854 406338
rect 480954 410614 481574 446058
rect 488394 454054 489014 489498
rect 488394 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 489014 454054
rect 488394 453734 489014 453818
rect 488394 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 489014 453734
rect 481800 439174 482120 439206
rect 481800 438938 481842 439174
rect 482078 438938 482120 439174
rect 481800 438854 482120 438938
rect 481800 438618 481842 438854
rect 482078 438618 482120 438854
rect 481800 438586 482120 438618
rect 487228 439174 487548 439206
rect 487228 438938 487270 439174
rect 487506 438938 487548 439174
rect 487228 438854 487548 438938
rect 487228 438618 487270 438854
rect 487506 438618 487548 438854
rect 487228 438586 487548 438618
rect 484514 435454 484834 435486
rect 484514 435218 484556 435454
rect 484792 435218 484834 435454
rect 484514 435134 484834 435218
rect 484514 434898 484556 435134
rect 484792 434898 484834 435134
rect 484514 434866 484834 434898
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 378737 481574 410058
rect 488394 418054 489014 453498
rect 489942 435454 490262 435486
rect 489942 435218 489984 435454
rect 490220 435218 490262 435454
rect 489942 435134 490262 435218
rect 489942 434898 489984 435134
rect 490220 434898 490262 435134
rect 489942 434866 490262 434898
rect 488394 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 489014 418054
rect 488394 417734 489014 417818
rect 488394 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 489014 417734
rect 488394 382054 489014 417498
rect 490422 382397 490482 518059
rect 490696 511174 491016 511206
rect 490696 510938 490738 511174
rect 490974 510938 491016 511174
rect 490696 510854 491016 510938
rect 490696 510618 490738 510854
rect 490974 510618 491016 510854
rect 490696 510586 491016 510618
rect 491342 382397 491402 596803
rect 492114 565774 492734 601218
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 492114 493774 492734 529218
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 492114 455868 492734 457218
rect 495834 605494 496454 608991
rect 495834 605258 495866 605494
rect 496102 605258 496186 605494
rect 496422 605258 496454 605494
rect 495834 605174 496454 605258
rect 495834 604938 495866 605174
rect 496102 604938 496186 605174
rect 496422 604938 496454 605174
rect 495834 569494 496454 604938
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 495834 533494 496454 568938
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495834 497494 496454 532938
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 492656 439174 492976 439206
rect 492656 438938 492698 439174
rect 492934 438938 492976 439174
rect 492656 438854 492976 438938
rect 492656 438618 492698 438854
rect 492934 438618 492976 438854
rect 492656 438586 492976 438618
rect 492114 421774 492734 432068
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 492114 385774 492734 421218
rect 492114 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 492734 385774
rect 492114 385454 492734 385538
rect 492114 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 492734 385454
rect 490419 382396 490485 382397
rect 490419 382332 490420 382396
rect 490484 382332 490485 382396
rect 490419 382331 490485 382332
rect 491339 382396 491405 382397
rect 491339 382332 491340 382396
rect 491404 382332 491405 382396
rect 491339 382331 491405 382332
rect 488394 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 489014 382054
rect 488394 381734 489014 381818
rect 488394 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 489014 381734
rect 488394 378737 489014 381498
rect 492114 378737 492734 385218
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 495834 378737 496454 388938
rect 505794 579454 506414 608991
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 469568 331174 469888 331206
rect 469568 330938 469610 331174
rect 469846 330938 469888 331174
rect 469568 330854 469888 330938
rect 469568 330618 469610 330854
rect 469846 330618 469888 330854
rect 469568 330586 469888 330618
rect 473514 331174 474134 366618
rect 500288 367174 500608 367206
rect 500288 366938 500330 367174
rect 500566 366938 500608 367174
rect 500288 366854 500608 366938
rect 500288 366618 500330 366854
rect 500566 366618 500608 366854
rect 500288 366586 500608 366618
rect 484928 363454 485248 363486
rect 484928 363218 484970 363454
rect 485206 363218 485248 363454
rect 484928 363134 485248 363218
rect 484928 362898 484970 363134
rect 485206 362898 485248 363134
rect 484928 362866 485248 362898
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 463739 320380 463805 320381
rect 463739 320316 463740 320380
rect 463804 320316 463805 320380
rect 463739 320315 463805 320316
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 458771 307052 458837 307053
rect 458771 306988 458772 307052
rect 458836 306988 458837 307052
rect 458771 306987 458837 306988
rect 457299 301476 457365 301477
rect 457299 301412 457300 301476
rect 457364 301412 457365 301476
rect 457299 301411 457365 301412
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 205774 456734 241218
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 169774 456734 205218
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 457302 123725 457362 301411
rect 457483 278084 457549 278085
rect 457483 278020 457484 278084
rect 457548 278020 457549 278084
rect 457483 278019 457549 278020
rect 457486 126717 457546 278019
rect 457667 272508 457733 272509
rect 457667 272444 457668 272508
rect 457732 272444 457733 272508
rect 457667 272443 457733 272444
rect 457670 131205 457730 272443
rect 457667 131204 457733 131205
rect 457667 131140 457668 131204
rect 457732 131140 457733 131204
rect 457667 131139 457733 131140
rect 458774 129709 458834 306987
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 458955 268428 459021 268429
rect 458955 268364 458956 268428
rect 459020 268364 459021 268428
rect 458955 268363 459021 268364
rect 458958 135693 459018 268363
rect 459834 245494 460454 280938
rect 463742 276725 463802 320315
rect 473514 295174 474134 330618
rect 500288 331174 500608 331206
rect 500288 330938 500330 331174
rect 500566 330938 500608 331174
rect 500288 330854 500608 330938
rect 500288 330618 500330 330854
rect 500566 330618 500608 330854
rect 500288 330586 500608 330618
rect 484928 327454 485248 327486
rect 484928 327218 484970 327454
rect 485206 327218 485248 327454
rect 484928 327134 485248 327218
rect 484928 326898 484970 327134
rect 485206 326898 485248 327134
rect 484928 326866 485248 326898
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 463739 276724 463805 276725
rect 463739 276660 463740 276724
rect 463804 276660 463805 276724
rect 463739 276659 463805 276660
rect 473514 259417 474134 294618
rect 477234 298894 477854 320287
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 259417 477854 262338
rect 480954 302614 481574 320287
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 259417 481574 266058
rect 484674 306334 485294 320068
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 259417 485294 269778
rect 488394 310054 489014 320287
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 259417 489014 273498
rect 492114 313774 492734 320287
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 259417 492734 277218
rect 495834 317494 496454 320287
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 259417 496454 280938
rect 505794 291454 506414 326898
rect 509514 583174 510134 608991
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 513234 586894 513854 608991
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 509514 330854 510134 330938
rect 510659 330988 510725 330989
rect 510659 330924 510660 330988
rect 510724 330924 510725 330988
rect 510659 330923 510725 330924
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 507163 320652 507229 320653
rect 507163 320588 507164 320652
rect 507228 320588 507229 320652
rect 507163 320587 507229 320588
rect 506979 320380 507045 320381
rect 506979 320316 506980 320380
rect 507044 320316 507045 320380
rect 506979 320315 507045 320316
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 259417 506414 290898
rect 506982 289237 507042 320315
rect 506979 289236 507045 289237
rect 506979 289172 506980 289236
rect 507044 289172 507045 289236
rect 506979 289171 507045 289172
rect 507166 289101 507226 320587
rect 507347 320516 507413 320517
rect 507347 320452 507348 320516
rect 507412 320452 507413 320516
rect 507347 320451 507413 320452
rect 507350 294677 507410 320451
rect 509187 316708 509253 316709
rect 509187 316644 509188 316708
rect 509252 316644 509253 316708
rect 509187 316643 509253 316644
rect 509190 311910 509250 316643
rect 509006 311850 509250 311910
rect 507347 294676 507413 294677
rect 507347 294612 507348 294676
rect 507412 294612 507413 294676
rect 507347 294611 507413 294612
rect 509006 294541 509066 311850
rect 509514 295174 510134 330618
rect 510291 325276 510357 325277
rect 510291 325212 510292 325276
rect 510356 325212 510357 325276
rect 510291 325211 510357 325212
rect 510294 316709 510354 325211
rect 510475 320244 510541 320245
rect 510475 320180 510476 320244
rect 510540 320180 510541 320244
rect 510475 320179 510541 320180
rect 510291 316708 510357 316709
rect 510291 316644 510292 316708
rect 510356 316644 510357 316708
rect 510291 316643 510357 316644
rect 510478 302837 510538 320179
rect 510475 302836 510541 302837
rect 510475 302772 510476 302836
rect 510540 302772 510541 302836
rect 510475 302771 510541 302772
rect 510662 300253 510722 330923
rect 510843 323644 510909 323645
rect 510843 323580 510844 323644
rect 510908 323580 510909 323644
rect 510843 323579 510909 323580
rect 510846 305965 510906 323579
rect 511027 322012 511093 322013
rect 511027 321948 511028 322012
rect 511092 321948 511093 322012
rect 511027 321947 511093 321948
rect 510843 305964 510909 305965
rect 510843 305900 510844 305964
rect 510908 305900 510909 305964
rect 510843 305899 510909 305900
rect 511030 305693 511090 321947
rect 511211 321604 511277 321605
rect 511211 321540 511212 321604
rect 511276 321540 511277 321604
rect 511211 321539 511277 321540
rect 511214 305829 511274 321539
rect 511211 305828 511277 305829
rect 511211 305764 511212 305828
rect 511276 305764 511277 305828
rect 511211 305763 511277 305764
rect 511027 305692 511093 305693
rect 511027 305628 511028 305692
rect 511092 305628 511093 305692
rect 511027 305627 511093 305628
rect 510659 300252 510725 300253
rect 510659 300188 510660 300252
rect 510724 300188 510725 300252
rect 510659 300187 510725 300188
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509003 294540 509069 294541
rect 509003 294476 509004 294540
rect 509068 294476 509069 294540
rect 509003 294475 509069 294476
rect 507163 289100 507229 289101
rect 507163 289036 507164 289100
rect 507228 289036 507229 289100
rect 507163 289035 507229 289036
rect 509514 259417 510134 294618
rect 513234 298894 513854 334338
rect 516954 590614 517574 608991
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 514891 328540 514957 328541
rect 514891 328476 514892 328540
rect 514956 328476 514957 328540
rect 514891 328475 514957 328476
rect 514155 324052 514221 324053
rect 514155 323988 514156 324052
rect 514220 323988 514221 324052
rect 514155 323987 514221 323988
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 514158 297533 514218 323987
rect 514707 322420 514773 322421
rect 514707 322356 514708 322420
rect 514772 322356 514773 322420
rect 514707 322355 514773 322356
rect 514710 321570 514770 322355
rect 514526 321510 514770 321570
rect 514526 315349 514586 321510
rect 514523 315348 514589 315349
rect 514523 315284 514524 315348
rect 514588 315284 514589 315348
rect 514523 315283 514589 315284
rect 514894 300117 514954 328475
rect 515075 324460 515141 324461
rect 515075 324396 515076 324460
rect 515140 324396 515141 324460
rect 515075 324395 515141 324396
rect 514891 300116 514957 300117
rect 514891 300052 514892 300116
rect 514956 300052 514957 300116
rect 514891 300051 514957 300052
rect 514155 297532 514221 297533
rect 514155 297468 514156 297532
rect 514220 297468 514221 297532
rect 514155 297467 514221 297468
rect 515078 291957 515138 324395
rect 516954 302614 517574 338058
rect 520674 594334 521294 608991
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 524394 598054 525014 608991
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 464644 525014 489498
rect 528114 601774 528734 637218
rect 528114 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 528734 601774
rect 528114 601454 528734 601538
rect 528114 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 528734 601454
rect 528114 565774 528734 601218
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 524208 435454 524528 435486
rect 524208 435218 524250 435454
rect 524486 435218 524528 435454
rect 524208 435134 524528 435218
rect 524208 434898 524250 435134
rect 524486 434898 524528 435134
rect 524208 434866 524528 434898
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 518203 333436 518269 333437
rect 518203 333372 518204 333436
rect 518268 333372 518269 333436
rect 518203 333371 518269 333372
rect 517835 330172 517901 330173
rect 517835 330108 517836 330172
rect 517900 330108 517901 330172
rect 517835 330107 517901 330108
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 515075 291956 515141 291957
rect 515075 291892 515076 291956
rect 515140 291892 515141 291956
rect 515075 291891 515141 291892
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 259417 513854 262338
rect 516954 266614 517574 302058
rect 517838 291821 517898 330107
rect 518019 323236 518085 323237
rect 518019 323172 518020 323236
rect 518084 323172 518085 323236
rect 518019 323171 518085 323172
rect 517835 291820 517901 291821
rect 517835 291756 517836 291820
rect 517900 291756 517901 291820
rect 517835 291755 517901 291756
rect 518022 286381 518082 323171
rect 518206 297397 518266 333371
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 518203 297396 518269 297397
rect 518203 297332 518204 297396
rect 518268 297332 518269 297396
rect 518203 297331 518269 297332
rect 518019 286380 518085 286381
rect 518019 286316 518020 286380
rect 518084 286316 518085 286380
rect 518019 286315 518085 286316
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 259417 517574 266058
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 259417 521294 269778
rect 524394 418054 525014 425068
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 259417 525014 273498
rect 528114 421774 528734 457218
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 259417 528734 277218
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 641494 532454 676938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 542675 699820 542741 699821
rect 542675 699756 542676 699820
rect 542740 699756 542741 699820
rect 542675 699755 542741 699756
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541008 655174 541328 655206
rect 541008 654938 541050 655174
rect 541286 654938 541328 655174
rect 541008 654854 541328 654938
rect 541008 654618 541050 654854
rect 541286 654618 541328 654854
rect 541008 654586 541328 654618
rect 531834 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 532454 641494
rect 531834 641174 532454 641258
rect 531834 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 532454 641174
rect 531834 605494 532454 640938
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541008 619174 541328 619206
rect 541008 618938 541050 619174
rect 541286 618938 541328 619174
rect 541008 618854 541328 618938
rect 541008 618618 541050 618854
rect 541286 618618 541328 618854
rect 541008 618586 541328 618618
rect 531834 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 532454 605494
rect 531834 605174 532454 605258
rect 531834 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 532454 605174
rect 531834 569494 532454 604938
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 539568 439174 539888 439206
rect 539568 438938 539610 439174
rect 539846 438938 539888 439174
rect 539568 438854 539888 438938
rect 539568 438618 539610 438854
rect 539846 438618 539888 438854
rect 539568 438586 539888 438618
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 531834 317494 532454 352938
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 479568 259174 479888 259206
rect 479568 258938 479610 259174
rect 479846 258938 479888 259174
rect 479568 258854 479888 258938
rect 479568 258618 479610 258854
rect 479846 258618 479888 258854
rect 479568 258586 479888 258618
rect 510288 259174 510608 259206
rect 510288 258938 510330 259174
rect 510566 258938 510608 259174
rect 510288 258854 510608 258938
rect 510288 258618 510330 258854
rect 510566 258618 510608 258854
rect 510288 258586 510608 258618
rect 464208 255454 464528 255486
rect 464208 255218 464250 255454
rect 464486 255218 464528 255454
rect 464208 255134 464528 255218
rect 464208 254898 464250 255134
rect 464486 254898 464528 255134
rect 464208 254866 464528 254898
rect 494928 255454 495248 255486
rect 494928 255218 494970 255454
rect 495206 255218 495248 255454
rect 494928 255134 495248 255218
rect 494928 254898 494970 255134
rect 495206 254898 495248 255134
rect 494928 254866 495248 254898
rect 525648 255454 525968 255486
rect 525648 255218 525690 255454
rect 525926 255218 525968 255454
rect 525648 255134 525968 255218
rect 525648 254898 525690 255134
rect 525926 254898 525968 255134
rect 525648 254866 525968 254898
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 209494 460454 244938
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 479568 223174 479888 223206
rect 479568 222938 479610 223174
rect 479846 222938 479888 223174
rect 479568 222854 479888 222938
rect 479568 222618 479610 222854
rect 479846 222618 479888 222854
rect 479568 222586 479888 222618
rect 510288 223174 510608 223206
rect 510288 222938 510330 223174
rect 510566 222938 510608 223174
rect 510288 222854 510608 222938
rect 510288 222618 510330 222854
rect 510566 222618 510608 222854
rect 510288 222586 510608 222618
rect 464208 219454 464528 219486
rect 464208 219218 464250 219454
rect 464486 219218 464528 219454
rect 464208 219134 464528 219218
rect 464208 218898 464250 219134
rect 464486 218898 464528 219134
rect 464208 218866 464528 218898
rect 494928 219454 495248 219486
rect 494928 219218 494970 219454
rect 495206 219218 495248 219454
rect 494928 219134 495248 219218
rect 494928 218898 494970 219134
rect 495206 218898 495248 219134
rect 494928 218866 495248 218898
rect 525648 219454 525968 219486
rect 525648 219218 525690 219454
rect 525926 219218 525968 219454
rect 525648 219134 525968 219218
rect 525648 218898 525690 219134
rect 525926 218898 525968 219134
rect 525648 218866 525968 218898
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 458955 135692 459021 135693
rect 458955 135628 458956 135692
rect 459020 135628 459021 135692
rect 458955 135627 459021 135628
rect 458771 129708 458837 129709
rect 458771 129644 458772 129708
rect 458836 129644 458837 129708
rect 458771 129643 458837 129644
rect 457483 126716 457549 126717
rect 457483 126652 457484 126716
rect 457548 126652 457549 126716
rect 457483 126651 457549 126652
rect 457299 123724 457365 123725
rect 457299 123660 457300 123724
rect 457364 123660 457365 123724
rect 457299 123659 457365 123660
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 61774 456734 97218
rect 456114 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 456734 61774
rect 456114 61454 456734 61538
rect 456114 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 456734 61454
rect 456114 25774 456734 61218
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 454539 3364 454605 3365
rect 454539 3300 454540 3364
rect 454604 3300 454605 3364
rect 454539 3299 454605 3300
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 183454 470414 201919
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 187174 474134 201919
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 190894 477854 201919
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 194614 481574 201919
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 484674 198334 485294 201919
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 162334 485294 197778
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484208 147454 484528 147486
rect 484208 147218 484250 147454
rect 484486 147218 484528 147454
rect 484208 147134 484528 147218
rect 484208 146898 484250 147134
rect 484486 146898 484528 147134
rect 484208 146866 484528 146898
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 484674 126334 485294 161778
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484208 111454 484528 111486
rect 484208 111218 484250 111454
rect 484486 111218 484528 111454
rect 484208 111134 484528 111218
rect 484208 110898 484250 111134
rect 484486 110898 484528 111134
rect 484208 110866 484528 110898
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 90334 485294 125778
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 166054 489014 201919
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 130054 489014 165498
rect 488394 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 489014 130054
rect 488394 129734 489014 129818
rect 488394 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 489014 129734
rect 488394 94054 489014 129498
rect 488394 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 489014 94054
rect 488394 93734 489014 93818
rect 488394 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 489014 93734
rect 488394 58054 489014 93498
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 169774 492734 201919
rect 492114 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 492734 169774
rect 492114 169454 492734 169538
rect 492114 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 492734 169454
rect 492114 133774 492734 169218
rect 505794 183454 506414 201919
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147033 506414 182898
rect 509514 187174 510134 201919
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 147033 510134 150618
rect 513234 190894 513854 201919
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 147033 513854 154338
rect 516954 194614 517574 201919
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 514928 147454 515248 147486
rect 514928 147218 514970 147454
rect 515206 147218 515248 147454
rect 514928 147134 515248 147218
rect 514928 146898 514970 147134
rect 515206 146898 515248 147134
rect 516954 147033 517574 158058
rect 520674 198334 521294 201919
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 147033 521294 161778
rect 524394 166054 525014 201919
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 147033 525014 165498
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 147033 532454 172938
rect 541794 435454 542414 470898
rect 542678 467261 542738 699755
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 542675 467260 542741 467261
rect 542675 467196 542676 467260
rect 542740 467196 542741 467260
rect 542675 467195 542741 467196
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 545514 439174 546134 474618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 458849 549854 478338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 549234 442894 549854 445551
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 552954 410614 553574 446058
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 558867 699820 558933 699821
rect 558867 699756 558868 699820
rect 558932 699756 558933 699820
rect 558867 699755 558933 699756
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 554928 435454 555248 435486
rect 554928 435218 554970 435454
rect 555206 435218 555248 435454
rect 554928 435134 555248 435218
rect 554928 434898 554970 435134
rect 555206 434898 555248 435134
rect 554928 434866 555248 434898
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 379516 553574 410058
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 555382 367174 555702 367206
rect 555382 366938 555424 367174
rect 555660 366938 555702 367174
rect 555382 366854 555702 366938
rect 555382 366618 555424 366854
rect 555660 366618 555702 366854
rect 555382 366586 555702 366618
rect 553163 363454 553483 363486
rect 553163 363218 553205 363454
rect 553441 363218 553483 363454
rect 553163 363134 553483 363218
rect 553163 362898 553205 363134
rect 553441 362898 553483 363134
rect 553163 362866 553483 362898
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 547643 309772 547709 309773
rect 547643 309708 547644 309772
rect 547708 309708 547709 309772
rect 547643 309707 547709 309708
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 149564 546134 150618
rect 547646 148474 547706 309707
rect 548011 300388 548077 300389
rect 548011 300324 548012 300388
rect 548076 300324 548077 300388
rect 548011 300323 548077 300324
rect 548014 148613 548074 300323
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 548011 148612 548077 148613
rect 548011 148548 548012 148612
rect 548076 148548 548077 148612
rect 548011 148547 548077 148548
rect 547646 148414 548074 148474
rect 548014 148205 548074 148414
rect 548011 148204 548077 148205
rect 548011 148140 548012 148204
rect 548076 148140 548077 148204
rect 548011 148139 548077 148140
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 514928 146866 515248 146898
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 492114 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 492734 133774
rect 492114 133454 492734 133538
rect 492114 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 492734 133454
rect 492114 97774 492734 133218
rect 499568 115174 499888 115206
rect 499568 114938 499610 115174
rect 499846 114938 499888 115174
rect 499568 114854 499888 114938
rect 499568 114618 499610 114854
rect 499846 114618 499888 114854
rect 499568 114586 499888 114618
rect 530288 115174 530608 115206
rect 530288 114938 530330 115174
rect 530566 114938 530608 115174
rect 530288 114854 530608 114938
rect 530288 114618 530330 114854
rect 530566 114618 530608 114854
rect 530288 114586 530608 114618
rect 514928 111454 515248 111486
rect 514928 111218 514970 111454
rect 515206 111218 515248 111454
rect 514928 111134 515248 111218
rect 514928 110898 514970 111134
rect 515206 110898 515248 111134
rect 514928 110866 515248 110898
rect 541794 111454 542414 146898
rect 545648 147454 545968 147486
rect 545648 147218 545690 147454
rect 545926 147218 545968 147454
rect 545648 147134 545968 147218
rect 545648 146898 545690 147134
rect 545926 146898 545968 147134
rect 545648 146866 545968 146898
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 492114 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 492734 97774
rect 492114 97454 492734 97538
rect 492114 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 492734 97454
rect 492114 61774 492734 97218
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 65494 496454 87495
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 75454 506414 87495
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 79174 510134 87495
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 82894 513854 87495
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 86614 517574 87495
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 54334 521294 87495
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 58054 525014 87495
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 61774 528734 87495
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 65494 532454 87495
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 75454 542414 110898
rect 545648 111454 545968 111486
rect 545648 111218 545690 111454
rect 545926 111218 545968 111454
rect 545648 111134 545968 111218
rect 545648 110898 545690 111134
rect 545926 110898 545968 111134
rect 545648 110866 545968 110898
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 545514 79174 546134 80068
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 549234 53868 549854 82338
rect 552954 338614 553574 360068
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 556674 342334 557294 377778
rect 557602 363454 557922 363486
rect 557602 363218 557644 363454
rect 557880 363218 557922 363454
rect 557602 363134 557922 363218
rect 557602 362898 557644 363134
rect 557880 362898 557922 363134
rect 557602 362866 557922 362898
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 558870 320109 558930 699755
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 559821 367174 560141 367206
rect 559821 366938 559863 367174
rect 560099 366938 560141 367174
rect 559821 366854 560141 366938
rect 559821 366618 559863 366854
rect 560099 366618 560141 366854
rect 559821 366586 560141 366618
rect 560394 346054 561014 381498
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 379516 564734 385218
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 564260 367174 564580 367206
rect 564260 366938 564302 367174
rect 564538 366938 564580 367174
rect 564260 366854 564580 366938
rect 564260 366618 564302 366854
rect 564538 366618 564580 366854
rect 564260 366586 564580 366618
rect 562041 363454 562361 363486
rect 562041 363218 562083 363454
rect 562319 363218 562361 363454
rect 562041 363134 562361 363218
rect 562041 362898 562083 363134
rect 562319 362898 562361 363134
rect 562041 362866 562361 362898
rect 566480 363454 566800 363486
rect 566480 363218 566522 363454
rect 566758 363218 566800 363454
rect 566480 363134 566800 363218
rect 566480 362898 566522 363134
rect 566758 362898 566800 363134
rect 566480 362866 566800 362898
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 558867 320108 558933 320109
rect 558867 320044 558868 320108
rect 558932 320044 558933 320108
rect 558867 320043 558933 320044
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54235 557294 89778
rect 556674 53999 556706 54235
rect 556942 53999 557026 54235
rect 557262 53999 557294 54235
rect 556674 53868 557294 53999
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 543658 39454 543978 39486
rect 543658 39218 543700 39454
rect 543936 39218 543978 39454
rect 543658 39134 543978 39218
rect 543658 38898 543700 39134
rect 543936 38898 543978 39134
rect 543658 38866 543978 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 42618
rect 546372 43174 546692 43206
rect 546372 42938 546414 43174
rect 546650 42938 546692 43174
rect 546372 42854 546692 42938
rect 546372 42618 546414 42854
rect 546650 42618 546692 42854
rect 546372 42586 546692 42618
rect 551800 43174 552120 43206
rect 552954 43177 553574 50058
rect 551800 42938 551842 43174
rect 552078 42938 552120 43174
rect 551800 42854 552120 42938
rect 551800 42618 551842 42854
rect 552078 42618 552120 42854
rect 551800 42586 552120 42618
rect 557228 43174 557548 43206
rect 557228 42938 557270 43174
rect 557506 42938 557548 43174
rect 557228 42854 557548 42938
rect 557228 42618 557270 42854
rect 557506 42618 557548 42854
rect 557228 42586 557548 42618
rect 549086 39454 549406 39486
rect 549086 39218 549128 39454
rect 549364 39218 549406 39454
rect 549086 39134 549406 39218
rect 549086 38898 549128 39134
rect 549364 38898 549406 39134
rect 549086 38866 549406 38898
rect 554514 39454 554834 39486
rect 554514 39218 554556 39454
rect 554792 39218 554834 39454
rect 554514 39134 554834 39218
rect 554514 38898 554556 39134
rect 554792 38898 554834 39134
rect 554514 38866 554834 38898
rect 559942 39454 560262 39486
rect 559942 39218 559984 39454
rect 560220 39218 560262 39454
rect 559942 39134 560262 39218
rect 559942 38898 559984 39134
rect 560220 38898 560262 39134
rect 559942 38866 560262 38898
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 30068
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 35319
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 18334 557294 30068
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 22054 561014 57498
rect 564114 349774 564734 360068
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 562656 43174 562976 43206
rect 562656 42938 562698 43174
rect 562934 42938 562976 43174
rect 562656 42854 562976 42938
rect 562656 42618 562698 42854
rect 562934 42618 562976 42854
rect 562656 42586 562976 42618
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 353494 568454 388938
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 568699 367174 569019 367206
rect 568699 366938 568741 367174
rect 568977 366938 569019 367174
rect 568699 366854 569019 366938
rect 568699 366618 568741 366854
rect 568977 366618 569019 366854
rect 568699 366586 569019 366618
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 24146 673538 24382 673774
rect 24466 673538 24702 673774
rect 24146 673218 24382 673454
rect 24466 673218 24702 673454
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 24250 651218 24486 651454
rect 24250 650898 24486 651134
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 24250 615218 24486 615454
rect 24250 614898 24486 615134
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 24250 579218 24486 579454
rect 24250 578898 24486 579134
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 24250 543218 24486 543454
rect 24250 542898 24486 543134
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 24250 507218 24486 507454
rect 24250 506898 24486 507134
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 24250 471218 24486 471454
rect 24250 470898 24486 471134
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 24250 435218 24486 435454
rect 24250 434898 24486 435134
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 24250 399218 24486 399454
rect 24250 398898 24486 399134
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 24250 363218 24486 363454
rect 24250 362898 24486 363134
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 24250 327218 24486 327454
rect 24250 326898 24486 327134
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 24250 291218 24486 291454
rect 24250 290898 24486 291134
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 24250 255218 24486 255454
rect 24250 254898 24486 255134
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 24250 219218 24486 219454
rect 24250 218898 24486 219134
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 24250 183218 24486 183454
rect 24250 182898 24486 183134
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 24250 147218 24486 147454
rect 24250 146898 24486 147134
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 24250 111218 24486 111454
rect 24250 110898 24486 111134
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 24250 75218 24486 75454
rect 24250 74898 24486 75134
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 39610 654938 39846 655174
rect 39610 654618 39846 654854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 39610 618938 39846 619174
rect 39610 618618 39846 618854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 39610 582938 39846 583174
rect 39610 582618 39846 582854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 39610 546938 39846 547174
rect 39610 546618 39846 546854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 39610 510938 39846 511174
rect 39610 510618 39846 510854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 39610 474938 39846 475174
rect 39610 474618 39846 474854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 39610 438938 39846 439174
rect 39610 438618 39846 438854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 39610 402938 39846 403174
rect 39610 402618 39846 402854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 39610 366938 39846 367174
rect 39610 366618 39846 366854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 39610 330938 39846 331174
rect 39610 330618 39846 330854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 39610 294938 39846 295174
rect 39610 294618 39846 294854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 39610 258938 39846 259174
rect 39610 258618 39846 258854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 39610 222938 39846 223174
rect 39610 222618 39846 222854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 39610 186938 39846 187174
rect 39610 186618 39846 186854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 39610 150938 39846 151174
rect 39610 150618 39846 150854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 39610 114938 39846 115174
rect 39610 114618 39846 114854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 39610 78938 39846 79174
rect 39610 78618 39846 78854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 708442 52942 708678
rect 53026 708442 53262 708678
rect 52706 708122 52942 708358
rect 53026 708122 53262 708358
rect 52706 666098 52942 666334
rect 53026 666098 53262 666334
rect 52706 665778 52942 666014
rect 53026 665778 53262 666014
rect 56426 709402 56662 709638
rect 56746 709402 56982 709638
rect 56426 709082 56662 709318
rect 56746 709082 56982 709318
rect 56426 669818 56662 670054
rect 56746 669818 56982 670054
rect 56426 669498 56662 669734
rect 56746 669498 56982 669734
rect 54970 651218 55206 651454
rect 54970 650898 55206 651134
rect 52706 630098 52942 630334
rect 53026 630098 53262 630334
rect 52706 629778 52942 630014
rect 53026 629778 53262 630014
rect 56426 633818 56662 634054
rect 56746 633818 56982 634054
rect 56426 633498 56662 633734
rect 56746 633498 56982 633734
rect 54970 615218 55206 615454
rect 54970 614898 55206 615134
rect 52706 594098 52942 594334
rect 53026 594098 53262 594334
rect 52706 593778 52942 594014
rect 53026 593778 53262 594014
rect 56426 597818 56662 598054
rect 56746 597818 56982 598054
rect 56426 597498 56662 597734
rect 56746 597498 56982 597734
rect 54970 579218 55206 579454
rect 54970 578898 55206 579134
rect 52706 558098 52942 558334
rect 53026 558098 53262 558334
rect 52706 557778 52942 558014
rect 53026 557778 53262 558014
rect 56426 561818 56662 562054
rect 56746 561818 56982 562054
rect 56426 561498 56662 561734
rect 56746 561498 56982 561734
rect 54970 543218 55206 543454
rect 54970 542898 55206 543134
rect 52706 522098 52942 522334
rect 53026 522098 53262 522334
rect 52706 521778 52942 522014
rect 53026 521778 53262 522014
rect 56426 525818 56662 526054
rect 56746 525818 56982 526054
rect 56426 525498 56662 525734
rect 56746 525498 56982 525734
rect 54970 507218 55206 507454
rect 54970 506898 55206 507134
rect 52706 486098 52942 486334
rect 53026 486098 53262 486334
rect 52706 485778 52942 486014
rect 53026 485778 53262 486014
rect 56426 489818 56662 490054
rect 56746 489818 56982 490054
rect 56426 489498 56662 489734
rect 56746 489498 56982 489734
rect 54970 471218 55206 471454
rect 54970 470898 55206 471134
rect 52706 450098 52942 450334
rect 53026 450098 53262 450334
rect 52706 449778 52942 450014
rect 53026 449778 53262 450014
rect 56426 453818 56662 454054
rect 56746 453818 56982 454054
rect 56426 453498 56662 453734
rect 56746 453498 56982 453734
rect 54970 435218 55206 435454
rect 54970 434898 55206 435134
rect 52706 414098 52942 414334
rect 53026 414098 53262 414334
rect 52706 413778 52942 414014
rect 53026 413778 53262 414014
rect 56426 417818 56662 418054
rect 56746 417818 56982 418054
rect 56426 417498 56662 417734
rect 56746 417498 56982 417734
rect 54970 399218 55206 399454
rect 54970 398898 55206 399134
rect 52706 378098 52942 378334
rect 53026 378098 53262 378334
rect 52706 377778 52942 378014
rect 53026 377778 53262 378014
rect 56426 381818 56662 382054
rect 56746 381818 56982 382054
rect 56426 381498 56662 381734
rect 56746 381498 56982 381734
rect 54970 363218 55206 363454
rect 54970 362898 55206 363134
rect 52706 342098 52942 342334
rect 53026 342098 53262 342334
rect 52706 341778 52942 342014
rect 53026 341778 53262 342014
rect 56426 345818 56662 346054
rect 56746 345818 56982 346054
rect 56426 345498 56662 345734
rect 56746 345498 56982 345734
rect 54970 327218 55206 327454
rect 54970 326898 55206 327134
rect 52706 306098 52942 306334
rect 53026 306098 53262 306334
rect 52706 305778 52942 306014
rect 53026 305778 53262 306014
rect 56426 309818 56662 310054
rect 56746 309818 56982 310054
rect 56426 309498 56662 309734
rect 56746 309498 56982 309734
rect 54970 291218 55206 291454
rect 54970 290898 55206 291134
rect 52706 270098 52942 270334
rect 53026 270098 53262 270334
rect 52706 269778 52942 270014
rect 53026 269778 53262 270014
rect 56426 273818 56662 274054
rect 56746 273818 56982 274054
rect 56426 273498 56662 273734
rect 56746 273498 56982 273734
rect 54970 255218 55206 255454
rect 54970 254898 55206 255134
rect 52706 234098 52942 234334
rect 53026 234098 53262 234334
rect 52706 233778 52942 234014
rect 53026 233778 53262 234014
rect 56426 237818 56662 238054
rect 56746 237818 56982 238054
rect 56426 237498 56662 237734
rect 56746 237498 56982 237734
rect 54970 219218 55206 219454
rect 54970 218898 55206 219134
rect 52706 198098 52942 198334
rect 53026 198098 53262 198334
rect 52706 197778 52942 198014
rect 53026 197778 53262 198014
rect 56426 201818 56662 202054
rect 56746 201818 56982 202054
rect 56426 201498 56662 201734
rect 56746 201498 56982 201734
rect 54970 183218 55206 183454
rect 54970 182898 55206 183134
rect 52706 162098 52942 162334
rect 53026 162098 53262 162334
rect 52706 161778 52942 162014
rect 53026 161778 53262 162014
rect 56426 165818 56662 166054
rect 56746 165818 56982 166054
rect 56426 165498 56662 165734
rect 56746 165498 56982 165734
rect 54970 147218 55206 147454
rect 54970 146898 55206 147134
rect 52706 126098 52942 126334
rect 53026 126098 53262 126334
rect 52706 125778 52942 126014
rect 53026 125778 53262 126014
rect 56426 129818 56662 130054
rect 56746 129818 56982 130054
rect 56426 129498 56662 129734
rect 56746 129498 56982 129734
rect 54970 111218 55206 111454
rect 54970 110898 55206 111134
rect 52706 90098 52942 90334
rect 53026 90098 53262 90334
rect 52706 89778 52942 90014
rect 53026 89778 53262 90014
rect 56426 93818 56662 94054
rect 56746 93818 56982 94054
rect 56426 93498 56662 93734
rect 56746 93498 56982 93734
rect 54970 75218 55206 75454
rect 54970 74898 55206 75134
rect 52706 54098 52942 54334
rect 53026 54098 53262 54334
rect 52706 53778 52942 54014
rect 53026 53778 53262 54014
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 57818 56662 58054
rect 56746 57818 56982 58054
rect 56426 57498 56662 57734
rect 56746 57498 56982 57734
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 710362 60382 710598
rect 60466 710362 60702 710598
rect 60146 710042 60382 710278
rect 60466 710042 60702 710278
rect 60146 673538 60382 673774
rect 60466 673538 60702 673774
rect 60146 673218 60382 673454
rect 60466 673218 60702 673454
rect 60146 637538 60382 637774
rect 60466 637538 60702 637774
rect 60146 637218 60382 637454
rect 60466 637218 60702 637454
rect 60146 601538 60382 601774
rect 60466 601538 60702 601774
rect 60146 601218 60382 601454
rect 60466 601218 60702 601454
rect 60146 565538 60382 565774
rect 60466 565538 60702 565774
rect 60146 565218 60382 565454
rect 60466 565218 60702 565454
rect 60146 529538 60382 529774
rect 60466 529538 60702 529774
rect 60146 529218 60382 529454
rect 60466 529218 60702 529454
rect 60146 493538 60382 493774
rect 60466 493538 60702 493774
rect 60146 493218 60382 493454
rect 60466 493218 60702 493454
rect 60146 457538 60382 457774
rect 60466 457538 60702 457774
rect 60146 457218 60382 457454
rect 60466 457218 60702 457454
rect 60146 421538 60382 421774
rect 60466 421538 60702 421774
rect 60146 421218 60382 421454
rect 60466 421218 60702 421454
rect 60146 385538 60382 385774
rect 60466 385538 60702 385774
rect 60146 385218 60382 385454
rect 60466 385218 60702 385454
rect 60146 349538 60382 349774
rect 60466 349538 60702 349774
rect 60146 349218 60382 349454
rect 60466 349218 60702 349454
rect 60146 313538 60382 313774
rect 60466 313538 60702 313774
rect 60146 313218 60382 313454
rect 60466 313218 60702 313454
rect 60146 277538 60382 277774
rect 60466 277538 60702 277774
rect 60146 277218 60382 277454
rect 60466 277218 60702 277454
rect 60146 241538 60382 241774
rect 60466 241538 60702 241774
rect 60146 241218 60382 241454
rect 60466 241218 60702 241454
rect 60146 205538 60382 205774
rect 60466 205538 60702 205774
rect 60146 205218 60382 205454
rect 60466 205218 60702 205454
rect 60146 169538 60382 169774
rect 60466 169538 60702 169774
rect 60146 169218 60382 169454
rect 60466 169218 60702 169454
rect 60146 133538 60382 133774
rect 60466 133538 60702 133774
rect 60146 133218 60382 133454
rect 60466 133218 60702 133454
rect 60146 97538 60382 97774
rect 60466 97538 60702 97774
rect 60146 97218 60382 97454
rect 60466 97218 60702 97454
rect 60146 61538 60382 61774
rect 60466 61538 60702 61774
rect 60146 61218 60382 61454
rect 60466 61218 60702 61454
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 92426 709402 92662 709638
rect 92746 709402 92982 709638
rect 92426 709082 92662 709318
rect 92746 709082 92982 709318
rect 92426 669818 92662 670054
rect 92746 669818 92982 670054
rect 92426 669498 92662 669734
rect 92746 669498 92982 669734
rect 96146 710362 96382 710598
rect 96466 710362 96702 710598
rect 96146 710042 96382 710278
rect 96466 710042 96702 710278
rect 96146 673538 96382 673774
rect 96466 673538 96702 673774
rect 96146 673218 96382 673454
rect 96466 673218 96702 673454
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 128426 709402 128662 709638
rect 128746 709402 128982 709638
rect 128426 709082 128662 709318
rect 128746 709082 128982 709318
rect 128426 669818 128662 670054
rect 128746 669818 128982 670054
rect 128426 669498 128662 669734
rect 128746 669498 128982 669734
rect 132146 710362 132382 710598
rect 132466 710362 132702 710598
rect 132146 710042 132382 710278
rect 132466 710042 132702 710278
rect 132146 673538 132382 673774
rect 132466 673538 132702 673774
rect 132146 673218 132382 673454
rect 132466 673218 132702 673454
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 164426 709402 164662 709638
rect 164746 709402 164982 709638
rect 164426 709082 164662 709318
rect 164746 709082 164982 709318
rect 164426 669818 164662 670054
rect 164746 669818 164982 670054
rect 164426 669498 164662 669734
rect 164746 669498 164982 669734
rect 168146 710362 168382 710598
rect 168466 710362 168702 710598
rect 168146 710042 168382 710278
rect 168466 710042 168702 710278
rect 168146 673538 168382 673774
rect 168466 673538 168702 673774
rect 168146 673218 168382 673454
rect 168466 673218 168702 673454
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 204146 710362 204382 710598
rect 204466 710362 204702 710598
rect 204146 710042 204382 710278
rect 204466 710042 204702 710278
rect 204146 673538 204382 673774
rect 204466 673538 204702 673774
rect 204146 673218 204382 673454
rect 204466 673218 204702 673454
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 236426 709402 236662 709638
rect 236746 709402 236982 709638
rect 236426 709082 236662 709318
rect 236746 709082 236982 709318
rect 236426 669818 236662 670054
rect 236746 669818 236982 670054
rect 236426 669498 236662 669734
rect 236746 669498 236982 669734
rect 240146 710362 240382 710598
rect 240466 710362 240702 710598
rect 240146 710042 240382 710278
rect 240466 710042 240702 710278
rect 240146 673538 240382 673774
rect 240466 673538 240702 673774
rect 240146 673218 240382 673454
rect 240466 673218 240702 673454
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 272426 709402 272662 709638
rect 272746 709402 272982 709638
rect 272426 709082 272662 709318
rect 272746 709082 272982 709318
rect 272426 669818 272662 670054
rect 272746 669818 272982 670054
rect 272426 669498 272662 669734
rect 272746 669498 272982 669734
rect 276146 710362 276382 710598
rect 276466 710362 276702 710598
rect 276146 710042 276382 710278
rect 276466 710042 276702 710278
rect 276146 673538 276382 673774
rect 276466 673538 276702 673774
rect 276146 673218 276382 673454
rect 276466 673218 276702 673454
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 308426 709402 308662 709638
rect 308746 709402 308982 709638
rect 308426 709082 308662 709318
rect 308746 709082 308982 709318
rect 308426 669818 308662 670054
rect 308746 669818 308982 670054
rect 308426 669498 308662 669734
rect 308746 669498 308982 669734
rect 312146 710362 312382 710598
rect 312466 710362 312702 710598
rect 312146 710042 312382 710278
rect 312466 710042 312702 710278
rect 312146 673538 312382 673774
rect 312466 673538 312702 673774
rect 312146 673218 312382 673454
rect 312466 673218 312702 673454
rect 315866 711322 316102 711558
rect 316186 711322 316422 711558
rect 315866 711002 316102 711238
rect 316186 711002 316422 711238
rect 315866 677258 316102 677494
rect 316186 677258 316422 677494
rect 315866 676938 316102 677174
rect 316186 676938 316422 677174
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 70330 654938 70566 655174
rect 70330 654618 70566 654854
rect 101050 654938 101286 655174
rect 101050 654618 101286 654854
rect 131770 654938 132006 655174
rect 131770 654618 132006 654854
rect 162490 654938 162726 655174
rect 162490 654618 162726 654854
rect 193210 654938 193446 655174
rect 193210 654618 193446 654854
rect 223930 654938 224166 655174
rect 223930 654618 224166 654854
rect 254650 654938 254886 655174
rect 254650 654618 254886 654854
rect 285370 654938 285606 655174
rect 285370 654618 285606 654854
rect 316090 654938 316326 655174
rect 316090 654618 316326 654854
rect 346810 654938 347046 655174
rect 346810 654618 347046 654854
rect 85690 651218 85926 651454
rect 85690 650898 85926 651134
rect 116410 651218 116646 651454
rect 116410 650898 116646 651134
rect 147130 651218 147366 651454
rect 147130 650898 147366 651134
rect 177850 651218 178086 651454
rect 177850 650898 178086 651134
rect 208570 651218 208806 651454
rect 208570 650898 208806 651134
rect 239290 651218 239526 651454
rect 239290 650898 239526 651134
rect 270010 651218 270246 651454
rect 270010 650898 270246 651134
rect 300730 651218 300966 651454
rect 300730 650898 300966 651134
rect 331450 651218 331686 651454
rect 331450 650898 331686 651134
rect 362170 651218 362406 651454
rect 362170 650898 362406 651134
rect 63866 641258 64102 641494
rect 64186 641258 64422 641494
rect 63866 640938 64102 641174
rect 64186 640938 64422 641174
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 377530 654938 377766 655174
rect 377530 654618 377766 654854
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 70330 618938 70566 619174
rect 70330 618618 70566 618854
rect 101050 618938 101286 619174
rect 101050 618618 101286 618854
rect 131770 618938 132006 619174
rect 131770 618618 132006 618854
rect 162490 618938 162726 619174
rect 162490 618618 162726 618854
rect 193210 618938 193446 619174
rect 193210 618618 193446 618854
rect 223930 618938 224166 619174
rect 223930 618618 224166 618854
rect 254650 618938 254886 619174
rect 254650 618618 254886 618854
rect 285370 618938 285606 619174
rect 285370 618618 285606 618854
rect 316090 618938 316326 619174
rect 316090 618618 316326 618854
rect 346810 618938 347046 619174
rect 346810 618618 347046 618854
rect 85690 615218 85926 615454
rect 85690 614898 85926 615134
rect 116410 615218 116646 615454
rect 116410 614898 116646 615134
rect 147130 615218 147366 615454
rect 147130 614898 147366 615134
rect 177850 615218 178086 615454
rect 177850 614898 178086 615134
rect 208570 615218 208806 615454
rect 208570 614898 208806 615134
rect 239290 615218 239526 615454
rect 239290 614898 239526 615134
rect 270010 615218 270246 615454
rect 270010 614898 270246 615134
rect 300730 615218 300966 615454
rect 300730 614898 300966 615134
rect 331450 615218 331686 615454
rect 331450 614898 331686 615134
rect 362170 615218 362406 615454
rect 362170 614898 362406 615134
rect 63866 605258 64102 605494
rect 64186 605258 64422 605494
rect 63866 604938 64102 605174
rect 64186 604938 64422 605174
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 377530 618938 377766 619174
rect 377530 618618 377766 618854
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 70330 582938 70566 583174
rect 70330 582618 70566 582854
rect 101050 582938 101286 583174
rect 101050 582618 101286 582854
rect 131770 582938 132006 583174
rect 131770 582618 132006 582854
rect 162490 582938 162726 583174
rect 162490 582618 162726 582854
rect 193210 582938 193446 583174
rect 193210 582618 193446 582854
rect 223930 582938 224166 583174
rect 223930 582618 224166 582854
rect 254650 582938 254886 583174
rect 254650 582618 254886 582854
rect 285370 582938 285606 583174
rect 285370 582618 285606 582854
rect 316090 582938 316326 583174
rect 316090 582618 316326 582854
rect 346810 582938 347046 583174
rect 346810 582618 347046 582854
rect 85690 579218 85926 579454
rect 85690 578898 85926 579134
rect 116410 579218 116646 579454
rect 116410 578898 116646 579134
rect 147130 579218 147366 579454
rect 147130 578898 147366 579134
rect 177850 579218 178086 579454
rect 177850 578898 178086 579134
rect 208570 579218 208806 579454
rect 208570 578898 208806 579134
rect 239290 579218 239526 579454
rect 239290 578898 239526 579134
rect 270010 579218 270246 579454
rect 270010 578898 270246 579134
rect 300730 579218 300966 579454
rect 300730 578898 300966 579134
rect 331450 579218 331686 579454
rect 331450 578898 331686 579134
rect 362170 579218 362406 579454
rect 362170 578898 362406 579134
rect 63866 569258 64102 569494
rect 64186 569258 64422 569494
rect 63866 568938 64102 569174
rect 64186 568938 64422 569174
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 377530 582938 377766 583174
rect 377530 582618 377766 582854
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 70330 546938 70566 547174
rect 70330 546618 70566 546854
rect 101050 546938 101286 547174
rect 101050 546618 101286 546854
rect 131770 546938 132006 547174
rect 131770 546618 132006 546854
rect 162490 546938 162726 547174
rect 162490 546618 162726 546854
rect 193210 546938 193446 547174
rect 193210 546618 193446 546854
rect 223930 546938 224166 547174
rect 223930 546618 224166 546854
rect 254650 546938 254886 547174
rect 254650 546618 254886 546854
rect 285370 546938 285606 547174
rect 285370 546618 285606 546854
rect 316090 546938 316326 547174
rect 316090 546618 316326 546854
rect 346810 546938 347046 547174
rect 346810 546618 347046 546854
rect 85690 543218 85926 543454
rect 85690 542898 85926 543134
rect 116410 543218 116646 543454
rect 116410 542898 116646 543134
rect 147130 543218 147366 543454
rect 147130 542898 147366 543134
rect 177850 543218 178086 543454
rect 177850 542898 178086 543134
rect 208570 543218 208806 543454
rect 208570 542898 208806 543134
rect 239290 543218 239526 543454
rect 239290 542898 239526 543134
rect 270010 543218 270246 543454
rect 270010 542898 270246 543134
rect 300730 543218 300966 543454
rect 300730 542898 300966 543134
rect 331450 543218 331686 543454
rect 331450 542898 331686 543134
rect 362170 543218 362406 543454
rect 362170 542898 362406 543134
rect 63866 533258 64102 533494
rect 64186 533258 64422 533494
rect 63866 532938 64102 533174
rect 64186 532938 64422 533174
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 377530 546938 377766 547174
rect 377530 546618 377766 546854
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 70330 510938 70566 511174
rect 70330 510618 70566 510854
rect 101050 510938 101286 511174
rect 101050 510618 101286 510854
rect 131770 510938 132006 511174
rect 131770 510618 132006 510854
rect 162490 510938 162726 511174
rect 162490 510618 162726 510854
rect 193210 510938 193446 511174
rect 193210 510618 193446 510854
rect 223930 510938 224166 511174
rect 223930 510618 224166 510854
rect 254650 510938 254886 511174
rect 254650 510618 254886 510854
rect 285370 510938 285606 511174
rect 285370 510618 285606 510854
rect 316090 510938 316326 511174
rect 316090 510618 316326 510854
rect 346810 510938 347046 511174
rect 346810 510618 347046 510854
rect 85690 507218 85926 507454
rect 85690 506898 85926 507134
rect 116410 507218 116646 507454
rect 116410 506898 116646 507134
rect 147130 507218 147366 507454
rect 147130 506898 147366 507134
rect 177850 507218 178086 507454
rect 177850 506898 178086 507134
rect 208570 507218 208806 507454
rect 208570 506898 208806 507134
rect 239290 507218 239526 507454
rect 239290 506898 239526 507134
rect 270010 507218 270246 507454
rect 270010 506898 270246 507134
rect 300730 507218 300966 507454
rect 300730 506898 300966 507134
rect 331450 507218 331686 507454
rect 331450 506898 331686 507134
rect 362170 507218 362406 507454
rect 362170 506898 362406 507134
rect 63866 497258 64102 497494
rect 64186 497258 64422 497494
rect 63866 496938 64102 497174
rect 64186 496938 64422 497174
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 377530 510938 377766 511174
rect 377530 510618 377766 510854
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 70330 474938 70566 475174
rect 70330 474618 70566 474854
rect 101050 474938 101286 475174
rect 101050 474618 101286 474854
rect 131770 474938 132006 475174
rect 131770 474618 132006 474854
rect 162490 474938 162726 475174
rect 162490 474618 162726 474854
rect 193210 474938 193446 475174
rect 193210 474618 193446 474854
rect 223930 474938 224166 475174
rect 223930 474618 224166 474854
rect 254650 474938 254886 475174
rect 254650 474618 254886 474854
rect 285370 474938 285606 475174
rect 285370 474618 285606 474854
rect 316090 474938 316326 475174
rect 316090 474618 316326 474854
rect 346810 474938 347046 475174
rect 346810 474618 347046 474854
rect 85690 471218 85926 471454
rect 85690 470898 85926 471134
rect 116410 471218 116646 471454
rect 116410 470898 116646 471134
rect 147130 471218 147366 471454
rect 147130 470898 147366 471134
rect 177850 471218 178086 471454
rect 177850 470898 178086 471134
rect 208570 471218 208806 471454
rect 208570 470898 208806 471134
rect 239290 471218 239526 471454
rect 239290 470898 239526 471134
rect 270010 471218 270246 471454
rect 270010 470898 270246 471134
rect 300730 471218 300966 471454
rect 300730 470898 300966 471134
rect 331450 471218 331686 471454
rect 331450 470898 331686 471134
rect 362170 471218 362406 471454
rect 362170 470898 362406 471134
rect 63866 461258 64102 461494
rect 64186 461258 64422 461494
rect 63866 460938 64102 461174
rect 64186 460938 64422 461174
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 377530 474938 377766 475174
rect 377530 474618 377766 474854
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 70330 438938 70566 439174
rect 70330 438618 70566 438854
rect 101050 438938 101286 439174
rect 101050 438618 101286 438854
rect 131770 438938 132006 439174
rect 131770 438618 132006 438854
rect 162490 438938 162726 439174
rect 162490 438618 162726 438854
rect 193210 438938 193446 439174
rect 193210 438618 193446 438854
rect 223930 438938 224166 439174
rect 223930 438618 224166 438854
rect 254650 438938 254886 439174
rect 254650 438618 254886 438854
rect 285370 438938 285606 439174
rect 285370 438618 285606 438854
rect 316090 438938 316326 439174
rect 316090 438618 316326 438854
rect 346810 438938 347046 439174
rect 346810 438618 347046 438854
rect 85690 435218 85926 435454
rect 85690 434898 85926 435134
rect 116410 435218 116646 435454
rect 116410 434898 116646 435134
rect 147130 435218 147366 435454
rect 147130 434898 147366 435134
rect 177850 435218 178086 435454
rect 177850 434898 178086 435134
rect 208570 435218 208806 435454
rect 208570 434898 208806 435134
rect 239290 435218 239526 435454
rect 239290 434898 239526 435134
rect 270010 435218 270246 435454
rect 270010 434898 270246 435134
rect 300730 435218 300966 435454
rect 300730 434898 300966 435134
rect 331450 435218 331686 435454
rect 331450 434898 331686 435134
rect 362170 435218 362406 435454
rect 362170 434898 362406 435134
rect 63866 425258 64102 425494
rect 64186 425258 64422 425494
rect 63866 424938 64102 425174
rect 64186 424938 64422 425174
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 377530 438938 377766 439174
rect 377530 438618 377766 438854
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 70330 402938 70566 403174
rect 70330 402618 70566 402854
rect 101050 402938 101286 403174
rect 101050 402618 101286 402854
rect 131770 402938 132006 403174
rect 131770 402618 132006 402854
rect 162490 402938 162726 403174
rect 162490 402618 162726 402854
rect 193210 402938 193446 403174
rect 193210 402618 193446 402854
rect 223930 402938 224166 403174
rect 223930 402618 224166 402854
rect 254650 402938 254886 403174
rect 254650 402618 254886 402854
rect 285370 402938 285606 403174
rect 285370 402618 285606 402854
rect 316090 402938 316326 403174
rect 316090 402618 316326 402854
rect 346810 402938 347046 403174
rect 346810 402618 347046 402854
rect 85690 399218 85926 399454
rect 85690 398898 85926 399134
rect 116410 399218 116646 399454
rect 116410 398898 116646 399134
rect 147130 399218 147366 399454
rect 147130 398898 147366 399134
rect 177850 399218 178086 399454
rect 177850 398898 178086 399134
rect 208570 399218 208806 399454
rect 208570 398898 208806 399134
rect 239290 399218 239526 399454
rect 239290 398898 239526 399134
rect 270010 399218 270246 399454
rect 270010 398898 270246 399134
rect 300730 399218 300966 399454
rect 300730 398898 300966 399134
rect 331450 399218 331686 399454
rect 331450 398898 331686 399134
rect 362170 399218 362406 399454
rect 362170 398898 362406 399134
rect 63866 389258 64102 389494
rect 64186 389258 64422 389494
rect 63866 388938 64102 389174
rect 64186 388938 64422 389174
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 377530 402938 377766 403174
rect 377530 402618 377766 402854
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 70330 366938 70566 367174
rect 70330 366618 70566 366854
rect 101050 366938 101286 367174
rect 101050 366618 101286 366854
rect 131770 366938 132006 367174
rect 131770 366618 132006 366854
rect 162490 366938 162726 367174
rect 162490 366618 162726 366854
rect 193210 366938 193446 367174
rect 193210 366618 193446 366854
rect 223930 366938 224166 367174
rect 223930 366618 224166 366854
rect 254650 366938 254886 367174
rect 254650 366618 254886 366854
rect 285370 366938 285606 367174
rect 285370 366618 285606 366854
rect 316090 366938 316326 367174
rect 316090 366618 316326 366854
rect 346810 366938 347046 367174
rect 346810 366618 347046 366854
rect 85690 363218 85926 363454
rect 85690 362898 85926 363134
rect 116410 363218 116646 363454
rect 116410 362898 116646 363134
rect 147130 363218 147366 363454
rect 147130 362898 147366 363134
rect 177850 363218 178086 363454
rect 177850 362898 178086 363134
rect 208570 363218 208806 363454
rect 208570 362898 208806 363134
rect 239290 363218 239526 363454
rect 239290 362898 239526 363134
rect 270010 363218 270246 363454
rect 270010 362898 270246 363134
rect 300730 363218 300966 363454
rect 300730 362898 300966 363134
rect 331450 363218 331686 363454
rect 331450 362898 331686 363134
rect 362170 363218 362406 363454
rect 362170 362898 362406 363134
rect 63866 353258 64102 353494
rect 64186 353258 64422 353494
rect 63866 352938 64102 353174
rect 64186 352938 64422 353174
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 377530 366938 377766 367174
rect 377530 366618 377766 366854
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 70330 330938 70566 331174
rect 70330 330618 70566 330854
rect 101050 330938 101286 331174
rect 101050 330618 101286 330854
rect 131770 330938 132006 331174
rect 131770 330618 132006 330854
rect 162490 330938 162726 331174
rect 162490 330618 162726 330854
rect 193210 330938 193446 331174
rect 193210 330618 193446 330854
rect 223930 330938 224166 331174
rect 223930 330618 224166 330854
rect 254650 330938 254886 331174
rect 254650 330618 254886 330854
rect 285370 330938 285606 331174
rect 285370 330618 285606 330854
rect 316090 330938 316326 331174
rect 316090 330618 316326 330854
rect 346810 330938 347046 331174
rect 346810 330618 347046 330854
rect 85690 327218 85926 327454
rect 85690 326898 85926 327134
rect 116410 327218 116646 327454
rect 116410 326898 116646 327134
rect 147130 327218 147366 327454
rect 147130 326898 147366 327134
rect 177850 327218 178086 327454
rect 177850 326898 178086 327134
rect 208570 327218 208806 327454
rect 208570 326898 208806 327134
rect 239290 327218 239526 327454
rect 239290 326898 239526 327134
rect 270010 327218 270246 327454
rect 270010 326898 270246 327134
rect 300730 327218 300966 327454
rect 300730 326898 300966 327134
rect 331450 327218 331686 327454
rect 331450 326898 331686 327134
rect 362170 327218 362406 327454
rect 362170 326898 362406 327134
rect 63866 317258 64102 317494
rect 64186 317258 64422 317494
rect 63866 316938 64102 317174
rect 64186 316938 64422 317174
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 377530 330938 377766 331174
rect 377530 330618 377766 330854
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 70330 294938 70566 295174
rect 70330 294618 70566 294854
rect 101050 294938 101286 295174
rect 101050 294618 101286 294854
rect 131770 294938 132006 295174
rect 131770 294618 132006 294854
rect 162490 294938 162726 295174
rect 162490 294618 162726 294854
rect 193210 294938 193446 295174
rect 193210 294618 193446 294854
rect 223930 294938 224166 295174
rect 223930 294618 224166 294854
rect 254650 294938 254886 295174
rect 254650 294618 254886 294854
rect 285370 294938 285606 295174
rect 285370 294618 285606 294854
rect 316090 294938 316326 295174
rect 316090 294618 316326 294854
rect 346810 294938 347046 295174
rect 346810 294618 347046 294854
rect 85690 291218 85926 291454
rect 85690 290898 85926 291134
rect 116410 291218 116646 291454
rect 116410 290898 116646 291134
rect 147130 291218 147366 291454
rect 147130 290898 147366 291134
rect 177850 291218 178086 291454
rect 177850 290898 178086 291134
rect 208570 291218 208806 291454
rect 208570 290898 208806 291134
rect 239290 291218 239526 291454
rect 239290 290898 239526 291134
rect 270010 291218 270246 291454
rect 270010 290898 270246 291134
rect 300730 291218 300966 291454
rect 300730 290898 300966 291134
rect 331450 291218 331686 291454
rect 331450 290898 331686 291134
rect 362170 291218 362406 291454
rect 362170 290898 362406 291134
rect 63866 281258 64102 281494
rect 64186 281258 64422 281494
rect 63866 280938 64102 281174
rect 64186 280938 64422 281174
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 377530 294938 377766 295174
rect 377530 294618 377766 294854
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 70330 258938 70566 259174
rect 70330 258618 70566 258854
rect 101050 258938 101286 259174
rect 101050 258618 101286 258854
rect 131770 258938 132006 259174
rect 131770 258618 132006 258854
rect 162490 258938 162726 259174
rect 162490 258618 162726 258854
rect 193210 258938 193446 259174
rect 193210 258618 193446 258854
rect 223930 258938 224166 259174
rect 223930 258618 224166 258854
rect 254650 258938 254886 259174
rect 254650 258618 254886 258854
rect 285370 258938 285606 259174
rect 285370 258618 285606 258854
rect 316090 258938 316326 259174
rect 316090 258618 316326 258854
rect 346810 258938 347046 259174
rect 346810 258618 347046 258854
rect 85690 255218 85926 255454
rect 85690 254898 85926 255134
rect 116410 255218 116646 255454
rect 116410 254898 116646 255134
rect 147130 255218 147366 255454
rect 147130 254898 147366 255134
rect 177850 255218 178086 255454
rect 177850 254898 178086 255134
rect 208570 255218 208806 255454
rect 208570 254898 208806 255134
rect 239290 255218 239526 255454
rect 239290 254898 239526 255134
rect 270010 255218 270246 255454
rect 270010 254898 270246 255134
rect 300730 255218 300966 255454
rect 300730 254898 300966 255134
rect 331450 255218 331686 255454
rect 331450 254898 331686 255134
rect 362170 255218 362406 255454
rect 362170 254898 362406 255134
rect 63866 245258 64102 245494
rect 64186 245258 64422 245494
rect 63866 244938 64102 245174
rect 64186 244938 64422 245174
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 377530 258938 377766 259174
rect 377530 258618 377766 258854
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 70330 222938 70566 223174
rect 70330 222618 70566 222854
rect 101050 222938 101286 223174
rect 101050 222618 101286 222854
rect 131770 222938 132006 223174
rect 131770 222618 132006 222854
rect 162490 222938 162726 223174
rect 162490 222618 162726 222854
rect 193210 222938 193446 223174
rect 193210 222618 193446 222854
rect 223930 222938 224166 223174
rect 223930 222618 224166 222854
rect 254650 222938 254886 223174
rect 254650 222618 254886 222854
rect 285370 222938 285606 223174
rect 285370 222618 285606 222854
rect 316090 222938 316326 223174
rect 316090 222618 316326 222854
rect 346810 222938 347046 223174
rect 346810 222618 347046 222854
rect 85690 219218 85926 219454
rect 85690 218898 85926 219134
rect 116410 219218 116646 219454
rect 116410 218898 116646 219134
rect 147130 219218 147366 219454
rect 147130 218898 147366 219134
rect 177850 219218 178086 219454
rect 177850 218898 178086 219134
rect 208570 219218 208806 219454
rect 208570 218898 208806 219134
rect 239290 219218 239526 219454
rect 239290 218898 239526 219134
rect 270010 219218 270246 219454
rect 270010 218898 270246 219134
rect 300730 219218 300966 219454
rect 300730 218898 300966 219134
rect 331450 219218 331686 219454
rect 331450 218898 331686 219134
rect 362170 219218 362406 219454
rect 362170 218898 362406 219134
rect 63866 209258 64102 209494
rect 64186 209258 64422 209494
rect 63866 208938 64102 209174
rect 64186 208938 64422 209174
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 377530 222938 377766 223174
rect 377530 222618 377766 222854
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 70330 186938 70566 187174
rect 70330 186618 70566 186854
rect 101050 186938 101286 187174
rect 101050 186618 101286 186854
rect 131770 186938 132006 187174
rect 131770 186618 132006 186854
rect 162490 186938 162726 187174
rect 162490 186618 162726 186854
rect 193210 186938 193446 187174
rect 193210 186618 193446 186854
rect 223930 186938 224166 187174
rect 223930 186618 224166 186854
rect 254650 186938 254886 187174
rect 254650 186618 254886 186854
rect 285370 186938 285606 187174
rect 285370 186618 285606 186854
rect 316090 186938 316326 187174
rect 316090 186618 316326 186854
rect 346810 186938 347046 187174
rect 346810 186618 347046 186854
rect 85690 183218 85926 183454
rect 85690 182898 85926 183134
rect 116410 183218 116646 183454
rect 116410 182898 116646 183134
rect 147130 183218 147366 183454
rect 147130 182898 147366 183134
rect 177850 183218 178086 183454
rect 177850 182898 178086 183134
rect 208570 183218 208806 183454
rect 208570 182898 208806 183134
rect 239290 183218 239526 183454
rect 239290 182898 239526 183134
rect 270010 183218 270246 183454
rect 270010 182898 270246 183134
rect 300730 183218 300966 183454
rect 300730 182898 300966 183134
rect 331450 183218 331686 183454
rect 331450 182898 331686 183134
rect 362170 183218 362406 183454
rect 362170 182898 362406 183134
rect 63866 173258 64102 173494
rect 64186 173258 64422 173494
rect 63866 172938 64102 173174
rect 64186 172938 64422 173174
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 377530 186938 377766 187174
rect 377530 186618 377766 186854
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 70330 150938 70566 151174
rect 70330 150618 70566 150854
rect 101050 150938 101286 151174
rect 101050 150618 101286 150854
rect 131770 150938 132006 151174
rect 131770 150618 132006 150854
rect 162490 150938 162726 151174
rect 162490 150618 162726 150854
rect 193210 150938 193446 151174
rect 193210 150618 193446 150854
rect 223930 150938 224166 151174
rect 223930 150618 224166 150854
rect 254650 150938 254886 151174
rect 254650 150618 254886 150854
rect 285370 150938 285606 151174
rect 285370 150618 285606 150854
rect 316090 150938 316326 151174
rect 316090 150618 316326 150854
rect 346810 150938 347046 151174
rect 346810 150618 347046 150854
rect 85690 147218 85926 147454
rect 85690 146898 85926 147134
rect 116410 147218 116646 147454
rect 116410 146898 116646 147134
rect 147130 147218 147366 147454
rect 147130 146898 147366 147134
rect 177850 147218 178086 147454
rect 177850 146898 178086 147134
rect 208570 147218 208806 147454
rect 208570 146898 208806 147134
rect 239290 147218 239526 147454
rect 239290 146898 239526 147134
rect 270010 147218 270246 147454
rect 270010 146898 270246 147134
rect 300730 147218 300966 147454
rect 300730 146898 300966 147134
rect 331450 147218 331686 147454
rect 331450 146898 331686 147134
rect 362170 147218 362406 147454
rect 362170 146898 362406 147134
rect 63866 137258 64102 137494
rect 64186 137258 64422 137494
rect 63866 136938 64102 137174
rect 64186 136938 64422 137174
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 377530 150938 377766 151174
rect 377530 150618 377766 150854
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 70330 114938 70566 115174
rect 70330 114618 70566 114854
rect 101050 114938 101286 115174
rect 101050 114618 101286 114854
rect 131770 114938 132006 115174
rect 131770 114618 132006 114854
rect 162490 114938 162726 115174
rect 162490 114618 162726 114854
rect 193210 114938 193446 115174
rect 193210 114618 193446 114854
rect 223930 114938 224166 115174
rect 223930 114618 224166 114854
rect 254650 114938 254886 115174
rect 254650 114618 254886 114854
rect 285370 114938 285606 115174
rect 285370 114618 285606 114854
rect 316090 114938 316326 115174
rect 316090 114618 316326 114854
rect 346810 114938 347046 115174
rect 346810 114618 347046 114854
rect 85690 111218 85926 111454
rect 85690 110898 85926 111134
rect 116410 111218 116646 111454
rect 116410 110898 116646 111134
rect 147130 111218 147366 111454
rect 147130 110898 147366 111134
rect 177850 111218 178086 111454
rect 177850 110898 178086 111134
rect 208570 111218 208806 111454
rect 208570 110898 208806 111134
rect 239290 111218 239526 111454
rect 239290 110898 239526 111134
rect 270010 111218 270246 111454
rect 270010 110898 270246 111134
rect 300730 111218 300966 111454
rect 300730 110898 300966 111134
rect 331450 111218 331686 111454
rect 331450 110898 331686 111134
rect 362170 111218 362406 111454
rect 362170 110898 362406 111134
rect 63866 101258 64102 101494
rect 64186 101258 64422 101494
rect 63866 100938 64102 101174
rect 64186 100938 64422 101174
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 377530 114938 377766 115174
rect 377530 114618 377766 114854
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 70330 78938 70566 79174
rect 70330 78618 70566 78854
rect 101050 78938 101286 79174
rect 101050 78618 101286 78854
rect 131770 78938 132006 79174
rect 131770 78618 132006 78854
rect 162490 78938 162726 79174
rect 162490 78618 162726 78854
rect 193210 78938 193446 79174
rect 193210 78618 193446 78854
rect 223930 78938 224166 79174
rect 223930 78618 224166 78854
rect 254650 78938 254886 79174
rect 254650 78618 254886 78854
rect 285370 78938 285606 79174
rect 285370 78618 285606 78854
rect 316090 78938 316326 79174
rect 316090 78618 316326 78854
rect 346810 78938 347046 79174
rect 346810 78618 347046 78854
rect 85690 75218 85926 75454
rect 85690 74898 85926 75134
rect 116410 75218 116646 75454
rect 116410 74898 116646 75134
rect 147130 75218 147366 75454
rect 147130 74898 147366 75134
rect 177850 75218 178086 75454
rect 177850 74898 178086 75134
rect 208570 75218 208806 75454
rect 208570 74898 208806 75134
rect 239290 75218 239526 75454
rect 239290 74898 239526 75134
rect 270010 75218 270246 75454
rect 270010 74898 270246 75134
rect 300730 75218 300966 75454
rect 300730 74898 300966 75134
rect 331450 75218 331686 75454
rect 331450 74898 331686 75134
rect 362170 75218 362406 75454
rect 362170 74898 362406 75134
rect 63866 65258 64102 65494
rect 64186 65258 64422 65494
rect 63866 64938 64102 65174
rect 64186 64938 64422 65174
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 54098 88942 54334
rect 89026 54098 89262 54334
rect 88706 53778 88942 54014
rect 89026 53778 89262 54014
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 57818 92662 58054
rect 92746 57818 92982 58054
rect 92426 57498 92662 57734
rect 92746 57498 92982 57734
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 54098 124942 54334
rect 125026 54098 125262 54334
rect 124706 53778 124942 54014
rect 125026 53778 125262 54014
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 57818 128662 58054
rect 128746 57818 128982 58054
rect 128426 57498 128662 57734
rect 128746 57498 128982 57734
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 54098 160942 54334
rect 161026 54098 161262 54334
rect 160706 53778 160942 54014
rect 161026 53778 161262 54014
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 57818 164662 58054
rect 164746 57818 164982 58054
rect 164426 57498 164662 57734
rect 164746 57498 164982 57734
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 57818 200662 58054
rect 200746 57818 200982 58054
rect 200426 57498 200662 57734
rect 200746 57498 200982 57734
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 54098 232942 54334
rect 233026 54098 233262 54334
rect 232706 53778 232942 54014
rect 233026 53778 233262 54014
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 57818 236662 58054
rect 236746 57818 236982 58054
rect 236426 57498 236662 57734
rect 236746 57498 236982 57734
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 54098 268942 54334
rect 269026 54098 269262 54334
rect 268706 53778 268942 54014
rect 269026 53778 269262 54014
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 57818 272662 58054
rect 272746 57818 272982 58054
rect 272426 57498 272662 57734
rect 272746 57498 272982 57734
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 304706 54098 304942 54334
rect 305026 54098 305262 54334
rect 304706 53778 304942 54014
rect 305026 53778 305262 54014
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 57818 308662 58054
rect 308746 57818 308982 58054
rect 308426 57498 308662 57734
rect 308746 57498 308982 57734
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 54098 340942 54334
rect 341026 54098 341262 54334
rect 340706 53778 340942 54014
rect 341026 53778 341262 54014
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 57818 344662 58054
rect 344746 57818 344982 58054
rect 344426 57498 344662 57734
rect 344746 57498 344982 57734
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 377530 78938 377766 79174
rect 377530 78618 377766 78854
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 387866 65258 388102 65494
rect 388186 65258 388422 65494
rect 387866 64938 388102 65174
rect 388186 64938 388422 65174
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 404700 327218 404936 327454
rect 404700 326898 404936 327134
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408414 330938 408650 331174
rect 408414 330618 408650 330854
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 412128 327218 412364 327454
rect 412128 326898 412364 327134
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 415842 330938 416078 331174
rect 415842 330618 416078 330854
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 426666 438938 426902 439174
rect 426666 438618 426902 438854
rect 432347 438938 432583 439174
rect 432347 438618 432583 438854
rect 438028 438938 438264 439174
rect 438028 438618 438264 438854
rect 443709 438938 443945 439174
rect 443709 438618 443945 438854
rect 423826 435218 424062 435454
rect 423826 434898 424062 435134
rect 429507 435218 429743 435454
rect 429507 434898 429743 435134
rect 435188 435218 435424 435454
rect 435188 434898 435424 435134
rect 440869 435218 441105 435454
rect 440869 434898 441105 435134
rect 420146 421538 420382 421774
rect 420466 421538 420702 421774
rect 420146 421218 420382 421454
rect 420466 421218 420702 421454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 419556 327218 419792 327454
rect 419556 326898 419792 327134
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 423270 330938 423506 331174
rect 423270 330618 423506 330854
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 430698 330938 430934 331174
rect 430698 330618 430934 330854
rect 426984 327218 427220 327454
rect 426984 326898 427220 327134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 484706 708442 484942 708678
rect 485026 708442 485262 708678
rect 484706 708122 484942 708358
rect 485026 708122 485262 708358
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 479610 654938 479846 655174
rect 479610 654618 479846 654854
rect 510330 654938 510566 655174
rect 510330 654618 510566 654854
rect 464250 651218 464486 651454
rect 464250 650898 464486 651134
rect 494970 651218 495206 651454
rect 494970 650898 495206 651134
rect 525690 651218 525926 651454
rect 525690 650898 525926 651134
rect 528146 637538 528382 637774
rect 528466 637538 528702 637774
rect 528146 637218 528382 637454
rect 528466 637218 528702 637454
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 453424 510938 453660 511174
rect 453424 510618 453660 510854
rect 455862 510938 456098 511174
rect 455862 510618 456098 510854
rect 458300 510938 458536 511174
rect 458300 510618 458536 510854
rect 452205 507218 452441 507454
rect 452205 506898 452441 507134
rect 454643 507218 454879 507454
rect 454643 506898 454879 507134
rect 457081 507218 457317 507454
rect 457081 506898 457317 507134
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 456146 421538 456382 421774
rect 456466 421538 456702 421774
rect 456146 421218 456382 421454
rect 456466 421218 456702 421454
rect 479610 618938 479846 619174
rect 479610 618618 479846 618854
rect 510330 618938 510566 619174
rect 510330 618618 510566 618854
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 525690 615218 525926 615454
rect 525690 614898 525926 615134
rect 459866 605258 460102 605494
rect 460186 605258 460422 605494
rect 459866 604938 460102 605174
rect 460186 604938 460422 605174
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 460738 510938 460974 511174
rect 460738 510618 460974 510854
rect 459519 507218 459755 507454
rect 459519 506898 459755 507134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 454250 363218 454486 363454
rect 454250 362898 454486 363134
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 454250 327218 454486 327454
rect 454250 326898 454486 327134
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 429610 150938 429846 151174
rect 429610 150618 429846 150854
rect 414250 147218 414486 147454
rect 414250 146898 414486 147134
rect 444970 147218 445206 147454
rect 444970 146898 445206 147134
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 412706 90098 412942 90334
rect 413026 90098 413262 90334
rect 412706 89778 412942 90014
rect 413026 89778 413262 90014
rect 412706 54098 412942 54334
rect 413026 54098 413262 54334
rect 412706 53778 412942 54014
rect 413026 53778 413262 54014
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 129818 416662 130054
rect 416746 129818 416982 130054
rect 416426 129498 416662 129734
rect 416746 129498 416982 129734
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 416426 57818 416662 58054
rect 416746 57818 416982 58054
rect 416426 57498 416662 57734
rect 416746 57498 416982 57734
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 133538 420382 133774
rect 420466 133538 420702 133774
rect 420146 133218 420382 133454
rect 420466 133218 420702 133454
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 420146 61538 420382 61774
rect 420466 61538 420702 61774
rect 420146 61218 420382 61454
rect 420466 61218 420702 61454
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 423866 65258 424102 65494
rect 424186 65258 424422 65494
rect 423866 64938 424102 65174
rect 424186 64938 424422 65174
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 90098 448942 90334
rect 449026 90098 449262 90334
rect 448706 89778 448942 90014
rect 449026 89778 449262 90014
rect 448706 54098 448942 54334
rect 449026 54098 449262 54334
rect 448706 53778 448942 54014
rect 449026 53778 449262 54014
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 452426 57818 452662 58054
rect 452746 57818 452982 58054
rect 452426 57498 452662 57734
rect 452746 57498 452982 57734
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473700 435218 473936 435454
rect 473700 434898 473936 435134
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 469610 366938 469846 367174
rect 469610 366618 469846 366854
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 476414 438938 476650 439174
rect 476414 438618 476650 438854
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 492146 601538 492382 601774
rect 492466 601538 492702 601774
rect 492146 601218 492382 601454
rect 492466 601218 492702 601454
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 482205 507218 482441 507454
rect 482205 506898 482441 507134
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 483424 510938 483660 511174
rect 483424 510618 483660 510854
rect 485862 510938 486098 511174
rect 485862 510618 486098 510854
rect 488300 510938 488536 511174
rect 488300 510618 488536 510854
rect 484643 507218 484879 507454
rect 484643 506898 484879 507134
rect 487081 507218 487317 507454
rect 487081 506898 487317 507134
rect 489519 507218 489755 507454
rect 489519 506898 489755 507134
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 479128 435218 479364 435454
rect 479128 434898 479364 435134
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 488426 453818 488662 454054
rect 488746 453818 488982 454054
rect 488426 453498 488662 453734
rect 488746 453498 488982 453734
rect 481842 438938 482078 439174
rect 481842 438618 482078 438854
rect 487270 438938 487506 439174
rect 487270 438618 487506 438854
rect 484556 435218 484792 435454
rect 484556 434898 484792 435134
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 489984 435218 490220 435454
rect 489984 434898 490220 435134
rect 488426 417818 488662 418054
rect 488746 417818 488982 418054
rect 488426 417498 488662 417734
rect 488746 417498 488982 417734
rect 490738 510938 490974 511174
rect 490738 510618 490974 510854
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 495866 605258 496102 605494
rect 496186 605258 496422 605494
rect 495866 604938 496102 605174
rect 496186 604938 496422 605174
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 492698 438938 492934 439174
rect 492698 438618 492934 438854
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 492146 385538 492382 385774
rect 492466 385538 492702 385774
rect 492146 385218 492382 385454
rect 492466 385218 492702 385454
rect 488426 381818 488662 382054
rect 488746 381818 488982 382054
rect 488426 381498 488662 381734
rect 488746 381498 488982 381734
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 469610 330938 469846 331174
rect 469610 330618 469846 330854
rect 500330 366938 500566 367174
rect 500330 366618 500566 366854
rect 484970 363218 485206 363454
rect 484970 362898 485206 363134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 500330 330938 500566 331174
rect 500330 330618 500566 330854
rect 484970 327218 485206 327454
rect 484970 326898 485206 327134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 528146 601538 528382 601774
rect 528466 601538 528702 601774
rect 528146 601218 528382 601454
rect 528466 601218 528702 601454
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 524250 435218 524486 435454
rect 524250 434898 524486 435134
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541050 654938 541286 655174
rect 541050 654618 541286 654854
rect 531866 641258 532102 641494
rect 532186 641258 532422 641494
rect 531866 640938 532102 641174
rect 532186 640938 532422 641174
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541050 618938 541286 619174
rect 541050 618618 541286 618854
rect 531866 605258 532102 605494
rect 532186 605258 532422 605494
rect 531866 604938 532102 605174
rect 532186 604938 532422 605174
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 539610 438938 539846 439174
rect 539610 438618 539846 438854
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 479610 258938 479846 259174
rect 479610 258618 479846 258854
rect 510330 258938 510566 259174
rect 510330 258618 510566 258854
rect 464250 255218 464486 255454
rect 464250 254898 464486 255134
rect 494970 255218 495206 255454
rect 494970 254898 495206 255134
rect 525690 255218 525926 255454
rect 525690 254898 525926 255134
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 479610 222938 479846 223174
rect 479610 222618 479846 222854
rect 510330 222938 510566 223174
rect 510330 222618 510566 222854
rect 464250 219218 464486 219454
rect 464250 218898 464486 219134
rect 494970 219218 495206 219454
rect 494970 218898 495206 219134
rect 525690 219218 525926 219454
rect 525690 218898 525926 219134
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 456146 61538 456382 61774
rect 456466 61538 456702 61774
rect 456146 61218 456382 61454
rect 456466 61218 456702 61454
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 484250 147218 484486 147454
rect 484250 146898 484486 147134
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484250 111218 484486 111454
rect 484250 110898 484486 111134
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 488426 129818 488662 130054
rect 488746 129818 488982 130054
rect 488426 129498 488662 129734
rect 488746 129498 488982 129734
rect 488426 93818 488662 94054
rect 488746 93818 488982 94054
rect 488426 93498 488662 93734
rect 488746 93498 488982 93734
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 169538 492382 169774
rect 492466 169538 492702 169774
rect 492146 169218 492382 169454
rect 492466 169218 492702 169454
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 514970 147218 515206 147454
rect 514970 146898 515206 147134
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 554970 435218 555206 435454
rect 554970 434898 555206 435134
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 555424 366938 555660 367174
rect 555424 366618 555660 366854
rect 553205 363218 553441 363454
rect 553205 362898 553441 363134
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 492146 133538 492382 133774
rect 492466 133538 492702 133774
rect 492146 133218 492382 133454
rect 492466 133218 492702 133454
rect 499610 114938 499846 115174
rect 499610 114618 499846 114854
rect 530330 114938 530566 115174
rect 530330 114618 530566 114854
rect 514970 111218 515206 111454
rect 514970 110898 515206 111134
rect 545690 147218 545926 147454
rect 545690 146898 545926 147134
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 492146 97538 492382 97774
rect 492466 97538 492702 97774
rect 492146 97218 492382 97454
rect 492466 97218 492702 97454
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 545690 111218 545926 111454
rect 545690 110898 545926 111134
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 557644 363218 557880 363454
rect 557644 362898 557880 363134
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 559863 366938 560099 367174
rect 559863 366618 560099 366854
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 564302 366938 564538 367174
rect 564302 366618 564538 366854
rect 562083 363218 562319 363454
rect 562083 362898 562319 363134
rect 566522 363218 566758 363454
rect 566522 362898 566758 363134
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 53999 556942 54235
rect 557026 53999 557262 54235
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 543700 39218 543936 39454
rect 543700 38898 543936 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546414 42938 546650 43174
rect 546414 42618 546650 42854
rect 551842 42938 552078 43174
rect 551842 42618 552078 42854
rect 557270 42938 557506 43174
rect 557270 42618 557506 42854
rect 549128 39218 549364 39454
rect 549128 38898 549364 39134
rect 554556 39218 554792 39454
rect 554556 38898 554792 39134
rect 559984 39218 560220 39454
rect 559984 38898 560220 39134
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 562698 42938 562934 43174
rect 562698 42618 562934 42854
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 568741 366938 568977 367174
rect 568741 366618 568977 366854
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 39610 655174
rect 39846 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 70330 655174
rect 70566 654938 101050 655174
rect 101286 654938 131770 655174
rect 132006 654938 162490 655174
rect 162726 654938 193210 655174
rect 193446 654938 223930 655174
rect 224166 654938 254650 655174
rect 254886 654938 285370 655174
rect 285606 654938 316090 655174
rect 316326 654938 346810 655174
rect 347046 654938 377530 655174
rect 377766 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 479610 655174
rect 479846 654938 510330 655174
rect 510566 654938 541050 655174
rect 541286 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 39610 654854
rect 39846 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 70330 654854
rect 70566 654618 101050 654854
rect 101286 654618 131770 654854
rect 132006 654618 162490 654854
rect 162726 654618 193210 654854
rect 193446 654618 223930 654854
rect 224166 654618 254650 654854
rect 254886 654618 285370 654854
rect 285606 654618 316090 654854
rect 316326 654618 346810 654854
rect 347046 654618 377530 654854
rect 377766 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 479610 654854
rect 479846 654618 510330 654854
rect 510566 654618 541050 654854
rect 541286 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 24250 651454
rect 24486 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 54970 651454
rect 55206 651218 85690 651454
rect 85926 651218 116410 651454
rect 116646 651218 147130 651454
rect 147366 651218 177850 651454
rect 178086 651218 208570 651454
rect 208806 651218 239290 651454
rect 239526 651218 270010 651454
rect 270246 651218 300730 651454
rect 300966 651218 331450 651454
rect 331686 651218 362170 651454
rect 362406 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 464250 651454
rect 464486 651218 494970 651454
rect 495206 651218 525690 651454
rect 525926 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 24250 651134
rect 24486 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 54970 651134
rect 55206 650898 85690 651134
rect 85926 650898 116410 651134
rect 116646 650898 147130 651134
rect 147366 650898 177850 651134
rect 178086 650898 208570 651134
rect 208806 650898 239290 651134
rect 239526 650898 270010 651134
rect 270246 650898 300730 651134
rect 300966 650898 331450 651134
rect 331686 650898 362170 651134
rect 362406 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 464250 651134
rect 464486 650898 494970 651134
rect 495206 650898 525690 651134
rect 525926 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 39610 619174
rect 39846 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 70330 619174
rect 70566 618938 101050 619174
rect 101286 618938 131770 619174
rect 132006 618938 162490 619174
rect 162726 618938 193210 619174
rect 193446 618938 223930 619174
rect 224166 618938 254650 619174
rect 254886 618938 285370 619174
rect 285606 618938 316090 619174
rect 316326 618938 346810 619174
rect 347046 618938 377530 619174
rect 377766 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 479610 619174
rect 479846 618938 510330 619174
rect 510566 618938 541050 619174
rect 541286 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 39610 618854
rect 39846 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 70330 618854
rect 70566 618618 101050 618854
rect 101286 618618 131770 618854
rect 132006 618618 162490 618854
rect 162726 618618 193210 618854
rect 193446 618618 223930 618854
rect 224166 618618 254650 618854
rect 254886 618618 285370 618854
rect 285606 618618 316090 618854
rect 316326 618618 346810 618854
rect 347046 618618 377530 618854
rect 377766 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 479610 618854
rect 479846 618618 510330 618854
rect 510566 618618 541050 618854
rect 541286 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 24250 615454
rect 24486 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 54970 615454
rect 55206 615218 85690 615454
rect 85926 615218 116410 615454
rect 116646 615218 147130 615454
rect 147366 615218 177850 615454
rect 178086 615218 208570 615454
rect 208806 615218 239290 615454
rect 239526 615218 270010 615454
rect 270246 615218 300730 615454
rect 300966 615218 331450 615454
rect 331686 615218 362170 615454
rect 362406 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 525690 615454
rect 525926 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 24250 615134
rect 24486 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 54970 615134
rect 55206 614898 85690 615134
rect 85926 614898 116410 615134
rect 116646 614898 147130 615134
rect 147366 614898 177850 615134
rect 178086 614898 208570 615134
rect 208806 614898 239290 615134
rect 239526 614898 270010 615134
rect 270246 614898 300730 615134
rect 300966 614898 331450 615134
rect 331686 614898 362170 615134
rect 362406 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 525690 615134
rect 525926 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 495866 605494
rect 496102 605258 496186 605494
rect 496422 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 495866 605174
rect 496102 604938 496186 605174
rect 496422 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 39610 583174
rect 39846 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 70330 583174
rect 70566 582938 101050 583174
rect 101286 582938 131770 583174
rect 132006 582938 162490 583174
rect 162726 582938 193210 583174
rect 193446 582938 223930 583174
rect 224166 582938 254650 583174
rect 254886 582938 285370 583174
rect 285606 582938 316090 583174
rect 316326 582938 346810 583174
rect 347046 582938 377530 583174
rect 377766 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 39610 582854
rect 39846 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 70330 582854
rect 70566 582618 101050 582854
rect 101286 582618 131770 582854
rect 132006 582618 162490 582854
rect 162726 582618 193210 582854
rect 193446 582618 223930 582854
rect 224166 582618 254650 582854
rect 254886 582618 285370 582854
rect 285606 582618 316090 582854
rect 316326 582618 346810 582854
rect 347046 582618 377530 582854
rect 377766 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 24250 579454
rect 24486 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 54970 579454
rect 55206 579218 85690 579454
rect 85926 579218 116410 579454
rect 116646 579218 147130 579454
rect 147366 579218 177850 579454
rect 178086 579218 208570 579454
rect 208806 579218 239290 579454
rect 239526 579218 270010 579454
rect 270246 579218 300730 579454
rect 300966 579218 331450 579454
rect 331686 579218 362170 579454
rect 362406 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 24250 579134
rect 24486 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 54970 579134
rect 55206 578898 85690 579134
rect 85926 578898 116410 579134
rect 116646 578898 147130 579134
rect 147366 578898 177850 579134
rect 178086 578898 208570 579134
rect 208806 578898 239290 579134
rect 239526 578898 270010 579134
rect 270246 578898 300730 579134
rect 300966 578898 331450 579134
rect 331686 578898 362170 579134
rect 362406 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 63866 569494
rect 64102 569258 64186 569494
rect 64422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 63866 569174
rect 64102 568938 64186 569174
rect 64422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 39610 547174
rect 39846 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 70330 547174
rect 70566 546938 101050 547174
rect 101286 546938 131770 547174
rect 132006 546938 162490 547174
rect 162726 546938 193210 547174
rect 193446 546938 223930 547174
rect 224166 546938 254650 547174
rect 254886 546938 285370 547174
rect 285606 546938 316090 547174
rect 316326 546938 346810 547174
rect 347046 546938 377530 547174
rect 377766 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 39610 546854
rect 39846 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 70330 546854
rect 70566 546618 101050 546854
rect 101286 546618 131770 546854
rect 132006 546618 162490 546854
rect 162726 546618 193210 546854
rect 193446 546618 223930 546854
rect 224166 546618 254650 546854
rect 254886 546618 285370 546854
rect 285606 546618 316090 546854
rect 316326 546618 346810 546854
rect 347046 546618 377530 546854
rect 377766 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 24250 543454
rect 24486 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 54970 543454
rect 55206 543218 85690 543454
rect 85926 543218 116410 543454
rect 116646 543218 147130 543454
rect 147366 543218 177850 543454
rect 178086 543218 208570 543454
rect 208806 543218 239290 543454
rect 239526 543218 270010 543454
rect 270246 543218 300730 543454
rect 300966 543218 331450 543454
rect 331686 543218 362170 543454
rect 362406 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 24250 543134
rect 24486 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 54970 543134
rect 55206 542898 85690 543134
rect 85926 542898 116410 543134
rect 116646 542898 147130 543134
rect 147366 542898 177850 543134
rect 178086 542898 208570 543134
rect 208806 542898 239290 543134
rect 239526 542898 270010 543134
rect 270246 542898 300730 543134
rect 300966 542898 331450 543134
rect 331686 542898 362170 543134
rect 362406 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 63866 533494
rect 64102 533258 64186 533494
rect 64422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 63866 533174
rect 64102 532938 64186 533174
rect 64422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 39610 511174
rect 39846 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 70330 511174
rect 70566 510938 101050 511174
rect 101286 510938 131770 511174
rect 132006 510938 162490 511174
rect 162726 510938 193210 511174
rect 193446 510938 223930 511174
rect 224166 510938 254650 511174
rect 254886 510938 285370 511174
rect 285606 510938 316090 511174
rect 316326 510938 346810 511174
rect 347046 510938 377530 511174
rect 377766 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 453424 511174
rect 453660 510938 455862 511174
rect 456098 510938 458300 511174
rect 458536 510938 460738 511174
rect 460974 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 483424 511174
rect 483660 510938 485862 511174
rect 486098 510938 488300 511174
rect 488536 510938 490738 511174
rect 490974 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 39610 510854
rect 39846 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 70330 510854
rect 70566 510618 101050 510854
rect 101286 510618 131770 510854
rect 132006 510618 162490 510854
rect 162726 510618 193210 510854
rect 193446 510618 223930 510854
rect 224166 510618 254650 510854
rect 254886 510618 285370 510854
rect 285606 510618 316090 510854
rect 316326 510618 346810 510854
rect 347046 510618 377530 510854
rect 377766 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 453424 510854
rect 453660 510618 455862 510854
rect 456098 510618 458300 510854
rect 458536 510618 460738 510854
rect 460974 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 483424 510854
rect 483660 510618 485862 510854
rect 486098 510618 488300 510854
rect 488536 510618 490738 510854
rect 490974 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 24250 507454
rect 24486 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 54970 507454
rect 55206 507218 85690 507454
rect 85926 507218 116410 507454
rect 116646 507218 147130 507454
rect 147366 507218 177850 507454
rect 178086 507218 208570 507454
rect 208806 507218 239290 507454
rect 239526 507218 270010 507454
rect 270246 507218 300730 507454
rect 300966 507218 331450 507454
rect 331686 507218 362170 507454
rect 362406 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 452205 507454
rect 452441 507218 454643 507454
rect 454879 507218 457081 507454
rect 457317 507218 459519 507454
rect 459755 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 482205 507454
rect 482441 507218 484643 507454
rect 484879 507218 487081 507454
rect 487317 507218 489519 507454
rect 489755 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 24250 507134
rect 24486 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 54970 507134
rect 55206 506898 85690 507134
rect 85926 506898 116410 507134
rect 116646 506898 147130 507134
rect 147366 506898 177850 507134
rect 178086 506898 208570 507134
rect 208806 506898 239290 507134
rect 239526 506898 270010 507134
rect 270246 506898 300730 507134
rect 300966 506898 331450 507134
rect 331686 506898 362170 507134
rect 362406 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 452205 507134
rect 452441 506898 454643 507134
rect 454879 506898 457081 507134
rect 457317 506898 459519 507134
rect 459755 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 482205 507134
rect 482441 506898 484643 507134
rect 484879 506898 487081 507134
rect 487317 506898 489519 507134
rect 489755 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 39610 475174
rect 39846 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 70330 475174
rect 70566 474938 101050 475174
rect 101286 474938 131770 475174
rect 132006 474938 162490 475174
rect 162726 474938 193210 475174
rect 193446 474938 223930 475174
rect 224166 474938 254650 475174
rect 254886 474938 285370 475174
rect 285606 474938 316090 475174
rect 316326 474938 346810 475174
rect 347046 474938 377530 475174
rect 377766 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 39610 474854
rect 39846 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 70330 474854
rect 70566 474618 101050 474854
rect 101286 474618 131770 474854
rect 132006 474618 162490 474854
rect 162726 474618 193210 474854
rect 193446 474618 223930 474854
rect 224166 474618 254650 474854
rect 254886 474618 285370 474854
rect 285606 474618 316090 474854
rect 316326 474618 346810 474854
rect 347046 474618 377530 474854
rect 377766 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 24250 471454
rect 24486 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 54970 471454
rect 55206 471218 85690 471454
rect 85926 471218 116410 471454
rect 116646 471218 147130 471454
rect 147366 471218 177850 471454
rect 178086 471218 208570 471454
rect 208806 471218 239290 471454
rect 239526 471218 270010 471454
rect 270246 471218 300730 471454
rect 300966 471218 331450 471454
rect 331686 471218 362170 471454
rect 362406 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 24250 471134
rect 24486 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 54970 471134
rect 55206 470898 85690 471134
rect 85926 470898 116410 471134
rect 116646 470898 147130 471134
rect 147366 470898 177850 471134
rect 178086 470898 208570 471134
rect 208806 470898 239290 471134
rect 239526 470898 270010 471134
rect 270246 470898 300730 471134
rect 300966 470898 331450 471134
rect 331686 470898 362170 471134
rect 362406 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 39610 439174
rect 39846 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 70330 439174
rect 70566 438938 101050 439174
rect 101286 438938 131770 439174
rect 132006 438938 162490 439174
rect 162726 438938 193210 439174
rect 193446 438938 223930 439174
rect 224166 438938 254650 439174
rect 254886 438938 285370 439174
rect 285606 438938 316090 439174
rect 316326 438938 346810 439174
rect 347046 438938 377530 439174
rect 377766 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 426666 439174
rect 426902 438938 432347 439174
rect 432583 438938 438028 439174
rect 438264 438938 443709 439174
rect 443945 438938 476414 439174
rect 476650 438938 481842 439174
rect 482078 438938 487270 439174
rect 487506 438938 492698 439174
rect 492934 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 539610 439174
rect 539846 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 39610 438854
rect 39846 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 70330 438854
rect 70566 438618 101050 438854
rect 101286 438618 131770 438854
rect 132006 438618 162490 438854
rect 162726 438618 193210 438854
rect 193446 438618 223930 438854
rect 224166 438618 254650 438854
rect 254886 438618 285370 438854
rect 285606 438618 316090 438854
rect 316326 438618 346810 438854
rect 347046 438618 377530 438854
rect 377766 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 426666 438854
rect 426902 438618 432347 438854
rect 432583 438618 438028 438854
rect 438264 438618 443709 438854
rect 443945 438618 476414 438854
rect 476650 438618 481842 438854
rect 482078 438618 487270 438854
rect 487506 438618 492698 438854
rect 492934 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 539610 438854
rect 539846 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 24250 435454
rect 24486 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 54970 435454
rect 55206 435218 85690 435454
rect 85926 435218 116410 435454
rect 116646 435218 147130 435454
rect 147366 435218 177850 435454
rect 178086 435218 208570 435454
rect 208806 435218 239290 435454
rect 239526 435218 270010 435454
rect 270246 435218 300730 435454
rect 300966 435218 331450 435454
rect 331686 435218 362170 435454
rect 362406 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 423826 435454
rect 424062 435218 429507 435454
rect 429743 435218 435188 435454
rect 435424 435218 440869 435454
rect 441105 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 473700 435454
rect 473936 435218 479128 435454
rect 479364 435218 484556 435454
rect 484792 435218 489984 435454
rect 490220 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 524250 435454
rect 524486 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 554970 435454
rect 555206 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 24250 435134
rect 24486 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 54970 435134
rect 55206 434898 85690 435134
rect 85926 434898 116410 435134
rect 116646 434898 147130 435134
rect 147366 434898 177850 435134
rect 178086 434898 208570 435134
rect 208806 434898 239290 435134
rect 239526 434898 270010 435134
rect 270246 434898 300730 435134
rect 300966 434898 331450 435134
rect 331686 434898 362170 435134
rect 362406 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 423826 435134
rect 424062 434898 429507 435134
rect 429743 434898 435188 435134
rect 435424 434898 440869 435134
rect 441105 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 473700 435134
rect 473936 434898 479128 435134
rect 479364 434898 484556 435134
rect 484792 434898 489984 435134
rect 490220 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 524250 435134
rect 524486 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 554970 435134
rect 555206 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 39610 403174
rect 39846 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 70330 403174
rect 70566 402938 101050 403174
rect 101286 402938 131770 403174
rect 132006 402938 162490 403174
rect 162726 402938 193210 403174
rect 193446 402938 223930 403174
rect 224166 402938 254650 403174
rect 254886 402938 285370 403174
rect 285606 402938 316090 403174
rect 316326 402938 346810 403174
rect 347046 402938 377530 403174
rect 377766 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 39610 402854
rect 39846 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 70330 402854
rect 70566 402618 101050 402854
rect 101286 402618 131770 402854
rect 132006 402618 162490 402854
rect 162726 402618 193210 402854
rect 193446 402618 223930 402854
rect 224166 402618 254650 402854
rect 254886 402618 285370 402854
rect 285606 402618 316090 402854
rect 316326 402618 346810 402854
rect 347046 402618 377530 402854
rect 377766 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 24250 399454
rect 24486 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 54970 399454
rect 55206 399218 85690 399454
rect 85926 399218 116410 399454
rect 116646 399218 147130 399454
rect 147366 399218 177850 399454
rect 178086 399218 208570 399454
rect 208806 399218 239290 399454
rect 239526 399218 270010 399454
rect 270246 399218 300730 399454
rect 300966 399218 331450 399454
rect 331686 399218 362170 399454
rect 362406 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 24250 399134
rect 24486 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 54970 399134
rect 55206 398898 85690 399134
rect 85926 398898 116410 399134
rect 116646 398898 147130 399134
rect 147366 398898 177850 399134
rect 178086 398898 208570 399134
rect 208806 398898 239290 399134
rect 239526 398898 270010 399134
rect 270246 398898 300730 399134
rect 300966 398898 331450 399134
rect 331686 398898 362170 399134
rect 362406 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 39610 367174
rect 39846 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 70330 367174
rect 70566 366938 101050 367174
rect 101286 366938 131770 367174
rect 132006 366938 162490 367174
rect 162726 366938 193210 367174
rect 193446 366938 223930 367174
rect 224166 366938 254650 367174
rect 254886 366938 285370 367174
rect 285606 366938 316090 367174
rect 316326 366938 346810 367174
rect 347046 366938 377530 367174
rect 377766 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 469610 367174
rect 469846 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 500330 367174
rect 500566 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 555424 367174
rect 555660 366938 559863 367174
rect 560099 366938 564302 367174
rect 564538 366938 568741 367174
rect 568977 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 39610 366854
rect 39846 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 70330 366854
rect 70566 366618 101050 366854
rect 101286 366618 131770 366854
rect 132006 366618 162490 366854
rect 162726 366618 193210 366854
rect 193446 366618 223930 366854
rect 224166 366618 254650 366854
rect 254886 366618 285370 366854
rect 285606 366618 316090 366854
rect 316326 366618 346810 366854
rect 347046 366618 377530 366854
rect 377766 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 469610 366854
rect 469846 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 500330 366854
rect 500566 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 555424 366854
rect 555660 366618 559863 366854
rect 560099 366618 564302 366854
rect 564538 366618 568741 366854
rect 568977 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 24250 363454
rect 24486 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 54970 363454
rect 55206 363218 85690 363454
rect 85926 363218 116410 363454
rect 116646 363218 147130 363454
rect 147366 363218 177850 363454
rect 178086 363218 208570 363454
rect 208806 363218 239290 363454
rect 239526 363218 270010 363454
rect 270246 363218 300730 363454
rect 300966 363218 331450 363454
rect 331686 363218 362170 363454
rect 362406 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 454250 363454
rect 454486 363218 484970 363454
rect 485206 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 553205 363454
rect 553441 363218 557644 363454
rect 557880 363218 562083 363454
rect 562319 363218 566522 363454
rect 566758 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 24250 363134
rect 24486 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 54970 363134
rect 55206 362898 85690 363134
rect 85926 362898 116410 363134
rect 116646 362898 147130 363134
rect 147366 362898 177850 363134
rect 178086 362898 208570 363134
rect 208806 362898 239290 363134
rect 239526 362898 270010 363134
rect 270246 362898 300730 363134
rect 300966 362898 331450 363134
rect 331686 362898 362170 363134
rect 362406 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 454250 363134
rect 454486 362898 484970 363134
rect 485206 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 553205 363134
rect 553441 362898 557644 363134
rect 557880 362898 562083 363134
rect 562319 362898 566522 363134
rect 566758 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 39610 331174
rect 39846 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 70330 331174
rect 70566 330938 101050 331174
rect 101286 330938 131770 331174
rect 132006 330938 162490 331174
rect 162726 330938 193210 331174
rect 193446 330938 223930 331174
rect 224166 330938 254650 331174
rect 254886 330938 285370 331174
rect 285606 330938 316090 331174
rect 316326 330938 346810 331174
rect 347046 330938 377530 331174
rect 377766 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 408414 331174
rect 408650 330938 415842 331174
rect 416078 330938 423270 331174
rect 423506 330938 430698 331174
rect 430934 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 469610 331174
rect 469846 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 500330 331174
rect 500566 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 39610 330854
rect 39846 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 70330 330854
rect 70566 330618 101050 330854
rect 101286 330618 131770 330854
rect 132006 330618 162490 330854
rect 162726 330618 193210 330854
rect 193446 330618 223930 330854
rect 224166 330618 254650 330854
rect 254886 330618 285370 330854
rect 285606 330618 316090 330854
rect 316326 330618 346810 330854
rect 347046 330618 377530 330854
rect 377766 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 408414 330854
rect 408650 330618 415842 330854
rect 416078 330618 423270 330854
rect 423506 330618 430698 330854
rect 430934 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 469610 330854
rect 469846 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 500330 330854
rect 500566 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 24250 327454
rect 24486 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 54970 327454
rect 55206 327218 85690 327454
rect 85926 327218 116410 327454
rect 116646 327218 147130 327454
rect 147366 327218 177850 327454
rect 178086 327218 208570 327454
rect 208806 327218 239290 327454
rect 239526 327218 270010 327454
rect 270246 327218 300730 327454
rect 300966 327218 331450 327454
rect 331686 327218 362170 327454
rect 362406 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 404700 327454
rect 404936 327218 412128 327454
rect 412364 327218 419556 327454
rect 419792 327218 426984 327454
rect 427220 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 454250 327454
rect 454486 327218 484970 327454
rect 485206 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 24250 327134
rect 24486 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 54970 327134
rect 55206 326898 85690 327134
rect 85926 326898 116410 327134
rect 116646 326898 147130 327134
rect 147366 326898 177850 327134
rect 178086 326898 208570 327134
rect 208806 326898 239290 327134
rect 239526 326898 270010 327134
rect 270246 326898 300730 327134
rect 300966 326898 331450 327134
rect 331686 326898 362170 327134
rect 362406 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 404700 327134
rect 404936 326898 412128 327134
rect 412364 326898 419556 327134
rect 419792 326898 426984 327134
rect 427220 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 454250 327134
rect 454486 326898 484970 327134
rect 485206 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 39610 295174
rect 39846 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 70330 295174
rect 70566 294938 101050 295174
rect 101286 294938 131770 295174
rect 132006 294938 162490 295174
rect 162726 294938 193210 295174
rect 193446 294938 223930 295174
rect 224166 294938 254650 295174
rect 254886 294938 285370 295174
rect 285606 294938 316090 295174
rect 316326 294938 346810 295174
rect 347046 294938 377530 295174
rect 377766 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 39610 294854
rect 39846 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 70330 294854
rect 70566 294618 101050 294854
rect 101286 294618 131770 294854
rect 132006 294618 162490 294854
rect 162726 294618 193210 294854
rect 193446 294618 223930 294854
rect 224166 294618 254650 294854
rect 254886 294618 285370 294854
rect 285606 294618 316090 294854
rect 316326 294618 346810 294854
rect 347046 294618 377530 294854
rect 377766 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 24250 291454
rect 24486 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 54970 291454
rect 55206 291218 85690 291454
rect 85926 291218 116410 291454
rect 116646 291218 147130 291454
rect 147366 291218 177850 291454
rect 178086 291218 208570 291454
rect 208806 291218 239290 291454
rect 239526 291218 270010 291454
rect 270246 291218 300730 291454
rect 300966 291218 331450 291454
rect 331686 291218 362170 291454
rect 362406 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 24250 291134
rect 24486 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 54970 291134
rect 55206 290898 85690 291134
rect 85926 290898 116410 291134
rect 116646 290898 147130 291134
rect 147366 290898 177850 291134
rect 178086 290898 208570 291134
rect 208806 290898 239290 291134
rect 239526 290898 270010 291134
rect 270246 290898 300730 291134
rect 300966 290898 331450 291134
rect 331686 290898 362170 291134
rect 362406 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 39610 259174
rect 39846 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 70330 259174
rect 70566 258938 101050 259174
rect 101286 258938 131770 259174
rect 132006 258938 162490 259174
rect 162726 258938 193210 259174
rect 193446 258938 223930 259174
rect 224166 258938 254650 259174
rect 254886 258938 285370 259174
rect 285606 258938 316090 259174
rect 316326 258938 346810 259174
rect 347046 258938 377530 259174
rect 377766 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 479610 259174
rect 479846 258938 510330 259174
rect 510566 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 39610 258854
rect 39846 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 70330 258854
rect 70566 258618 101050 258854
rect 101286 258618 131770 258854
rect 132006 258618 162490 258854
rect 162726 258618 193210 258854
rect 193446 258618 223930 258854
rect 224166 258618 254650 258854
rect 254886 258618 285370 258854
rect 285606 258618 316090 258854
rect 316326 258618 346810 258854
rect 347046 258618 377530 258854
rect 377766 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 479610 258854
rect 479846 258618 510330 258854
rect 510566 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 24250 255454
rect 24486 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 54970 255454
rect 55206 255218 85690 255454
rect 85926 255218 116410 255454
rect 116646 255218 147130 255454
rect 147366 255218 177850 255454
rect 178086 255218 208570 255454
rect 208806 255218 239290 255454
rect 239526 255218 270010 255454
rect 270246 255218 300730 255454
rect 300966 255218 331450 255454
rect 331686 255218 362170 255454
rect 362406 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 464250 255454
rect 464486 255218 494970 255454
rect 495206 255218 525690 255454
rect 525926 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 24250 255134
rect 24486 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 54970 255134
rect 55206 254898 85690 255134
rect 85926 254898 116410 255134
rect 116646 254898 147130 255134
rect 147366 254898 177850 255134
rect 178086 254898 208570 255134
rect 208806 254898 239290 255134
rect 239526 254898 270010 255134
rect 270246 254898 300730 255134
rect 300966 254898 331450 255134
rect 331686 254898 362170 255134
rect 362406 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 464250 255134
rect 464486 254898 494970 255134
rect 495206 254898 525690 255134
rect 525926 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 39610 223174
rect 39846 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 70330 223174
rect 70566 222938 101050 223174
rect 101286 222938 131770 223174
rect 132006 222938 162490 223174
rect 162726 222938 193210 223174
rect 193446 222938 223930 223174
rect 224166 222938 254650 223174
rect 254886 222938 285370 223174
rect 285606 222938 316090 223174
rect 316326 222938 346810 223174
rect 347046 222938 377530 223174
rect 377766 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 479610 223174
rect 479846 222938 510330 223174
rect 510566 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 39610 222854
rect 39846 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 70330 222854
rect 70566 222618 101050 222854
rect 101286 222618 131770 222854
rect 132006 222618 162490 222854
rect 162726 222618 193210 222854
rect 193446 222618 223930 222854
rect 224166 222618 254650 222854
rect 254886 222618 285370 222854
rect 285606 222618 316090 222854
rect 316326 222618 346810 222854
rect 347046 222618 377530 222854
rect 377766 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 479610 222854
rect 479846 222618 510330 222854
rect 510566 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 24250 219454
rect 24486 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 54970 219454
rect 55206 219218 85690 219454
rect 85926 219218 116410 219454
rect 116646 219218 147130 219454
rect 147366 219218 177850 219454
rect 178086 219218 208570 219454
rect 208806 219218 239290 219454
rect 239526 219218 270010 219454
rect 270246 219218 300730 219454
rect 300966 219218 331450 219454
rect 331686 219218 362170 219454
rect 362406 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 464250 219454
rect 464486 219218 494970 219454
rect 495206 219218 525690 219454
rect 525926 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 24250 219134
rect 24486 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 54970 219134
rect 55206 218898 85690 219134
rect 85926 218898 116410 219134
rect 116646 218898 147130 219134
rect 147366 218898 177850 219134
rect 178086 218898 208570 219134
rect 208806 218898 239290 219134
rect 239526 218898 270010 219134
rect 270246 218898 300730 219134
rect 300966 218898 331450 219134
rect 331686 218898 362170 219134
rect 362406 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 464250 219134
rect 464486 218898 494970 219134
rect 495206 218898 525690 219134
rect 525926 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 39610 187174
rect 39846 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 70330 187174
rect 70566 186938 101050 187174
rect 101286 186938 131770 187174
rect 132006 186938 162490 187174
rect 162726 186938 193210 187174
rect 193446 186938 223930 187174
rect 224166 186938 254650 187174
rect 254886 186938 285370 187174
rect 285606 186938 316090 187174
rect 316326 186938 346810 187174
rect 347046 186938 377530 187174
rect 377766 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 39610 186854
rect 39846 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 70330 186854
rect 70566 186618 101050 186854
rect 101286 186618 131770 186854
rect 132006 186618 162490 186854
rect 162726 186618 193210 186854
rect 193446 186618 223930 186854
rect 224166 186618 254650 186854
rect 254886 186618 285370 186854
rect 285606 186618 316090 186854
rect 316326 186618 346810 186854
rect 347046 186618 377530 186854
rect 377766 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 24250 183454
rect 24486 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 54970 183454
rect 55206 183218 85690 183454
rect 85926 183218 116410 183454
rect 116646 183218 147130 183454
rect 147366 183218 177850 183454
rect 178086 183218 208570 183454
rect 208806 183218 239290 183454
rect 239526 183218 270010 183454
rect 270246 183218 300730 183454
rect 300966 183218 331450 183454
rect 331686 183218 362170 183454
rect 362406 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 24250 183134
rect 24486 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 54970 183134
rect 55206 182898 85690 183134
rect 85926 182898 116410 183134
rect 116646 182898 147130 183134
rect 147366 182898 177850 183134
rect 178086 182898 208570 183134
rect 208806 182898 239290 183134
rect 239526 182898 270010 183134
rect 270246 182898 300730 183134
rect 300966 182898 331450 183134
rect 331686 182898 362170 183134
rect 362406 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 39610 151174
rect 39846 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 70330 151174
rect 70566 150938 101050 151174
rect 101286 150938 131770 151174
rect 132006 150938 162490 151174
rect 162726 150938 193210 151174
rect 193446 150938 223930 151174
rect 224166 150938 254650 151174
rect 254886 150938 285370 151174
rect 285606 150938 316090 151174
rect 316326 150938 346810 151174
rect 347046 150938 377530 151174
rect 377766 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 429610 151174
rect 429846 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 39610 150854
rect 39846 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 70330 150854
rect 70566 150618 101050 150854
rect 101286 150618 131770 150854
rect 132006 150618 162490 150854
rect 162726 150618 193210 150854
rect 193446 150618 223930 150854
rect 224166 150618 254650 150854
rect 254886 150618 285370 150854
rect 285606 150618 316090 150854
rect 316326 150618 346810 150854
rect 347046 150618 377530 150854
rect 377766 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 429610 150854
rect 429846 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 24250 147454
rect 24486 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 54970 147454
rect 55206 147218 85690 147454
rect 85926 147218 116410 147454
rect 116646 147218 147130 147454
rect 147366 147218 177850 147454
rect 178086 147218 208570 147454
rect 208806 147218 239290 147454
rect 239526 147218 270010 147454
rect 270246 147218 300730 147454
rect 300966 147218 331450 147454
rect 331686 147218 362170 147454
rect 362406 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 414250 147454
rect 414486 147218 444970 147454
rect 445206 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 484250 147454
rect 484486 147218 514970 147454
rect 515206 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 545690 147454
rect 545926 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 24250 147134
rect 24486 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 54970 147134
rect 55206 146898 85690 147134
rect 85926 146898 116410 147134
rect 116646 146898 147130 147134
rect 147366 146898 177850 147134
rect 178086 146898 208570 147134
rect 208806 146898 239290 147134
rect 239526 146898 270010 147134
rect 270246 146898 300730 147134
rect 300966 146898 331450 147134
rect 331686 146898 362170 147134
rect 362406 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 414250 147134
rect 414486 146898 444970 147134
rect 445206 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 484250 147134
rect 484486 146898 514970 147134
rect 515206 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 545690 147134
rect 545926 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 39610 115174
rect 39846 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 70330 115174
rect 70566 114938 101050 115174
rect 101286 114938 131770 115174
rect 132006 114938 162490 115174
rect 162726 114938 193210 115174
rect 193446 114938 223930 115174
rect 224166 114938 254650 115174
rect 254886 114938 285370 115174
rect 285606 114938 316090 115174
rect 316326 114938 346810 115174
rect 347046 114938 377530 115174
rect 377766 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 499610 115174
rect 499846 114938 530330 115174
rect 530566 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 39610 114854
rect 39846 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 70330 114854
rect 70566 114618 101050 114854
rect 101286 114618 131770 114854
rect 132006 114618 162490 114854
rect 162726 114618 193210 114854
rect 193446 114618 223930 114854
rect 224166 114618 254650 114854
rect 254886 114618 285370 114854
rect 285606 114618 316090 114854
rect 316326 114618 346810 114854
rect 347046 114618 377530 114854
rect 377766 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 499610 114854
rect 499846 114618 530330 114854
rect 530566 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 24250 111454
rect 24486 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 54970 111454
rect 55206 111218 85690 111454
rect 85926 111218 116410 111454
rect 116646 111218 147130 111454
rect 147366 111218 177850 111454
rect 178086 111218 208570 111454
rect 208806 111218 239290 111454
rect 239526 111218 270010 111454
rect 270246 111218 300730 111454
rect 300966 111218 331450 111454
rect 331686 111218 362170 111454
rect 362406 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 484250 111454
rect 484486 111218 514970 111454
rect 515206 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 545690 111454
rect 545926 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 24250 111134
rect 24486 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 54970 111134
rect 55206 110898 85690 111134
rect 85926 110898 116410 111134
rect 116646 110898 147130 111134
rect 147366 110898 177850 111134
rect 178086 110898 208570 111134
rect 208806 110898 239290 111134
rect 239526 110898 270010 111134
rect 270246 110898 300730 111134
rect 300966 110898 331450 111134
rect 331686 110898 362170 111134
rect 362406 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 484250 111134
rect 484486 110898 514970 111134
rect 515206 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 545690 111134
rect 545926 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 39610 79174
rect 39846 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 70330 79174
rect 70566 78938 101050 79174
rect 101286 78938 131770 79174
rect 132006 78938 162490 79174
rect 162726 78938 193210 79174
rect 193446 78938 223930 79174
rect 224166 78938 254650 79174
rect 254886 78938 285370 79174
rect 285606 78938 316090 79174
rect 316326 78938 346810 79174
rect 347046 78938 377530 79174
rect 377766 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 39610 78854
rect 39846 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 70330 78854
rect 70566 78618 101050 78854
rect 101286 78618 131770 78854
rect 132006 78618 162490 78854
rect 162726 78618 193210 78854
rect 193446 78618 223930 78854
rect 224166 78618 254650 78854
rect 254886 78618 285370 78854
rect 285606 78618 316090 78854
rect 316326 78618 346810 78854
rect 347046 78618 377530 78854
rect 377766 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 24250 75454
rect 24486 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 54970 75454
rect 55206 75218 85690 75454
rect 85926 75218 116410 75454
rect 116646 75218 147130 75454
rect 147366 75218 177850 75454
rect 178086 75218 208570 75454
rect 208806 75218 239290 75454
rect 239526 75218 270010 75454
rect 270246 75218 300730 75454
rect 300966 75218 331450 75454
rect 331686 75218 362170 75454
rect 362406 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 24250 75134
rect 24486 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 54970 75134
rect 55206 74898 85690 75134
rect 85926 74898 116410 75134
rect 116646 74898 147130 75134
rect 147366 74898 177850 75134
rect 178086 74898 208570 75134
rect 208806 74898 239290 75134
rect 239526 74898 270010 75134
rect 270246 74898 300730 75134
rect 300966 74898 331450 75134
rect 331686 74898 362170 75134
rect 362406 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54235 589182 54334
rect 521262 54098 556706 54235
rect -8726 54014 556706 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53999 556706 54014
rect 556942 53999 557026 54235
rect 557262 54098 589182 54235
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect 557262 54014 592650 54098
rect 557262 53999 589182 54014
rect 521262 53778 589182 53999
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546414 43174
rect 546650 42938 551842 43174
rect 552078 42938 557270 43174
rect 557506 42938 562698 43174
rect 562934 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546414 42854
rect 546650 42618 551842 42854
rect 552078 42618 557270 42854
rect 557506 42618 562698 42854
rect 562934 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 543700 39454
rect 543936 39218 549128 39454
rect 549364 39218 554556 39454
rect 554792 39218 559984 39454
rect 560220 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 543700 39134
rect 543936 38898 549128 39134
rect 549364 38898 554556 39134
rect 554792 38898 559984 39134
rect 560220 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use posit_unit  posit_unit
timestamp 0
transform 1 0 460000 0 1 200000
box 0 2128 70000 67504
use multiplexer  proj_multiplexer
timestamp 0
transform 1 0 450000 0 1 320000
box 0 0 60000 60000
use tholin_avalonsemi_5401  tholin_avalonsemi_5401
timestamp 0
transform 1 0 520000 0 1 425000
box 842 0 40000 40000
use tholin_avalonsemi_tbb1143  tholin_avalonsemi_tbb1143
timestamp 0
transform 1 0 400000 0 1 305000
box 1066 1935 32000 32000
use tt2_tholin_diceroll  tt2_tholin_diceroll
timestamp 0
transform 1 0 470000 0 1 432000
box 1066 0 22976 24000
use tt2_tholin_multiplexed_counter  tt2_tholin_multiplexed_counter
timestamp 0
transform 1 0 550000 0 1 360000
box 842 0 19122 20000
use tt2_tholin_multiplier  tt2_tholin_multiplier
timestamp 0
transform 1 0 450000 0 1 500000
box 0 0 11118 16584
use tt2_tholin_namebadge  tt2_tholin_namebadge
timestamp 0
transform 1 0 420000 0 1 420000
box 1066 0 23987 25000
use tune_player  tune_player
timestamp 0
transform 1 0 540000 0 1 30000
box 0 2128 22976 21808
use wrapped_6502  wrapped_6502
timestamp 0
transform 1 0 410000 0 1 120000
box 1066 2128 45000 45000
use wrapped_MC14500  wrapped_MC14500
timestamp 0
transform 1 0 480000 0 1 500000
box 566 0 12000 18000
use wrapped_as1802  wrapped_as1802
timestamp 0
transform 1 0 480000 0 1 80000
box 1066 1776 70000 70000
use wrapped_as2650  wrapped_as2650
timestamp 0
transform 1 0 460000 0 1 600000
box 0 0 83812 78600
use wrapped_as512512512  wrapped_as512512512
timestamp 0
transform 1 0 20000 0 1 50000
box 1066 2128 360000 617488
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 58855 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 667017 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 58855 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 667017 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 58855 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 667017 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 58855 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 667017 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 58855 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 667017 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 58855 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 667017 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 58855 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 667017 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 58855 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 667017 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 50068 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 669548 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 135791 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 163505 434414 422599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 442833 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 379772 470414 608991 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 665809 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 87495 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 147033 506414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 259417 506414 608991 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 665809 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 58855 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 667017 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 58855 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 667017 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 58855 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 667017 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 58855 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 667017 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 58855 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 667017 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 58855 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 667017 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 58855 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 667017 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 58855 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 667017 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 58855 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 667017 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 135791 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 163505 441854 422599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 442833 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 259417 477854 320287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 378737 477854 608991 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 665809 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 87495 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 147033 513854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 259417 513854 608991 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 665809 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 30068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 53868 549854 445551 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 458849 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 58855 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 58855 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 58855 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 58855 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 58855 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 58855 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 58855 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 58855 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 135791 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 163505 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 259417 485294 320068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 517884 485294 608991 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 665809 485294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 87495 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 147033 521294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 259417 521294 608991 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 665809 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 30068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 53868 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 50068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 669548 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 58855 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 667017 96734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 58855 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 667017 132734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 58855 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 667017 168734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 58855 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 667017 204734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 58855 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 667017 240734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 58855 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 667017 276734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 58855 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 667017 312734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 58855 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 667017 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 135791 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 163505 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 500068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 517884 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 201919 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 259417 492734 320287 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 378737 492734 432068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 455868 492734 608991 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 665809 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 87495 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 259417 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 360068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 379516 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 58855 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 667017 93014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 58855 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 667017 129014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 58855 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 667017 165014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 58855 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 667017 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 58855 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 667017 237014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 58855 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 667017 273014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 58855 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 667017 309014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 58855 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 667017 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 135791 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 163505 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 517884 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 259417 489014 320287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 378737 489014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 517884 489014 608991 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 665809 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 87495 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 147033 525014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 259417 525014 425068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 464644 525014 608991 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 665809 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 58855 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 667017 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 58855 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 667017 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 58855 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 667017 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 58855 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 667017 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 58855 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 667017 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 58855 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 667017 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 50068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 669548 316454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 58855 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 667017 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 135791 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 163505 424454 420068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 444412 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 500068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 517884 460454 608991 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 665809 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 87495 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 259417 496454 320287 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 378737 496454 608991 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 665809 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 87495 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 147033 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 58855 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 667017 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 58855 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 667017 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 58855 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 667017 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 58855 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 667017 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 58855 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 667017 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 58855 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 667017 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 58855 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 667017 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 58855 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 667017 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 58855 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 667017 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 135791 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 163505 438134 420068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 444412 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 259417 474134 432068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 455868 474134 608991 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 665809 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 87495 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 147033 510134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 259417 510134 608991 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 665809 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 80068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 149564 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 58855 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 667017 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 58855 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 667017 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 58855 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 667017 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 50068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 669548 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 58855 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 667017 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 58855 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 667017 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 50068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 669548 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 58855 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 667017 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 58855 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 667017 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 120068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 164540 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 259417 481574 320287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 378737 481574 608991 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 665809 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 87495 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 147033 517574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 259417 517574 608991 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 665809 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 35319 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 43177 553574 360068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 379516 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 362288 651336 362288 651336 0 vccd1
rlabel via4 45704 658776 45704 658776 0 vccd2
rlabel via4 377144 666216 377144 666216 0 vdda1
rlabel via4 60584 637656 60584 637656 0 vdda2
rlabel via4 344864 669936 344864 669936 0 vssa1
rlabel via4 64304 641376 64304 641376 0 vssa2
rlabel via4 377648 655056 377648 655056 0 vssd1
rlabel via4 373424 50496 373424 50496 0 vssd2
rlabel metal2 422510 446036 422510 446036 0 design_clk
rlabel metal3 450708 501179 450708 501179 0 dsi_all\[0\]
rlabel metal1 444498 444414 444498 444414 0 dsi_all\[10\]
rlabel metal2 447166 174862 447166 174862 0 dsi_all\[11\]
rlabel metal2 447166 185946 447166 185946 0 dsi_all\[12\]
rlabel metal1 445464 331330 445464 331330 0 dsi_all\[13\]
rlabel metal2 447166 331517 447166 331517 0 dsi_all\[14\]
rlabel metal1 445648 331398 445648 331398 0 dsi_all\[15\]
rlabel metal3 448738 332860 448738 332860 0 dsi_all\[16\]
rlabel metal2 447166 333047 447166 333047 0 dsi_all\[17\]
rlabel metal2 447258 333285 447258 333285 0 dsi_all\[18\]
rlabel metal2 447166 334237 447166 334237 0 dsi_all\[19\]
rlabel metal2 450570 502095 450570 502095 0 dsi_all\[1\]
rlabel metal2 447258 334543 447258 334543 0 dsi_all\[20\]
rlabel metal3 448738 335580 448738 335580 0 dsi_all\[21\]
rlabel metal1 445556 335750 445556 335750 0 dsi_all\[22\]
rlabel metal1 444774 335818 444774 335818 0 dsi_all\[23\]
rlabel metal2 447166 337025 447166 337025 0 dsi_all\[24\]
rlabel metal2 447258 337263 447258 337263 0 dsi_all\[25\]
rlabel metal2 447166 338419 447166 338419 0 dsi_all\[26\]
rlabel metal3 450156 505531 450156 505531 0 dsi_all\[2\]
rlabel metal3 450340 507707 450340 507707 0 dsi_all\[3\]
rlabel metal2 541459 464916 541459 464916 0 dsi_all\[4\]
rlabel metal1 504942 153170 504942 153170 0 dsi_all\[5\]
rlabel metal2 450570 166668 450570 166668 0 dsi_all\[6\]
rlabel metal2 523671 600100 523671 600100 0 dsi_all\[7\]
rlabel metal2 447166 447576 447166 447576 0 dsi_all\[8\]
rlabel metal2 447902 447644 447902 447644 0 dsi_all\[9\]
rlabel metal2 488658 318274 488658 318274 0 dso_6502\[0\]
rlabel metal3 456128 137156 456128 137156 0 dso_6502\[10\]
rlabel metal3 456128 138652 456128 138652 0 dso_6502\[11\]
rlabel metal3 455898 140148 455898 140148 0 dso_6502\[12\]
rlabel metal3 456128 141644 456128 141644 0 dso_6502\[13\]
rlabel metal1 475502 268430 475502 268430 0 dso_6502\[14\]
rlabel metal3 455898 144636 455898 144636 0 dso_6502\[15\]
rlabel metal1 475272 276658 475272 276658 0 dso_6502\[16\]
rlabel metal1 475226 294474 475226 294474 0 dso_6502\[17\]
rlabel metal1 476284 269858 476284 269858 0 dso_6502\[18\]
rlabel metal1 476100 271218 476100 271218 0 dso_6502\[19\]
rlabel metal2 488888 318138 488888 318138 0 dso_6502\[1\]
rlabel metal3 456358 152116 456358 152116 0 dso_6502\[20\]
rlabel metal3 455898 153612 455898 153612 0 dso_6502\[21\]
rlabel metal3 455898 155108 455898 155108 0 dso_6502\[22\]
rlabel metal3 455898 156604 455898 156604 0 dso_6502\[23\]
rlabel metal3 456404 158100 456404 158100 0 dso_6502\[24\]
rlabel metal3 455898 159596 455898 159596 0 dso_6502\[25\]
rlabel metal3 455898 161092 455898 161092 0 dso_6502\[26\]
rlabel metal2 489072 318036 489072 318036 0 dso_6502\[2\]
rlabel metal1 489118 317934 489118 317934 0 dso_6502\[3\]
rlabel metal2 488934 295013 488934 295013 0 dso_6502\[4\]
rlabel metal3 474559 307020 474559 307020 0 dso_6502\[5\]
rlabel metal3 473869 272476 473869 272476 0 dso_6502\[6\]
rlabel metal3 456036 132668 456036 132668 0 dso_6502\[7\]
rlabel metal3 456266 134164 456266 134164 0 dso_6502\[8\]
rlabel metal3 456979 135660 456979 135660 0 dso_6502\[9\]
rlabel metal2 447350 347055 447350 347055 0 dso_LCD\[0\]
rlabel metal2 447258 347361 447258 347361 0 dso_LCD\[1\]
rlabel metal2 423568 354076 423568 354076 0 dso_LCD\[2\]
rlabel metal2 423430 354212 423430 354212 0 dso_LCD\[3\]
rlabel metal1 445464 349010 445464 349010 0 dso_LCD\[4\]
rlabel metal2 447350 349843 447350 349843 0 dso_LCD\[5\]
rlabel metal2 447258 350047 447258 350047 0 dso_LCD\[6\]
rlabel metal2 447166 350353 447166 350353 0 dso_LCD\[7\]
rlabel metal3 550290 81804 550290 81804 0 dso_as1802\[0\]
rlabel metal3 550336 106284 550336 106284 0 dso_as1802\[10\]
rlabel metal1 525136 268362 525136 268362 0 dso_as1802\[11\]
rlabel metal3 550382 111180 550382 111180 0 dso_as1802\[12\]
rlabel metal3 550428 113628 550428 113628 0 dso_as1802\[13\]
rlabel metal3 550474 116076 550474 116076 0 dso_as1802\[14\]
rlabel metal3 550612 118524 550612 118524 0 dso_as1802\[15\]
rlabel metal3 550658 120972 550658 120972 0 dso_as1802\[16\]
rlabel metal3 550566 123420 550566 123420 0 dso_as1802\[17\]
rlabel metal1 527390 309842 527390 309842 0 dso_as1802\[18\]
rlabel metal1 527206 308550 527206 308550 0 dso_as1802\[19\]
rlabel metal1 522974 307122 522974 307122 0 dso_as1802\[1\]
rlabel metal1 526010 269994 526010 269994 0 dso_as1802\[20\]
rlabel metal3 551210 133212 551210 133212 0 dso_as1802\[21\]
rlabel via2 549861 136204 549861 136204 0 dso_as1802\[22\]
rlabel via2 549539 138652 549539 138652 0 dso_as1802\[23\]
rlabel metal3 551256 140556 551256 140556 0 dso_as1802\[24\]
rlabel metal1 550344 149430 550344 149430 0 dso_as1802\[25\]
rlabel metal4 547676 229092 547676 229092 0 dso_as1802\[26\]
rlabel metal1 524400 271150 524400 271150 0 dso_as1802\[2\]
rlabel metal1 524998 271218 524998 271218 0 dso_as1802\[3\]
rlabel metal3 551302 91596 551302 91596 0 dso_as1802\[4\]
rlabel metal3 551164 94044 551164 94044 0 dso_as1802\[5\]
rlabel via2 549355 96764 549355 96764 0 dso_as1802\[6\]
rlabel via2 549493 99348 549493 99348 0 dso_as1802\[7\]
rlabel metal2 543030 233954 543030 233954 0 dso_as1802\[8\]
rlabel metal1 524538 272578 524538 272578 0 dso_as1802\[9\]
rlabel metal2 461610 503540 461610 503540 0 dso_as2650\[0\]
rlabel metal2 487002 381640 487002 381640 0 dso_as2650\[10\]
rlabel metal2 464370 491368 464370 491368 0 dso_as2650\[11\]
rlabel metal2 489387 379916 489387 379916 0 dso_as2650\[12\]
rlabel metal3 459778 638588 459778 638588 0 dso_as2650\[13\]
rlabel metal3 459456 641444 459456 641444 0 dso_as2650\[14\]
rlabel metal3 460276 644013 460276 644013 0 dso_as2650\[15\]
rlabel metal3 459502 647156 459502 647156 0 dso_as2650\[16\]
rlabel metal1 477894 598230 477894 598230 0 dso_as2650\[17\]
rlabel metal1 477940 596802 477940 596802 0 dso_as2650\[18\]
rlabel metal3 460460 655807 460460 655807 0 dso_as2650\[19\]
rlabel metal3 459732 604316 459732 604316 0 dso_as2650\[1\]
rlabel metal2 499737 379916 499737 379916 0 dso_as2650\[20\]
rlabel metal2 501071 379916 501071 379916 0 dso_as2650\[21\]
rlabel metal2 502405 379916 502405 379916 0 dso_as2650\[22\]
rlabel metal2 503746 489760 503746 489760 0 dso_as2650\[23\]
rlabel metal2 504843 379916 504843 379916 0 dso_as2650\[24\]
rlabel metal2 506322 381470 506322 381470 0 dso_as2650\[25\]
rlabel metal2 507419 379916 507419 379916 0 dso_as2650\[26\]
rlabel metal2 462990 491844 462990 491844 0 dso_as2650\[2\]
rlabel metal2 468510 491028 468510 491028 0 dso_as2650\[3\]
rlabel metal2 467130 491606 467130 491606 0 dso_as2650\[4\]
rlabel metal2 463082 491674 463082 491674 0 dso_as2650\[5\]
rlabel metal2 469890 450840 469890 450840 0 dso_as2650\[6\]
rlabel metal2 467222 490042 467222 490042 0 dso_as2650\[7\]
rlabel metal2 467314 452676 467314 452676 0 dso_as2650\[8\]
rlabel metal2 468602 489396 468602 489396 0 dso_as2650\[9\]
rlabel metal2 443946 362542 443946 362542 0 dso_as512512512\[0\]
rlabel metal2 447258 366503 447258 366503 0 dso_as512512512\[10\]
rlabel metal2 447166 366809 447166 366809 0 dso_as512512512\[11\]
rlabel metal2 447350 367727 447350 367727 0 dso_as512512512\[12\]
rlabel metal2 447258 368033 447258 368033 0 dso_as512512512\[13\]
rlabel metal2 447166 368339 447166 368339 0 dso_as512512512\[14\]
rlabel metal2 447258 369291 447258 369291 0 dso_as512512512\[15\]
rlabel metal2 447166 369529 447166 369529 0 dso_as512512512\[16\]
rlabel metal2 447350 370515 447350 370515 0 dso_as512512512\[17\]
rlabel metal2 447258 370753 447258 370753 0 dso_as512512512\[18\]
rlabel metal2 447166 370991 447166 370991 0 dso_as512512512\[19\]
rlabel metal2 447166 361335 447166 361335 0 dso_as512512512\[1\]
rlabel metal2 447258 371943 447258 371943 0 dso_as512512512\[20\]
rlabel metal2 447350 372283 447350 372283 0 dso_as512512512\[21\]
rlabel metal2 447166 372521 447166 372521 0 dso_as512512512\[22\]
rlabel metal2 447258 373541 447258 373541 0 dso_as512512512\[23\]
rlabel metal2 447166 373779 447166 373779 0 dso_as512512512\[24\]
rlabel metal2 447350 374765 447350 374765 0 dso_as512512512\[25\]
rlabel metal2 447258 374969 447258 374969 0 dso_as512512512\[26\]
rlabel via2 447166 375275 447166 375275 0 dso_as512512512\[27\]
rlabel metal1 445556 362746 445556 362746 0 dso_as512512512\[2\]
rlabel metal2 447258 362525 447258 362525 0 dso_as512512512\[3\]
rlabel metal2 447166 362831 447166 362831 0 dso_as512512512\[4\]
rlabel metal2 447258 363817 447258 363817 0 dso_as512512512\[5\]
rlabel metal2 447166 364055 447166 364055 0 dso_as512512512\[6\]
rlabel metal2 447350 365041 447350 365041 0 dso_as512512512\[7\]
rlabel metal2 447258 365279 447258 365279 0 dso_as512512512\[8\]
rlabel via2 447166 365517 447166 365517 0 dso_as512512512\[9\]
rlabel metal2 520858 423480 520858 423480 0 dso_as5401\[0\]
rlabel metal3 511236 371756 511236 371756 0 dso_as5401\[10\]
rlabel metal3 511374 372164 511374 372164 0 dso_as5401\[11\]
rlabel metal2 538377 425068 538377 425068 0 dso_as5401\[12\]
rlabel metal2 539803 425068 539803 425068 0 dso_as5401\[13\]
rlabel metal2 541466 422630 541466 422630 0 dso_as5401\[14\]
rlabel metal2 542747 425068 542747 425068 0 dso_as5401\[15\]
rlabel metal2 544410 424160 544410 424160 0 dso_as5401\[16\]
rlabel metal2 545882 424228 545882 424228 0 dso_as5401\[17\]
rlabel metal2 547354 424194 547354 424194 0 dso_as5401\[18\]
rlabel metal1 531806 385662 531806 385662 0 dso_as5401\[19\]
rlabel metal2 522139 425068 522139 425068 0 dso_as5401\[1\]
rlabel metal2 538890 399840 538890 399840 0 dso_as5401\[20\]
rlabel metal2 540270 399908 540270 399908 0 dso_as5401\[21\]
rlabel metal2 544410 394551 544410 394551 0 dso_as5401\[22\]
rlabel metal2 547170 399840 547170 399840 0 dso_as5401\[23\]
rlabel metal2 556186 424058 556186 424058 0 dso_as5401\[24\]
rlabel metal2 557658 424024 557658 424024 0 dso_as5401\[25\]
rlabel metal2 559130 423990 559130 423990 0 dso_as5401\[26\]
rlabel metal2 523611 425068 523611 425068 0 dso_as5401\[2\]
rlabel metal1 522468 422382 522468 422382 0 dso_as5401\[3\]
rlabel metal2 526555 425068 526555 425068 0 dso_as5401\[4\]
rlabel metal2 528218 424092 528218 424092 0 dso_as5401\[5\]
rlabel metal2 522422 396916 522422 396916 0 dso_as5401\[6\]
rlabel metal3 511604 370532 511604 370532 0 dso_as5401\[7\]
rlabel metal2 523710 397154 523710 397154 0 dso_as5401\[8\]
rlabel metal3 511604 371348 511604 371348 0 dso_as5401\[9\]
rlabel metal3 511328 362780 511328 362780 0 dso_counter\[0\]
rlabel metal3 511512 366860 511512 366860 0 dso_counter\[10\]
rlabel metal2 547170 363562 547170 363562 0 dso_counter\[11\]
rlabel metal3 511512 363188 511512 363188 0 dso_counter\[1\]
rlabel metal3 511650 363596 511650 363596 0 dso_counter\[2\]
rlabel metal3 511052 364004 511052 364004 0 dso_counter\[3\]
rlabel metal3 511650 364412 511650 364412 0 dso_counter\[4\]
rlabel metal2 559130 359390 559130 359390 0 dso_counter\[5\]
rlabel metal2 560786 359288 560786 359288 0 dso_counter\[6\]
rlabel metal2 562442 359322 562442 359322 0 dso_counter\[7\]
rlabel metal2 564098 359220 564098 359220 0 dso_counter\[8\]
rlabel metal2 518926 362372 518926 362372 0 dso_counter\[9\]
rlabel metal2 462767 379916 462767 379916 0 dso_diceroll\[0\]
rlabel metal2 464055 379916 464055 379916 0 dso_diceroll\[1\]
rlabel metal2 465343 379916 465343 379916 0 dso_diceroll\[2\]
rlabel metal2 466394 404896 466394 404896 0 dso_diceroll\[3\]
rlabel metal2 467682 382116 467682 382116 0 dso_diceroll\[4\]
rlabel metal1 485760 429182 485760 429182 0 dso_diceroll\[5\]
rlabel metal2 470258 382150 470258 382150 0 dso_diceroll\[6\]
rlabel metal1 481252 387090 481252 387090 0 dso_diceroll\[7\]
rlabel metal3 449796 350812 449796 350812 0 dso_mc14500\[0\]
rlabel metal3 449934 351356 449934 351356 0 dso_mc14500\[1\]
rlabel metal3 449842 351900 449842 351900 0 dso_mc14500\[2\]
rlabel metal3 449750 352444 449750 352444 0 dso_mc14500\[3\]
rlabel metal3 449014 352988 449014 352988 0 dso_mc14500\[4\]
rlabel metal3 448784 353532 448784 353532 0 dso_mc14500\[5\]
rlabel metal3 449612 354076 449612 354076 0 dso_mc14500\[6\]
rlabel metal3 449888 354620 449888 354620 0 dso_mc14500\[7\]
rlabel metal3 449244 355164 449244 355164 0 dso_mc14500\[8\]
rlabel metal2 450991 500140 450991 500140 0 dso_multiplier\[0\]
rlabel metal2 452417 500140 452417 500140 0 dso_multiplier\[1\]
rlabel metal2 454611 379916 454611 379916 0 dso_multiplier\[2\]
rlabel metal2 455269 500140 455269 500140 0 dso_multiplier\[3\]
rlabel metal2 457187 379916 457187 379916 0 dso_multiplier\[4\]
rlabel metal2 458475 379916 458475 379916 0 dso_multiplier\[5\]
rlabel metal2 459915 500140 459915 500140 0 dso_multiplier\[6\]
rlabel metal2 461249 500140 461249 500140 0 dso_multiplier\[7\]
rlabel metal2 488198 311605 488198 311605 0 dso_posit\[0\]
rlabel metal1 488014 318070 488014 318070 0 dso_posit\[1\]
rlabel metal1 488198 318002 488198 318002 0 dso_posit\[2\]
rlabel metal2 488244 318036 488244 318036 0 dso_posit\[3\]
rlabel metal2 447166 356201 447166 356201 0 dso_tbb1143\[0\]
rlabel metal1 445556 356218 445556 356218 0 dso_tbb1143\[1\]
rlabel metal2 447258 356711 447258 356711 0 dso_tbb1143\[2\]
rlabel metal2 447166 357663 447166 357663 0 dso_tbb1143\[3\]
rlabel metal2 447258 357969 447258 357969 0 dso_tbb1143\[4\]
rlabel metal1 445694 358938 445694 358938 0 dso_tbb1143\[5\]
rlabel metal2 447166 359193 447166 359193 0 dso_tbb1143\[6\]
rlabel metal2 447258 359431 447258 359431 0 dso_tbb1143\[7\]
rlabel metal3 540684 50131 540684 50131 0 dso_tune
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel metal2 580198 457453 580198 457453 0 io_in[10]
rlabel metal2 519570 413916 519570 413916 0 io_in[11]
rlabel metal2 580198 563703 580198 563703 0 io_in[12]
rlabel metal2 580198 617185 580198 617185 0 io_in[13]
rlabel via2 580198 670701 580198 670701 0 io_in[14]
rlabel metal3 559291 699788 559291 699788 0 io_in[15]
rlabel metal2 444222 509524 444222 509524 0 io_in[16]
rlabel metal2 429870 574304 429870 574304 0 io_in[17]
rlabel metal2 365010 702110 365010 702110 0 io_in[18]
rlabel metal3 374049 700604 374049 700604 0 io_in[19]
rlabel metal2 580198 46597 580198 46597 0 io_in[1]
rlabel metal2 235198 702008 235198 702008 0 io_in[20]
rlabel metal1 309764 700366 309764 700366 0 io_in[21]
rlabel metal4 444268 510068 444268 510068 0 io_in[22]
rlabel metal2 40526 701957 40526 701957 0 io_in[23]
rlabel metal3 1878 684284 1878 684284 0 io_in[24]
rlabel metal3 2016 632060 2016 632060 0 io_in[25]
rlabel metal3 1970 579972 1970 579972 0 io_in[26]
rlabel metal3 1924 527884 1924 527884 0 io_in[27]
rlabel metal1 4508 565862 4508 565862 0 io_in[28]
rlabel metal3 1924 423572 1924 423572 0 io_in[29]
rlabel metal2 580198 86547 580198 86547 0 io_in[2]
rlabel metal1 5980 115906 5980 115906 0 io_in[30]
rlabel metal1 5750 140114 5750 140114 0 io_in[31]
rlabel metal2 445786 272204 445786 272204 0 io_in[32]
rlabel metal1 4324 102170 4324 102170 0 io_in[33]
rlabel metal1 4646 89726 4646 89726 0 io_in[34]
rlabel metal3 1924 110636 1924 110636 0 io_in[35]
rlabel metal3 1878 71604 1878 71604 0 io_in[36]
rlabel metal3 1924 32436 1924 32436 0 io_in[37]
rlabel metal2 558210 219028 558210 219028 0 io_in[3]
rlabel metal2 580198 166413 580198 166413 0 io_in[4]
rlabel metal2 579830 206329 579830 206329 0 io_in[5]
rlabel via2 580198 245565 580198 245565 0 io_in[6]
rlabel metal2 580198 299081 580198 299081 0 io_in[7]
rlabel metal3 582138 351900 582138 351900 0 io_in[8]
rlabel metal3 582000 404940 582000 404940 0 io_in[9]
rlabel via2 580198 33099 580198 33099 0 io_oeb[0]
rlabel metal3 582046 484636 582046 484636 0 io_oeb[10]
rlabel metal2 580198 537319 580198 537319 0 io_oeb[11]
rlabel metal2 522330 365194 522330 365194 0 io_oeb[12]
rlabel metal3 581954 644028 581954 644028 0 io_oeb[13]
rlabel metal3 581908 697204 581908 697204 0 io_oeb[14]
rlabel metal1 488566 317968 488566 317968 0 io_oeb[15]
rlabel metal2 462346 691604 462346 691604 0 io_oeb[16]
rlabel metal1 480976 317934 480976 317934 0 io_oeb[17]
rlabel metal2 332534 702076 332534 702076 0 io_oeb[18]
rlabel metal2 445326 493272 445326 493272 0 io_oeb[19]
rlabel metal2 559590 186558 559590 186558 0 io_oeb[1]
rlabel metal2 482402 319253 482402 319253 0 io_oeb[20]
rlabel metal2 137862 701940 137862 701940 0 io_oeb[21]
rlabel metal2 442382 326808 442382 326808 0 io_oeb[22]
rlabel metal2 445418 493612 445418 493612 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal3 2062 606084 2062 606084 0 io_oeb[25]
rlabel metal2 4094 622404 4094 622404 0 io_oeb[26]
rlabel metal3 1878 501772 1878 501772 0 io_oeb[27]
rlabel metal3 2062 449548 2062 449548 0 io_oeb[28]
rlabel metal1 4370 253946 4370 253946 0 io_oeb[29]
rlabel metal2 562350 211446 562350 211446 0 io_oeb[2]
rlabel metal3 2016 345372 2016 345372 0 io_oeb[30]
rlabel metal3 1970 293148 1970 293148 0 io_oeb[31]
rlabel metal1 5566 83198 5566 83198 0 io_oeb[32]
rlabel metal1 4600 115906 4600 115906 0 io_oeb[33]
rlabel metal3 2016 136748 2016 136748 0 io_oeb[34]
rlabel metal3 1832 84660 1832 84660 0 io_oeb[35]
rlabel metal3 1878 45492 1878 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 580198 152915 580198 152915 0 io_oeb[3]
rlabel metal2 580198 192831 580198 192831 0 io_oeb[4]
rlabel metal2 580198 232781 580198 232781 0 io_oeb[5]
rlabel metal3 581954 272204 581954 272204 0 io_oeb[6]
rlabel metal2 481482 319124 481482 319124 0 io_oeb[7]
rlabel metal2 485070 319532 485070 319532 0 io_oeb[8]
rlabel metal3 581908 431596 581908 431596 0 io_oeb[9]
rlabel metal2 580014 20213 580014 20213 0 io_out[0]
rlabel metal2 580014 471019 580014 471019 0 io_out[10]
rlabel metal3 581954 524484 581954 524484 0 io_out[11]
rlabel metal2 579646 577269 579646 577269 0 io_out[12]
rlabel metal1 579002 630666 579002 630666 0 io_out[13]
rlabel metal2 579646 683519 579646 683519 0 io_out[14]
rlabel metal3 543099 699788 543099 699788 0 io_out[15]
rlabel metal2 444314 509184 444314 509184 0 io_out[16]
rlabel metal2 413678 521876 413678 521876 0 io_out[17]
rlabel metal2 348818 686912 348818 686912 0 io_out[18]
rlabel metal2 445234 494054 445234 494054 0 io_out[19]
rlabel metal2 580198 60163 580198 60163 0 io_out[1]
rlabel metal2 219006 702042 219006 702042 0 io_out[20]
rlabel metal2 154146 686844 154146 686844 0 io_out[21]
rlabel metal2 89194 686810 89194 686810 0 io_out[22]
rlabel metal2 24334 686113 24334 686113 0 io_out[23]
rlabel metal3 1924 671228 1924 671228 0 io_out[24]
rlabel metal3 1740 619140 1740 619140 0 io_out[25]
rlabel metal3 2062 566916 2062 566916 0 io_out[26]
rlabel metal2 385066 467806 385066 467806 0 io_out[27]
rlabel metal3 1970 462604 1970 462604 0 io_out[28]
rlabel metal3 2016 410516 2016 410516 0 io_out[29]
rlabel metal2 580198 100079 580198 100079 0 io_out[2]
rlabel metal1 388562 80070 388562 80070 0 io_out[30]
rlabel metal1 4462 212466 4462 212466 0 io_out[31]
rlabel metal3 2016 254116 2016 254116 0 io_out[32]
rlabel metal1 4462 101558 4462 101558 0 io_out[33]
rlabel metal2 424166 255952 424166 255952 0 io_out[34]
rlabel metal3 1878 97580 1878 97580 0 io_out[35]
rlabel metal3 1970 58548 1970 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel via2 580198 139349 580198 139349 0 io_out[3]
rlabel metal2 580198 179265 580198 179265 0 io_out[4]
rlabel metal3 581908 219028 581908 219028 0 io_out[5]
rlabel metal3 581954 258876 581954 258876 0 io_out[6]
rlabel metal2 580198 312647 580198 312647 0 io_out[7]
rlabel metal2 580198 364735 580198 364735 0 io_out[8]
rlabel metal3 582092 418268 582092 418268 0 io_out[9]
rlabel metal1 487830 318206 487830 318206 0 oeb_6502
rlabel metal3 548688 148580 548688 148580 0 oeb_as1802
rlabel metal3 459410 678572 459410 678572 0 oeb_as2650
rlabel metal2 403650 518840 403650 518840 0 oeb_as512512512
rlabel metal3 560778 444924 560778 444924 0 oeb_as5401
rlabel metal3 449704 355708 449704 355708 0 oeb_mc14500
rlabel metal3 449980 339932 449980 339932 0 rst_6502
rlabel metal2 427478 446070 427478 446070 0 rst_LCD
rlabel metal3 449106 341020 449106 341020 0 rst_as1802
rlabel metal2 540546 599158 540546 599158 0 rst_as2650
rlabel metal2 447166 343111 447166 343111 0 rst_as512512512
rlabel metal2 525090 465688 525090 465688 0 rst_as5401
rlabel metal3 449980 343196 449980 343196 0 rst_counter
rlabel metal3 449106 343740 449106 343740 0 rst_diceroll
rlabel metal3 449060 344284 449060 344284 0 rst_mc14500
rlabel metal3 449934 344828 449934 344828 0 rst_posit
rlabel metal2 447166 345219 447166 345219 0 rst_tbb1143
rlabel metal3 449244 345916 449244 345916 0 rst_tune
rlabel metal2 598 1843 598 1843 0 wb_clk_i
rlabel metal2 1702 1979 1702 1979 0 wb_rst_i
rlabel metal2 2898 25371 2898 25371 0 wbs_ack_o
rlabel metal2 406778 178228 406778 178228 0 wbs_adr_i[0]
rlabel metal2 403926 178245 403926 178245 0 wbs_adr_i[10]
rlabel metal2 403742 178279 403742 178279 0 wbs_adr_i[11]
rlabel metal2 403834 176868 403834 176868 0 wbs_adr_i[12]
rlabel metal2 58466 25388 58466 25388 0 wbs_adr_i[13]
rlabel metal2 62054 25422 62054 25422 0 wbs_adr_i[14]
rlabel metal2 65550 25456 65550 25456 0 wbs_adr_i[15]
rlabel metal2 69138 23994 69138 23994 0 wbs_adr_i[16]
rlabel metal2 72634 24028 72634 24028 0 wbs_adr_i[17]
rlabel metal2 76222 24062 76222 24062 0 wbs_adr_i[18]
rlabel metal2 79718 24096 79718 24096 0 wbs_adr_i[19]
rlabel metal2 12374 23960 12374 23960 0 wbs_adr_i[1]
rlabel metal2 83306 24130 83306 24130 0 wbs_adr_i[20]
rlabel metal3 511098 349316 511098 349316 0 wbs_adr_i[21]
rlabel metal3 511650 350540 511650 350540 0 wbs_adr_i[22]
rlabel metal2 93978 25286 93978 25286 0 wbs_adr_i[23]
rlabel metal2 97474 24232 97474 24232 0 wbs_adr_i[24]
rlabel metal2 101062 24300 101062 24300 0 wbs_adr_i[25]
rlabel metal2 104558 23926 104558 23926 0 wbs_adr_i[26]
rlabel metal2 407974 174556 407974 174556 0 wbs_adr_i[27]
rlabel metal2 410550 174590 410550 174590 0 wbs_adr_i[28]
rlabel metal2 115230 25252 115230 25252 0 wbs_adr_i[29]
rlabel metal2 17066 2030 17066 2030 0 wbs_adr_i[2]
rlabel metal2 118818 22838 118818 22838 0 wbs_adr_i[30]
rlabel metal2 122314 22872 122314 22872 0 wbs_adr_i[31]
rlabel metal2 21850 2064 21850 2064 0 wbs_adr_i[3]
rlabel metal2 392886 172465 392886 172465 0 wbs_adr_i[4]
rlabel metal2 392610 151198 392610 151198 0 wbs_adr_i[5]
rlabel metal2 393070 172567 393070 172567 0 wbs_adr_i[6]
rlabel metal2 37214 22668 37214 22668 0 wbs_adr_i[7]
rlabel metal2 40710 22702 40710 22702 0 wbs_adr_i[8]
rlabel metal2 44298 22736 44298 22736 0 wbs_adr_i[9]
rlabel metal2 4094 1911 4094 1911 0 wbs_cyc_i
rlabel metal2 389850 150535 389850 150535 0 wbs_dat_i[0]
rlabel metal2 390310 171530 390310 171530 0 wbs_dat_i[10]
rlabel metal2 390126 170068 390126 170068 0 wbs_dat_i[11]
rlabel metal2 56074 21274 56074 21274 0 wbs_dat_i[12]
rlabel metal2 59662 21308 59662 21308 0 wbs_dat_i[13]
rlabel metal2 63250 21342 63250 21342 0 wbs_dat_i[14]
rlabel metal2 387458 171768 387458 171768 0 wbs_dat_i[15]
rlabel metal2 387550 173978 387550 173978 0 wbs_dat_i[16]
rlabel metal2 387090 169898 387090 169898 0 wbs_dat_i[17]
rlabel metal2 77418 21410 77418 21410 0 wbs_dat_i[18]
rlabel metal2 80914 21444 80914 21444 0 wbs_dat_i[19]
rlabel metal2 384330 149175 384330 149175 0 wbs_dat_i[1]
rlabel metal2 384514 168708 384514 168708 0 wbs_dat_i[20]
rlabel metal2 384606 171530 384606 171530 0 wbs_dat_i[21]
rlabel metal2 384422 168878 384422 168878 0 wbs_dat_i[22]
rlabel metal2 95174 21172 95174 21172 0 wbs_dat_i[23]
rlabel metal2 98670 21512 98670 21512 0 wbs_dat_i[24]
rlabel metal2 102258 21138 102258 21138 0 wbs_dat_i[25]
rlabel metal2 391506 167229 391506 167229 0 wbs_dat_i[26]
rlabel metal1 245594 39270 245594 39270 0 wbs_dat_i[27]
rlabel metal2 520398 326332 520398 326332 0 wbs_dat_i[28]
rlabel metal2 116426 20152 116426 20152 0 wbs_dat_i[29]
rlabel metal2 18262 19846 18262 19846 0 wbs_dat_i[2]
rlabel metal2 119922 20118 119922 20118 0 wbs_dat_i[30]
rlabel metal1 260314 40018 260314 40018 0 wbs_dat_i[31]
rlabel metal2 23046 19880 23046 19880 0 wbs_dat_i[3]
rlabel metal1 205436 39474 205436 39474 0 wbs_dat_i[4]
rlabel metal2 385894 165665 385894 165665 0 wbs_dat_i[5]
rlabel metal2 385710 165716 385710 165716 0 wbs_dat_i[6]
rlabel metal2 38410 20016 38410 20016 0 wbs_dat_i[7]
rlabel metal2 41906 21206 41906 21206 0 wbs_dat_i[8]
rlabel metal2 45494 20050 45494 20050 0 wbs_dat_i[9]
rlabel metal2 388470 147900 388470 147900 0 wbs_dat_o[0]
rlabel metal2 388654 168708 388654 168708 0 wbs_dat_o[10]
rlabel metal2 391322 164322 391322 164322 0 wbs_dat_o[11]
rlabel metal2 57270 18520 57270 18520 0 wbs_dat_o[12]
rlabel metal2 60858 18452 60858 18452 0 wbs_dat_o[13]
rlabel metal2 64354 18554 64354 18554 0 wbs_dat_o[14]
rlabel metal2 67942 2234 67942 2234 0 wbs_dat_o[15]
rlabel metal2 521962 316438 521962 316438 0 wbs_dat_o[16]
rlabel metal2 75026 18622 75026 18622 0 wbs_dat_o[17]
rlabel metal2 78614 1860 78614 1860 0 wbs_dat_o[18]
rlabel metal2 82110 18656 82110 18656 0 wbs_dat_o[19]
rlabel metal2 14766 2132 14766 2132 0 wbs_dat_o[1]
rlabel metal2 521686 318546 521686 318546 0 wbs_dat_o[20]
rlabel metal2 520582 319396 520582 319396 0 wbs_dat_o[21]
rlabel metal2 520490 320314 520490 320314 0 wbs_dat_o[22]
rlabel metal2 96278 18792 96278 18792 0 wbs_dat_o[23]
rlabel metal2 99866 2166 99866 2166 0 wbs_dat_o[24]
rlabel metal2 103362 18418 103362 18418 0 wbs_dat_o[25]
rlabel metal2 106950 1826 106950 1826 0 wbs_dat_o[26]
rlabel metal2 523250 323544 523250 323544 0 wbs_dat_o[27]
rlabel metal2 114034 1792 114034 1792 0 wbs_dat_o[28]
rlabel metal2 117622 17160 117622 17160 0 wbs_dat_o[29]
rlabel metal2 19458 17058 19458 17058 0 wbs_dat_o[2]
rlabel metal2 121118 17194 121118 17194 0 wbs_dat_o[30]
rlabel metal2 405122 161942 405122 161942 0 wbs_dat_o[31]
rlabel metal2 24242 17092 24242 17092 0 wbs_dat_o[3]
rlabel metal2 407882 145010 407882 145010 0 wbs_dat_o[4]
rlabel metal2 32430 2200 32430 2200 0 wbs_dat_o[5]
rlabel metal2 36018 1894 36018 1894 0 wbs_dat_o[6]
rlabel metal2 39606 17126 39606 17126 0 wbs_dat_o[7]
rlabel metal2 43102 1928 43102 1928 0 wbs_dat_o[8]
rlabel metal2 46690 25303 46690 25303 0 wbs_dat_o[9]
rlabel metal2 5290 2183 5290 2183 0 wbs_stb_i
rlabel metal2 6486 2047 6486 2047 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
