magic
tech sky130B
magscale 1 2
timestamp 1683542783
<< viali >>
rect 2053 18717 2087 18751
rect 1777 18649 1811 18683
rect 3709 17153 3743 17187
rect 5273 17153 5307 17187
rect 5457 17153 5491 17187
rect 7481 17153 7515 17187
rect 7665 17153 7699 17187
rect 3433 17085 3467 17119
rect 3617 17085 3651 17119
rect 3525 16949 3559 16983
rect 5457 16949 5491 16983
rect 7573 16949 7607 16983
rect 7297 16677 7331 16711
rect 4445 16609 4479 16643
rect 5641 16609 5675 16643
rect 5733 16609 5767 16643
rect 5917 16609 5951 16643
rect 6561 16609 6595 16643
rect 3157 16541 3191 16575
rect 3249 16541 3283 16575
rect 4629 16541 4663 16575
rect 5825 16541 5859 16575
rect 8033 16541 8067 16575
rect 11713 16541 11747 16575
rect 3433 16473 3467 16507
rect 6745 16473 6779 16507
rect 7297 16473 7331 16507
rect 7849 16473 7883 16507
rect 8217 16473 8251 16507
rect 3157 16405 3191 16439
rect 4813 16405 4847 16439
rect 5457 16405 5491 16439
rect 6837 16405 6871 16439
rect 11621 16405 11655 16439
rect 9597 16201 9631 16235
rect 3157 16133 3191 16167
rect 3341 16133 3375 16167
rect 14933 16133 14967 16167
rect 5457 16065 5491 16099
rect 7297 16065 7331 16099
rect 7481 16065 7515 16099
rect 7573 16065 7607 16099
rect 9321 16065 9355 16099
rect 11161 16065 11195 16099
rect 12173 16065 12207 16099
rect 13001 16065 13035 16099
rect 13093 16065 13127 16099
rect 13277 16065 13311 16099
rect 13369 16065 13403 16099
rect 14565 16065 14599 16099
rect 14658 16065 14692 16099
rect 14841 16065 14875 16099
rect 15030 16065 15064 16099
rect 5549 15997 5583 16031
rect 5733 15997 5767 16031
rect 7205 15997 7239 16031
rect 10977 15997 11011 16031
rect 11897 15997 11931 16031
rect 3525 15861 3559 15895
rect 5641 15861 5675 15895
rect 7205 15861 7239 15895
rect 12817 15861 12851 15895
rect 15209 15861 15243 15895
rect 5641 15657 5675 15691
rect 6745 15657 6779 15691
rect 6837 15657 6871 15691
rect 7389 15657 7423 15691
rect 14749 15657 14783 15691
rect 16865 15657 16899 15691
rect 12265 15589 12299 15623
rect 16681 15589 16715 15623
rect 16773 15589 16807 15623
rect 6929 15521 6963 15555
rect 10333 15521 10367 15555
rect 13369 15521 13403 15555
rect 2329 15453 2363 15487
rect 2513 15453 2547 15487
rect 3065 15453 3099 15487
rect 3157 15453 3191 15487
rect 3249 15453 3283 15487
rect 4537 15453 4571 15487
rect 4629 15453 4663 15487
rect 4813 15453 4847 15487
rect 4905 15453 4939 15487
rect 6653 15453 6687 15487
rect 7389 15453 7423 15487
rect 7573 15453 7607 15487
rect 10057 15453 10091 15487
rect 10149 15453 10183 15487
rect 10425 15453 10459 15487
rect 11253 15453 11287 15487
rect 11345 15453 11379 15487
rect 11529 15453 11563 15487
rect 11621 15453 11655 15487
rect 12265 15453 12299 15487
rect 14565 15453 14599 15487
rect 14749 15453 14783 15487
rect 15301 15453 15335 15487
rect 15485 15453 15519 15487
rect 15577 15453 15611 15487
rect 15669 15453 15703 15487
rect 17141 15453 17175 15487
rect 2421 15385 2455 15419
rect 5917 15385 5951 15419
rect 13277 15385 13311 15419
rect 16405 15385 16439 15419
rect 3433 15317 3467 15351
rect 5089 15317 5123 15351
rect 9873 15317 9907 15351
rect 11069 15317 11103 15351
rect 12817 15317 12851 15351
rect 13185 15317 13219 15351
rect 15945 15317 15979 15351
rect 17049 15317 17083 15351
rect 2145 15113 2179 15147
rect 10425 15113 10459 15147
rect 10793 15113 10827 15147
rect 11713 15113 11747 15147
rect 13001 15113 13035 15147
rect 14749 15113 14783 15147
rect 2053 15045 2087 15079
rect 3893 15045 3927 15079
rect 7205 15045 7239 15079
rect 8033 15045 8067 15079
rect 9321 15045 9355 15079
rect 19165 15045 19199 15079
rect 3709 14977 3743 15011
rect 3985 14977 4019 15011
rect 4077 14977 4111 15011
rect 4721 14977 4755 15011
rect 5825 14977 5859 15011
rect 5917 14977 5951 15011
rect 6837 14977 6871 15011
rect 8217 14977 8251 15011
rect 8309 14977 8343 15011
rect 9045 14977 9079 15011
rect 10885 14977 10919 15011
rect 11897 14977 11931 15011
rect 12265 14977 12299 15011
rect 12461 14977 12495 15011
rect 13277 14977 13311 15011
rect 14657 14977 14691 15011
rect 14841 14977 14875 15011
rect 15485 14977 15519 15011
rect 15761 14977 15795 15011
rect 18337 14977 18371 15011
rect 18981 14977 19015 15011
rect 19257 14977 19291 15011
rect 2329 14909 2363 14943
rect 4997 14909 5031 14943
rect 6745 14909 6779 14943
rect 8953 14909 8987 14943
rect 9413 14909 9447 14943
rect 11069 14909 11103 14943
rect 12081 14909 12115 14943
rect 12173 14909 12207 14943
rect 13001 14909 13035 14943
rect 15577 14909 15611 14943
rect 15669 14909 15703 14943
rect 17141 14909 17175 14943
rect 17601 14909 17635 14943
rect 18061 14909 18095 14943
rect 18245 14909 18279 14943
rect 4813 14841 4847 14875
rect 6561 14841 6595 14875
rect 8033 14841 8067 14875
rect 17417 14841 17451 14875
rect 18981 14841 19015 14875
rect 1685 14773 1719 14807
rect 4261 14773 4295 14807
rect 4905 14773 4939 14807
rect 8769 14773 8803 14807
rect 13185 14773 13219 14807
rect 15301 14773 15335 14807
rect 18153 14773 18187 14807
rect 12357 14569 12391 14603
rect 14473 14569 14507 14603
rect 15577 14569 15611 14603
rect 19441 14569 19475 14603
rect 14565 14501 14599 14535
rect 18337 14501 18371 14535
rect 17509 14433 17543 14467
rect 18245 14433 18279 14467
rect 20085 14433 20119 14467
rect 7849 14365 7883 14399
rect 8125 14365 8159 14399
rect 9262 14365 9296 14399
rect 9689 14365 9723 14399
rect 9781 14365 9815 14399
rect 12265 14365 12299 14399
rect 12449 14365 12483 14399
rect 13093 14365 13127 14399
rect 13369 14365 13403 14399
rect 14289 14365 14323 14399
rect 14657 14365 14691 14399
rect 14749 14365 14783 14399
rect 15485 14365 15519 14399
rect 15669 14365 15703 14399
rect 17417 14365 17451 14399
rect 17601 14365 17635 14399
rect 18153 14365 18187 14399
rect 18429 14365 18463 14399
rect 19566 14365 19600 14399
rect 19993 14365 20027 14399
rect 7113 14297 7147 14331
rect 7297 14297 7331 14331
rect 7757 14297 7791 14331
rect 11253 14297 11287 14331
rect 6929 14229 6963 14263
rect 9137 14229 9171 14263
rect 9321 14229 9355 14263
rect 11161 14229 11195 14263
rect 12909 14229 12943 14263
rect 13277 14229 13311 14263
rect 15025 14229 15059 14263
rect 18613 14229 18647 14263
rect 19625 14229 19659 14263
rect 1593 14025 1627 14059
rect 2053 14025 2087 14059
rect 8585 14025 8619 14059
rect 14657 14025 14691 14059
rect 15761 14025 15795 14059
rect 3617 13957 3651 13991
rect 10609 13957 10643 13991
rect 18061 13957 18095 13991
rect 18153 13957 18187 13991
rect 1961 13889 1995 13923
rect 3525 13889 3559 13923
rect 3709 13889 3743 13923
rect 3893 13889 3927 13923
rect 3985 13889 4019 13923
rect 5089 13889 5123 13923
rect 5273 13889 5307 13923
rect 8401 13889 8435 13923
rect 8585 13889 8619 13923
rect 10793 13889 10827 13923
rect 11989 13889 12023 13923
rect 12081 13889 12115 13923
rect 12173 13889 12207 13923
rect 12357 13889 12391 13923
rect 13185 13889 13219 13923
rect 13369 13889 13403 13923
rect 14565 13889 14599 13923
rect 14749 13889 14783 13923
rect 15945 13889 15979 13923
rect 16037 13889 16071 13923
rect 16221 13889 16255 13923
rect 16313 13889 16347 13923
rect 17785 13889 17819 13923
rect 2237 13821 2271 13855
rect 5181 13821 5215 13855
rect 11161 13821 11195 13855
rect 17693 13821 17727 13855
rect 3341 13685 3375 13719
rect 11713 13685 11747 13719
rect 13277 13685 13311 13719
rect 17509 13685 17543 13719
rect 3065 13481 3099 13515
rect 16497 13481 16531 13515
rect 17693 13481 17727 13515
rect 19901 13481 19935 13515
rect 6469 13413 6503 13447
rect 9689 13413 9723 13447
rect 10701 13413 10735 13447
rect 13277 13413 13311 13447
rect 2329 13345 2363 13379
rect 2421 13345 2455 13379
rect 5365 13345 5399 13379
rect 5457 13345 5491 13379
rect 9229 13345 9263 13379
rect 11621 13345 11655 13379
rect 17969 13345 18003 13379
rect 18153 13345 18187 13379
rect 3341 13277 3375 13311
rect 3985 13277 4019 13311
rect 4169 13277 4203 13311
rect 6653 13277 6687 13311
rect 6745 13277 6779 13311
rect 6837 13277 6871 13311
rect 7113 13277 7147 13311
rect 9321 13277 9355 13311
rect 10333 13277 10367 13311
rect 10487 13277 10521 13311
rect 11161 13277 11195 13311
rect 11713 13277 11747 13311
rect 13001 13277 13035 13311
rect 13093 13277 13127 13311
rect 15209 13277 15243 13311
rect 15577 13277 15611 13311
rect 16313 13277 16347 13311
rect 16589 13277 16623 13311
rect 17877 13277 17911 13311
rect 18061 13277 18095 13311
rect 19993 13277 20027 13311
rect 3065 13209 3099 13243
rect 4077 13209 4111 13243
rect 6955 13209 6989 13243
rect 13277 13209 13311 13243
rect 15301 13209 15335 13243
rect 15393 13209 15427 13243
rect 1869 13141 1903 13175
rect 2237 13141 2271 13175
rect 3249 13141 3283 13175
rect 4905 13141 4939 13175
rect 5273 13141 5307 13175
rect 11345 13141 11379 13175
rect 15025 13141 15059 13175
rect 16037 13141 16071 13175
rect 2145 12937 2179 12971
rect 5089 12937 5123 12971
rect 8493 12937 8527 12971
rect 16865 12937 16899 12971
rect 18153 12937 18187 12971
rect 19809 12937 19843 12971
rect 1961 12869 1995 12903
rect 4997 12869 5031 12903
rect 9045 12869 9079 12903
rect 13461 12869 13495 12903
rect 17017 12869 17051 12903
rect 17233 12869 17267 12903
rect 19073 12869 19107 12903
rect 1777 12801 1811 12835
rect 2697 12801 2731 12835
rect 6561 12801 6595 12835
rect 6929 12801 6963 12835
rect 7297 12801 7331 12835
rect 8033 12801 8067 12835
rect 8769 12801 8803 12835
rect 10609 12801 10643 12835
rect 10885 12801 10919 12835
rect 18245 12801 18279 12835
rect 18429 12801 18463 12835
rect 18981 12801 19015 12835
rect 19257 12801 19291 12835
rect 19993 12801 20027 12835
rect 20171 12801 20205 12835
rect 3249 12733 3283 12767
rect 5181 12733 5215 12767
rect 7389 12733 7423 12767
rect 8677 12733 8711 12767
rect 9137 12733 9171 12767
rect 13093 12733 13127 12767
rect 10793 12665 10827 12699
rect 19257 12665 19291 12699
rect 4629 12597 4663 12631
rect 10701 12597 10735 12631
rect 13461 12597 13495 12631
rect 13645 12597 13679 12631
rect 17049 12597 17083 12631
rect 20085 12597 20119 12631
rect 6745 12393 6779 12427
rect 13553 12393 13587 12427
rect 15301 12393 15335 12427
rect 17693 12393 17727 12427
rect 14289 12325 14323 12359
rect 4813 12257 4847 12291
rect 4905 12257 4939 12291
rect 11253 12257 11287 12291
rect 14749 12257 14783 12291
rect 19717 12257 19751 12291
rect 2697 12189 2731 12223
rect 6377 12189 6411 12223
rect 6745 12189 6779 12223
rect 6929 12189 6963 12223
rect 10885 12189 10919 12223
rect 11345 12189 11379 12223
rect 12081 12189 12115 12223
rect 13369 12189 13403 12223
rect 13553 12189 13587 12223
rect 14473 12189 14507 12223
rect 14566 12189 14600 12223
rect 14841 12189 14875 12223
rect 15301 12189 15335 12223
rect 15485 12189 15519 12223
rect 17141 12189 17175 12223
rect 17233 12189 17267 12223
rect 17969 12189 18003 12223
rect 18061 12189 18095 12223
rect 18153 12189 18187 12223
rect 18337 12189 18371 12223
rect 20085 12189 20119 12223
rect 2881 12121 2915 12155
rect 10977 12121 11011 12155
rect 20269 12121 20303 12155
rect 4353 12053 4387 12087
rect 4721 12053 4755 12087
rect 6561 12053 6595 12087
rect 10609 12053 10643 12087
rect 11069 12053 11103 12087
rect 11989 12053 12023 12087
rect 13737 12053 13771 12087
rect 3525 11849 3559 11883
rect 4445 11849 4479 11883
rect 7297 11849 7331 11883
rect 11805 11849 11839 11883
rect 13553 11849 13587 11883
rect 18689 11849 18723 11883
rect 19717 11849 19751 11883
rect 5365 11781 5399 11815
rect 8309 11781 8343 11815
rect 12081 11781 12115 11815
rect 15945 11781 15979 11815
rect 17693 11781 17727 11815
rect 18889 11781 18923 11815
rect 2329 11713 2363 11747
rect 4353 11713 4387 11747
rect 5181 11713 5215 11747
rect 5457 11713 5491 11747
rect 5549 11713 5583 11747
rect 7205 11713 7239 11747
rect 8033 11713 8067 11747
rect 8125 11713 8159 11747
rect 8769 11713 8803 11747
rect 8953 11713 8987 11747
rect 9321 11713 9355 11747
rect 10425 11713 10459 11747
rect 10517 11713 10551 11747
rect 10609 11713 10643 11747
rect 10701 11713 10735 11747
rect 11989 11713 12023 11747
rect 12173 11713 12207 11747
rect 13185 11713 13219 11747
rect 13369 11713 13403 11747
rect 15025 11713 15059 11747
rect 15209 11713 15243 11747
rect 15669 11713 15703 11747
rect 15817 11713 15851 11747
rect 16037 11713 16071 11747
rect 16134 11713 16168 11747
rect 16865 11713 16899 11747
rect 17877 11713 17911 11747
rect 17969 11713 18003 11747
rect 19349 11713 19383 11747
rect 2053 11645 2087 11679
rect 3065 11645 3099 11679
rect 3157 11645 3191 11679
rect 4537 11645 4571 11679
rect 7389 11645 7423 11679
rect 17141 11645 17175 11679
rect 19441 11645 19475 11679
rect 8309 11577 8343 11611
rect 12357 11577 12391 11611
rect 17049 11577 17083 11611
rect 2145 11509 2179 11543
rect 2237 11509 2271 11543
rect 2881 11509 2915 11543
rect 3985 11509 4019 11543
rect 5733 11509 5767 11543
rect 6837 11509 6871 11543
rect 10241 11509 10275 11543
rect 15209 11509 15243 11543
rect 16313 11509 16347 11543
rect 16957 11509 16991 11543
rect 18521 11509 18555 11543
rect 18705 11509 18739 11543
rect 19349 11509 19383 11543
rect 1961 11305 1995 11339
rect 2513 11305 2547 11339
rect 4997 11305 5031 11339
rect 9137 11305 9171 11339
rect 11437 11305 11471 11339
rect 15945 11305 15979 11339
rect 18245 11305 18279 11339
rect 18724 11305 18758 11339
rect 18613 11237 18647 11271
rect 5365 11169 5399 11203
rect 7021 11169 7055 11203
rect 7205 11169 7239 11203
rect 9597 11169 9631 11203
rect 11621 11169 11655 11203
rect 18521 11169 18555 11203
rect 2697 11101 2731 11135
rect 2881 11101 2915 11135
rect 5181 11101 5215 11135
rect 5457 11101 5491 11135
rect 9321 11101 9355 11135
rect 9413 11101 9447 11135
rect 9505 11101 9539 11135
rect 11713 11101 11747 11135
rect 11805 11101 11839 11135
rect 11897 11101 11931 11135
rect 14473 11101 14507 11135
rect 16129 11101 16163 11135
rect 16221 11101 16255 11135
rect 1685 11033 1719 11067
rect 6929 11033 6963 11067
rect 14381 11033 14415 11067
rect 18889 11033 18923 11067
rect 6561 10965 6595 10999
rect 1961 10761 1995 10795
rect 13737 10761 13771 10795
rect 19809 10761 19843 10795
rect 1777 10693 1811 10727
rect 18061 10693 18095 10727
rect 2053 10625 2087 10659
rect 12909 10625 12943 10659
rect 13093 10625 13127 10659
rect 14013 10625 14047 10659
rect 15761 10625 15795 10659
rect 16037 10625 16071 10659
rect 16221 10625 16255 10659
rect 17877 10625 17911 10659
rect 18521 10625 18555 10659
rect 18613 10625 18647 10659
rect 18797 10625 18831 10659
rect 19717 10625 19751 10659
rect 20085 10625 20119 10659
rect 20269 10625 20303 10659
rect 13921 10557 13955 10591
rect 14105 10557 14139 10591
rect 14197 10557 14231 10591
rect 15577 10557 15611 10591
rect 17509 10557 17543 10591
rect 18981 10557 19015 10591
rect 15853 10489 15887 10523
rect 15945 10489 15979 10523
rect 1777 10421 1811 10455
rect 13001 10421 13035 10455
rect 2973 10217 3007 10251
rect 8585 10217 8619 10251
rect 11713 10217 11747 10251
rect 14381 10217 14415 10251
rect 14611 10217 14645 10251
rect 15853 10217 15887 10251
rect 16037 10217 16071 10251
rect 16497 10217 16531 10251
rect 13737 10149 13771 10183
rect 14473 10149 14507 10183
rect 1593 10013 1627 10047
rect 1860 10013 1894 10047
rect 7205 10013 7239 10047
rect 10333 10013 10367 10047
rect 10609 10013 10643 10047
rect 13553 10013 13587 10047
rect 13737 10013 13771 10047
rect 14289 10013 14323 10047
rect 14749 10013 14783 10047
rect 16497 10013 16531 10047
rect 16773 10013 16807 10047
rect 18153 10013 18187 10047
rect 18705 10013 18739 10047
rect 18889 10013 18923 10047
rect 7472 9945 7506 9979
rect 15669 9945 15703 9979
rect 15885 9945 15919 9979
rect 16681 9945 16715 9979
rect 17601 9945 17635 9979
rect 2964 9605 2998 9639
rect 4782 9605 4816 9639
rect 15301 9605 15335 9639
rect 15945 9605 15979 9639
rect 8217 9537 8251 9571
rect 9781 9537 9815 9571
rect 10048 9537 10082 9571
rect 15209 9537 15243 9571
rect 15853 9537 15887 9571
rect 16037 9537 16071 9571
rect 18981 9537 19015 9571
rect 19901 9537 19935 9571
rect 2697 9469 2731 9503
rect 4537 9469 4571 9503
rect 6837 9469 6871 9503
rect 7941 9469 7975 9503
rect 4077 9401 4111 9435
rect 19073 9401 19107 9435
rect 5917 9333 5951 9367
rect 11161 9333 11195 9367
rect 3433 9129 3467 9163
rect 5825 9129 5859 9163
rect 6469 9129 6503 9163
rect 11897 9129 11931 9163
rect 15945 9129 15979 9163
rect 18797 9129 18831 9163
rect 18705 9061 18739 9095
rect 2053 8993 2087 9027
rect 7849 8993 7883 9027
rect 10609 8993 10643 9027
rect 17049 8993 17083 9027
rect 18337 8993 18371 9027
rect 2320 8925 2354 8959
rect 4445 8925 4479 8959
rect 4712 8925 4746 8959
rect 7593 8925 7627 8959
rect 10333 8925 10367 8959
rect 13553 8925 13587 8959
rect 13737 8925 13771 8959
rect 14657 8925 14691 8959
rect 16313 8925 16347 8959
rect 16405 8925 16439 8959
rect 16865 8925 16899 8959
rect 17233 8925 17267 8959
rect 14289 8857 14323 8891
rect 14473 8857 14507 8891
rect 13737 8789 13771 8823
rect 9873 8585 9907 8619
rect 16221 8585 16255 8619
rect 18797 8585 18831 8619
rect 13921 8517 13955 8551
rect 14013 8517 14047 8551
rect 8493 8449 8527 8483
rect 8760 8449 8794 8483
rect 13829 8449 13863 8483
rect 14131 8449 14165 8483
rect 14749 8449 14783 8483
rect 14933 8449 14967 8483
rect 16129 8449 16163 8483
rect 16313 8449 16347 8483
rect 16957 8449 16991 8483
rect 17141 8449 17175 8483
rect 18153 8449 18187 8483
rect 18245 8449 18279 8483
rect 18429 8449 18463 8483
rect 18521 8449 18555 8483
rect 18613 8449 18647 8483
rect 19257 8449 19291 8483
rect 14289 8381 14323 8415
rect 19349 8381 19383 8415
rect 17141 8313 17175 8347
rect 13645 8245 13679 8279
rect 14841 8245 14875 8279
rect 2973 8041 3007 8075
rect 5917 8041 5951 8075
rect 8217 8041 8251 8075
rect 11805 8041 11839 8075
rect 1593 7905 1627 7939
rect 4537 7905 4571 7939
rect 13553 7905 13587 7939
rect 16313 7905 16347 7939
rect 18521 7905 18555 7939
rect 18705 7905 18739 7939
rect 1849 7837 1883 7871
rect 6837 7837 6871 7871
rect 10425 7837 10459 7871
rect 10681 7837 10715 7871
rect 13461 7837 13495 7871
rect 17693 7837 17727 7871
rect 18429 7837 18463 7871
rect 18613 7837 18647 7871
rect 4804 7769 4838 7803
rect 7104 7769 7138 7803
rect 16037 7769 16071 7803
rect 17785 7769 17819 7803
rect 13001 7701 13035 7735
rect 13369 7701 13403 7735
rect 15669 7701 15703 7735
rect 16129 7701 16163 7735
rect 18889 7701 18923 7735
rect 16129 7497 16163 7531
rect 16865 7497 16899 7531
rect 2605 7429 2639 7463
rect 9597 7429 9631 7463
rect 17877 7429 17911 7463
rect 4353 7361 4387 7395
rect 7849 7361 7883 7395
rect 14013 7361 14047 7395
rect 17049 7361 17083 7395
rect 17141 7361 17175 7395
rect 17417 7361 17451 7395
rect 18153 7361 18187 7395
rect 18889 7361 18923 7395
rect 19073 7361 19107 7395
rect 14289 7293 14323 7327
rect 15945 7293 15979 7327
rect 16313 7293 16347 7327
rect 18061 7293 18095 7327
rect 17325 7225 17359 7259
rect 13829 7157 13863 7191
rect 14197 7157 14231 7191
rect 15761 7157 15795 7191
rect 18153 7157 18187 7191
rect 18337 7157 18371 7191
rect 18889 7157 18923 7191
rect 15853 6953 15887 6987
rect 11713 6885 11747 6919
rect 4537 6817 4571 6851
rect 13645 6817 13679 6851
rect 14565 6817 14599 6851
rect 14933 6817 14967 6851
rect 1593 6749 1627 6783
rect 1860 6749 1894 6783
rect 4804 6749 4838 6783
rect 10333 6749 10367 6783
rect 10600 6749 10634 6783
rect 13369 6749 13403 6783
rect 14657 6749 14691 6783
rect 15669 6749 15703 6783
rect 18245 6749 18279 6783
rect 18797 6749 18831 6783
rect 19625 6749 19659 6783
rect 19901 6749 19935 6783
rect 20085 6749 20119 6783
rect 6377 6681 6411 6715
rect 15025 6681 15059 6715
rect 15485 6681 15519 6715
rect 18061 6681 18095 6715
rect 2973 6613 3007 6647
rect 5917 6613 5951 6647
rect 7665 6613 7699 6647
rect 13001 6613 13035 6647
rect 13461 6613 13495 6647
rect 14381 6613 14415 6647
rect 19441 6613 19475 6647
rect 9321 6409 9355 6443
rect 11161 6409 11195 6443
rect 13645 6409 13679 6443
rect 15301 6409 15335 6443
rect 18705 6409 18739 6443
rect 19809 6409 19843 6443
rect 2964 6341 2998 6375
rect 4804 6341 4838 6375
rect 8208 6341 8242 6375
rect 10048 6341 10082 6375
rect 15117 6341 15151 6375
rect 2697 6273 2731 6307
rect 7941 6273 7975 6307
rect 9781 6273 9815 6307
rect 13553 6273 13587 6307
rect 15393 6273 15427 6307
rect 16957 6273 16991 6307
rect 17049 6273 17083 6307
rect 18705 6273 18739 6307
rect 18889 6273 18923 6307
rect 19073 6273 19107 6307
rect 19717 6273 19751 6307
rect 19901 6273 19935 6307
rect 4537 6205 4571 6239
rect 13737 6205 13771 6239
rect 15117 6137 15151 6171
rect 4077 6069 4111 6103
rect 5917 6069 5951 6103
rect 13185 6069 13219 6103
rect 17233 6069 17267 6103
rect 5641 5865 5675 5899
rect 16405 5865 16439 5899
rect 11161 5797 11195 5831
rect 13185 5729 13219 5763
rect 17049 5729 17083 5763
rect 4261 5661 4295 5695
rect 4537 5661 4571 5695
rect 7113 5661 7147 5695
rect 7380 5661 7414 5695
rect 9781 5661 9815 5695
rect 10048 5661 10082 5695
rect 17601 5661 17635 5695
rect 17785 5661 17819 5695
rect 16773 5593 16807 5627
rect 8493 5525 8527 5559
rect 12541 5525 12575 5559
rect 12909 5525 12943 5559
rect 13001 5525 13035 5559
rect 16865 5525 16899 5559
rect 17693 5525 17727 5559
rect 6009 5321 6043 5355
rect 14841 5321 14875 5355
rect 10048 5253 10082 5287
rect 13645 5253 13679 5287
rect 15945 5253 15979 5287
rect 17693 5253 17727 5287
rect 1593 5185 1627 5219
rect 1860 5185 1894 5219
rect 4896 5185 4930 5219
rect 7113 5185 7147 5219
rect 7380 5185 7414 5219
rect 13093 5185 13127 5219
rect 14197 5185 14231 5219
rect 14381 5185 14415 5219
rect 14473 5185 14507 5219
rect 14565 5185 14599 5219
rect 15301 5185 15335 5219
rect 15485 5185 15519 5219
rect 15577 5185 15611 5219
rect 15670 5185 15704 5219
rect 17417 5185 17451 5219
rect 4629 5117 4663 5151
rect 9781 5117 9815 5151
rect 17325 5117 17359 5151
rect 17785 5117 17819 5151
rect 11161 5049 11195 5083
rect 2973 4981 3007 5015
rect 8493 4981 8527 5015
rect 17141 4981 17175 5015
rect 14381 4777 14415 4811
rect 16681 4777 16715 4811
rect 17693 4777 17727 4811
rect 18337 4777 18371 4811
rect 11713 4709 11747 4743
rect 15117 4709 15151 4743
rect 10333 4573 10367 4607
rect 14289 4573 14323 4607
rect 15209 4573 15243 4607
rect 16589 4573 16623 4607
rect 16773 4573 16807 4607
rect 17141 4573 17175 4607
rect 17601 4573 17635 4607
rect 18245 4573 18279 4607
rect 10600 4505 10634 4539
rect 16957 4437 16991 4471
rect 1869 4233 1903 4267
rect 1777 4097 1811 4131
rect 1961 4097 1995 4131
rect 3056 4097 3090 4131
rect 4629 4097 4663 4131
rect 4896 4097 4930 4131
rect 7113 4097 7147 4131
rect 7380 4097 7414 4131
rect 10048 4097 10082 4131
rect 13921 4097 13955 4131
rect 14105 4097 14139 4131
rect 14381 4097 14415 4131
rect 14473 4097 14507 4131
rect 14657 4097 14691 4131
rect 2789 4029 2823 4063
rect 9781 4029 9815 4063
rect 11161 3961 11195 3995
rect 4169 3893 4203 3927
rect 6009 3893 6043 3927
rect 8493 3893 8527 3927
rect 4077 3689 4111 3723
rect 8217 3689 8251 3723
rect 14289 3689 14323 3723
rect 16681 3689 16715 3723
rect 17141 3689 17175 3723
rect 17785 3689 17819 3723
rect 12449 3621 12483 3655
rect 1777 3553 1811 3587
rect 4169 3553 4203 3587
rect 13001 3553 13035 3587
rect 13369 3553 13403 3587
rect 14841 3553 14875 3587
rect 4261 3485 4295 3519
rect 6837 3485 6871 3519
rect 9137 3485 9171 3519
rect 11069 3485 11103 3519
rect 13173 3485 13207 3519
rect 14473 3485 14507 3519
rect 14565 3485 14599 3519
rect 14933 3485 14967 3519
rect 15393 3485 15427 3519
rect 15577 3485 15611 3519
rect 16865 3485 16899 3519
rect 16957 3485 16991 3519
rect 17233 3485 17267 3519
rect 17693 3485 17727 3519
rect 17969 3485 18003 3519
rect 18061 3485 18095 3519
rect 2044 3417 2078 3451
rect 3985 3417 4019 3451
rect 7104 3417 7138 3451
rect 9404 3417 9438 3451
rect 11336 3417 11370 3451
rect 18245 3417 18279 3451
rect 3157 3349 3191 3383
rect 10517 3349 10551 3383
rect 14657 3349 14691 3383
rect 15485 3349 15519 3383
rect 7021 3145 7055 3179
rect 9137 3145 9171 3179
rect 10057 3145 10091 3179
rect 12265 3145 12299 3179
rect 2605 3077 2639 3111
rect 4353 3077 4387 3111
rect 5641 3077 5675 3111
rect 7849 3077 7883 3111
rect 13553 3077 13587 3111
rect 5457 3009 5491 3043
rect 5549 3009 5583 3043
rect 6561 3009 6595 3043
rect 6837 3009 6871 3043
rect 10241 3009 10275 3043
rect 12265 3009 12299 3043
rect 12541 3009 12575 3043
rect 13737 3009 13771 3043
rect 14657 3009 14691 3043
rect 14841 3009 14875 3043
rect 15669 3009 15703 3043
rect 15945 3009 15979 3043
rect 16129 3009 16163 3043
rect 17141 3009 17175 3043
rect 5273 2941 5307 2975
rect 6009 2941 6043 2975
rect 10517 2941 10551 2975
rect 14013 2941 14047 2975
rect 17233 2941 17267 2975
rect 17509 2941 17543 2975
rect 6653 2873 6687 2907
rect 12357 2873 12391 2907
rect 13921 2873 13955 2907
rect 14473 2873 14507 2907
rect 10425 2805 10459 2839
rect 15485 2805 15519 2839
rect 2421 2601 2455 2635
rect 4353 2601 4387 2635
rect 5365 2601 5399 2635
rect 5549 2601 5583 2635
rect 6745 2601 6779 2635
rect 8585 2601 8619 2635
rect 12449 2601 12483 2635
rect 14841 2601 14875 2635
rect 15577 2601 15611 2635
rect 1685 2533 1719 2567
rect 11161 2533 11195 2567
rect 2789 2465 2823 2499
rect 9781 2465 9815 2499
rect 1685 2397 1719 2431
rect 1961 2397 1995 2431
rect 2605 2397 2639 2431
rect 2881 2397 2915 2431
rect 4077 2397 4111 2431
rect 4353 2397 4387 2431
rect 6561 2397 6595 2431
rect 6745 2397 6779 2431
rect 8309 2397 8343 2431
rect 8401 2397 8435 2431
rect 10048 2397 10082 2431
rect 12449 2397 12483 2431
rect 12633 2397 12667 2431
rect 12725 2397 12759 2431
rect 15761 2397 15795 2431
rect 16037 2397 16071 2431
rect 5181 2329 5215 2363
rect 5381 2329 5415 2363
rect 8585 2329 8619 2363
rect 14657 2329 14691 2363
rect 14857 2329 14891 2363
rect 1869 2261 1903 2295
rect 4169 2261 4203 2295
rect 15025 2261 15059 2295
rect 15945 2261 15979 2295
<< metal1 >>
rect 1104 19610 21043 19632
rect 1104 19558 5894 19610
rect 5946 19558 5958 19610
rect 6010 19558 6022 19610
rect 6074 19558 6086 19610
rect 6138 19558 6150 19610
rect 6202 19558 10839 19610
rect 10891 19558 10903 19610
rect 10955 19558 10967 19610
rect 11019 19558 11031 19610
rect 11083 19558 11095 19610
rect 11147 19558 15784 19610
rect 15836 19558 15848 19610
rect 15900 19558 15912 19610
rect 15964 19558 15976 19610
rect 16028 19558 16040 19610
rect 16092 19558 20729 19610
rect 20781 19558 20793 19610
rect 20845 19558 20857 19610
rect 20909 19558 20921 19610
rect 20973 19558 20985 19610
rect 21037 19558 21043 19610
rect 1104 19536 21043 19558
rect 1104 19066 20884 19088
rect 1104 19014 3422 19066
rect 3474 19014 3486 19066
rect 3538 19014 3550 19066
rect 3602 19014 3614 19066
rect 3666 19014 3678 19066
rect 3730 19014 8367 19066
rect 8419 19014 8431 19066
rect 8483 19014 8495 19066
rect 8547 19014 8559 19066
rect 8611 19014 8623 19066
rect 8675 19014 13312 19066
rect 13364 19014 13376 19066
rect 13428 19014 13440 19066
rect 13492 19014 13504 19066
rect 13556 19014 13568 19066
rect 13620 19014 18257 19066
rect 18309 19014 18321 19066
rect 18373 19014 18385 19066
rect 18437 19014 18449 19066
rect 18501 19014 18513 19066
rect 18565 19014 20884 19066
rect 1104 18992 20884 19014
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18748 2099 18751
rect 2498 18748 2504 18760
rect 2087 18720 2504 18748
rect 2087 18717 2099 18720
rect 2041 18711 2099 18717
rect 2498 18708 2504 18720
rect 2556 18708 2562 18760
rect 934 18640 940 18692
rect 992 18680 998 18692
rect 1765 18683 1823 18689
rect 1765 18680 1777 18683
rect 992 18652 1777 18680
rect 992 18640 998 18652
rect 1765 18649 1777 18652
rect 1811 18649 1823 18683
rect 1765 18643 1823 18649
rect 1104 18522 21043 18544
rect 1104 18470 5894 18522
rect 5946 18470 5958 18522
rect 6010 18470 6022 18522
rect 6074 18470 6086 18522
rect 6138 18470 6150 18522
rect 6202 18470 10839 18522
rect 10891 18470 10903 18522
rect 10955 18470 10967 18522
rect 11019 18470 11031 18522
rect 11083 18470 11095 18522
rect 11147 18470 15784 18522
rect 15836 18470 15848 18522
rect 15900 18470 15912 18522
rect 15964 18470 15976 18522
rect 16028 18470 16040 18522
rect 16092 18470 20729 18522
rect 20781 18470 20793 18522
rect 20845 18470 20857 18522
rect 20909 18470 20921 18522
rect 20973 18470 20985 18522
rect 21037 18470 21043 18522
rect 1104 18448 21043 18470
rect 1104 17978 20884 18000
rect 1104 17926 3422 17978
rect 3474 17926 3486 17978
rect 3538 17926 3550 17978
rect 3602 17926 3614 17978
rect 3666 17926 3678 17978
rect 3730 17926 8367 17978
rect 8419 17926 8431 17978
rect 8483 17926 8495 17978
rect 8547 17926 8559 17978
rect 8611 17926 8623 17978
rect 8675 17926 13312 17978
rect 13364 17926 13376 17978
rect 13428 17926 13440 17978
rect 13492 17926 13504 17978
rect 13556 17926 13568 17978
rect 13620 17926 18257 17978
rect 18309 17926 18321 17978
rect 18373 17926 18385 17978
rect 18437 17926 18449 17978
rect 18501 17926 18513 17978
rect 18565 17926 20884 17978
rect 1104 17904 20884 17926
rect 1104 17434 21043 17456
rect 1104 17382 5894 17434
rect 5946 17382 5958 17434
rect 6010 17382 6022 17434
rect 6074 17382 6086 17434
rect 6138 17382 6150 17434
rect 6202 17382 10839 17434
rect 10891 17382 10903 17434
rect 10955 17382 10967 17434
rect 11019 17382 11031 17434
rect 11083 17382 11095 17434
rect 11147 17382 15784 17434
rect 15836 17382 15848 17434
rect 15900 17382 15912 17434
rect 15964 17382 15976 17434
rect 16028 17382 16040 17434
rect 16092 17382 20729 17434
rect 20781 17382 20793 17434
rect 20845 17382 20857 17434
rect 20909 17382 20921 17434
rect 20973 17382 20985 17434
rect 21037 17382 21043 17434
rect 1104 17360 21043 17382
rect 5276 17224 7512 17252
rect 3050 17144 3056 17196
rect 3108 17184 3114 17196
rect 3697 17187 3755 17193
rect 3697 17184 3709 17187
rect 3108 17156 3709 17184
rect 3108 17144 3114 17156
rect 3697 17153 3709 17156
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 4062 17144 4068 17196
rect 4120 17184 4126 17196
rect 5276 17193 5304 17224
rect 5261 17187 5319 17193
rect 5261 17184 5273 17187
rect 4120 17156 5273 17184
rect 4120 17144 4126 17156
rect 5261 17153 5273 17156
rect 5307 17153 5319 17187
rect 5261 17147 5319 17153
rect 5445 17187 5503 17193
rect 5445 17153 5457 17187
rect 5491 17184 5503 17187
rect 5994 17184 6000 17196
rect 5491 17156 6000 17184
rect 5491 17153 5503 17156
rect 5445 17147 5503 17153
rect 3421 17119 3479 17125
rect 3421 17085 3433 17119
rect 3467 17085 3479 17119
rect 3421 17079 3479 17085
rect 3605 17119 3663 17125
rect 3605 17085 3617 17119
rect 3651 17116 3663 17119
rect 5460 17116 5488 17147
rect 5994 17144 6000 17156
rect 6052 17144 6058 17196
rect 7484 17193 7512 17224
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17153 7527 17187
rect 7469 17147 7527 17153
rect 7653 17187 7711 17193
rect 7653 17153 7665 17187
rect 7699 17184 7711 17187
rect 8110 17184 8116 17196
rect 7699 17156 8116 17184
rect 7699 17153 7711 17156
rect 7653 17147 7711 17153
rect 3651 17088 5488 17116
rect 7484 17116 7512 17147
rect 8110 17144 8116 17156
rect 8168 17144 8174 17196
rect 7742 17116 7748 17128
rect 7484 17088 7748 17116
rect 3651 17085 3663 17088
rect 3605 17079 3663 17085
rect 3326 17008 3332 17060
rect 3384 17048 3390 17060
rect 3436 17048 3464 17079
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 4062 17048 4068 17060
rect 3384 17020 4068 17048
rect 3384 17008 3390 17020
rect 4062 17008 4068 17020
rect 4120 17008 4126 17060
rect 3142 16940 3148 16992
rect 3200 16980 3206 16992
rect 3513 16983 3571 16989
rect 3513 16980 3525 16983
rect 3200 16952 3525 16980
rect 3200 16940 3206 16952
rect 3513 16949 3525 16952
rect 3559 16949 3571 16983
rect 3513 16943 3571 16949
rect 5442 16940 5448 16992
rect 5500 16940 5506 16992
rect 7282 16940 7288 16992
rect 7340 16980 7346 16992
rect 7561 16983 7619 16989
rect 7561 16980 7573 16983
rect 7340 16952 7573 16980
rect 7340 16940 7346 16952
rect 7561 16949 7573 16952
rect 7607 16949 7619 16983
rect 7561 16943 7619 16949
rect 1104 16890 20884 16912
rect 1104 16838 3422 16890
rect 3474 16838 3486 16890
rect 3538 16838 3550 16890
rect 3602 16838 3614 16890
rect 3666 16838 3678 16890
rect 3730 16838 8367 16890
rect 8419 16838 8431 16890
rect 8483 16838 8495 16890
rect 8547 16838 8559 16890
rect 8611 16838 8623 16890
rect 8675 16838 13312 16890
rect 13364 16838 13376 16890
rect 13428 16838 13440 16890
rect 13492 16838 13504 16890
rect 13556 16838 13568 16890
rect 13620 16838 18257 16890
rect 18309 16838 18321 16890
rect 18373 16838 18385 16890
rect 18437 16838 18449 16890
rect 18501 16838 18513 16890
rect 18565 16838 20884 16890
rect 1104 16816 20884 16838
rect 5810 16736 5816 16788
rect 5868 16776 5874 16788
rect 5868 16748 7328 16776
rect 5868 16736 5874 16748
rect 4062 16668 4068 16720
rect 4120 16708 4126 16720
rect 5994 16708 6000 16720
rect 4120 16680 4476 16708
rect 4120 16668 4126 16680
rect 4448 16649 4476 16680
rect 4632 16680 6000 16708
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16609 4491 16643
rect 4433 16603 4491 16609
rect 3142 16532 3148 16584
rect 3200 16532 3206 16584
rect 3234 16532 3240 16584
rect 3292 16572 3298 16584
rect 4062 16572 4068 16584
rect 3292 16544 4068 16572
rect 3292 16532 3298 16544
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 4632 16581 4660 16680
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 7300 16717 7328 16748
rect 7285 16711 7343 16717
rect 7285 16677 7297 16711
rect 7331 16708 7343 16711
rect 7558 16708 7564 16720
rect 7331 16680 7564 16708
rect 7331 16677 7343 16680
rect 7285 16671 7343 16677
rect 7558 16668 7564 16680
rect 7616 16668 7622 16720
rect 5442 16600 5448 16652
rect 5500 16640 5506 16652
rect 5629 16643 5687 16649
rect 5629 16640 5641 16643
rect 5500 16612 5641 16640
rect 5500 16600 5506 16612
rect 5629 16609 5641 16612
rect 5675 16609 5687 16643
rect 5629 16603 5687 16609
rect 5718 16600 5724 16652
rect 5776 16600 5782 16652
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16640 5963 16643
rect 6549 16643 6607 16649
rect 6549 16640 6561 16643
rect 5951 16612 6561 16640
rect 5951 16609 5963 16612
rect 5905 16603 5963 16609
rect 6549 16609 6561 16612
rect 6595 16609 6607 16643
rect 6549 16603 6607 16609
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 5810 16532 5816 16584
rect 5868 16532 5874 16584
rect 5994 16532 6000 16584
rect 6052 16572 6058 16584
rect 6052 16544 7328 16572
rect 6052 16532 6058 16544
rect 3421 16507 3479 16513
rect 3421 16473 3433 16507
rect 3467 16504 3479 16507
rect 4338 16504 4344 16516
rect 3467 16476 4344 16504
rect 3467 16473 3479 16476
rect 3421 16467 3479 16473
rect 4338 16464 4344 16476
rect 4396 16504 4402 16516
rect 6733 16507 6791 16513
rect 4396 16476 6132 16504
rect 4396 16464 4402 16476
rect 3142 16396 3148 16448
rect 3200 16396 3206 16448
rect 4798 16396 4804 16448
rect 4856 16396 4862 16448
rect 5258 16396 5264 16448
rect 5316 16436 5322 16448
rect 5445 16439 5503 16445
rect 5445 16436 5457 16439
rect 5316 16408 5457 16436
rect 5316 16396 5322 16408
rect 5445 16405 5457 16408
rect 5491 16405 5503 16439
rect 6104 16436 6132 16476
rect 6733 16473 6745 16507
rect 6779 16504 6791 16507
rect 7190 16504 7196 16516
rect 6779 16476 7196 16504
rect 6779 16473 6791 16476
rect 6733 16467 6791 16473
rect 7190 16464 7196 16476
rect 7248 16464 7254 16516
rect 7300 16513 7328 16544
rect 7742 16532 7748 16584
rect 7800 16572 7806 16584
rect 8021 16575 8079 16581
rect 8021 16572 8033 16575
rect 7800 16544 8033 16572
rect 7800 16532 7806 16544
rect 8021 16541 8033 16544
rect 8067 16541 8079 16575
rect 8021 16535 8079 16541
rect 11330 16532 11336 16584
rect 11388 16572 11394 16584
rect 11701 16575 11759 16581
rect 11701 16572 11713 16575
rect 11388 16544 11713 16572
rect 11388 16532 11394 16544
rect 11701 16541 11713 16544
rect 11747 16541 11759 16575
rect 11701 16535 11759 16541
rect 7285 16507 7343 16513
rect 7285 16473 7297 16507
rect 7331 16504 7343 16507
rect 7374 16504 7380 16516
rect 7331 16476 7380 16504
rect 7331 16473 7343 16476
rect 7285 16467 7343 16473
rect 7374 16464 7380 16476
rect 7432 16464 7438 16516
rect 7837 16507 7895 16513
rect 7837 16473 7849 16507
rect 7883 16473 7895 16507
rect 7837 16467 7895 16473
rect 6825 16439 6883 16445
rect 6825 16436 6837 16439
rect 6104 16408 6837 16436
rect 5445 16399 5503 16405
rect 6825 16405 6837 16408
rect 6871 16436 6883 16439
rect 7466 16436 7472 16448
rect 6871 16408 7472 16436
rect 6871 16405 6883 16408
rect 6825 16399 6883 16405
rect 7466 16396 7472 16408
rect 7524 16436 7530 16448
rect 7852 16436 7880 16467
rect 8110 16464 8116 16516
rect 8168 16504 8174 16516
rect 8205 16507 8263 16513
rect 8205 16504 8217 16507
rect 8168 16476 8217 16504
rect 8168 16464 8174 16476
rect 8205 16473 8217 16476
rect 8251 16473 8263 16507
rect 8205 16467 8263 16473
rect 7524 16408 7880 16436
rect 7524 16396 7530 16408
rect 11606 16396 11612 16448
rect 11664 16436 11670 16448
rect 13078 16436 13084 16448
rect 11664 16408 13084 16436
rect 11664 16396 11670 16408
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 1104 16346 21043 16368
rect 1104 16294 5894 16346
rect 5946 16294 5958 16346
rect 6010 16294 6022 16346
rect 6074 16294 6086 16346
rect 6138 16294 6150 16346
rect 6202 16294 10839 16346
rect 10891 16294 10903 16346
rect 10955 16294 10967 16346
rect 11019 16294 11031 16346
rect 11083 16294 11095 16346
rect 11147 16294 15784 16346
rect 15836 16294 15848 16346
rect 15900 16294 15912 16346
rect 15964 16294 15976 16346
rect 16028 16294 16040 16346
rect 16092 16294 20729 16346
rect 20781 16294 20793 16346
rect 20845 16294 20857 16346
rect 20909 16294 20921 16346
rect 20973 16294 20985 16346
rect 21037 16294 21043 16346
rect 1104 16272 21043 16294
rect 8018 16192 8024 16244
rect 8076 16232 8082 16244
rect 9585 16235 9643 16241
rect 9585 16232 9597 16235
rect 8076 16204 9597 16232
rect 8076 16192 8082 16204
rect 9585 16201 9597 16204
rect 9631 16232 9643 16235
rect 9631 16204 14412 16232
rect 9631 16201 9643 16204
rect 9585 16195 9643 16201
rect 3145 16167 3203 16173
rect 3145 16133 3157 16167
rect 3191 16164 3203 16167
rect 3234 16164 3240 16176
rect 3191 16136 3240 16164
rect 3191 16133 3203 16136
rect 3145 16127 3203 16133
rect 3234 16124 3240 16136
rect 3292 16124 3298 16176
rect 3326 16124 3332 16176
rect 3384 16124 3390 16176
rect 12710 16124 12716 16176
rect 12768 16164 12774 16176
rect 12768 16136 13400 16164
rect 12768 16124 12774 16136
rect 5442 16056 5448 16108
rect 5500 16056 5506 16108
rect 7282 16056 7288 16108
rect 7340 16056 7346 16108
rect 7466 16056 7472 16108
rect 7524 16056 7530 16108
rect 7558 16056 7564 16108
rect 7616 16056 7622 16108
rect 8938 16056 8944 16108
rect 8996 16096 9002 16108
rect 9309 16099 9367 16105
rect 9309 16096 9321 16099
rect 8996 16068 9321 16096
rect 8996 16056 9002 16068
rect 9309 16065 9321 16068
rect 9355 16065 9367 16099
rect 9309 16059 9367 16065
rect 11149 16099 11207 16105
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11606 16096 11612 16108
rect 11195 16068 11612 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 4798 15988 4804 16040
rect 4856 16028 4862 16040
rect 5537 16031 5595 16037
rect 5537 16028 5549 16031
rect 4856 16000 5549 16028
rect 4856 15988 4862 16000
rect 5537 15997 5549 16000
rect 5583 15997 5595 16031
rect 5537 15991 5595 15997
rect 5626 15988 5632 16040
rect 5684 16028 5690 16040
rect 5721 16031 5779 16037
rect 5721 16028 5733 16031
rect 5684 16000 5733 16028
rect 5684 15988 5690 16000
rect 5721 15997 5733 16000
rect 5767 16028 5779 16031
rect 5810 16028 5816 16040
rect 5767 16000 5816 16028
rect 5767 15997 5779 16000
rect 5721 15991 5779 15997
rect 5810 15988 5816 16000
rect 5868 15988 5874 16040
rect 6822 15988 6828 16040
rect 6880 16028 6886 16040
rect 7193 16031 7251 16037
rect 7193 16028 7205 16031
rect 6880 16000 7205 16028
rect 6880 15988 6886 16000
rect 7193 15997 7205 16000
rect 7239 15997 7251 16031
rect 7193 15991 7251 15997
rect 9324 15960 9352 16059
rect 11606 16056 11612 16068
rect 11664 16056 11670 16108
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12434 16096 12440 16108
rect 12207 16068 12440 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 10410 15988 10416 16040
rect 10468 16028 10474 16040
rect 10965 16031 11023 16037
rect 10965 16028 10977 16031
rect 10468 16000 10977 16028
rect 10468 15988 10474 16000
rect 10965 15997 10977 16000
rect 11011 16028 11023 16031
rect 11698 16028 11704 16040
rect 11011 16000 11704 16028
rect 11011 15997 11023 16000
rect 10965 15991 11023 15997
rect 11698 15988 11704 16000
rect 11756 15988 11762 16040
rect 11882 15988 11888 16040
rect 11940 15988 11946 16040
rect 13004 16028 13032 16059
rect 13078 16056 13084 16108
rect 13136 16056 13142 16108
rect 13372 16105 13400 16136
rect 14384 16108 14412 16204
rect 14458 16124 14464 16176
rect 14516 16164 14522 16176
rect 14921 16167 14979 16173
rect 14921 16164 14933 16167
rect 14516 16136 14933 16164
rect 14516 16124 14522 16136
rect 14921 16133 14933 16136
rect 14967 16133 14979 16167
rect 14921 16127 14979 16133
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 13170 16028 13176 16040
rect 13004 16000 13176 16028
rect 13170 15988 13176 16000
rect 13228 15988 13234 16040
rect 13280 16028 13308 16059
rect 14366 16056 14372 16108
rect 14424 16096 14430 16108
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 14424 16068 14565 16096
rect 14424 16056 14430 16068
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 13722 16028 13728 16040
rect 13280 16000 13728 16028
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 14568 16028 14596 16059
rect 14642 16056 14648 16108
rect 14700 16096 14706 16108
rect 14700 16068 14745 16096
rect 14700 16056 14706 16068
rect 14826 16056 14832 16108
rect 14884 16056 14890 16108
rect 15010 16056 15016 16108
rect 15068 16105 15074 16108
rect 15068 16059 15076 16105
rect 15068 16056 15074 16059
rect 15102 16028 15108 16040
rect 14568 16000 15108 16028
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 11606 15960 11612 15972
rect 9324 15932 11612 15960
rect 11606 15920 11612 15932
rect 11664 15960 11670 15972
rect 15654 15960 15660 15972
rect 11664 15932 15660 15960
rect 11664 15920 11670 15932
rect 15654 15920 15660 15932
rect 15712 15920 15718 15972
rect 3234 15852 3240 15904
rect 3292 15892 3298 15904
rect 3513 15895 3571 15901
rect 3513 15892 3525 15895
rect 3292 15864 3525 15892
rect 3292 15852 3298 15864
rect 3513 15861 3525 15864
rect 3559 15861 3571 15895
rect 3513 15855 3571 15861
rect 5629 15895 5687 15901
rect 5629 15861 5641 15895
rect 5675 15892 5687 15895
rect 6730 15892 6736 15904
rect 5675 15864 6736 15892
rect 5675 15861 5687 15864
rect 5629 15855 5687 15861
rect 6730 15852 6736 15864
rect 6788 15852 6794 15904
rect 7190 15852 7196 15904
rect 7248 15852 7254 15904
rect 12802 15852 12808 15904
rect 12860 15852 12866 15904
rect 15194 15852 15200 15904
rect 15252 15852 15258 15904
rect 1104 15802 20884 15824
rect 1104 15750 3422 15802
rect 3474 15750 3486 15802
rect 3538 15750 3550 15802
rect 3602 15750 3614 15802
rect 3666 15750 3678 15802
rect 3730 15750 8367 15802
rect 8419 15750 8431 15802
rect 8483 15750 8495 15802
rect 8547 15750 8559 15802
rect 8611 15750 8623 15802
rect 8675 15750 13312 15802
rect 13364 15750 13376 15802
rect 13428 15750 13440 15802
rect 13492 15750 13504 15802
rect 13556 15750 13568 15802
rect 13620 15750 18257 15802
rect 18309 15750 18321 15802
rect 18373 15750 18385 15802
rect 18437 15750 18449 15802
rect 18501 15750 18513 15802
rect 18565 15750 20884 15802
rect 1104 15728 20884 15750
rect 3970 15648 3976 15700
rect 4028 15688 4034 15700
rect 5626 15688 5632 15700
rect 4028 15660 5632 15688
rect 4028 15648 4034 15660
rect 5626 15648 5632 15660
rect 5684 15688 5690 15700
rect 6733 15691 6791 15697
rect 6733 15688 6745 15691
rect 5684 15660 6745 15688
rect 5684 15648 5690 15660
rect 6733 15657 6745 15660
rect 6779 15657 6791 15691
rect 6733 15651 6791 15657
rect 4062 15620 4068 15632
rect 2746 15592 4068 15620
rect 2746 15552 2774 15592
rect 4062 15580 4068 15592
rect 4120 15620 4126 15632
rect 5718 15620 5724 15632
rect 4120 15592 5724 15620
rect 4120 15580 4126 15592
rect 5718 15580 5724 15592
rect 5776 15580 5782 15632
rect 6748 15620 6776 15651
rect 6822 15648 6828 15700
rect 6880 15648 6886 15700
rect 7374 15648 7380 15700
rect 7432 15648 7438 15700
rect 11238 15648 11244 15700
rect 11296 15688 11302 15700
rect 14737 15691 14795 15697
rect 11296 15660 14136 15688
rect 11296 15648 11302 15660
rect 7098 15620 7104 15632
rect 6748 15592 7104 15620
rect 7098 15580 7104 15592
rect 7156 15580 7162 15632
rect 10060 15592 11008 15620
rect 3326 15552 3332 15564
rect 2332 15524 2774 15552
rect 2976 15524 3332 15552
rect 2332 15493 2360 15524
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15453 2375 15487
rect 2317 15447 2375 15453
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15484 2559 15487
rect 2976 15484 3004 15524
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 4338 15512 4344 15564
rect 4396 15552 4402 15564
rect 4396 15524 4844 15552
rect 4396 15512 4402 15524
rect 2547 15456 3004 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 3050 15444 3056 15496
rect 3108 15444 3114 15496
rect 3145 15487 3203 15493
rect 3145 15453 3157 15487
rect 3191 15453 3203 15487
rect 3145 15447 3203 15453
rect 2409 15419 2467 15425
rect 2409 15385 2421 15419
rect 2455 15416 2467 15419
rect 3160 15416 3188 15447
rect 3234 15444 3240 15496
rect 3292 15444 3298 15496
rect 3970 15444 3976 15496
rect 4028 15484 4034 15496
rect 4525 15487 4583 15493
rect 4525 15484 4537 15487
rect 4028 15456 4537 15484
rect 4028 15444 4034 15456
rect 4525 15453 4537 15456
rect 4571 15453 4583 15487
rect 4525 15447 4583 15453
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15484 4675 15487
rect 4706 15484 4712 15496
rect 4663 15456 4712 15484
rect 4663 15453 4675 15456
rect 4617 15447 4675 15453
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 4816 15493 4844 15524
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 6972 15524 7604 15552
rect 6972 15512 6978 15524
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15453 4859 15487
rect 4801 15447 4859 15453
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15453 4951 15487
rect 4893 15447 4951 15453
rect 3694 15416 3700 15428
rect 2455 15388 3700 15416
rect 2455 15385 2467 15388
rect 2409 15379 2467 15385
rect 3694 15376 3700 15388
rect 3752 15416 3758 15428
rect 4908 15416 4936 15447
rect 6638 15444 6644 15496
rect 6696 15444 6702 15496
rect 7576 15493 7604 15524
rect 10060 15493 10088 15592
rect 10318 15512 10324 15564
rect 10376 15512 10382 15564
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15453 7435 15487
rect 7377 15447 7435 15453
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15453 7619 15487
rect 7561 15447 7619 15453
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15453 10103 15487
rect 10045 15447 10103 15453
rect 10137 15487 10195 15493
rect 10137 15453 10149 15487
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 3752 15388 4936 15416
rect 5905 15419 5963 15425
rect 3752 15376 3758 15388
rect 5905 15385 5917 15419
rect 5951 15416 5963 15419
rect 6362 15416 6368 15428
rect 5951 15388 6368 15416
rect 5951 15385 5963 15388
rect 5905 15379 5963 15385
rect 6362 15376 6368 15388
rect 6420 15376 6426 15428
rect 7392 15416 7420 15447
rect 8110 15416 8116 15428
rect 7392 15388 8116 15416
rect 8110 15376 8116 15388
rect 8168 15376 8174 15428
rect 10152 15416 10180 15447
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 10410 15484 10416 15496
rect 10284 15456 10416 15484
rect 10284 15444 10290 15456
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 10980 15484 11008 15592
rect 11146 15580 11152 15632
rect 11204 15620 11210 15632
rect 11790 15620 11796 15632
rect 11204 15592 11796 15620
rect 11204 15580 11210 15592
rect 11790 15580 11796 15592
rect 11848 15580 11854 15632
rect 12253 15623 12311 15629
rect 12253 15589 12265 15623
rect 12299 15620 12311 15623
rect 12434 15620 12440 15632
rect 12299 15592 12440 15620
rect 12299 15589 12311 15592
rect 12253 15583 12311 15589
rect 12434 15580 12440 15592
rect 12492 15580 12498 15632
rect 13170 15580 13176 15632
rect 13228 15620 13234 15632
rect 14108 15620 14136 15660
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 15010 15688 15016 15700
rect 14783 15660 15016 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 15010 15648 15016 15660
rect 15068 15648 15074 15700
rect 15102 15648 15108 15700
rect 15160 15688 15166 15700
rect 16853 15691 16911 15697
rect 16853 15688 16865 15691
rect 15160 15660 16865 15688
rect 15160 15648 15166 15660
rect 16853 15657 16865 15660
rect 16899 15688 16911 15691
rect 18138 15688 18144 15700
rect 16899 15660 18144 15688
rect 16899 15657 16911 15660
rect 16853 15651 16911 15657
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 16669 15623 16727 15629
rect 16669 15620 16681 15623
rect 13228 15592 13400 15620
rect 14108 15592 14780 15620
rect 13228 15580 13234 15592
rect 13372 15561 13400 15592
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15521 13415 15555
rect 13357 15515 13415 15521
rect 11054 15484 11060 15496
rect 10980 15456 11060 15484
rect 11054 15444 11060 15456
rect 11112 15444 11118 15496
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 11146 15416 11152 15428
rect 10152 15388 11152 15416
rect 11146 15376 11152 15388
rect 11204 15376 11210 15428
rect 3326 15308 3332 15360
rect 3384 15348 3390 15360
rect 3421 15351 3479 15357
rect 3421 15348 3433 15351
rect 3384 15320 3433 15348
rect 3384 15308 3390 15320
rect 3421 15317 3433 15320
rect 3467 15317 3479 15351
rect 3421 15311 3479 15317
rect 4982 15308 4988 15360
rect 5040 15348 5046 15360
rect 5077 15351 5135 15357
rect 5077 15348 5089 15351
rect 5040 15320 5089 15348
rect 5040 15308 5046 15320
rect 5077 15317 5089 15320
rect 5123 15317 5135 15351
rect 5077 15311 5135 15317
rect 9858 15308 9864 15360
rect 9916 15308 9922 15360
rect 10686 15308 10692 15360
rect 10744 15348 10750 15360
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 10744 15320 11069 15348
rect 10744 15308 10750 15320
rect 11057 15317 11069 15320
rect 11103 15317 11115 15351
rect 11256 15348 11284 15447
rect 11330 15444 11336 15496
rect 11388 15444 11394 15496
rect 11514 15444 11520 15496
rect 11572 15444 11578 15496
rect 11606 15444 11612 15496
rect 11664 15444 11670 15496
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15484 12311 15487
rect 12894 15484 12900 15496
rect 12299 15456 12900 15484
rect 12299 15453 12311 15456
rect 12253 15447 12311 15453
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 14553 15487 14611 15493
rect 14553 15484 14565 15487
rect 13096 15456 14565 15484
rect 11882 15376 11888 15428
rect 11940 15416 11946 15428
rect 13096 15416 13124 15456
rect 14553 15453 14565 15456
rect 14599 15484 14611 15487
rect 14642 15484 14648 15496
rect 14599 15456 14648 15484
rect 14599 15453 14611 15456
rect 14553 15447 14611 15453
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 14752 15493 14780 15592
rect 15120 15592 16681 15620
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 15010 15484 15016 15496
rect 14783 15456 15016 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 15010 15444 15016 15456
rect 15068 15444 15074 15496
rect 11940 15388 13124 15416
rect 13265 15419 13323 15425
rect 11940 15376 11946 15388
rect 13265 15385 13277 15419
rect 13311 15416 13323 15419
rect 13814 15416 13820 15428
rect 13311 15388 13820 15416
rect 13311 15385 13323 15388
rect 13265 15379 13323 15385
rect 13814 15376 13820 15388
rect 13872 15376 13878 15428
rect 12805 15351 12863 15357
rect 12805 15348 12817 15351
rect 11256 15320 12817 15348
rect 11057 15311 11115 15317
rect 12805 15317 12817 15320
rect 12851 15317 12863 15351
rect 12805 15311 12863 15317
rect 12986 15308 12992 15360
rect 13044 15348 13050 15360
rect 13173 15351 13231 15357
rect 13173 15348 13185 15351
rect 13044 15320 13185 15348
rect 13044 15308 13050 15320
rect 13173 15317 13185 15320
rect 13219 15348 13231 15351
rect 15120 15348 15148 15592
rect 16669 15589 16681 15592
rect 16715 15589 16727 15623
rect 16669 15583 16727 15589
rect 16758 15580 16764 15632
rect 16816 15580 16822 15632
rect 18874 15552 18880 15564
rect 15580 15524 18880 15552
rect 15286 15444 15292 15496
rect 15344 15444 15350 15496
rect 15580 15493 15608 15524
rect 18874 15512 18880 15524
rect 18932 15512 18938 15564
rect 15473 15487 15531 15493
rect 15473 15453 15485 15487
rect 15519 15453 15531 15487
rect 15473 15447 15531 15453
rect 15565 15487 15623 15493
rect 15565 15453 15577 15487
rect 15611 15453 15623 15487
rect 15565 15447 15623 15453
rect 15488 15416 15516 15447
rect 15654 15444 15660 15496
rect 15712 15484 15718 15496
rect 16482 15484 16488 15496
rect 15712 15456 16488 15484
rect 15712 15444 15718 15456
rect 16482 15444 16488 15456
rect 16540 15444 16546 15496
rect 17129 15487 17187 15493
rect 17129 15453 17141 15487
rect 17175 15484 17187 15487
rect 17402 15484 17408 15496
rect 17175 15456 17408 15484
rect 17175 15453 17187 15456
rect 17129 15447 17187 15453
rect 17402 15444 17408 15456
rect 17460 15444 17466 15496
rect 16393 15419 16451 15425
rect 16393 15416 16405 15419
rect 15488 15388 16405 15416
rect 16393 15385 16405 15388
rect 16439 15385 16451 15419
rect 16393 15379 16451 15385
rect 13219 15320 15148 15348
rect 13219 15317 13231 15320
rect 13173 15311 13231 15317
rect 15654 15308 15660 15360
rect 15712 15348 15718 15360
rect 15933 15351 15991 15357
rect 15933 15348 15945 15351
rect 15712 15320 15945 15348
rect 15712 15308 15718 15320
rect 15933 15317 15945 15320
rect 15979 15317 15991 15351
rect 15933 15311 15991 15317
rect 17037 15351 17095 15357
rect 17037 15317 17049 15351
rect 17083 15348 17095 15351
rect 17862 15348 17868 15360
rect 17083 15320 17868 15348
rect 17083 15317 17095 15320
rect 17037 15311 17095 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 1104 15258 21043 15280
rect 1104 15206 5894 15258
rect 5946 15206 5958 15258
rect 6010 15206 6022 15258
rect 6074 15206 6086 15258
rect 6138 15206 6150 15258
rect 6202 15206 10839 15258
rect 10891 15206 10903 15258
rect 10955 15206 10967 15258
rect 11019 15206 11031 15258
rect 11083 15206 11095 15258
rect 11147 15206 15784 15258
rect 15836 15206 15848 15258
rect 15900 15206 15912 15258
rect 15964 15206 15976 15258
rect 16028 15206 16040 15258
rect 16092 15206 20729 15258
rect 20781 15206 20793 15258
rect 20845 15206 20857 15258
rect 20909 15206 20921 15258
rect 20973 15206 20985 15258
rect 21037 15206 21043 15258
rect 1104 15184 21043 15206
rect 2133 15147 2191 15153
rect 2133 15113 2145 15147
rect 2179 15144 2191 15147
rect 3142 15144 3148 15156
rect 2179 15116 3148 15144
rect 2179 15113 2191 15116
rect 2133 15107 2191 15113
rect 3142 15104 3148 15116
rect 3200 15104 3206 15156
rect 6822 15144 6828 15156
rect 5828 15116 6828 15144
rect 2041 15079 2099 15085
rect 2041 15045 2053 15079
rect 2087 15076 2099 15079
rect 2222 15076 2228 15088
rect 2087 15048 2228 15076
rect 2087 15045 2099 15048
rect 2041 15039 2099 15045
rect 2222 15036 2228 15048
rect 2280 15036 2286 15088
rect 3234 15036 3240 15088
rect 3292 15076 3298 15088
rect 3881 15079 3939 15085
rect 3881 15076 3893 15079
rect 3292 15048 3893 15076
rect 3292 15036 3298 15048
rect 3881 15045 3893 15048
rect 3927 15045 3939 15079
rect 3881 15039 3939 15045
rect 3694 14968 3700 15020
rect 3752 14968 3758 15020
rect 3970 14968 3976 15020
rect 4028 14968 4034 15020
rect 4062 14968 4068 15020
rect 4120 14968 4126 15020
rect 4706 14968 4712 15020
rect 4764 14968 4770 15020
rect 5828 15017 5856 15116
rect 6822 15104 6828 15116
rect 6880 15144 6886 15156
rect 7742 15144 7748 15156
rect 6880 15116 7748 15144
rect 6880 15104 6886 15116
rect 7742 15104 7748 15116
rect 7800 15104 7806 15156
rect 10226 15144 10232 15156
rect 8220 15116 10232 15144
rect 6362 15036 6368 15088
rect 6420 15076 6426 15088
rect 7193 15079 7251 15085
rect 7193 15076 7205 15079
rect 6420 15048 7205 15076
rect 6420 15036 6426 15048
rect 7193 15045 7205 15048
rect 7239 15045 7251 15079
rect 7193 15039 7251 15045
rect 8018 15036 8024 15088
rect 8076 15036 8082 15088
rect 5813 15011 5871 15017
rect 5813 14977 5825 15011
rect 5859 14977 5871 15011
rect 5813 14971 5871 14977
rect 5905 15011 5963 15017
rect 5905 14977 5917 15011
rect 5951 15008 5963 15011
rect 6638 15008 6644 15020
rect 5951 14980 6644 15008
rect 5951 14977 5963 14980
rect 5905 14971 5963 14977
rect 6638 14968 6644 14980
rect 6696 15008 6702 15020
rect 6825 15011 6883 15017
rect 6825 15008 6837 15011
rect 6696 14980 6837 15008
rect 6696 14968 6702 14980
rect 6825 14977 6837 14980
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 7834 14968 7840 15020
rect 7892 15008 7898 15020
rect 8220 15017 8248 15116
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 10318 15104 10324 15156
rect 10376 15144 10382 15156
rect 10413 15147 10471 15153
rect 10413 15144 10425 15147
rect 10376 15116 10425 15144
rect 10376 15104 10382 15116
rect 10413 15113 10425 15116
rect 10459 15113 10471 15147
rect 10413 15107 10471 15113
rect 10781 15147 10839 15153
rect 10781 15113 10793 15147
rect 10827 15144 10839 15147
rect 11422 15144 11428 15156
rect 10827 15116 11428 15144
rect 10827 15113 10839 15116
rect 10781 15107 10839 15113
rect 11422 15104 11428 15116
rect 11480 15104 11486 15156
rect 11514 15104 11520 15156
rect 11572 15144 11578 15156
rect 11701 15147 11759 15153
rect 11701 15144 11713 15147
rect 11572 15116 11713 15144
rect 11572 15104 11578 15116
rect 11701 15113 11713 15116
rect 11747 15113 11759 15147
rect 11701 15107 11759 15113
rect 11790 15104 11796 15156
rect 11848 15144 11854 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 11848 15116 13001 15144
rect 11848 15104 11854 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 14737 15147 14795 15153
rect 14737 15113 14749 15147
rect 14783 15144 14795 15147
rect 14826 15144 14832 15156
rect 14783 15116 14832 15144
rect 14783 15113 14795 15116
rect 14737 15107 14795 15113
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 16850 15144 16856 15156
rect 14936 15116 16856 15144
rect 9122 15076 9128 15088
rect 8312 15048 9128 15076
rect 8312 15017 8340 15048
rect 9122 15036 9128 15048
rect 9180 15036 9186 15088
rect 9309 15079 9367 15085
rect 9309 15045 9321 15079
rect 9355 15076 9367 15079
rect 12802 15076 12808 15088
rect 9355 15048 12808 15076
rect 9355 15045 9367 15048
rect 9309 15039 9367 15045
rect 12802 15036 12808 15048
rect 12860 15036 12866 15088
rect 14936 15076 14964 15116
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 19153 15079 19211 15085
rect 19153 15076 19165 15079
rect 14660 15048 14964 15076
rect 18616 15048 19165 15076
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 7892 14980 8217 15008
rect 7892 14968 7898 14980
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 8205 14971 8263 14977
rect 8297 15011 8355 15017
rect 8297 14977 8309 15011
rect 8343 14977 8355 15011
rect 8297 14971 8355 14977
rect 9033 15011 9091 15017
rect 9033 14977 9045 15011
rect 9079 15008 9091 15011
rect 9858 15008 9864 15020
rect 9079 14980 9864 15008
rect 9079 14977 9091 14980
rect 9033 14971 9091 14977
rect 9858 14968 9864 14980
rect 9916 14968 9922 15020
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 15008 10931 15011
rect 11790 15008 11796 15020
rect 10919 14980 11796 15008
rect 10919 14977 10931 14980
rect 10873 14971 10931 14977
rect 11790 14968 11796 14980
rect 11848 14968 11854 15020
rect 11882 14968 11888 15020
rect 11940 14968 11946 15020
rect 12250 14968 12256 15020
rect 12308 14968 12314 15020
rect 12449 15011 12507 15017
rect 12449 14977 12461 15011
rect 12495 15008 12507 15011
rect 12912 15008 13032 15014
rect 13265 15011 13323 15017
rect 13265 15008 13277 15011
rect 12495 14980 12756 15008
rect 12495 14977 12507 14980
rect 12449 14971 12507 14977
rect 2314 14900 2320 14952
rect 2372 14900 2378 14952
rect 3050 14900 3056 14952
rect 3108 14940 3114 14952
rect 3988 14940 4016 14968
rect 3108 14912 4016 14940
rect 3108 14900 3114 14912
rect 4982 14900 4988 14952
rect 5040 14900 5046 14952
rect 6454 14900 6460 14952
rect 6512 14940 6518 14952
rect 6733 14943 6791 14949
rect 6733 14940 6745 14943
rect 6512 14912 6745 14940
rect 6512 14900 6518 14912
rect 6733 14909 6745 14912
rect 6779 14940 6791 14943
rect 6914 14940 6920 14952
rect 6779 14912 6920 14940
rect 6779 14909 6791 14912
rect 6733 14903 6791 14909
rect 6914 14900 6920 14912
rect 6972 14900 6978 14952
rect 8938 14900 8944 14952
rect 8996 14900 9002 14952
rect 9401 14943 9459 14949
rect 9401 14909 9413 14943
rect 9447 14909 9459 14943
rect 9401 14903 9459 14909
rect 11057 14943 11115 14949
rect 11057 14909 11069 14943
rect 11103 14909 11115 14943
rect 11057 14903 11115 14909
rect 4798 14832 4804 14884
rect 4856 14872 4862 14884
rect 6549 14875 6607 14881
rect 6549 14872 6561 14875
rect 4856 14844 6561 14872
rect 4856 14832 4862 14844
rect 6549 14841 6561 14844
rect 6595 14841 6607 14875
rect 6549 14835 6607 14841
rect 8021 14875 8079 14881
rect 8021 14841 8033 14875
rect 8067 14872 8079 14875
rect 9214 14872 9220 14884
rect 8067 14844 9220 14872
rect 8067 14841 8079 14844
rect 8021 14835 8079 14841
rect 9214 14832 9220 14844
rect 9272 14872 9278 14884
rect 9416 14872 9444 14903
rect 9272 14844 9444 14872
rect 9272 14832 9278 14844
rect 1673 14807 1731 14813
rect 1673 14773 1685 14807
rect 1719 14804 1731 14807
rect 2038 14804 2044 14816
rect 1719 14776 2044 14804
rect 1719 14773 1731 14776
rect 1673 14767 1731 14773
rect 2038 14764 2044 14776
rect 2096 14764 2102 14816
rect 4246 14764 4252 14816
rect 4304 14764 4310 14816
rect 4890 14764 4896 14816
rect 4948 14764 4954 14816
rect 8757 14807 8815 14813
rect 8757 14773 8769 14807
rect 8803 14804 8815 14807
rect 8846 14804 8852 14816
rect 8803 14776 8852 14804
rect 8803 14773 8815 14776
rect 8757 14767 8815 14773
rect 8846 14764 8852 14776
rect 8904 14764 8910 14816
rect 11072 14804 11100 14903
rect 11238 14900 11244 14952
rect 11296 14940 11302 14952
rect 12069 14943 12127 14949
rect 12069 14940 12081 14943
rect 11296 14912 12081 14940
rect 11296 14900 11302 14912
rect 12069 14909 12081 14912
rect 12115 14909 12127 14943
rect 12069 14903 12127 14909
rect 12158 14900 12164 14952
rect 12216 14900 12222 14952
rect 11698 14832 11704 14884
rect 11756 14872 11762 14884
rect 12728 14872 12756 14980
rect 12912 14986 13277 15008
rect 12802 14900 12808 14952
rect 12860 14940 12866 14952
rect 12912 14940 12940 14986
rect 13004 14980 13277 14986
rect 13265 14977 13277 14980
rect 13311 14977 13323 15011
rect 13265 14971 13323 14977
rect 13630 14968 13636 15020
rect 13688 15008 13694 15020
rect 14660 15017 14688 15048
rect 18616 15020 18644 15048
rect 19153 15045 19165 15048
rect 19199 15045 19211 15079
rect 19153 15039 19211 15045
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 13688 14980 14657 15008
rect 13688 14968 13694 14980
rect 14645 14977 14657 14980
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 14826 14968 14832 15020
rect 14884 14968 14890 15020
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 15473 15011 15531 15017
rect 15473 15008 15485 15011
rect 15252 14980 15485 15008
rect 15252 14968 15258 14980
rect 15473 14977 15485 14980
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 15746 14968 15752 15020
rect 15804 14968 15810 15020
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 18325 15011 18383 15017
rect 18325 15008 18337 15011
rect 16816 14980 18337 15008
rect 16816 14968 16822 14980
rect 18325 14977 18337 14980
rect 18371 15008 18383 15011
rect 18598 15008 18604 15020
rect 18371 14980 18604 15008
rect 18371 14977 18383 14980
rect 18325 14971 18383 14977
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 18966 14968 18972 15020
rect 19024 14968 19030 15020
rect 19242 14968 19248 15020
rect 19300 14968 19306 15020
rect 12860 14912 12940 14940
rect 12989 14943 13047 14949
rect 12860 14900 12866 14912
rect 12989 14909 13001 14943
rect 13035 14940 13047 14943
rect 13078 14940 13084 14952
rect 13035 14912 13084 14940
rect 13035 14909 13047 14912
rect 12989 14903 13047 14909
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 15562 14900 15568 14952
rect 15620 14900 15626 14952
rect 15657 14943 15715 14949
rect 15657 14909 15669 14943
rect 15703 14909 15715 14943
rect 15657 14903 15715 14909
rect 15378 14872 15384 14884
rect 11756 14844 15384 14872
rect 11756 14832 11762 14844
rect 15378 14832 15384 14844
rect 15436 14872 15442 14884
rect 15672 14872 15700 14903
rect 17126 14900 17132 14952
rect 17184 14900 17190 14952
rect 17586 14900 17592 14952
rect 17644 14940 17650 14952
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 17644 14912 18061 14940
rect 17644 14900 17650 14912
rect 18049 14909 18061 14912
rect 18095 14909 18107 14943
rect 18049 14903 18107 14909
rect 18233 14943 18291 14949
rect 18233 14909 18245 14943
rect 18279 14940 18291 14943
rect 19260 14940 19288 14968
rect 18279 14912 19288 14940
rect 18279 14909 18291 14912
rect 18233 14903 18291 14909
rect 15436 14844 15700 14872
rect 15436 14832 15442 14844
rect 17402 14832 17408 14884
rect 17460 14832 17466 14884
rect 18874 14832 18880 14884
rect 18932 14872 18938 14884
rect 18969 14875 19027 14881
rect 18969 14872 18981 14875
rect 18932 14844 18981 14872
rect 18932 14832 18938 14844
rect 18969 14841 18981 14844
rect 19015 14841 19027 14875
rect 18969 14835 19027 14841
rect 12066 14804 12072 14816
rect 11072 14776 12072 14804
rect 12066 14764 12072 14776
rect 12124 14764 12130 14816
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 13078 14804 13084 14816
rect 12676 14776 13084 14804
rect 12676 14764 12682 14776
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 13170 14764 13176 14816
rect 13228 14764 13234 14816
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15654 14804 15660 14816
rect 15335 14776 15660 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 18046 14764 18052 14816
rect 18104 14804 18110 14816
rect 18141 14807 18199 14813
rect 18141 14804 18153 14807
rect 18104 14776 18153 14804
rect 18104 14764 18110 14776
rect 18141 14773 18153 14776
rect 18187 14773 18199 14807
rect 18141 14767 18199 14773
rect 1104 14714 20884 14736
rect 1104 14662 3422 14714
rect 3474 14662 3486 14714
rect 3538 14662 3550 14714
rect 3602 14662 3614 14714
rect 3666 14662 3678 14714
rect 3730 14662 8367 14714
rect 8419 14662 8431 14714
rect 8483 14662 8495 14714
rect 8547 14662 8559 14714
rect 8611 14662 8623 14714
rect 8675 14662 13312 14714
rect 13364 14662 13376 14714
rect 13428 14662 13440 14714
rect 13492 14662 13504 14714
rect 13556 14662 13568 14714
rect 13620 14662 18257 14714
rect 18309 14662 18321 14714
rect 18373 14662 18385 14714
rect 18437 14662 18449 14714
rect 18501 14662 18513 14714
rect 18565 14662 20884 14714
rect 1104 14640 20884 14662
rect 12345 14603 12403 14609
rect 12345 14569 12357 14603
rect 12391 14600 12403 14603
rect 13170 14600 13176 14612
rect 12391 14572 13176 14600
rect 12391 14569 12403 14572
rect 12345 14563 12403 14569
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 14366 14560 14372 14612
rect 14424 14600 14430 14612
rect 14461 14603 14519 14609
rect 14461 14600 14473 14603
rect 14424 14572 14473 14600
rect 14424 14560 14430 14572
rect 14461 14569 14473 14572
rect 14507 14600 14519 14603
rect 14507 14572 14780 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 12250 14492 12256 14544
rect 12308 14532 12314 14544
rect 14553 14535 14611 14541
rect 14553 14532 14565 14535
rect 12308 14504 14565 14532
rect 12308 14492 12314 14504
rect 14553 14501 14565 14504
rect 14599 14532 14611 14535
rect 14642 14532 14648 14544
rect 14599 14504 14648 14532
rect 14599 14501 14611 14504
rect 14553 14495 14611 14501
rect 14642 14492 14648 14504
rect 14700 14492 14706 14544
rect 14752 14532 14780 14572
rect 14826 14560 14832 14612
rect 14884 14600 14890 14612
rect 15565 14603 15623 14609
rect 15565 14600 15577 14603
rect 14884 14572 15577 14600
rect 14884 14560 14890 14572
rect 15565 14569 15577 14572
rect 15611 14569 15623 14603
rect 19242 14600 19248 14612
rect 15565 14563 15623 14569
rect 18340 14572 19248 14600
rect 14918 14532 14924 14544
rect 14752 14504 14924 14532
rect 14918 14492 14924 14504
rect 14976 14492 14982 14544
rect 18340 14541 18368 14572
rect 19242 14560 19248 14572
rect 19300 14600 19306 14612
rect 19429 14603 19487 14609
rect 19429 14600 19441 14603
rect 19300 14572 19441 14600
rect 19300 14560 19306 14572
rect 19429 14569 19441 14572
rect 19475 14569 19487 14603
rect 19429 14563 19487 14569
rect 18325 14535 18383 14541
rect 18325 14501 18337 14535
rect 18371 14501 18383 14535
rect 18325 14495 18383 14501
rect 8938 14424 8944 14476
rect 8996 14464 9002 14476
rect 8996 14436 9628 14464
rect 8996 14424 9002 14436
rect 9600 14408 9628 14436
rect 13722 14424 13728 14476
rect 13780 14464 13786 14476
rect 17497 14467 17555 14473
rect 17497 14464 17509 14467
rect 13780 14436 17509 14464
rect 13780 14424 13786 14436
rect 6454 14356 6460 14408
rect 6512 14396 6518 14408
rect 7837 14399 7895 14405
rect 7837 14396 7849 14399
rect 6512 14368 7849 14396
rect 6512 14356 6518 14368
rect 7837 14365 7849 14368
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 8110 14356 8116 14408
rect 8168 14356 8174 14408
rect 9214 14356 9220 14408
rect 9272 14405 9278 14408
rect 9272 14399 9308 14405
rect 9296 14365 9308 14399
rect 9272 14359 9308 14365
rect 9272 14356 9278 14359
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 9640 14368 9689 14396
rect 9640 14356 9646 14368
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 9677 14359 9735 14365
rect 9769 14399 9827 14405
rect 9769 14365 9781 14399
rect 9815 14396 9827 14399
rect 11698 14396 11704 14408
rect 9815 14368 11704 14396
rect 9815 14365 9827 14368
rect 9769 14359 9827 14365
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 11882 14356 11888 14408
rect 11940 14396 11946 14408
rect 12250 14396 12256 14408
rect 11940 14368 12256 14396
rect 11940 14356 11946 14368
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 12434 14356 12440 14408
rect 12492 14356 12498 14408
rect 12894 14356 12900 14408
rect 12952 14396 12958 14408
rect 13081 14399 13139 14405
rect 13081 14396 13093 14399
rect 12952 14368 13093 14396
rect 12952 14356 12958 14368
rect 13081 14365 13093 14368
rect 13127 14365 13139 14399
rect 13081 14359 13139 14365
rect 13354 14356 13360 14408
rect 13412 14356 13418 14408
rect 14274 14356 14280 14408
rect 14332 14356 14338 14408
rect 14660 14405 14688 14436
rect 17497 14433 17509 14436
rect 17543 14433 17555 14467
rect 18233 14467 18291 14473
rect 18233 14464 18245 14467
rect 17497 14427 17555 14433
rect 17604 14436 18245 14464
rect 17604 14408 17632 14436
rect 18233 14433 18245 14436
rect 18279 14433 18291 14467
rect 18598 14464 18604 14476
rect 18233 14427 18291 14433
rect 18432 14436 18604 14464
rect 14645 14399 14703 14405
rect 14645 14365 14657 14399
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14396 14795 14399
rect 14826 14396 14832 14408
rect 14783 14368 14832 14396
rect 14783 14365 14795 14368
rect 14737 14359 14795 14365
rect 14826 14356 14832 14368
rect 14884 14396 14890 14408
rect 15286 14396 15292 14408
rect 14884 14368 15292 14396
rect 14884 14356 14890 14368
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14365 15531 14399
rect 15473 14359 15531 14365
rect 15657 14399 15715 14405
rect 15657 14365 15669 14399
rect 15703 14396 15715 14399
rect 16574 14396 16580 14408
rect 15703 14368 16580 14396
rect 15703 14365 15715 14368
rect 15657 14359 15715 14365
rect 5718 14288 5724 14340
rect 5776 14328 5782 14340
rect 5776 14300 7052 14328
rect 5776 14288 5782 14300
rect 6914 14220 6920 14272
rect 6972 14220 6978 14272
rect 7024 14260 7052 14300
rect 7098 14288 7104 14340
rect 7156 14288 7162 14340
rect 7285 14331 7343 14337
rect 7285 14297 7297 14331
rect 7331 14328 7343 14331
rect 7745 14331 7803 14337
rect 7745 14328 7757 14331
rect 7331 14300 7757 14328
rect 7331 14297 7343 14300
rect 7285 14291 7343 14297
rect 7745 14297 7757 14300
rect 7791 14297 7803 14331
rect 7745 14291 7803 14297
rect 7300 14260 7328 14291
rect 11238 14288 11244 14340
rect 11296 14288 11302 14340
rect 14550 14288 14556 14340
rect 14608 14328 14614 14340
rect 15488 14328 15516 14359
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 14608 14300 16068 14328
rect 14608 14288 14614 14300
rect 7024 14232 7328 14260
rect 9125 14263 9183 14269
rect 9125 14229 9137 14263
rect 9171 14260 9183 14263
rect 9214 14260 9220 14272
rect 9171 14232 9220 14260
rect 9171 14229 9183 14232
rect 9125 14223 9183 14229
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 9306 14220 9312 14272
rect 9364 14220 9370 14272
rect 11149 14263 11207 14269
rect 11149 14229 11161 14263
rect 11195 14260 11207 14263
rect 11606 14260 11612 14272
rect 11195 14232 11612 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 12897 14263 12955 14269
rect 12897 14260 12909 14263
rect 11848 14232 12909 14260
rect 11848 14220 11854 14232
rect 12897 14229 12909 14232
rect 12943 14229 12955 14263
rect 12897 14223 12955 14229
rect 12986 14220 12992 14272
rect 13044 14260 13050 14272
rect 13265 14263 13323 14269
rect 13265 14260 13277 14263
rect 13044 14232 13277 14260
rect 13044 14220 13050 14232
rect 13265 14229 13277 14232
rect 13311 14229 13323 14263
rect 13265 14223 13323 14229
rect 15013 14263 15071 14269
rect 15013 14229 15025 14263
rect 15059 14260 15071 14263
rect 15470 14260 15476 14272
rect 15059 14232 15476 14260
rect 15059 14229 15071 14232
rect 15013 14223 15071 14229
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 16040 14260 16068 14300
rect 16114 14288 16120 14340
rect 16172 14328 16178 14340
rect 17420 14328 17448 14359
rect 17586 14356 17592 14408
rect 17644 14356 17650 14408
rect 18138 14356 18144 14408
rect 18196 14356 18202 14408
rect 18432 14405 18460 14436
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 19886 14424 19892 14476
rect 19944 14464 19950 14476
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 19944 14436 20085 14464
rect 19944 14424 19950 14436
rect 20073 14433 20085 14436
rect 20119 14433 20131 14467
rect 20073 14427 20131 14433
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14365 18475 14399
rect 19554 14399 19612 14405
rect 19554 14396 19566 14399
rect 18417 14359 18475 14365
rect 19306 14368 19566 14396
rect 19306 14328 19334 14368
rect 19554 14365 19566 14368
rect 19600 14365 19612 14399
rect 19554 14359 19612 14365
rect 19978 14356 19984 14408
rect 20036 14356 20042 14408
rect 16172 14300 17448 14328
rect 18064 14300 19334 14328
rect 16172 14288 16178 14300
rect 17402 14260 17408 14272
rect 16040 14232 17408 14260
rect 17402 14220 17408 14232
rect 17460 14260 17466 14272
rect 18064 14260 18092 14300
rect 17460 14232 18092 14260
rect 17460 14220 17466 14232
rect 18138 14220 18144 14272
rect 18196 14260 18202 14272
rect 18601 14263 18659 14269
rect 18601 14260 18613 14263
rect 18196 14232 18613 14260
rect 18196 14220 18202 14232
rect 18601 14229 18613 14232
rect 18647 14229 18659 14263
rect 18601 14223 18659 14229
rect 19610 14220 19616 14272
rect 19668 14220 19674 14272
rect 1104 14170 21043 14192
rect 1104 14118 5894 14170
rect 5946 14118 5958 14170
rect 6010 14118 6022 14170
rect 6074 14118 6086 14170
rect 6138 14118 6150 14170
rect 6202 14118 10839 14170
rect 10891 14118 10903 14170
rect 10955 14118 10967 14170
rect 11019 14118 11031 14170
rect 11083 14118 11095 14170
rect 11147 14118 15784 14170
rect 15836 14118 15848 14170
rect 15900 14118 15912 14170
rect 15964 14118 15976 14170
rect 16028 14118 16040 14170
rect 16092 14118 20729 14170
rect 20781 14118 20793 14170
rect 20845 14118 20857 14170
rect 20909 14118 20921 14170
rect 20973 14118 20985 14170
rect 21037 14118 21043 14170
rect 1104 14096 21043 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1762 14056 1768 14068
rect 1627 14028 1768 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 2038 14016 2044 14068
rect 2096 14016 2102 14068
rect 8573 14059 8631 14065
rect 8573 14025 8585 14059
rect 8619 14056 8631 14059
rect 9306 14056 9312 14068
rect 8619 14028 9312 14056
rect 8619 14025 8631 14028
rect 8573 14019 8631 14025
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 11882 14056 11888 14068
rect 9600 14028 11888 14056
rect 3605 13991 3663 13997
rect 3605 13957 3617 13991
rect 3651 13988 3663 13991
rect 4798 13988 4804 14000
rect 3651 13960 4804 13988
rect 3651 13957 3663 13960
rect 3605 13951 3663 13957
rect 4798 13948 4804 13960
rect 4856 13948 4862 14000
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13920 2007 13923
rect 2038 13920 2044 13932
rect 1995 13892 2044 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 2038 13880 2044 13892
rect 2096 13880 2102 13932
rect 3326 13880 3332 13932
rect 3384 13920 3390 13932
rect 3513 13923 3571 13929
rect 3513 13920 3525 13923
rect 3384 13892 3525 13920
rect 3384 13880 3390 13892
rect 3513 13889 3525 13892
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 3697 13923 3755 13929
rect 3697 13889 3709 13923
rect 3743 13889 3755 13923
rect 3697 13883 3755 13889
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13821 2283 13855
rect 2225 13815 2283 13821
rect 2240 13784 2268 13815
rect 2314 13812 2320 13864
rect 2372 13852 2378 13864
rect 2372 13824 2774 13852
rect 2372 13812 2378 13824
rect 2406 13784 2412 13796
rect 2240 13756 2412 13784
rect 2406 13744 2412 13756
rect 2464 13744 2470 13796
rect 2746 13784 2774 13824
rect 3712 13784 3740 13883
rect 3878 13880 3884 13932
rect 3936 13880 3942 13932
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 3786 13812 3792 13864
rect 3844 13852 3850 13864
rect 3988 13852 4016 13883
rect 3844 13824 4016 13852
rect 3844 13812 3850 13824
rect 5092 13784 5120 13883
rect 5258 13880 5264 13932
rect 5316 13880 5322 13932
rect 8389 13923 8447 13929
rect 8389 13889 8401 13923
rect 8435 13920 8447 13923
rect 8573 13923 8631 13929
rect 8435 13892 8524 13920
rect 8435 13889 8447 13892
rect 8389 13883 8447 13889
rect 5169 13855 5227 13861
rect 5169 13821 5181 13855
rect 5215 13852 5227 13855
rect 5350 13852 5356 13864
rect 5215 13824 5356 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 8496 13852 8524 13892
rect 8573 13889 8585 13923
rect 8619 13920 8631 13923
rect 9600 13920 9628 14028
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 12124 14028 12480 14056
rect 12124 14016 12130 14028
rect 9674 13948 9680 14000
rect 9732 13988 9738 14000
rect 10597 13991 10655 13997
rect 10597 13988 10609 13991
rect 9732 13960 10609 13988
rect 9732 13948 9738 13960
rect 10597 13957 10609 13960
rect 10643 13988 10655 13991
rect 10643 13960 12388 13988
rect 10643 13957 10655 13960
rect 10597 13951 10655 13957
rect 8619 13892 9628 13920
rect 10781 13923 10839 13929
rect 8619 13889 8631 13892
rect 8573 13883 8631 13889
rect 10781 13889 10793 13923
rect 10827 13920 10839 13923
rect 11606 13920 11612 13932
rect 10827 13892 11612 13920
rect 10827 13889 10839 13892
rect 10781 13883 10839 13889
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 11882 13920 11888 13932
rect 11716 13892 11888 13920
rect 8754 13852 8760 13864
rect 8496 13824 8760 13852
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 11330 13852 11336 13864
rect 11195 13824 11336 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 11422 13812 11428 13864
rect 11480 13852 11486 13864
rect 11716 13852 11744 13892
rect 11882 13880 11888 13892
rect 11940 13920 11946 13932
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 11940 13892 11989 13920
rect 11940 13880 11946 13892
rect 11977 13889 11989 13892
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 12066 13880 12072 13932
rect 12124 13880 12130 13932
rect 12360 13929 12388 13960
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13889 12403 13923
rect 12452 13920 12480 14028
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 12802 14056 12808 14068
rect 12584 14028 12808 14056
rect 12584 14016 12590 14028
rect 12802 14016 12808 14028
rect 12860 14056 12866 14068
rect 14458 14056 14464 14068
rect 12860 14028 14464 14056
rect 12860 14016 12866 14028
rect 14458 14016 14464 14028
rect 14516 14056 14522 14068
rect 14516 14028 14596 14056
rect 14516 14016 14522 14028
rect 12452 13892 12940 13920
rect 12345 13883 12403 13889
rect 11480 13824 11744 13852
rect 11480 13812 11486 13824
rect 11790 13812 11796 13864
rect 11848 13852 11854 13864
rect 12176 13852 12204 13883
rect 12802 13852 12808 13864
rect 11848 13824 12808 13852
rect 11848 13812 11854 13824
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 5442 13784 5448 13796
rect 2746 13756 5448 13784
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 9030 13744 9036 13796
rect 9088 13784 9094 13796
rect 12434 13784 12440 13796
rect 9088 13756 12440 13784
rect 9088 13744 9094 13756
rect 12434 13744 12440 13756
rect 12492 13744 12498 13796
rect 12912 13784 12940 13892
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 13173 13923 13231 13929
rect 13173 13920 13185 13923
rect 13044 13892 13185 13920
rect 13044 13880 13050 13892
rect 13173 13889 13185 13892
rect 13219 13889 13231 13923
rect 13173 13883 13231 13889
rect 13188 13852 13216 13883
rect 13354 13880 13360 13932
rect 13412 13920 13418 13932
rect 13722 13920 13728 13932
rect 13412 13892 13728 13920
rect 13412 13880 13418 13892
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 14568 13929 14596 14028
rect 14642 14016 14648 14068
rect 14700 14016 14706 14068
rect 15562 14016 15568 14068
rect 15620 14056 15626 14068
rect 15749 14059 15807 14065
rect 15749 14056 15761 14059
rect 15620 14028 15761 14056
rect 15620 14016 15626 14028
rect 15749 14025 15761 14028
rect 15795 14025 15807 14059
rect 15749 14019 15807 14025
rect 15948 14028 16252 14056
rect 15948 13988 15976 14028
rect 14752 13960 15976 13988
rect 16224 13988 16252 14028
rect 16224 13960 18000 13988
rect 14752 13929 14780 13960
rect 14553 13923 14611 13929
rect 14553 13889 14565 13923
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13889 15991 13923
rect 15933 13883 15991 13889
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 16071 13892 16160 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 14458 13852 14464 13864
rect 13188 13824 14464 13852
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 15948 13852 15976 13883
rect 15948 13824 16068 13852
rect 13630 13784 13636 13796
rect 12912 13756 13636 13784
rect 13630 13744 13636 13756
rect 13688 13744 13694 13796
rect 3326 13676 3332 13728
rect 3384 13676 3390 13728
rect 11698 13676 11704 13728
rect 11756 13676 11762 13728
rect 12986 13676 12992 13728
rect 13044 13716 13050 13728
rect 13265 13719 13323 13725
rect 13265 13716 13277 13719
rect 13044 13688 13277 13716
rect 13044 13676 13050 13688
rect 13265 13685 13277 13688
rect 13311 13685 13323 13719
rect 16040 13716 16068 13824
rect 16132 13784 16160 13892
rect 16206 13880 16212 13932
rect 16264 13880 16270 13932
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13920 16359 13923
rect 16482 13920 16488 13932
rect 16347 13892 16488 13920
rect 16347 13889 16359 13892
rect 16301 13883 16359 13889
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 17770 13880 17776 13932
rect 17828 13880 17834 13932
rect 17972 13920 18000 13960
rect 18046 13948 18052 14000
rect 18104 13948 18110 14000
rect 18138 13948 18144 14000
rect 18196 13948 18202 14000
rect 19886 13920 19892 13932
rect 17972 13892 19892 13920
rect 19886 13880 19892 13892
rect 19944 13880 19950 13932
rect 17678 13812 17684 13864
rect 17736 13812 17742 13864
rect 16850 13784 16856 13796
rect 16132 13756 16856 13784
rect 16850 13744 16856 13756
rect 16908 13784 16914 13796
rect 17586 13784 17592 13796
rect 16908 13756 17592 13784
rect 16908 13744 16914 13756
rect 17586 13744 17592 13756
rect 17644 13744 17650 13796
rect 16666 13716 16672 13728
rect 16040 13688 16672 13716
rect 13265 13679 13323 13685
rect 16666 13676 16672 13688
rect 16724 13676 16730 13728
rect 17494 13676 17500 13728
rect 17552 13676 17558 13728
rect 1104 13626 20884 13648
rect 1104 13574 3422 13626
rect 3474 13574 3486 13626
rect 3538 13574 3550 13626
rect 3602 13574 3614 13626
rect 3666 13574 3678 13626
rect 3730 13574 8367 13626
rect 8419 13574 8431 13626
rect 8483 13574 8495 13626
rect 8547 13574 8559 13626
rect 8611 13574 8623 13626
rect 8675 13574 13312 13626
rect 13364 13574 13376 13626
rect 13428 13574 13440 13626
rect 13492 13574 13504 13626
rect 13556 13574 13568 13626
rect 13620 13574 18257 13626
rect 18309 13574 18321 13626
rect 18373 13574 18385 13626
rect 18437 13574 18449 13626
rect 18501 13574 18513 13626
rect 18565 13574 20884 13626
rect 1104 13552 20884 13574
rect 3053 13515 3111 13521
rect 3053 13481 3065 13515
rect 3099 13512 3111 13515
rect 3878 13512 3884 13524
rect 3099 13484 3884 13512
rect 3099 13481 3111 13484
rect 3053 13475 3111 13481
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 13078 13472 13084 13524
rect 13136 13512 13142 13524
rect 16390 13512 16396 13524
rect 13136 13484 16396 13512
rect 13136 13472 13142 13484
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 16482 13472 16488 13524
rect 16540 13472 16546 13524
rect 17678 13472 17684 13524
rect 17736 13472 17742 13524
rect 19886 13472 19892 13524
rect 19944 13472 19950 13524
rect 6457 13447 6515 13453
rect 6457 13444 6469 13447
rect 2332 13416 6469 13444
rect 2332 13385 2360 13416
rect 6457 13413 6469 13416
rect 6503 13413 6515 13447
rect 6457 13407 6515 13413
rect 6564 13416 7052 13444
rect 2317 13379 2375 13385
rect 2317 13345 2329 13379
rect 2363 13345 2375 13379
rect 2317 13339 2375 13345
rect 2406 13336 2412 13388
rect 2464 13336 2470 13388
rect 4890 13336 4896 13388
rect 4948 13376 4954 13388
rect 5353 13379 5411 13385
rect 5353 13376 5365 13379
rect 4948 13348 5365 13376
rect 4948 13336 4954 13348
rect 5353 13345 5365 13348
rect 5399 13345 5411 13379
rect 5353 13339 5411 13345
rect 5442 13336 5448 13388
rect 5500 13376 5506 13388
rect 6564 13376 6592 13416
rect 6914 13376 6920 13388
rect 5500 13348 6592 13376
rect 6656 13348 6920 13376
rect 5500 13336 5506 13348
rect 3329 13311 3387 13317
rect 3329 13277 3341 13311
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 2314 13200 2320 13252
rect 2372 13240 2378 13252
rect 3053 13243 3111 13249
rect 3053 13240 3065 13243
rect 2372 13212 3065 13240
rect 2372 13200 2378 13212
rect 3053 13209 3065 13212
rect 3099 13209 3111 13243
rect 3344 13240 3372 13271
rect 3970 13268 3976 13320
rect 4028 13268 4034 13320
rect 4154 13268 4160 13320
rect 4212 13268 4218 13320
rect 6656 13317 6684 13348
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 7024 13376 7052 13416
rect 9674 13404 9680 13456
rect 9732 13404 9738 13456
rect 10689 13447 10747 13453
rect 10689 13413 10701 13447
rect 10735 13444 10747 13447
rect 12158 13444 12164 13456
rect 10735 13416 12164 13444
rect 10735 13413 10747 13416
rect 10689 13407 10747 13413
rect 12158 13404 12164 13416
rect 12216 13404 12222 13456
rect 13170 13404 13176 13456
rect 13228 13444 13234 13456
rect 13265 13447 13323 13453
rect 13265 13444 13277 13447
rect 13228 13416 13277 13444
rect 13228 13404 13234 13416
rect 13265 13413 13277 13416
rect 13311 13413 13323 13447
rect 18874 13444 18880 13456
rect 13265 13407 13323 13413
rect 15120 13416 18880 13444
rect 7374 13376 7380 13388
rect 7024 13348 7380 13376
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13277 6699 13311
rect 6641 13271 6699 13277
rect 6730 13268 6736 13320
rect 6788 13268 6794 13320
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13308 6883 13311
rect 7024 13308 7052 13348
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 8938 13336 8944 13388
rect 8996 13376 9002 13388
rect 9217 13379 9275 13385
rect 9217 13376 9229 13379
rect 8996 13348 9229 13376
rect 8996 13336 9002 13348
rect 9217 13345 9229 13348
rect 9263 13376 9275 13379
rect 9263 13348 11560 13376
rect 9263 13345 9275 13348
rect 9217 13339 9275 13345
rect 6871 13280 7052 13308
rect 7101 13311 7159 13317
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 7101 13277 7113 13311
rect 7147 13308 7159 13311
rect 8018 13308 8024 13320
rect 7147 13280 8024 13308
rect 7147 13277 7159 13280
rect 7101 13271 7159 13277
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 8294 13268 8300 13320
rect 8352 13308 8358 13320
rect 9306 13308 9312 13320
rect 8352 13280 9312 13308
rect 8352 13268 8358 13280
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 10336 13317 10364 13348
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13277 10379 13311
rect 10321 13271 10379 13277
rect 10475 13311 10533 13317
rect 10475 13277 10487 13311
rect 10521 13308 10533 13311
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 10521 13280 11161 13308
rect 10521 13277 10533 13280
rect 10475 13271 10533 13277
rect 11149 13277 11161 13280
rect 11195 13308 11207 13311
rect 11422 13308 11428 13320
rect 11195 13280 11428 13308
rect 11195 13277 11207 13280
rect 11149 13271 11207 13277
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 11532 13308 11560 13348
rect 11606 13336 11612 13388
rect 11664 13376 11670 13388
rect 15120 13376 15148 13416
rect 18874 13404 18880 13416
rect 18932 13404 18938 13456
rect 17494 13376 17500 13388
rect 11664 13348 15148 13376
rect 15212 13348 17500 13376
rect 11664 13336 11670 13348
rect 11701 13311 11759 13317
rect 11701 13308 11713 13311
rect 11532 13280 11713 13308
rect 11701 13277 11713 13280
rect 11747 13308 11759 13311
rect 11790 13308 11796 13320
rect 11747 13280 11796 13308
rect 11747 13277 11759 13280
rect 11701 13271 11759 13277
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 12986 13268 12992 13320
rect 13044 13268 13050 13320
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13308 13139 13311
rect 13630 13308 13636 13320
rect 13127 13280 13636 13308
rect 13127 13277 13139 13280
rect 13081 13271 13139 13277
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 15212 13317 15240 13348
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 17957 13379 18015 13385
rect 17957 13376 17969 13379
rect 17604 13348 17969 13376
rect 15197 13311 15255 13317
rect 15197 13277 15209 13311
rect 15243 13277 15255 13311
rect 15197 13271 15255 13277
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 15565 13311 15623 13317
rect 15565 13308 15577 13311
rect 15528 13280 15577 13308
rect 15528 13268 15534 13280
rect 15565 13277 15577 13280
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 16298 13268 16304 13320
rect 16356 13268 16362 13320
rect 16574 13268 16580 13320
rect 16632 13268 16638 13320
rect 17034 13268 17040 13320
rect 17092 13308 17098 13320
rect 17604 13308 17632 13348
rect 17957 13345 17969 13348
rect 18003 13345 18015 13379
rect 17957 13339 18015 13345
rect 18138 13336 18144 13388
rect 18196 13336 18202 13388
rect 17092 13280 17632 13308
rect 17092 13268 17098 13280
rect 17678 13268 17684 13320
rect 17736 13308 17742 13320
rect 17865 13311 17923 13317
rect 17865 13308 17877 13311
rect 17736 13280 17877 13308
rect 17736 13268 17742 13280
rect 17865 13277 17877 13280
rect 17911 13277 17923 13311
rect 17865 13271 17923 13277
rect 18046 13268 18052 13320
rect 18104 13268 18110 13320
rect 19702 13268 19708 13320
rect 19760 13308 19766 13320
rect 19981 13311 20039 13317
rect 19981 13308 19993 13311
rect 19760 13280 19993 13308
rect 19760 13268 19766 13280
rect 19981 13277 19993 13280
rect 20027 13277 20039 13311
rect 19981 13271 20039 13277
rect 4065 13243 4123 13249
rect 4065 13240 4077 13243
rect 3344 13212 4077 13240
rect 3053 13203 3111 13209
rect 4065 13209 4077 13212
rect 4111 13209 4123 13243
rect 4065 13203 4123 13209
rect 4264 13212 6776 13240
rect 1670 13132 1676 13184
rect 1728 13172 1734 13184
rect 1857 13175 1915 13181
rect 1857 13172 1869 13175
rect 1728 13144 1869 13172
rect 1728 13132 1734 13144
rect 1857 13141 1869 13144
rect 1903 13141 1915 13175
rect 1857 13135 1915 13141
rect 2222 13132 2228 13184
rect 2280 13132 2286 13184
rect 3142 13132 3148 13184
rect 3200 13172 3206 13184
rect 3237 13175 3295 13181
rect 3237 13172 3249 13175
rect 3200 13144 3249 13172
rect 3200 13132 3206 13144
rect 3237 13141 3249 13144
rect 3283 13172 3295 13175
rect 4264 13172 4292 13212
rect 6748 13184 6776 13212
rect 6914 13200 6920 13252
rect 6972 13249 6978 13252
rect 6972 13243 7001 13249
rect 6989 13209 7001 13243
rect 6972 13203 7001 13209
rect 6972 13200 6978 13203
rect 11514 13200 11520 13252
rect 11572 13240 11578 13252
rect 12250 13240 12256 13252
rect 11572 13212 12256 13240
rect 11572 13200 11578 13212
rect 12250 13200 12256 13212
rect 12308 13240 12314 13252
rect 13265 13243 13323 13249
rect 13265 13240 13277 13243
rect 12308 13212 13277 13240
rect 12308 13200 12314 13212
rect 13265 13209 13277 13212
rect 13311 13240 13323 13243
rect 13311 13212 15240 13240
rect 13311 13209 13323 13212
rect 13265 13203 13323 13209
rect 3283 13144 4292 13172
rect 4893 13175 4951 13181
rect 3283 13141 3295 13144
rect 3237 13135 3295 13141
rect 4893 13141 4905 13175
rect 4939 13172 4951 13175
rect 5074 13172 5080 13184
rect 4939 13144 5080 13172
rect 4939 13141 4951 13144
rect 4893 13135 4951 13141
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 5261 13175 5319 13181
rect 5261 13141 5273 13175
rect 5307 13172 5319 13175
rect 5810 13172 5816 13184
rect 5307 13144 5816 13172
rect 5307 13141 5319 13144
rect 5261 13135 5319 13141
rect 5810 13132 5816 13144
rect 5868 13172 5874 13184
rect 6270 13172 6276 13184
rect 5868 13144 6276 13172
rect 5868 13132 5874 13144
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 6730 13132 6736 13184
rect 6788 13132 6794 13184
rect 11330 13132 11336 13184
rect 11388 13172 11394 13184
rect 12894 13172 12900 13184
rect 11388 13144 12900 13172
rect 11388 13132 11394 13144
rect 12894 13132 12900 13144
rect 12952 13132 12958 13184
rect 14182 13132 14188 13184
rect 14240 13172 14246 13184
rect 15013 13175 15071 13181
rect 15013 13172 15025 13175
rect 14240 13144 15025 13172
rect 14240 13132 14246 13144
rect 15013 13141 15025 13144
rect 15059 13141 15071 13175
rect 15212 13172 15240 13212
rect 15286 13200 15292 13252
rect 15344 13200 15350 13252
rect 15381 13243 15439 13249
rect 15381 13209 15393 13243
rect 15427 13240 15439 13243
rect 16592 13240 16620 13268
rect 19610 13240 19616 13252
rect 15427 13212 16068 13240
rect 16592 13212 19616 13240
rect 15427 13209 15439 13212
rect 15381 13203 15439 13209
rect 15654 13172 15660 13184
rect 15212 13144 15660 13172
rect 15013 13135 15071 13141
rect 15654 13132 15660 13144
rect 15712 13172 15718 13184
rect 15930 13172 15936 13184
rect 15712 13144 15936 13172
rect 15712 13132 15718 13144
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 16040 13181 16068 13212
rect 19610 13200 19616 13212
rect 19668 13200 19674 13252
rect 16025 13175 16083 13181
rect 16025 13141 16037 13175
rect 16071 13141 16083 13175
rect 16025 13135 16083 13141
rect 1104 13082 21043 13104
rect 1104 13030 5894 13082
rect 5946 13030 5958 13082
rect 6010 13030 6022 13082
rect 6074 13030 6086 13082
rect 6138 13030 6150 13082
rect 6202 13030 10839 13082
rect 10891 13030 10903 13082
rect 10955 13030 10967 13082
rect 11019 13030 11031 13082
rect 11083 13030 11095 13082
rect 11147 13030 15784 13082
rect 15836 13030 15848 13082
rect 15900 13030 15912 13082
rect 15964 13030 15976 13082
rect 16028 13030 16040 13082
rect 16092 13030 20729 13082
rect 20781 13030 20793 13082
rect 20845 13030 20857 13082
rect 20909 13030 20921 13082
rect 20973 13030 20985 13082
rect 21037 13030 21043 13082
rect 1104 13008 21043 13030
rect 2133 12971 2191 12977
rect 2133 12937 2145 12971
rect 2179 12968 2191 12971
rect 3142 12968 3148 12980
rect 2179 12940 3148 12968
rect 2179 12937 2191 12940
rect 2133 12931 2191 12937
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 5074 12928 5080 12980
rect 5132 12928 5138 12980
rect 8481 12971 8539 12977
rect 8481 12937 8493 12971
rect 8527 12968 8539 12971
rect 8754 12968 8760 12980
rect 8527 12940 8760 12968
rect 8527 12937 8539 12940
rect 8481 12931 8539 12937
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9122 12968 9128 12980
rect 8864 12940 9128 12968
rect 1949 12903 2007 12909
rect 1949 12869 1961 12903
rect 1995 12900 2007 12903
rect 2222 12900 2228 12912
rect 1995 12872 2228 12900
rect 1995 12869 2007 12872
rect 1949 12863 2007 12869
rect 2222 12860 2228 12872
rect 2280 12900 2286 12912
rect 2774 12900 2780 12912
rect 2280 12872 2780 12900
rect 2280 12860 2286 12872
rect 2774 12860 2780 12872
rect 2832 12900 2838 12912
rect 3970 12900 3976 12912
rect 2832 12872 3976 12900
rect 2832 12860 2838 12872
rect 3970 12860 3976 12872
rect 4028 12860 4034 12912
rect 4798 12860 4804 12912
rect 4856 12900 4862 12912
rect 4985 12903 5043 12909
rect 4985 12900 4997 12903
rect 4856 12872 4997 12900
rect 4856 12860 4862 12872
rect 4985 12869 4997 12872
rect 5031 12900 5043 12903
rect 5031 12872 6960 12900
rect 5031 12869 5043 12872
rect 4985 12863 5043 12869
rect 1765 12835 1823 12841
rect 1765 12801 1777 12835
rect 1811 12832 1823 12835
rect 2038 12832 2044 12844
rect 1811 12804 2044 12832
rect 1811 12801 1823 12804
rect 1765 12795 1823 12801
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 2682 12792 2688 12844
rect 2740 12792 2746 12844
rect 4154 12832 4160 12844
rect 3160 12804 4160 12832
rect 2056 12764 2084 12792
rect 3160 12764 3188 12804
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6932 12841 6960 12872
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6328 12804 6561 12832
rect 6328 12792 6334 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 6917 12835 6975 12841
rect 6917 12801 6929 12835
rect 6963 12801 6975 12835
rect 6917 12795 6975 12801
rect 7282 12792 7288 12844
rect 7340 12792 7346 12844
rect 8018 12792 8024 12844
rect 8076 12792 8082 12844
rect 8757 12835 8815 12841
rect 8757 12801 8769 12835
rect 8803 12833 8815 12835
rect 8864 12833 8892 12940
rect 9122 12928 9128 12940
rect 9180 12968 9186 12980
rect 12710 12968 12716 12980
rect 9180 12940 12716 12968
rect 9180 12928 9186 12940
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 13004 12940 16252 12968
rect 9030 12860 9036 12912
rect 9088 12860 9094 12912
rect 12434 12860 12440 12912
rect 12492 12900 12498 12912
rect 13004 12900 13032 12940
rect 12492 12872 13032 12900
rect 12492 12860 12498 12872
rect 13078 12860 13084 12912
rect 13136 12900 13142 12912
rect 13449 12903 13507 12909
rect 13449 12900 13461 12903
rect 13136 12872 13461 12900
rect 13136 12860 13142 12872
rect 13449 12869 13461 12872
rect 13495 12869 13507 12903
rect 13449 12863 13507 12869
rect 14090 12860 14096 12912
rect 14148 12900 14154 12912
rect 15286 12900 15292 12912
rect 14148 12872 15292 12900
rect 14148 12860 14154 12872
rect 15286 12860 15292 12872
rect 15344 12860 15350 12912
rect 8803 12805 8892 12833
rect 8803 12801 8815 12805
rect 8757 12795 8815 12801
rect 9306 12792 9312 12844
rect 9364 12832 9370 12844
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 9364 12804 10609 12832
rect 9364 12792 9370 12804
rect 10597 12801 10609 12804
rect 10643 12832 10655 12835
rect 10778 12832 10784 12844
rect 10643 12804 10784 12832
rect 10643 12801 10655 12804
rect 10597 12795 10655 12801
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 12986 12832 12992 12844
rect 10919 12804 12992 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 2056 12736 3188 12764
rect 3237 12767 3295 12773
rect 3237 12733 3249 12767
rect 3283 12764 3295 12767
rect 3786 12764 3792 12776
rect 3283 12736 3792 12764
rect 3283 12733 3295 12736
rect 3237 12727 3295 12733
rect 3050 12656 3056 12708
rect 3108 12696 3114 12708
rect 3252 12696 3280 12727
rect 3786 12724 3792 12736
rect 3844 12724 3850 12776
rect 5166 12724 5172 12776
rect 5224 12724 5230 12776
rect 7374 12724 7380 12776
rect 7432 12724 7438 12776
rect 3108 12668 3280 12696
rect 8036 12696 8064 12792
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 8665 12767 8723 12773
rect 8665 12764 8677 12767
rect 8352 12736 8677 12764
rect 8352 12724 8358 12736
rect 8665 12733 8677 12736
rect 8711 12733 8723 12767
rect 8665 12727 8723 12733
rect 9122 12724 9128 12776
rect 9180 12724 9186 12776
rect 9232 12736 12434 12764
rect 9232 12696 9260 12736
rect 8036 12668 9260 12696
rect 10781 12699 10839 12705
rect 3108 12656 3114 12668
rect 10781 12665 10793 12699
rect 10827 12696 10839 12699
rect 11330 12696 11336 12708
rect 10827 12668 11336 12696
rect 10827 12665 10839 12668
rect 10781 12659 10839 12665
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 12406 12696 12434 12736
rect 12802 12724 12808 12776
rect 12860 12764 12866 12776
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 12860 12736 13093 12764
rect 12860 12724 12866 12736
rect 13081 12733 13093 12736
rect 13127 12733 13139 12767
rect 15102 12764 15108 12776
rect 13081 12727 13139 12733
rect 13372 12736 15108 12764
rect 13372 12696 13400 12736
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 16224 12764 16252 12940
rect 16298 12928 16304 12980
rect 16356 12968 16362 12980
rect 16853 12971 16911 12977
rect 16853 12968 16865 12971
rect 16356 12940 16865 12968
rect 16356 12928 16362 12940
rect 16853 12937 16865 12940
rect 16899 12937 16911 12971
rect 16853 12931 16911 12937
rect 17678 12928 17684 12980
rect 17736 12968 17742 12980
rect 18141 12971 18199 12977
rect 18141 12968 18153 12971
rect 17736 12940 18153 12968
rect 17736 12928 17742 12940
rect 18141 12937 18153 12940
rect 18187 12937 18199 12971
rect 18141 12931 18199 12937
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 19242 12968 19248 12980
rect 18748 12940 19248 12968
rect 18748 12928 18754 12940
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 19797 12971 19855 12977
rect 19797 12937 19809 12971
rect 19843 12937 19855 12971
rect 19797 12931 19855 12937
rect 16390 12860 16396 12912
rect 16448 12900 16454 12912
rect 17034 12909 17040 12912
rect 17005 12903 17040 12909
rect 17005 12900 17017 12903
rect 16448 12872 17017 12900
rect 16448 12860 16454 12872
rect 17005 12869 17017 12872
rect 17005 12863 17040 12869
rect 17034 12860 17040 12863
rect 17092 12860 17098 12912
rect 17126 12860 17132 12912
rect 17184 12900 17190 12912
rect 17221 12903 17279 12909
rect 17221 12900 17233 12903
rect 17184 12872 17233 12900
rect 17184 12860 17190 12872
rect 17221 12869 17233 12872
rect 17267 12869 17279 12903
rect 17221 12863 17279 12869
rect 18046 12860 18052 12912
rect 18104 12900 18110 12912
rect 19061 12903 19119 12909
rect 19061 12900 19073 12903
rect 18104 12872 19073 12900
rect 18104 12860 18110 12872
rect 19061 12869 19073 12872
rect 19107 12900 19119 12903
rect 19812 12900 19840 12931
rect 19107 12872 19840 12900
rect 19107 12869 19119 12872
rect 19061 12863 19119 12869
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 17862 12832 17868 12844
rect 17368 12804 17868 12832
rect 17368 12792 17374 12804
rect 17862 12792 17868 12804
rect 17920 12832 17926 12844
rect 18233 12835 18291 12841
rect 18233 12832 18245 12835
rect 17920 12804 18245 12832
rect 17920 12792 17926 12804
rect 18233 12801 18245 12804
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12832 18475 12835
rect 18598 12832 18604 12844
rect 18463 12804 18604 12832
rect 18463 12801 18475 12804
rect 18417 12795 18475 12801
rect 18598 12792 18604 12804
rect 18656 12832 18662 12844
rect 18969 12835 19027 12841
rect 18969 12832 18981 12835
rect 18656 12804 18981 12832
rect 18656 12792 18662 12804
rect 18969 12801 18981 12804
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 19242 12792 19248 12844
rect 19300 12792 19306 12844
rect 19702 12792 19708 12844
rect 19760 12832 19766 12844
rect 19981 12835 20039 12841
rect 19981 12832 19993 12835
rect 19760 12804 19993 12832
rect 19760 12792 19766 12804
rect 19981 12801 19993 12804
rect 20027 12801 20039 12835
rect 20159 12835 20217 12841
rect 20159 12832 20171 12835
rect 19981 12795 20039 12801
rect 20088 12804 20171 12832
rect 19334 12764 19340 12776
rect 16224 12736 19340 12764
rect 19334 12724 19340 12736
rect 19392 12764 19398 12776
rect 20088 12764 20116 12804
rect 20159 12801 20171 12804
rect 20205 12801 20217 12835
rect 20159 12795 20217 12801
rect 19392 12736 20116 12764
rect 19392 12724 19398 12736
rect 15286 12696 15292 12708
rect 12406 12668 13400 12696
rect 13464 12668 15292 12696
rect 4614 12588 4620 12640
rect 4672 12588 4678 12640
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 8110 12628 8116 12640
rect 7984 12600 8116 12628
rect 7984 12588 7990 12600
rect 8110 12588 8116 12600
rect 8168 12588 8174 12640
rect 10502 12588 10508 12640
rect 10560 12628 10566 12640
rect 10689 12631 10747 12637
rect 10689 12628 10701 12631
rect 10560 12600 10701 12628
rect 10560 12588 10566 12600
rect 10689 12597 10701 12600
rect 10735 12597 10747 12631
rect 10689 12591 10747 12597
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 12802 12628 12808 12640
rect 12584 12600 12808 12628
rect 12584 12588 12590 12600
rect 12802 12588 12808 12600
rect 12860 12588 12866 12640
rect 13464 12637 13492 12668
rect 15286 12656 15292 12668
rect 15344 12696 15350 12708
rect 15746 12696 15752 12708
rect 15344 12668 15752 12696
rect 15344 12656 15350 12668
rect 15746 12656 15752 12668
rect 15804 12656 15810 12708
rect 18966 12656 18972 12708
rect 19024 12696 19030 12708
rect 19245 12699 19303 12705
rect 19245 12696 19257 12699
rect 19024 12668 19257 12696
rect 19024 12656 19030 12668
rect 19245 12665 19257 12668
rect 19291 12665 19303 12699
rect 19245 12659 19303 12665
rect 13449 12631 13507 12637
rect 13449 12597 13461 12631
rect 13495 12597 13507 12631
rect 13449 12591 13507 12597
rect 13630 12588 13636 12640
rect 13688 12588 13694 12640
rect 17034 12588 17040 12640
rect 17092 12588 17098 12640
rect 20070 12588 20076 12640
rect 20128 12588 20134 12640
rect 1104 12538 20884 12560
rect 1104 12486 3422 12538
rect 3474 12486 3486 12538
rect 3538 12486 3550 12538
rect 3602 12486 3614 12538
rect 3666 12486 3678 12538
rect 3730 12486 8367 12538
rect 8419 12486 8431 12538
rect 8483 12486 8495 12538
rect 8547 12486 8559 12538
rect 8611 12486 8623 12538
rect 8675 12486 13312 12538
rect 13364 12486 13376 12538
rect 13428 12486 13440 12538
rect 13492 12486 13504 12538
rect 13556 12486 13568 12538
rect 13620 12486 18257 12538
rect 18309 12486 18321 12538
rect 18373 12486 18385 12538
rect 18437 12486 18449 12538
rect 18501 12486 18513 12538
rect 18565 12486 20884 12538
rect 1104 12464 20884 12486
rect 6730 12384 6736 12436
rect 6788 12384 6794 12436
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 7834 12424 7840 12436
rect 7156 12396 7840 12424
rect 7156 12384 7162 12396
rect 7834 12384 7840 12396
rect 7892 12424 7898 12436
rect 9122 12424 9128 12436
rect 7892 12396 9128 12424
rect 7892 12384 7898 12396
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 11238 12384 11244 12436
rect 11296 12424 11302 12436
rect 12526 12424 12532 12436
rect 11296 12396 12532 12424
rect 11296 12384 11302 12396
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 13541 12427 13599 12433
rect 13541 12393 13553 12427
rect 13587 12424 13599 12427
rect 13630 12424 13636 12436
rect 13587 12396 13636 12424
rect 13587 12393 13599 12396
rect 13541 12387 13599 12393
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 14366 12384 14372 12436
rect 14424 12424 14430 12436
rect 15010 12424 15016 12436
rect 14424 12396 15016 12424
rect 14424 12384 14430 12396
rect 15010 12384 15016 12396
rect 15068 12424 15074 12436
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 15068 12396 15301 12424
rect 15068 12384 15074 12396
rect 15289 12393 15301 12396
rect 15335 12393 15347 12427
rect 15289 12387 15347 12393
rect 15746 12384 15752 12436
rect 15804 12424 15810 12436
rect 17310 12424 17316 12436
rect 15804 12396 17316 12424
rect 15804 12384 15810 12396
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 17681 12427 17739 12433
rect 17681 12393 17693 12427
rect 17727 12424 17739 12427
rect 17770 12424 17776 12436
rect 17727 12396 17776 12424
rect 17727 12393 17739 12396
rect 17681 12387 17739 12393
rect 17770 12384 17776 12396
rect 17828 12384 17834 12436
rect 2314 12316 2320 12368
rect 2372 12356 2378 12368
rect 2372 12328 4936 12356
rect 2372 12316 2378 12328
rect 4246 12248 4252 12300
rect 4304 12288 4310 12300
rect 4908 12297 4936 12328
rect 12710 12316 12716 12368
rect 12768 12356 12774 12368
rect 14277 12359 14335 12365
rect 14277 12356 14289 12359
rect 12768 12328 14289 12356
rect 12768 12316 12774 12328
rect 14277 12325 14289 12328
rect 14323 12325 14335 12359
rect 17328 12356 17356 12384
rect 19978 12356 19984 12368
rect 17328 12328 19984 12356
rect 14277 12319 14335 12325
rect 4801 12291 4859 12297
rect 4801 12288 4813 12291
rect 4304 12260 4813 12288
rect 4304 12248 4310 12260
rect 4801 12257 4813 12260
rect 4847 12257 4859 12291
rect 4801 12251 4859 12257
rect 4893 12291 4951 12297
rect 4893 12257 4905 12291
rect 4939 12257 4951 12291
rect 4893 12251 4951 12257
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12288 11299 12291
rect 11514 12288 11520 12300
rect 11287 12260 11520 12288
rect 11287 12257 11299 12260
rect 11241 12251 11299 12257
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 14734 12248 14740 12300
rect 14792 12288 14798 12300
rect 16574 12288 16580 12300
rect 14792 12260 16580 12288
rect 14792 12248 14798 12260
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 18690 12288 18696 12300
rect 17144 12260 18000 12288
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12220 2743 12223
rect 3050 12220 3056 12232
rect 2731 12192 3056 12220
rect 2731 12189 2743 12192
rect 2685 12183 2743 12189
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 6365 12223 6423 12229
rect 6365 12220 6377 12223
rect 4120 12192 6377 12220
rect 4120 12180 4126 12192
rect 6365 12189 6377 12192
rect 6411 12189 6423 12223
rect 6365 12183 6423 12189
rect 6730 12180 6736 12232
rect 6788 12180 6794 12232
rect 6914 12180 6920 12232
rect 6972 12180 6978 12232
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 10873 12223 10931 12229
rect 10873 12220 10885 12223
rect 10468 12192 10885 12220
rect 10468 12180 10474 12192
rect 10873 12189 10885 12192
rect 10919 12189 10931 12223
rect 10873 12183 10931 12189
rect 11330 12180 11336 12232
rect 11388 12180 11394 12232
rect 12066 12180 12072 12232
rect 12124 12180 12130 12232
rect 13170 12180 13176 12232
rect 13228 12220 13234 12232
rect 13357 12223 13415 12229
rect 13357 12220 13369 12223
rect 13228 12192 13369 12220
rect 13228 12180 13234 12192
rect 13357 12189 13369 12192
rect 13403 12189 13415 12223
rect 13357 12183 13415 12189
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 14090 12220 14096 12232
rect 13587 12192 14096 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 14090 12180 14096 12192
rect 14148 12220 14154 12232
rect 14274 12220 14280 12232
rect 14148 12192 14280 12220
rect 14148 12180 14154 12192
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14458 12180 14464 12232
rect 14516 12180 14522 12232
rect 14550 12180 14556 12232
rect 14608 12220 14614 12232
rect 14829 12223 14887 12229
rect 14608 12192 14653 12220
rect 14608 12180 14614 12192
rect 14829 12189 14841 12223
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 2130 12112 2136 12164
rect 2188 12152 2194 12164
rect 2406 12152 2412 12164
rect 2188 12124 2412 12152
rect 2188 12112 2194 12124
rect 2406 12112 2412 12124
rect 2464 12152 2470 12164
rect 2869 12155 2927 12161
rect 2869 12152 2881 12155
rect 2464 12124 2881 12152
rect 2464 12112 2470 12124
rect 2869 12121 2881 12124
rect 2915 12152 2927 12155
rect 4522 12152 4528 12164
rect 2915 12124 4528 12152
rect 2915 12121 2927 12124
rect 2869 12115 2927 12121
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 10778 12112 10784 12164
rect 10836 12152 10842 12164
rect 10965 12155 11023 12161
rect 10965 12152 10977 12155
rect 10836 12124 10977 12152
rect 10836 12112 10842 12124
rect 10965 12121 10977 12124
rect 11011 12121 11023 12155
rect 10965 12115 11023 12121
rect 14642 12112 14648 12164
rect 14700 12152 14706 12164
rect 14844 12152 14872 12183
rect 15286 12180 15292 12232
rect 15344 12180 15350 12232
rect 15470 12180 15476 12232
rect 15528 12180 15534 12232
rect 17144 12229 17172 12260
rect 17972 12232 18000 12260
rect 18156 12260 18696 12288
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 15580 12192 17141 12220
rect 15580 12152 15608 12192
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 17221 12223 17279 12229
rect 17221 12189 17233 12223
rect 17267 12220 17279 12223
rect 17310 12220 17316 12232
rect 17267 12192 17316 12220
rect 17267 12189 17279 12192
rect 17221 12183 17279 12189
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17954 12180 17960 12232
rect 18012 12180 18018 12232
rect 18156 12229 18184 12260
rect 18690 12248 18696 12260
rect 18748 12248 18754 12300
rect 19720 12297 19748 12328
rect 19978 12316 19984 12328
rect 20036 12316 20042 12368
rect 19705 12291 19763 12297
rect 19705 12257 19717 12291
rect 19751 12257 19763 12291
rect 19705 12251 19763 12257
rect 18049 12223 18107 12229
rect 18049 12189 18061 12223
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 18141 12223 18199 12229
rect 18141 12189 18153 12223
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 18064 12152 18092 12183
rect 18230 12180 18236 12232
rect 18288 12220 18294 12232
rect 18325 12223 18383 12229
rect 18325 12220 18337 12223
rect 18288 12192 18337 12220
rect 18288 12180 18294 12192
rect 18325 12189 18337 12192
rect 18371 12220 18383 12223
rect 18598 12220 18604 12232
rect 18371 12192 18604 12220
rect 18371 12189 18383 12192
rect 18325 12183 18383 12189
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 19058 12180 19064 12232
rect 19116 12220 19122 12232
rect 20070 12220 20076 12232
rect 19116 12192 20076 12220
rect 19116 12180 19122 12192
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 14700 12124 15608 12152
rect 17052 12124 18092 12152
rect 14700 12112 14706 12124
rect 4341 12087 4399 12093
rect 4341 12053 4353 12087
rect 4387 12084 4399 12087
rect 4430 12084 4436 12096
rect 4387 12056 4436 12084
rect 4387 12053 4399 12056
rect 4341 12047 4399 12053
rect 4430 12044 4436 12056
rect 4488 12044 4494 12096
rect 4709 12087 4767 12093
rect 4709 12053 4721 12087
rect 4755 12084 4767 12087
rect 4798 12084 4804 12096
rect 4755 12056 4804 12084
rect 4755 12053 4767 12056
rect 4709 12047 4767 12053
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 7282 12084 7288 12096
rect 6595 12056 7288 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 10594 12044 10600 12096
rect 10652 12044 10658 12096
rect 11057 12087 11115 12093
rect 11057 12053 11069 12087
rect 11103 12084 11115 12087
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11103 12056 11989 12084
rect 11103 12053 11115 12056
rect 11057 12047 11115 12053
rect 11977 12053 11989 12056
rect 12023 12084 12035 12087
rect 13170 12084 13176 12096
rect 12023 12056 13176 12084
rect 12023 12053 12035 12056
rect 11977 12047 12035 12053
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 13725 12087 13783 12093
rect 13725 12053 13737 12087
rect 13771 12084 13783 12087
rect 13998 12084 14004 12096
rect 13771 12056 14004 12084
rect 13771 12053 13783 12056
rect 13725 12047 13783 12053
rect 13998 12044 14004 12056
rect 14056 12044 14062 12096
rect 15194 12044 15200 12096
rect 15252 12084 15258 12096
rect 16482 12084 16488 12096
rect 15252 12056 16488 12084
rect 15252 12044 15258 12056
rect 16482 12044 16488 12056
rect 16540 12044 16546 12096
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 17052 12084 17080 12124
rect 19334 12112 19340 12164
rect 19392 12152 19398 12164
rect 20257 12155 20315 12161
rect 20257 12152 20269 12155
rect 19392 12124 20269 12152
rect 19392 12112 19398 12124
rect 20257 12121 20269 12124
rect 20303 12121 20315 12155
rect 20257 12115 20315 12121
rect 16632 12056 17080 12084
rect 16632 12044 16638 12056
rect 1104 11994 21043 12016
rect 1104 11942 5894 11994
rect 5946 11942 5958 11994
rect 6010 11942 6022 11994
rect 6074 11942 6086 11994
rect 6138 11942 6150 11994
rect 6202 11942 10839 11994
rect 10891 11942 10903 11994
rect 10955 11942 10967 11994
rect 11019 11942 11031 11994
rect 11083 11942 11095 11994
rect 11147 11942 15784 11994
rect 15836 11942 15848 11994
rect 15900 11942 15912 11994
rect 15964 11942 15976 11994
rect 16028 11942 16040 11994
rect 16092 11942 20729 11994
rect 20781 11942 20793 11994
rect 20845 11942 20857 11994
rect 20909 11942 20921 11994
rect 20973 11942 20985 11994
rect 21037 11942 21043 11994
rect 1104 11920 21043 11942
rect 3326 11840 3332 11892
rect 3384 11880 3390 11892
rect 3513 11883 3571 11889
rect 3513 11880 3525 11883
rect 3384 11852 3525 11880
rect 3384 11840 3390 11852
rect 3513 11849 3525 11852
rect 3559 11849 3571 11883
rect 3513 11843 3571 11849
rect 4430 11840 4436 11892
rect 4488 11840 4494 11892
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 7285 11883 7343 11889
rect 7285 11880 7297 11883
rect 7248 11852 7297 11880
rect 7248 11840 7254 11852
rect 7285 11849 7297 11852
rect 7331 11849 7343 11883
rect 11238 11880 11244 11892
rect 7285 11843 7343 11849
rect 7944 11852 11244 11880
rect 3050 11772 3056 11824
rect 3108 11812 3114 11824
rect 4890 11812 4896 11824
rect 3108 11784 4896 11812
rect 3108 11772 3114 11784
rect 4890 11772 4896 11784
rect 4948 11812 4954 11824
rect 4948 11784 5304 11812
rect 4948 11772 4954 11784
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11744 2375 11747
rect 2958 11744 2964 11756
rect 2363 11716 2964 11744
rect 2363 11713 2375 11716
rect 2317 11707 2375 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 3878 11704 3884 11756
rect 3936 11744 3942 11756
rect 4341 11747 4399 11753
rect 4341 11744 4353 11747
rect 3936 11716 4353 11744
rect 3936 11704 3942 11716
rect 4341 11713 4353 11716
rect 4387 11744 4399 11747
rect 4387 11716 4936 11744
rect 4387 11713 4399 11716
rect 4341 11707 4399 11713
rect 2041 11679 2099 11685
rect 2041 11645 2053 11679
rect 2087 11676 2099 11679
rect 2130 11676 2136 11688
rect 2087 11648 2136 11676
rect 2087 11645 2099 11648
rect 2041 11639 2099 11645
rect 2130 11636 2136 11648
rect 2188 11636 2194 11688
rect 3050 11636 3056 11688
rect 3108 11636 3114 11688
rect 3145 11679 3203 11685
rect 3145 11645 3157 11679
rect 3191 11645 3203 11679
rect 3145 11639 3203 11645
rect 1946 11568 1952 11620
rect 2004 11608 2010 11620
rect 2682 11608 2688 11620
rect 2004 11580 2688 11608
rect 2004 11568 2010 11580
rect 2682 11568 2688 11580
rect 2740 11608 2746 11620
rect 3160 11608 3188 11639
rect 4522 11636 4528 11688
rect 4580 11636 4586 11688
rect 4908 11676 4936 11716
rect 4982 11704 4988 11756
rect 5040 11744 5046 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 5040 11716 5181 11744
rect 5040 11704 5046 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 5276 11744 5304 11784
rect 5350 11772 5356 11824
rect 5408 11772 5414 11824
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5276 11716 5457 11744
rect 5169 11707 5227 11713
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11744 5595 11747
rect 5810 11744 5816 11756
rect 5583 11716 5816 11744
rect 5583 11713 5595 11716
rect 5537 11707 5595 11713
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 6886 11716 7205 11744
rect 6730 11676 6736 11688
rect 4908 11648 6736 11676
rect 6730 11636 6736 11648
rect 6788 11676 6794 11688
rect 6886 11676 6914 11716
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 6788 11648 6914 11676
rect 6788 11636 6794 11648
rect 7374 11636 7380 11688
rect 7432 11636 7438 11688
rect 7944 11608 7972 11852
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 11790 11840 11796 11892
rect 11848 11840 11854 11892
rect 13541 11883 13599 11889
rect 13541 11849 13553 11883
rect 13587 11880 13599 11883
rect 13814 11880 13820 11892
rect 13587 11852 13820 11880
rect 13587 11849 13599 11852
rect 13541 11843 13599 11849
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 16022 11840 16028 11892
rect 16080 11880 16086 11892
rect 18677 11883 18735 11889
rect 16080 11852 18276 11880
rect 16080 11840 16086 11852
rect 8297 11815 8355 11821
rect 8297 11781 8309 11815
rect 8343 11812 8355 11815
rect 9490 11812 9496 11824
rect 8343 11784 9496 11812
rect 8343 11781 8355 11784
rect 8297 11775 8355 11781
rect 9490 11772 9496 11784
rect 9548 11772 9554 11824
rect 11698 11772 11704 11824
rect 11756 11812 11762 11824
rect 12066 11812 12072 11824
rect 11756 11784 12072 11812
rect 11756 11772 11762 11784
rect 12066 11772 12072 11784
rect 12124 11772 12130 11824
rect 13832 11812 13860 11840
rect 13832 11784 15240 11812
rect 8021 11747 8079 11753
rect 8021 11713 8033 11747
rect 8067 11713 8079 11747
rect 8021 11707 8079 11713
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11744 8171 11747
rect 8202 11744 8208 11756
rect 8159 11716 8208 11744
rect 8159 11713 8171 11716
rect 8113 11707 8171 11713
rect 2740 11580 7972 11608
rect 2740 11568 2746 11580
rect 2130 11500 2136 11552
rect 2188 11500 2194 11552
rect 2222 11500 2228 11552
rect 2280 11500 2286 11552
rect 2866 11500 2872 11552
rect 2924 11500 2930 11552
rect 3970 11500 3976 11552
rect 4028 11500 4034 11552
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 5721 11543 5779 11549
rect 5721 11540 5733 11543
rect 4764 11512 5733 11540
rect 4764 11500 4770 11512
rect 5721 11509 5733 11512
rect 5767 11509 5779 11543
rect 5721 11503 5779 11509
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11540 6883 11543
rect 7006 11540 7012 11552
rect 6871 11512 7012 11540
rect 6871 11509 6883 11512
rect 6825 11503 6883 11509
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 8036 11540 8064 11707
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 8754 11704 8760 11756
rect 8812 11704 8818 11756
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 9309 11747 9367 11753
rect 9309 11713 9321 11747
rect 9355 11744 9367 11747
rect 9582 11744 9588 11756
rect 9355 11716 9588 11744
rect 9355 11713 9367 11716
rect 9309 11707 9367 11713
rect 8956 11676 8984 11707
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 10318 11704 10324 11756
rect 10376 11744 10382 11756
rect 10413 11747 10471 11753
rect 10413 11744 10425 11747
rect 10376 11716 10425 11744
rect 10376 11704 10382 11716
rect 10413 11713 10425 11716
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 10502 11704 10508 11756
rect 10560 11704 10566 11756
rect 10594 11704 10600 11756
rect 10652 11704 10658 11756
rect 10686 11704 10692 11756
rect 10744 11704 10750 11756
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 11664 11716 11989 11744
rect 11664 11704 11670 11716
rect 11977 11713 11989 11716
rect 12023 11713 12035 11747
rect 11977 11707 12035 11713
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 8312 11648 8984 11676
rect 8312 11617 8340 11648
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 11790 11676 11796 11688
rect 11388 11648 11796 11676
rect 11388 11636 11394 11648
rect 11790 11636 11796 11648
rect 11848 11676 11854 11688
rect 12176 11676 12204 11707
rect 13170 11704 13176 11756
rect 13228 11704 13234 11756
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11744 13415 11747
rect 14734 11744 14740 11756
rect 13403 11716 14740 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 11848 11648 12664 11676
rect 11848 11636 11854 11648
rect 8297 11611 8355 11617
rect 8297 11577 8309 11611
rect 8343 11577 8355 11611
rect 8297 11571 8355 11577
rect 11882 11568 11888 11620
rect 11940 11608 11946 11620
rect 12345 11611 12403 11617
rect 12345 11608 12357 11611
rect 11940 11580 12357 11608
rect 11940 11568 11946 11580
rect 12345 11577 12357 11580
rect 12391 11577 12403 11611
rect 12636 11608 12664 11648
rect 12710 11636 12716 11688
rect 12768 11676 12774 11688
rect 13372 11676 13400 11707
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 15010 11704 15016 11756
rect 15068 11704 15074 11756
rect 15212 11753 15240 11784
rect 15930 11772 15936 11824
rect 15988 11772 15994 11824
rect 16482 11772 16488 11824
rect 16540 11812 16546 11824
rect 17681 11815 17739 11821
rect 17681 11812 17693 11815
rect 16540 11784 17693 11812
rect 16540 11772 16546 11784
rect 17681 11781 17693 11784
rect 17727 11781 17739 11815
rect 18138 11812 18144 11824
rect 17681 11775 17739 11781
rect 17880 11784 18144 11812
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11744 15255 11747
rect 15286 11744 15292 11756
rect 15243 11716 15292 11744
rect 15243 11713 15255 11716
rect 15197 11707 15255 11713
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 15657 11747 15715 11753
rect 15657 11713 15669 11747
rect 15703 11713 15715 11747
rect 15657 11707 15715 11713
rect 15805 11747 15863 11753
rect 15805 11713 15817 11747
rect 15851 11744 15863 11747
rect 15851 11713 15884 11744
rect 15805 11707 15884 11713
rect 12768 11648 13400 11676
rect 12768 11636 12774 11648
rect 14826 11636 14832 11688
rect 14884 11676 14890 11688
rect 15672 11676 15700 11707
rect 14884 11648 15700 11676
rect 15856 11676 15884 11707
rect 16022 11704 16028 11756
rect 16080 11704 16086 11756
rect 16114 11704 16120 11756
rect 16172 11753 16178 11756
rect 16172 11744 16180 11753
rect 16172 11716 16217 11744
rect 16172 11707 16180 11716
rect 16172 11704 16178 11707
rect 16850 11704 16856 11756
rect 16908 11704 16914 11756
rect 17880 11753 17908 11784
rect 18138 11772 18144 11784
rect 18196 11772 18202 11824
rect 18248 11812 18276 11852
rect 18677 11849 18689 11883
rect 18723 11880 18735 11883
rect 18966 11880 18972 11892
rect 18723 11852 18972 11880
rect 18723 11849 18735 11852
rect 18677 11843 18735 11849
rect 18966 11840 18972 11852
rect 19024 11840 19030 11892
rect 19610 11840 19616 11892
rect 19668 11880 19674 11892
rect 19705 11883 19763 11889
rect 19705 11880 19717 11883
rect 19668 11852 19717 11880
rect 19668 11840 19674 11852
rect 19705 11849 19717 11852
rect 19751 11849 19763 11883
rect 19705 11843 19763 11849
rect 18877 11815 18935 11821
rect 18877 11812 18889 11815
rect 18248 11784 18889 11812
rect 18877 11781 18889 11784
rect 18923 11812 18935 11815
rect 19518 11812 19524 11824
rect 18923 11784 19524 11812
rect 18923 11781 18935 11784
rect 18877 11775 18935 11781
rect 19518 11772 19524 11784
rect 19576 11772 19582 11824
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11713 17923 11747
rect 17865 11707 17923 11713
rect 17954 11704 17960 11756
rect 18012 11704 18018 11756
rect 18782 11704 18788 11756
rect 18840 11744 18846 11756
rect 19337 11747 19395 11753
rect 19337 11744 19349 11747
rect 18840 11716 19349 11744
rect 18840 11704 18846 11716
rect 19337 11713 19349 11716
rect 19383 11713 19395 11747
rect 19337 11707 19395 11713
rect 17129 11679 17187 11685
rect 15856 11648 17080 11676
rect 14884 11636 14890 11648
rect 15470 11608 15476 11620
rect 12636 11580 15476 11608
rect 12345 11571 12403 11577
rect 15470 11568 15476 11580
rect 15528 11608 15534 11620
rect 16022 11608 16028 11620
rect 15528 11580 16028 11608
rect 15528 11568 15534 11580
rect 16022 11568 16028 11580
rect 16080 11568 16086 11620
rect 17052 11617 17080 11648
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 18046 11676 18052 11688
rect 17175 11648 18052 11676
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 18874 11636 18880 11688
rect 18932 11676 18938 11688
rect 19429 11679 19487 11685
rect 19429 11676 19441 11679
rect 18932 11648 19441 11676
rect 18932 11636 18938 11648
rect 19429 11645 19441 11648
rect 19475 11645 19487 11679
rect 19429 11639 19487 11645
rect 17037 11611 17095 11617
rect 17037 11577 17049 11611
rect 17083 11577 17095 11611
rect 17037 11571 17095 11577
rect 17954 11568 17960 11620
rect 18012 11608 18018 11620
rect 20070 11608 20076 11620
rect 18012 11580 20076 11608
rect 18012 11568 18018 11580
rect 8938 11540 8944 11552
rect 8036 11512 8944 11540
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 10229 11543 10287 11549
rect 10229 11540 10241 11543
rect 10100 11512 10241 11540
rect 10100 11500 10106 11512
rect 10229 11509 10241 11512
rect 10275 11509 10287 11543
rect 10229 11503 10287 11509
rect 15194 11500 15200 11552
rect 15252 11500 15258 11552
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 16114 11540 16120 11552
rect 15344 11512 16120 11540
rect 15344 11500 15350 11512
rect 16114 11500 16120 11512
rect 16172 11500 16178 11552
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 16264 11512 16313 11540
rect 16264 11500 16270 11512
rect 16301 11509 16313 11512
rect 16347 11509 16359 11543
rect 16301 11503 16359 11509
rect 16942 11500 16948 11552
rect 17000 11500 17006 11552
rect 18509 11543 18567 11549
rect 18509 11509 18521 11543
rect 18555 11540 18567 11543
rect 18598 11540 18604 11552
rect 18555 11512 18604 11540
rect 18555 11509 18567 11512
rect 18509 11503 18567 11509
rect 18598 11500 18604 11512
rect 18656 11500 18662 11552
rect 18708 11549 18736 11580
rect 20070 11568 20076 11580
rect 20128 11568 20134 11620
rect 18693 11543 18751 11549
rect 18693 11509 18705 11543
rect 18739 11509 18751 11543
rect 18693 11503 18751 11509
rect 19334 11500 19340 11552
rect 19392 11500 19398 11552
rect 1104 11450 20884 11472
rect 1104 11398 3422 11450
rect 3474 11398 3486 11450
rect 3538 11398 3550 11450
rect 3602 11398 3614 11450
rect 3666 11398 3678 11450
rect 3730 11398 8367 11450
rect 8419 11398 8431 11450
rect 8483 11398 8495 11450
rect 8547 11398 8559 11450
rect 8611 11398 8623 11450
rect 8675 11398 13312 11450
rect 13364 11398 13376 11450
rect 13428 11398 13440 11450
rect 13492 11398 13504 11450
rect 13556 11398 13568 11450
rect 13620 11398 18257 11450
rect 18309 11398 18321 11450
rect 18373 11398 18385 11450
rect 18437 11398 18449 11450
rect 18501 11398 18513 11450
rect 18565 11398 20884 11450
rect 1104 11376 20884 11398
rect 1946 11296 1952 11348
rect 2004 11296 2010 11348
rect 2498 11296 2504 11348
rect 2556 11296 2562 11348
rect 4982 11296 4988 11348
rect 5040 11296 5046 11348
rect 5166 11296 5172 11348
rect 5224 11336 5230 11348
rect 5224 11308 6914 11336
rect 5224 11296 5230 11308
rect 4890 11228 4896 11280
rect 4948 11268 4954 11280
rect 6886 11268 6914 11308
rect 8754 11296 8760 11348
rect 8812 11336 8818 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 8812 11308 9137 11336
rect 8812 11296 8818 11308
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 9125 11299 9183 11305
rect 11422 11296 11428 11348
rect 11480 11296 11486 11348
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 15933 11339 15991 11345
rect 15933 11336 15945 11339
rect 14516 11308 15945 11336
rect 14516 11296 14522 11308
rect 15933 11305 15945 11308
rect 15979 11336 15991 11339
rect 16850 11336 16856 11348
rect 15979 11308 16856 11336
rect 15979 11305 15991 11308
rect 15933 11299 15991 11305
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 18138 11296 18144 11348
rect 18196 11336 18202 11348
rect 18233 11339 18291 11345
rect 18233 11336 18245 11339
rect 18196 11308 18245 11336
rect 18196 11296 18202 11308
rect 18233 11305 18245 11308
rect 18279 11305 18291 11339
rect 18233 11299 18291 11305
rect 18690 11296 18696 11348
rect 18748 11345 18754 11348
rect 18748 11339 18770 11345
rect 18758 11305 18770 11339
rect 18748 11299 18770 11305
rect 18748 11296 18754 11299
rect 14366 11268 14372 11280
rect 4948 11240 5856 11268
rect 6886 11240 14372 11268
rect 4948 11228 4954 11240
rect 3050 11160 3056 11212
rect 3108 11200 3114 11212
rect 4062 11200 4068 11212
rect 3108 11172 4068 11200
rect 3108 11160 3114 11172
rect 4062 11160 4068 11172
rect 4120 11200 4126 11212
rect 5353 11203 5411 11209
rect 5353 11200 5365 11203
rect 4120 11172 5365 11200
rect 4120 11160 4126 11172
rect 5353 11169 5365 11172
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 2590 11092 2596 11144
rect 2648 11132 2654 11144
rect 2685 11135 2743 11141
rect 2685 11132 2697 11135
rect 2648 11104 2697 11132
rect 2648 11092 2654 11104
rect 2685 11101 2697 11104
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 2958 11132 2964 11144
rect 2915 11104 2964 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 4522 11092 4528 11144
rect 4580 11132 4586 11144
rect 5166 11132 5172 11144
rect 4580 11104 5172 11132
rect 4580 11092 4586 11104
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 5626 11132 5632 11144
rect 5491 11104 5632 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 5828 11132 5856 11240
rect 7006 11160 7012 11212
rect 7064 11160 7070 11212
rect 7208 11209 7236 11240
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 16574 11268 16580 11280
rect 16132 11240 16580 11268
rect 7193 11203 7251 11209
rect 7193 11169 7205 11203
rect 7239 11169 7251 11203
rect 9585 11203 9643 11209
rect 9585 11200 9597 11203
rect 7193 11163 7251 11169
rect 8220 11172 9597 11200
rect 8220 11132 8248 11172
rect 9585 11169 9597 11172
rect 9631 11169 9643 11203
rect 9585 11163 9643 11169
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 14090 11200 14096 11212
rect 11664 11172 14096 11200
rect 11664 11160 11670 11172
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 5828 11104 8248 11132
rect 8938 11092 8944 11144
rect 8996 11132 9002 11144
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 8996 11104 9321 11132
rect 8996 11092 9002 11104
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 934 11024 940 11076
rect 992 11064 998 11076
rect 1673 11067 1731 11073
rect 1673 11064 1685 11067
rect 992 11036 1685 11064
rect 992 11024 998 11036
rect 1673 11033 1685 11036
rect 1719 11033 1731 11067
rect 1673 11027 1731 11033
rect 6914 11024 6920 11076
rect 6972 11024 6978 11076
rect 8202 11024 8208 11076
rect 8260 11064 8266 11076
rect 9416 11064 9444 11095
rect 9490 11092 9496 11144
rect 9548 11092 9554 11144
rect 11698 11092 11704 11144
rect 11756 11092 11762 11144
rect 11790 11092 11796 11144
rect 11848 11092 11854 11144
rect 11882 11092 11888 11144
rect 11940 11092 11946 11144
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11132 14519 11135
rect 14550 11132 14556 11144
rect 14507 11104 14556 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 10318 11064 10324 11076
rect 8260 11036 9444 11064
rect 9600 11036 10324 11064
rect 8260 11024 8266 11036
rect 6546 10956 6552 11008
rect 6604 10956 6610 11008
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 9600 10996 9628 11036
rect 10318 11024 10324 11036
rect 10376 11024 10382 11076
rect 10410 11024 10416 11076
rect 10468 11064 10474 11076
rect 12710 11064 12716 11076
rect 10468 11036 12716 11064
rect 10468 11024 10474 11036
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 13078 11024 13084 11076
rect 13136 11064 13142 11076
rect 14369 11067 14427 11073
rect 14369 11064 14381 11067
rect 13136 11036 14381 11064
rect 13136 11024 13142 11036
rect 14369 11033 14381 11036
rect 14415 11033 14427 11067
rect 14369 11027 14427 11033
rect 8168 10968 9628 10996
rect 14476 10996 14504 11095
rect 14550 11092 14556 11104
rect 14608 11092 14614 11144
rect 16132 11141 16160 11240
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 18601 11271 18659 11277
rect 18601 11237 18613 11271
rect 18647 11237 18659 11271
rect 18601 11231 18659 11237
rect 18509 11203 18567 11209
rect 18509 11169 18521 11203
rect 18555 11169 18567 11203
rect 18616 11200 18644 11231
rect 18782 11200 18788 11212
rect 18616 11172 18788 11200
rect 18509 11163 18567 11169
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 16209 11135 16267 11141
rect 16209 11101 16221 11135
rect 16255 11132 16267 11135
rect 17954 11132 17960 11144
rect 16255 11104 17960 11132
rect 16255 11101 16267 11104
rect 16209 11095 16267 11101
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 16224 11064 16252 11095
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 18524 11132 18552 11163
rect 18782 11160 18788 11172
rect 18840 11160 18846 11212
rect 18874 11160 18880 11212
rect 18932 11160 18938 11212
rect 18690 11132 18696 11144
rect 18524 11104 18696 11132
rect 18690 11092 18696 11104
rect 18748 11132 18754 11144
rect 18892 11132 18920 11160
rect 18748 11104 18920 11132
rect 18748 11092 18754 11104
rect 14884 11036 16252 11064
rect 14884 11024 14890 11036
rect 18874 11024 18880 11076
rect 18932 11024 18938 11076
rect 16942 10996 16948 11008
rect 14476 10968 16948 10996
rect 8168 10956 8174 10968
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 1104 10906 21043 10928
rect 1104 10854 5894 10906
rect 5946 10854 5958 10906
rect 6010 10854 6022 10906
rect 6074 10854 6086 10906
rect 6138 10854 6150 10906
rect 6202 10854 10839 10906
rect 10891 10854 10903 10906
rect 10955 10854 10967 10906
rect 11019 10854 11031 10906
rect 11083 10854 11095 10906
rect 11147 10854 15784 10906
rect 15836 10854 15848 10906
rect 15900 10854 15912 10906
rect 15964 10854 15976 10906
rect 16028 10854 16040 10906
rect 16092 10854 20729 10906
rect 20781 10854 20793 10906
rect 20845 10854 20857 10906
rect 20909 10854 20921 10906
rect 20973 10854 20985 10906
rect 21037 10854 21043 10906
rect 1104 10832 21043 10854
rect 1949 10795 2007 10801
rect 1949 10761 1961 10795
rect 1995 10792 2007 10795
rect 2958 10792 2964 10804
rect 1995 10764 2964 10792
rect 1995 10761 2007 10764
rect 1949 10755 2007 10761
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 13725 10795 13783 10801
rect 13725 10792 13737 10795
rect 12492 10764 13737 10792
rect 12492 10752 12498 10764
rect 13725 10761 13737 10764
rect 13771 10761 13783 10795
rect 13725 10755 13783 10761
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 18932 10764 19809 10792
rect 18932 10752 18938 10764
rect 19797 10761 19809 10764
rect 19843 10761 19855 10795
rect 19797 10755 19855 10761
rect 1765 10727 1823 10733
rect 1765 10693 1777 10727
rect 1811 10724 1823 10727
rect 2130 10724 2136 10736
rect 1811 10696 2136 10724
rect 1811 10693 1823 10696
rect 1765 10687 1823 10693
rect 2130 10684 2136 10696
rect 2188 10684 2194 10736
rect 11698 10684 11704 10736
rect 11756 10724 11762 10736
rect 14826 10724 14832 10736
rect 11756 10696 14832 10724
rect 11756 10684 11762 10696
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2222 10656 2228 10668
rect 2087 10628 2228 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 12710 10616 12716 10668
rect 12768 10656 12774 10668
rect 13096 10665 13124 10696
rect 14826 10684 14832 10696
rect 14884 10684 14890 10736
rect 14918 10684 14924 10736
rect 14976 10724 14982 10736
rect 18049 10727 18107 10733
rect 14976 10696 16068 10724
rect 14976 10684 14982 10696
rect 12897 10659 12955 10665
rect 12897 10656 12909 10659
rect 12768 10628 12909 10656
rect 12768 10616 12774 10628
rect 12897 10625 12909 10628
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 15252 10628 15761 10656
rect 15252 10616 15258 10628
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 15838 10616 15844 10668
rect 15896 10656 15902 10668
rect 16040 10665 16068 10696
rect 18049 10693 18061 10727
rect 18095 10724 18107 10727
rect 18892 10724 18920 10752
rect 18095 10696 18920 10724
rect 18095 10693 18107 10696
rect 18049 10687 18107 10693
rect 16025 10659 16083 10665
rect 15896 10616 15916 10656
rect 16025 10625 16037 10659
rect 16071 10625 16083 10659
rect 16025 10619 16083 10625
rect 16206 10616 16212 10668
rect 16264 10616 16270 10668
rect 18524 10665 18552 10696
rect 18966 10684 18972 10736
rect 19024 10724 19030 10736
rect 19024 10696 20300 10724
rect 19024 10684 19030 10696
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 18509 10659 18567 10665
rect 18509 10625 18521 10659
rect 18555 10625 18567 10659
rect 18509 10619 18567 10625
rect 12820 10560 13032 10588
rect 10594 10480 10600 10532
rect 10652 10520 10658 10532
rect 12434 10520 12440 10532
rect 10652 10492 12440 10520
rect 10652 10480 10658 10492
rect 12434 10480 12440 10492
rect 12492 10480 12498 10532
rect 1765 10455 1823 10461
rect 1765 10421 1777 10455
rect 1811 10452 1823 10455
rect 1854 10452 1860 10464
rect 1811 10424 1860 10452
rect 1811 10421 1823 10424
rect 1765 10415 1823 10421
rect 1854 10412 1860 10424
rect 1912 10412 1918 10464
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 12820 10452 12848 10560
rect 13004 10520 13032 10560
rect 13906 10548 13912 10600
rect 13964 10548 13970 10600
rect 14093 10591 14151 10597
rect 14093 10557 14105 10591
rect 14139 10557 14151 10591
rect 14093 10551 14151 10557
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10588 14243 10591
rect 15565 10591 15623 10597
rect 15565 10588 15577 10591
rect 14231 10560 15577 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 15565 10557 15577 10560
rect 15611 10557 15623 10591
rect 15888 10588 15916 10616
rect 17034 10588 17040 10600
rect 15888 10560 17040 10588
rect 15565 10551 15623 10557
rect 14108 10520 14136 10551
rect 17034 10548 17040 10560
rect 17092 10588 17098 10600
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 17092 10560 17509 10588
rect 17092 10548 17098 10560
rect 17497 10557 17509 10560
rect 17543 10557 17555 10591
rect 17880 10588 17908 10619
rect 18598 10616 18604 10668
rect 18656 10616 18662 10668
rect 18690 10616 18696 10668
rect 18748 10656 18754 10668
rect 18785 10659 18843 10665
rect 18785 10656 18797 10659
rect 18748 10628 18797 10656
rect 18748 10616 18754 10628
rect 18785 10625 18797 10628
rect 18831 10625 18843 10659
rect 18785 10619 18843 10625
rect 19518 10616 19524 10668
rect 19576 10656 19582 10668
rect 19705 10659 19763 10665
rect 19705 10656 19717 10659
rect 19576 10628 19717 10656
rect 19576 10616 19582 10628
rect 19705 10625 19717 10628
rect 19751 10625 19763 10659
rect 19705 10619 19763 10625
rect 20070 10616 20076 10668
rect 20128 10616 20134 10668
rect 20272 10665 20300 10696
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10625 20315 10659
rect 20257 10619 20315 10625
rect 18616 10588 18644 10616
rect 17880 10560 18644 10588
rect 18969 10591 19027 10597
rect 17497 10551 17555 10557
rect 18969 10557 18981 10591
rect 19015 10557 19027 10591
rect 18969 10551 19027 10557
rect 13004 10492 14136 10520
rect 14274 10480 14280 10532
rect 14332 10520 14338 10532
rect 15841 10523 15899 10529
rect 15841 10520 15853 10523
rect 14332 10492 15853 10520
rect 14332 10480 14338 10492
rect 15841 10489 15853 10492
rect 15887 10489 15899 10523
rect 15841 10483 15899 10489
rect 15933 10523 15991 10529
rect 15933 10489 15945 10523
rect 15979 10520 15991 10523
rect 16022 10520 16028 10532
rect 15979 10492 16028 10520
rect 15979 10489 15991 10492
rect 15933 10483 15991 10489
rect 16022 10480 16028 10492
rect 16080 10480 16086 10532
rect 16942 10480 16948 10532
rect 17000 10520 17006 10532
rect 18984 10520 19012 10551
rect 17000 10492 19012 10520
rect 17000 10480 17006 10492
rect 9640 10424 12848 10452
rect 9640 10412 9646 10424
rect 12986 10412 12992 10464
rect 13044 10412 13050 10464
rect 1104 10362 20884 10384
rect 1104 10310 3422 10362
rect 3474 10310 3486 10362
rect 3538 10310 3550 10362
rect 3602 10310 3614 10362
rect 3666 10310 3678 10362
rect 3730 10310 8367 10362
rect 8419 10310 8431 10362
rect 8483 10310 8495 10362
rect 8547 10310 8559 10362
rect 8611 10310 8623 10362
rect 8675 10310 13312 10362
rect 13364 10310 13376 10362
rect 13428 10310 13440 10362
rect 13492 10310 13504 10362
rect 13556 10310 13568 10362
rect 13620 10310 18257 10362
rect 18309 10310 18321 10362
rect 18373 10310 18385 10362
rect 18437 10310 18449 10362
rect 18501 10310 18513 10362
rect 18565 10310 20884 10362
rect 1104 10288 20884 10310
rect 2958 10208 2964 10260
rect 3016 10208 3022 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 9490 10248 9496 10260
rect 8619 10220 9496 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 11698 10208 11704 10260
rect 11756 10208 11762 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 14369 10251 14427 10257
rect 14369 10248 14381 10251
rect 13964 10220 14381 10248
rect 13964 10208 13970 10220
rect 14369 10217 14381 10220
rect 14415 10217 14427 10251
rect 14369 10211 14427 10217
rect 14599 10251 14657 10257
rect 14599 10217 14611 10251
rect 14645 10248 14657 10251
rect 14734 10248 14740 10260
rect 14645 10220 14740 10248
rect 14645 10217 14657 10220
rect 14599 10211 14657 10217
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 15838 10208 15844 10260
rect 15896 10208 15902 10260
rect 16022 10208 16028 10260
rect 16080 10208 16086 10260
rect 16485 10251 16543 10257
rect 16485 10217 16497 10251
rect 16531 10248 16543 10251
rect 16666 10248 16672 10260
rect 16531 10220 16672 10248
rect 16531 10217 16543 10220
rect 16485 10211 16543 10217
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 13725 10183 13783 10189
rect 13725 10149 13737 10183
rect 13771 10180 13783 10183
rect 14461 10183 14519 10189
rect 14461 10180 14473 10183
rect 13771 10152 14473 10180
rect 13771 10149 13783 10152
rect 13725 10143 13783 10149
rect 14461 10149 14473 10152
rect 14507 10149 14519 10183
rect 14461 10143 14519 10149
rect 13740 10084 15792 10112
rect 1578 10004 1584 10056
rect 1636 10004 1642 10056
rect 1854 10053 1860 10056
rect 1848 10044 1860 10053
rect 1815 10016 1860 10044
rect 1848 10007 1860 10016
rect 1854 10004 1860 10007
rect 1912 10004 1918 10056
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 7834 10044 7840 10056
rect 7239 10016 7840 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 7834 10004 7840 10016
rect 7892 10004 7898 10056
rect 10318 10004 10324 10056
rect 10376 10004 10382 10056
rect 10597 10047 10655 10053
rect 10597 10013 10609 10047
rect 10643 10044 10655 10047
rect 10643 10016 12940 10044
rect 10643 10013 10655 10016
rect 10597 10007 10655 10013
rect 7460 9979 7518 9985
rect 7460 9945 7472 9979
rect 7506 9976 7518 9979
rect 8110 9976 8116 9988
rect 7506 9948 8116 9976
rect 7506 9945 7518 9948
rect 7460 9939 7518 9945
rect 8110 9936 8116 9948
rect 8168 9936 8174 9988
rect 12912 9908 12940 10016
rect 13538 10004 13544 10056
rect 13596 10004 13602 10056
rect 13740 10053 13768 10084
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 14274 10004 14280 10056
rect 14332 10004 14338 10056
rect 14734 10004 14740 10056
rect 14792 10004 14798 10056
rect 12986 9936 12992 9988
rect 13044 9976 13050 9988
rect 15657 9979 15715 9985
rect 15657 9976 15669 9979
rect 13044 9948 15669 9976
rect 13044 9936 13050 9948
rect 15657 9945 15669 9948
rect 15703 9945 15715 9979
rect 15764 9976 15792 10084
rect 16040 10044 16068 10208
rect 19058 10112 19064 10124
rect 18708 10084 19064 10112
rect 16485 10047 16543 10053
rect 16485 10044 16497 10047
rect 16040 10016 16497 10044
rect 16485 10013 16497 10016
rect 16531 10013 16543 10047
rect 16485 10007 16543 10013
rect 16758 10004 16764 10056
rect 16816 10004 16822 10056
rect 18138 10004 18144 10056
rect 18196 10004 18202 10056
rect 18708 10053 18736 10084
rect 19058 10072 19064 10084
rect 19116 10072 19122 10124
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10013 18751 10047
rect 18693 10007 18751 10013
rect 18874 10004 18880 10056
rect 18932 10004 18938 10056
rect 15873 9979 15931 9985
rect 15873 9976 15885 9979
rect 15764 9948 15885 9976
rect 15657 9939 15715 9945
rect 15873 9945 15885 9948
rect 15919 9976 15931 9979
rect 16390 9976 16396 9988
rect 15919 9948 16396 9976
rect 15919 9945 15931 9948
rect 15873 9939 15931 9945
rect 16390 9936 16396 9948
rect 16448 9936 16454 9988
rect 16574 9936 16580 9988
rect 16632 9976 16638 9988
rect 16669 9979 16727 9985
rect 16669 9976 16681 9979
rect 16632 9948 16681 9976
rect 16632 9936 16638 9948
rect 16669 9945 16681 9948
rect 16715 9976 16727 9979
rect 17589 9979 17647 9985
rect 17589 9976 17601 9979
rect 16715 9948 17601 9976
rect 16715 9945 16727 9948
rect 16669 9939 16727 9945
rect 17589 9945 17601 9948
rect 17635 9945 17647 9979
rect 17589 9939 17647 9945
rect 14734 9908 14740 9920
rect 12912 9880 14740 9908
rect 14734 9868 14740 9880
rect 14792 9868 14798 9920
rect 1104 9818 21043 9840
rect 1104 9766 5894 9818
rect 5946 9766 5958 9818
rect 6010 9766 6022 9818
rect 6074 9766 6086 9818
rect 6138 9766 6150 9818
rect 6202 9766 10839 9818
rect 10891 9766 10903 9818
rect 10955 9766 10967 9818
rect 11019 9766 11031 9818
rect 11083 9766 11095 9818
rect 11147 9766 15784 9818
rect 15836 9766 15848 9818
rect 15900 9766 15912 9818
rect 15964 9766 15976 9818
rect 16028 9766 16040 9818
rect 16092 9766 20729 9818
rect 20781 9766 20793 9818
rect 20845 9766 20857 9818
rect 20909 9766 20921 9818
rect 20973 9766 20985 9818
rect 21037 9766 21043 9818
rect 1104 9744 21043 9766
rect 2952 9639 3010 9645
rect 2952 9605 2964 9639
rect 2998 9636 3010 9639
rect 3970 9636 3976 9648
rect 2998 9608 3976 9636
rect 2998 9605 3010 9608
rect 2952 9599 3010 9605
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 4614 9596 4620 9648
rect 4672 9636 4678 9648
rect 4770 9639 4828 9645
rect 4770 9636 4782 9639
rect 4672 9608 4782 9636
rect 4672 9596 4678 9608
rect 4770 9605 4782 9608
rect 4816 9605 4828 9639
rect 10318 9636 10324 9648
rect 4770 9599 4828 9605
rect 9784 9608 10324 9636
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 9784 9577 9812 9608
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 15102 9596 15108 9648
rect 15160 9636 15166 9648
rect 15289 9639 15347 9645
rect 15289 9636 15301 9639
rect 15160 9608 15301 9636
rect 15160 9596 15166 9608
rect 15289 9605 15301 9608
rect 15335 9605 15347 9639
rect 15289 9599 15347 9605
rect 15933 9639 15991 9645
rect 15933 9605 15945 9639
rect 15979 9636 15991 9639
rect 16758 9636 16764 9648
rect 15979 9608 16764 9636
rect 15979 9605 15991 9608
rect 15933 9599 15991 9605
rect 16758 9596 16764 9608
rect 16816 9596 16822 9648
rect 10042 9577 10048 9580
rect 8205 9571 8263 9577
rect 8205 9568 8217 9571
rect 7892 9540 8217 9568
rect 7892 9528 7898 9540
rect 8205 9537 8217 9540
rect 8251 9568 8263 9571
rect 9769 9571 9827 9577
rect 9769 9568 9781 9571
rect 8251 9540 9781 9568
rect 8251 9537 8263 9540
rect 8205 9531 8263 9537
rect 9769 9537 9781 9540
rect 9815 9537 9827 9571
rect 10036 9568 10048 9577
rect 10003 9540 10048 9568
rect 9769 9531 9827 9537
rect 10036 9531 10048 9540
rect 10042 9528 10048 9531
rect 10100 9528 10106 9580
rect 15194 9528 15200 9580
rect 15252 9528 15258 9580
rect 15841 9571 15899 9577
rect 15841 9537 15853 9571
rect 15887 9537 15899 9571
rect 15841 9531 15899 9537
rect 16025 9571 16083 9577
rect 16025 9537 16037 9571
rect 16071 9568 16083 9571
rect 16114 9568 16120 9580
rect 16071 9540 16120 9568
rect 16071 9537 16083 9540
rect 16025 9531 16083 9537
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 1636 9472 2697 9500
rect 1636 9460 1642 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 4430 9460 4436 9512
rect 4488 9500 4494 9512
rect 4525 9503 4583 9509
rect 4525 9500 4537 9503
rect 4488 9472 4537 9500
rect 4488 9460 4494 9472
rect 4525 9469 4537 9472
rect 4571 9469 4583 9503
rect 4525 9463 4583 9469
rect 6822 9460 6828 9512
rect 6880 9460 6886 9512
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9500 7987 9503
rect 8846 9500 8852 9512
rect 7975 9472 8852 9500
rect 7975 9469 7987 9472
rect 7929 9463 7987 9469
rect 8846 9460 8852 9472
rect 8904 9460 8910 9512
rect 3878 9392 3884 9444
rect 3936 9432 3942 9444
rect 4065 9435 4123 9441
rect 4065 9432 4077 9435
rect 3936 9404 4077 9432
rect 3936 9392 3942 9404
rect 4065 9401 4077 9404
rect 4111 9401 4123 9435
rect 4065 9395 4123 9401
rect 14734 9392 14740 9444
rect 14792 9432 14798 9444
rect 15856 9432 15884 9531
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 18138 9528 18144 9580
rect 18196 9568 18202 9580
rect 18966 9568 18972 9580
rect 18196 9540 18972 9568
rect 18196 9528 18202 9540
rect 18966 9528 18972 9540
rect 19024 9528 19030 9580
rect 19889 9571 19947 9577
rect 19889 9537 19901 9571
rect 19935 9568 19947 9571
rect 20070 9568 20076 9580
rect 19935 9540 20076 9568
rect 19935 9537 19947 9540
rect 19889 9531 19947 9537
rect 20070 9528 20076 9540
rect 20128 9528 20134 9580
rect 14792 9404 15884 9432
rect 19061 9435 19119 9441
rect 14792 9392 14798 9404
rect 19061 9401 19073 9435
rect 19107 9432 19119 9435
rect 19334 9432 19340 9444
rect 19107 9404 19340 9432
rect 19107 9401 19119 9404
rect 19061 9395 19119 9401
rect 19334 9392 19340 9404
rect 19392 9392 19398 9444
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 4856 9336 5917 9364
rect 4856 9324 4862 9336
rect 5905 9333 5917 9336
rect 5951 9333 5963 9367
rect 5905 9327 5963 9333
rect 11149 9367 11207 9373
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 13170 9364 13176 9376
rect 11195 9336 13176 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 15194 9324 15200 9376
rect 15252 9364 15258 9376
rect 16666 9364 16672 9376
rect 15252 9336 16672 9364
rect 15252 9324 15258 9336
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 1104 9274 20884 9296
rect 1104 9222 3422 9274
rect 3474 9222 3486 9274
rect 3538 9222 3550 9274
rect 3602 9222 3614 9274
rect 3666 9222 3678 9274
rect 3730 9222 8367 9274
rect 8419 9222 8431 9274
rect 8483 9222 8495 9274
rect 8547 9222 8559 9274
rect 8611 9222 8623 9274
rect 8675 9222 13312 9274
rect 13364 9222 13376 9274
rect 13428 9222 13440 9274
rect 13492 9222 13504 9274
rect 13556 9222 13568 9274
rect 13620 9222 18257 9274
rect 18309 9222 18321 9274
rect 18373 9222 18385 9274
rect 18437 9222 18449 9274
rect 18501 9222 18513 9274
rect 18565 9222 20884 9274
rect 1104 9200 20884 9222
rect 3050 9120 3056 9172
rect 3108 9160 3114 9172
rect 3421 9163 3479 9169
rect 3421 9160 3433 9163
rect 3108 9132 3433 9160
rect 3108 9120 3114 9132
rect 3421 9129 3433 9132
rect 3467 9129 3479 9163
rect 3421 9123 3479 9129
rect 5810 9120 5816 9172
rect 5868 9120 5874 9172
rect 6457 9163 6515 9169
rect 6457 9129 6469 9163
rect 6503 9160 6515 9163
rect 8018 9160 8024 9172
rect 6503 9132 8024 9160
rect 6503 9129 6515 9132
rect 6457 9123 6515 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 10244 9132 11284 9160
rect 1578 8984 1584 9036
rect 1636 9024 1642 9036
rect 2041 9027 2099 9033
rect 2041 9024 2053 9027
rect 1636 8996 2053 9024
rect 1636 8984 1642 8996
rect 2041 8993 2053 8996
rect 2087 8993 2099 9027
rect 2041 8987 2099 8993
rect 7834 8984 7840 9036
rect 7892 8984 7898 9036
rect 2308 8959 2366 8965
rect 2308 8925 2320 8959
rect 2354 8956 2366 8959
rect 2866 8956 2872 8968
rect 2354 8928 2872 8956
rect 2354 8925 2366 8928
rect 2308 8919 2366 8925
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 4430 8916 4436 8968
rect 4488 8916 4494 8968
rect 4706 8965 4712 8968
rect 4700 8956 4712 8965
rect 4667 8928 4712 8956
rect 4700 8919 4712 8928
rect 4706 8916 4712 8919
rect 4764 8916 4770 8968
rect 7581 8959 7639 8965
rect 7581 8925 7593 8959
rect 7627 8956 7639 8959
rect 10244 8956 10272 9132
rect 11256 9092 11284 9132
rect 11790 9120 11796 9172
rect 11848 9160 11854 9172
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 11848 9132 11897 9160
rect 11848 9120 11854 9132
rect 11885 9129 11897 9132
rect 11931 9129 11943 9163
rect 11885 9123 11943 9129
rect 14090 9120 14096 9172
rect 14148 9160 14154 9172
rect 15933 9163 15991 9169
rect 15933 9160 15945 9163
rect 14148 9132 15945 9160
rect 14148 9120 14154 9132
rect 15933 9129 15945 9132
rect 15979 9160 15991 9163
rect 18138 9160 18144 9172
rect 15979 9132 18144 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 18782 9120 18788 9172
rect 18840 9120 18846 9172
rect 14182 9092 14188 9104
rect 11256 9064 14188 9092
rect 14182 9052 14188 9064
rect 14240 9052 14246 9104
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 9024 10655 9027
rect 13078 9024 13084 9036
rect 10643 8996 13084 9024
rect 10643 8993 10655 8996
rect 10597 8987 10655 8993
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 13556 8996 14688 9024
rect 7627 8928 10272 8956
rect 7627 8925 7639 8928
rect 7581 8919 7639 8925
rect 10318 8916 10324 8968
rect 10376 8916 10382 8968
rect 13170 8916 13176 8968
rect 13228 8956 13234 8968
rect 13556 8965 13584 8996
rect 14660 8965 14688 8996
rect 14918 8984 14924 9036
rect 14976 9024 14982 9036
rect 14976 8996 16896 9024
rect 14976 8984 14982 8996
rect 13541 8959 13599 8965
rect 13541 8956 13553 8959
rect 13228 8928 13553 8956
rect 13228 8916 13234 8928
rect 13541 8925 13553 8928
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8956 13783 8959
rect 14645 8959 14703 8965
rect 13771 8928 14504 8956
rect 13771 8925 13783 8928
rect 13725 8919 13783 8925
rect 14476 8900 14504 8928
rect 14645 8925 14657 8959
rect 14691 8956 14703 8959
rect 14734 8956 14740 8968
rect 14691 8928 14740 8956
rect 14691 8925 14703 8928
rect 14645 8919 14703 8925
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 16298 8916 16304 8968
rect 16356 8916 16362 8968
rect 16393 8959 16451 8965
rect 16393 8925 16405 8959
rect 16439 8956 16451 8959
rect 16666 8956 16672 8968
rect 16439 8928 16672 8956
rect 16439 8925 16451 8928
rect 16393 8919 16451 8925
rect 16666 8916 16672 8928
rect 16724 8916 16730 8968
rect 16868 8965 16896 8996
rect 17034 8984 17040 9036
rect 17092 9024 17098 9036
rect 17862 9024 17868 9036
rect 17092 8996 17868 9024
rect 17092 8984 17098 8996
rect 17862 8984 17868 8996
rect 17920 8984 17926 9036
rect 18156 9024 18184 9120
rect 18693 9095 18751 9101
rect 18693 9061 18705 9095
rect 18739 9092 18751 9095
rect 18874 9092 18880 9104
rect 18739 9064 18880 9092
rect 18739 9061 18751 9064
rect 18693 9055 18751 9061
rect 18874 9052 18880 9064
rect 18932 9052 18938 9104
rect 18325 9027 18383 9033
rect 18325 9024 18337 9027
rect 18156 8996 18337 9024
rect 18325 8993 18337 8996
rect 18371 8993 18383 9027
rect 18325 8987 18383 8993
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8956 16911 8959
rect 16942 8956 16948 8968
rect 16899 8928 16948 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 16942 8916 16948 8928
rect 17000 8916 17006 8968
rect 17221 8959 17279 8965
rect 17221 8925 17233 8959
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 13814 8848 13820 8900
rect 13872 8888 13878 8900
rect 14277 8891 14335 8897
rect 14277 8888 14289 8891
rect 13872 8860 14289 8888
rect 13872 8848 13878 8860
rect 14277 8857 14289 8860
rect 14323 8857 14335 8891
rect 14277 8851 14335 8857
rect 14458 8848 14464 8900
rect 14516 8848 14522 8900
rect 15654 8848 15660 8900
rect 15712 8888 15718 8900
rect 17236 8888 17264 8919
rect 18138 8888 18144 8900
rect 15712 8860 18144 8888
rect 15712 8848 15718 8860
rect 18138 8848 18144 8860
rect 18196 8848 18202 8900
rect 13725 8823 13783 8829
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 13906 8820 13912 8832
rect 13771 8792 13912 8820
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 13906 8780 13912 8792
rect 13964 8780 13970 8832
rect 16298 8780 16304 8832
rect 16356 8820 16362 8832
rect 18046 8820 18052 8832
rect 16356 8792 18052 8820
rect 16356 8780 16362 8792
rect 18046 8780 18052 8792
rect 18104 8820 18110 8832
rect 18414 8820 18420 8832
rect 18104 8792 18420 8820
rect 18104 8780 18110 8792
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 1104 8730 21043 8752
rect 1104 8678 5894 8730
rect 5946 8678 5958 8730
rect 6010 8678 6022 8730
rect 6074 8678 6086 8730
rect 6138 8678 6150 8730
rect 6202 8678 10839 8730
rect 10891 8678 10903 8730
rect 10955 8678 10967 8730
rect 11019 8678 11031 8730
rect 11083 8678 11095 8730
rect 11147 8678 15784 8730
rect 15836 8678 15848 8730
rect 15900 8678 15912 8730
rect 15964 8678 15976 8730
rect 16028 8678 16040 8730
rect 16092 8678 20729 8730
rect 20781 8678 20793 8730
rect 20845 8678 20857 8730
rect 20909 8678 20921 8730
rect 20973 8678 20985 8730
rect 21037 8678 21043 8730
rect 1104 8656 21043 8678
rect 9861 8619 9919 8625
rect 9861 8585 9873 8619
rect 9907 8616 9919 8619
rect 11882 8616 11888 8628
rect 9907 8588 11888 8616
rect 9907 8585 9919 8588
rect 9861 8579 9919 8585
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 16209 8619 16267 8625
rect 16209 8585 16221 8619
rect 16255 8616 16267 8619
rect 17034 8616 17040 8628
rect 16255 8588 17040 8616
rect 16255 8585 16267 8588
rect 16209 8579 16267 8585
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 18785 8619 18843 8625
rect 18785 8585 18797 8619
rect 18831 8616 18843 8619
rect 18874 8616 18880 8628
rect 18831 8588 18880 8616
rect 18831 8585 18843 8588
rect 18785 8579 18843 8585
rect 18874 8576 18880 8588
rect 18932 8576 18938 8628
rect 10318 8548 10324 8560
rect 8496 8520 10324 8548
rect 8496 8489 8524 8520
rect 10318 8508 10324 8520
rect 10376 8508 10382 8560
rect 13906 8508 13912 8560
rect 13964 8508 13970 8560
rect 13998 8508 14004 8560
rect 14056 8548 14062 8560
rect 14056 8520 14964 8548
rect 14056 8508 14062 8520
rect 14936 8492 14964 8520
rect 16592 8520 19288 8548
rect 16592 8492 16620 8520
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 8748 8483 8806 8489
rect 8748 8449 8760 8483
rect 8794 8480 8806 8483
rect 11514 8480 11520 8492
rect 8794 8452 11520 8480
rect 8794 8449 8806 8452
rect 8748 8443 8806 8449
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 14090 8440 14096 8492
rect 14148 8489 14154 8492
rect 14148 8483 14177 8489
rect 14165 8449 14177 8483
rect 14148 8443 14177 8449
rect 14148 8440 14154 8443
rect 14734 8440 14740 8492
rect 14792 8440 14798 8492
rect 14918 8440 14924 8492
rect 14976 8440 14982 8492
rect 15102 8440 15108 8492
rect 15160 8480 15166 8492
rect 16117 8483 16175 8489
rect 16117 8480 16129 8483
rect 15160 8452 16129 8480
rect 15160 8440 15166 8452
rect 16117 8449 16129 8452
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 16574 8480 16580 8492
rect 16347 8452 16580 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8412 14335 8415
rect 15120 8412 15148 8440
rect 14323 8384 15148 8412
rect 16132 8412 16160 8443
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16684 8452 16957 8480
rect 16684 8412 16712 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17126 8440 17132 8492
rect 17184 8440 17190 8492
rect 18138 8440 18144 8492
rect 18196 8440 18202 8492
rect 18230 8440 18236 8492
rect 18288 8440 18294 8492
rect 18414 8440 18420 8492
rect 18472 8440 18478 8492
rect 18506 8440 18512 8492
rect 18564 8440 18570 8492
rect 19260 8489 19288 8520
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8449 18659 8483
rect 18601 8443 18659 8449
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8449 19303 8483
rect 19245 8443 19303 8449
rect 16132 8384 16712 8412
rect 18616 8412 18644 8443
rect 18690 8412 18696 8424
rect 18616 8384 18696 8412
rect 14323 8381 14335 8384
rect 14277 8375 14335 8381
rect 18690 8372 18696 8384
rect 18748 8412 18754 8424
rect 19337 8415 19395 8421
rect 19337 8412 19349 8415
rect 18748 8384 19349 8412
rect 18748 8372 18754 8384
rect 19337 8381 19349 8384
rect 19383 8381 19395 8415
rect 19337 8375 19395 8381
rect 16942 8304 16948 8356
rect 17000 8344 17006 8356
rect 17129 8347 17187 8353
rect 17129 8344 17141 8347
rect 17000 8316 17141 8344
rect 17000 8304 17006 8316
rect 17129 8313 17141 8316
rect 17175 8313 17187 8347
rect 17129 8307 17187 8313
rect 13630 8236 13636 8288
rect 13688 8236 13694 8288
rect 14826 8236 14832 8288
rect 14884 8236 14890 8288
rect 1104 8186 20884 8208
rect 1104 8134 3422 8186
rect 3474 8134 3486 8186
rect 3538 8134 3550 8186
rect 3602 8134 3614 8186
rect 3666 8134 3678 8186
rect 3730 8134 8367 8186
rect 8419 8134 8431 8186
rect 8483 8134 8495 8186
rect 8547 8134 8559 8186
rect 8611 8134 8623 8186
rect 8675 8134 13312 8186
rect 13364 8134 13376 8186
rect 13428 8134 13440 8186
rect 13492 8134 13504 8186
rect 13556 8134 13568 8186
rect 13620 8134 18257 8186
rect 18309 8134 18321 8186
rect 18373 8134 18385 8186
rect 18437 8134 18449 8186
rect 18501 8134 18513 8186
rect 18565 8134 20884 8186
rect 1104 8112 20884 8134
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2832 8044 2973 8072
rect 2832 8032 2838 8044
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 2961 8035 3019 8041
rect 5905 8075 5963 8081
rect 5905 8041 5917 8075
rect 5951 8072 5963 8075
rect 6454 8072 6460 8084
rect 5951 8044 6460 8072
rect 5951 8041 5963 8044
rect 5905 8035 5963 8041
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 8202 8032 8208 8084
rect 8260 8032 8266 8084
rect 11793 8075 11851 8081
rect 11793 8041 11805 8075
rect 11839 8072 11851 8075
rect 15654 8072 15660 8084
rect 11839 8044 15660 8072
rect 11839 8041 11851 8044
rect 11793 8035 11851 8041
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 16666 7964 16672 8016
rect 16724 8004 16730 8016
rect 16724 7976 17448 8004
rect 16724 7964 16730 7976
rect 17420 7948 17448 7976
rect 1578 7896 1584 7948
rect 1636 7896 1642 7948
rect 2682 7896 2688 7948
rect 2740 7936 2746 7948
rect 4430 7936 4436 7948
rect 2740 7908 4436 7936
rect 2740 7896 2746 7908
rect 4430 7896 4436 7908
rect 4488 7936 4494 7948
rect 4525 7939 4583 7945
rect 4525 7936 4537 7939
rect 4488 7908 4537 7936
rect 4488 7896 4494 7908
rect 4525 7905 4537 7908
rect 4571 7905 4583 7939
rect 4525 7899 4583 7905
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 13722 7936 13728 7948
rect 13587 7908 13728 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 13722 7896 13728 7908
rect 13780 7936 13786 7948
rect 16301 7939 16359 7945
rect 16301 7936 16313 7939
rect 13780 7908 16313 7936
rect 13780 7896 13786 7908
rect 16301 7905 16313 7908
rect 16347 7936 16359 7939
rect 17034 7936 17040 7948
rect 16347 7908 17040 7936
rect 16347 7905 16359 7908
rect 16301 7899 16359 7905
rect 17034 7896 17040 7908
rect 17092 7896 17098 7948
rect 17402 7896 17408 7948
rect 17460 7936 17466 7948
rect 17460 7908 17816 7936
rect 17460 7896 17466 7908
rect 1670 7828 1676 7880
rect 1728 7868 1734 7880
rect 1837 7871 1895 7877
rect 1837 7868 1849 7871
rect 1728 7840 1849 7868
rect 1728 7828 1734 7840
rect 1837 7837 1849 7840
rect 1883 7837 1895 7871
rect 1837 7831 1895 7837
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7834 7868 7840 7880
rect 6871 7840 7840 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 10376 7840 10425 7868
rect 10376 7828 10382 7840
rect 10413 7837 10425 7840
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 10502 7828 10508 7880
rect 10560 7868 10566 7880
rect 10669 7871 10727 7877
rect 10669 7868 10681 7871
rect 10560 7840 10681 7868
rect 10560 7828 10566 7840
rect 10669 7837 10681 7840
rect 10715 7837 10727 7871
rect 10669 7831 10727 7837
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7868 13507 7871
rect 13630 7868 13636 7880
rect 13495 7840 13636 7868
rect 13495 7837 13507 7840
rect 13449 7831 13507 7837
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 15562 7868 15568 7880
rect 14016 7840 15568 7868
rect 7098 7809 7104 7812
rect 4792 7803 4850 7809
rect 4792 7769 4804 7803
rect 4838 7800 4850 7803
rect 4838 7772 6914 7800
rect 4838 7769 4850 7772
rect 4792 7763 4850 7769
rect 6886 7732 6914 7772
rect 7092 7763 7104 7809
rect 7098 7760 7104 7763
rect 7156 7760 7162 7812
rect 14016 7800 14044 7840
rect 15562 7828 15568 7840
rect 15620 7828 15626 7880
rect 16758 7828 16764 7880
rect 16816 7868 16822 7880
rect 17126 7868 17132 7880
rect 16816 7840 17132 7868
rect 16816 7828 16822 7840
rect 17126 7828 17132 7840
rect 17184 7868 17190 7880
rect 17681 7871 17739 7877
rect 17681 7868 17693 7871
rect 17184 7840 17693 7868
rect 17184 7828 17190 7840
rect 17681 7837 17693 7840
rect 17727 7837 17739 7871
rect 17788 7868 17816 7908
rect 18046 7896 18052 7948
rect 18104 7936 18110 7948
rect 18509 7939 18567 7945
rect 18509 7936 18521 7939
rect 18104 7908 18521 7936
rect 18104 7896 18110 7908
rect 18509 7905 18521 7908
rect 18555 7905 18567 7939
rect 18509 7899 18567 7905
rect 18690 7896 18696 7948
rect 18748 7896 18754 7948
rect 18138 7868 18144 7880
rect 17788 7840 18144 7868
rect 17681 7831 17739 7837
rect 18138 7828 18144 7840
rect 18196 7868 18202 7880
rect 18414 7868 18420 7880
rect 18196 7840 18420 7868
rect 18196 7828 18202 7840
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 18598 7828 18604 7880
rect 18656 7828 18662 7880
rect 7208 7772 14044 7800
rect 7208 7732 7236 7772
rect 15102 7760 15108 7812
rect 15160 7800 15166 7812
rect 16025 7803 16083 7809
rect 16025 7800 16037 7803
rect 15160 7772 16037 7800
rect 15160 7760 15166 7772
rect 16025 7769 16037 7772
rect 16071 7769 16083 7803
rect 16025 7763 16083 7769
rect 17773 7803 17831 7809
rect 17773 7769 17785 7803
rect 17819 7800 17831 7803
rect 18616 7800 18644 7828
rect 17819 7772 18644 7800
rect 17819 7769 17831 7772
rect 17773 7763 17831 7769
rect 6886 7704 7236 7732
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 12989 7735 13047 7741
rect 12989 7732 13001 7735
rect 11940 7704 13001 7732
rect 11940 7692 11946 7704
rect 12989 7701 13001 7704
rect 13035 7701 13047 7735
rect 12989 7695 13047 7701
rect 13170 7692 13176 7744
rect 13228 7732 13234 7744
rect 13357 7735 13415 7741
rect 13357 7732 13369 7735
rect 13228 7704 13369 7732
rect 13228 7692 13234 7704
rect 13357 7701 13369 7704
rect 13403 7701 13415 7735
rect 13357 7695 13415 7701
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 15657 7735 15715 7741
rect 15657 7732 15669 7735
rect 15252 7704 15669 7732
rect 15252 7692 15258 7704
rect 15657 7701 15669 7704
rect 15703 7701 15715 7735
rect 15657 7695 15715 7701
rect 16117 7735 16175 7741
rect 16117 7701 16129 7735
rect 16163 7732 16175 7735
rect 16850 7732 16856 7744
rect 16163 7704 16856 7732
rect 16163 7701 16175 7704
rect 16117 7695 16175 7701
rect 16850 7692 16856 7704
rect 16908 7692 16914 7744
rect 18874 7692 18880 7744
rect 18932 7692 18938 7744
rect 1104 7642 21043 7664
rect 1104 7590 5894 7642
rect 5946 7590 5958 7642
rect 6010 7590 6022 7642
rect 6074 7590 6086 7642
rect 6138 7590 6150 7642
rect 6202 7590 10839 7642
rect 10891 7590 10903 7642
rect 10955 7590 10967 7642
rect 11019 7590 11031 7642
rect 11083 7590 11095 7642
rect 11147 7590 15784 7642
rect 15836 7590 15848 7642
rect 15900 7590 15912 7642
rect 15964 7590 15976 7642
rect 16028 7590 16040 7642
rect 16092 7590 20729 7642
rect 20781 7590 20793 7642
rect 20845 7590 20857 7642
rect 20909 7590 20921 7642
rect 20973 7590 20985 7642
rect 21037 7590 21043 7642
rect 1104 7568 21043 7590
rect 16117 7531 16175 7537
rect 16117 7497 16129 7531
rect 16163 7528 16175 7531
rect 16758 7528 16764 7540
rect 16163 7500 16764 7528
rect 16163 7497 16175 7500
rect 16117 7491 16175 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 16850 7488 16856 7540
rect 16908 7488 16914 7540
rect 19058 7528 19064 7540
rect 18248 7500 19064 7528
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 2593 7463 2651 7469
rect 2593 7460 2605 7463
rect 1636 7432 2605 7460
rect 1636 7420 1642 7432
rect 2593 7429 2605 7432
rect 2639 7460 2651 7463
rect 2682 7460 2688 7472
rect 2639 7432 2688 7460
rect 2639 7429 2651 7432
rect 2593 7423 2651 7429
rect 2682 7420 2688 7432
rect 2740 7420 2746 7472
rect 9585 7463 9643 7469
rect 9585 7429 9597 7463
rect 9631 7460 9643 7463
rect 10318 7460 10324 7472
rect 9631 7432 10324 7460
rect 9631 7429 9643 7432
rect 9585 7423 9643 7429
rect 10318 7420 10324 7432
rect 10376 7420 10382 7472
rect 14458 7420 14464 7472
rect 14516 7460 14522 7472
rect 14516 7432 17080 7460
rect 14516 7420 14522 7432
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 7650 7392 7656 7404
rect 4387 7364 7656 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 7650 7352 7656 7364
rect 7708 7392 7714 7404
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 7708 7364 7849 7392
rect 7708 7352 7714 7364
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7392 14059 7395
rect 14826 7392 14832 7404
rect 14047 7364 14832 7392
rect 14047 7361 14059 7364
rect 14001 7355 14059 7361
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 17052 7401 17080 7432
rect 17862 7420 17868 7472
rect 17920 7420 17926 7472
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7361 17187 7395
rect 17129 7355 17187 7361
rect 13170 7284 13176 7336
rect 13228 7324 13234 7336
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 13228 7296 14289 7324
rect 13228 7284 13234 7296
rect 14277 7293 14289 7296
rect 14323 7324 14335 7327
rect 15286 7324 15292 7336
rect 14323 7296 15292 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 15930 7284 15936 7336
rect 15988 7284 15994 7336
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7293 16359 7327
rect 17144 7324 17172 7355
rect 17402 7352 17408 7404
rect 17460 7352 17466 7404
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7392 18199 7395
rect 18248 7392 18276 7500
rect 19058 7488 19064 7500
rect 19116 7488 19122 7540
rect 18414 7420 18420 7472
rect 18472 7460 18478 7472
rect 18472 7432 19104 7460
rect 18472 7420 18478 7432
rect 18187 7364 18276 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 18598 7352 18604 7404
rect 18656 7392 18662 7404
rect 19076 7401 19104 7432
rect 18877 7395 18935 7401
rect 18877 7392 18889 7395
rect 18656 7364 18889 7392
rect 18656 7352 18662 7364
rect 18877 7361 18889 7364
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 19061 7395 19119 7401
rect 19061 7361 19073 7395
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17144 7296 18061 7324
rect 16301 7287 16359 7293
rect 18049 7293 18061 7296
rect 18095 7324 18107 7327
rect 18095 7296 18920 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 13906 7216 13912 7268
rect 13964 7256 13970 7268
rect 16316 7256 16344 7287
rect 17313 7259 17371 7265
rect 17313 7256 17325 7259
rect 13964 7228 17325 7256
rect 13964 7216 13970 7228
rect 17313 7225 17325 7228
rect 17359 7225 17371 7259
rect 17313 7219 17371 7225
rect 13814 7148 13820 7200
rect 13872 7148 13878 7200
rect 13998 7148 14004 7200
rect 14056 7188 14062 7200
rect 14185 7191 14243 7197
rect 14185 7188 14197 7191
rect 14056 7160 14197 7188
rect 14056 7148 14062 7160
rect 14185 7157 14197 7160
rect 14231 7157 14243 7191
rect 14185 7151 14243 7157
rect 14274 7148 14280 7200
rect 14332 7188 14338 7200
rect 15102 7188 15108 7200
rect 14332 7160 15108 7188
rect 14332 7148 14338 7160
rect 15102 7148 15108 7160
rect 15160 7188 15166 7200
rect 15749 7191 15807 7197
rect 15749 7188 15761 7191
rect 15160 7160 15761 7188
rect 15160 7148 15166 7160
rect 15749 7157 15761 7160
rect 15795 7157 15807 7191
rect 15749 7151 15807 7157
rect 18138 7148 18144 7200
rect 18196 7148 18202 7200
rect 18325 7191 18383 7197
rect 18325 7157 18337 7191
rect 18371 7188 18383 7191
rect 18598 7188 18604 7200
rect 18371 7160 18604 7188
rect 18371 7157 18383 7160
rect 18325 7151 18383 7157
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 18892 7197 18920 7296
rect 18877 7191 18935 7197
rect 18877 7157 18889 7191
rect 18923 7188 18935 7191
rect 19886 7188 19892 7200
rect 18923 7160 19892 7188
rect 18923 7157 18935 7160
rect 18877 7151 18935 7157
rect 19886 7148 19892 7160
rect 19944 7148 19950 7200
rect 1104 7098 20884 7120
rect 1104 7046 3422 7098
rect 3474 7046 3486 7098
rect 3538 7046 3550 7098
rect 3602 7046 3614 7098
rect 3666 7046 3678 7098
rect 3730 7046 8367 7098
rect 8419 7046 8431 7098
rect 8483 7046 8495 7098
rect 8547 7046 8559 7098
rect 8611 7046 8623 7098
rect 8675 7046 13312 7098
rect 13364 7046 13376 7098
rect 13428 7046 13440 7098
rect 13492 7046 13504 7098
rect 13556 7046 13568 7098
rect 13620 7046 18257 7098
rect 18309 7046 18321 7098
rect 18373 7046 18385 7098
rect 18437 7046 18449 7098
rect 18501 7046 18513 7098
rect 18565 7046 20884 7098
rect 1104 7024 20884 7046
rect 15841 6987 15899 6993
rect 15841 6953 15853 6987
rect 15887 6984 15899 6987
rect 15930 6984 15936 6996
rect 15887 6956 15936 6984
rect 15887 6953 15899 6956
rect 15841 6947 15899 6953
rect 11701 6919 11759 6925
rect 11701 6885 11713 6919
rect 11747 6914 11759 6919
rect 14458 6916 14464 6928
rect 11747 6886 11781 6914
rect 13556 6888 14464 6916
rect 11747 6885 11759 6886
rect 11701 6879 11759 6885
rect 4430 6808 4436 6860
rect 4488 6848 4494 6860
rect 4525 6851 4583 6857
rect 4525 6848 4537 6851
rect 4488 6820 4537 6848
rect 4488 6808 4494 6820
rect 4525 6817 4537 6820
rect 4571 6817 4583 6851
rect 11716 6848 11744 6879
rect 13556 6848 13584 6888
rect 14458 6876 14464 6888
rect 14516 6916 14522 6928
rect 14516 6888 14596 6916
rect 14516 6876 14522 6888
rect 11716 6820 13584 6848
rect 13633 6851 13691 6857
rect 4525 6811 4583 6817
rect 13633 6817 13645 6851
rect 13679 6848 13691 6851
rect 13722 6848 13728 6860
rect 13679 6820 13728 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 14568 6857 14596 6888
rect 14553 6851 14611 6857
rect 14553 6817 14565 6851
rect 14599 6817 14611 6851
rect 14553 6811 14611 6817
rect 14921 6851 14979 6857
rect 14921 6817 14933 6851
rect 14967 6848 14979 6851
rect 15856 6848 15884 6947
rect 15930 6944 15936 6956
rect 15988 6944 15994 6996
rect 19242 6848 19248 6860
rect 14967 6820 15884 6848
rect 18248 6820 19248 6848
rect 14967 6817 14979 6820
rect 14921 6811 14979 6817
rect 1578 6740 1584 6792
rect 1636 6740 1642 6792
rect 1854 6789 1860 6792
rect 1848 6743 1860 6789
rect 1854 6740 1860 6743
rect 1912 6740 1918 6792
rect 4792 6783 4850 6789
rect 4792 6749 4804 6783
rect 4838 6780 4850 6783
rect 6546 6780 6552 6792
rect 4838 6752 6552 6780
rect 4838 6749 4850 6752
rect 4792 6743 4850 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 9766 6740 9772 6792
rect 9824 6780 9830 6792
rect 10318 6780 10324 6792
rect 9824 6752 10324 6780
rect 9824 6740 9830 6752
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 10594 6789 10600 6792
rect 10588 6743 10600 6789
rect 10594 6740 10600 6743
rect 10652 6740 10658 6792
rect 13357 6783 13415 6789
rect 10704 6752 12434 6780
rect 6362 6672 6368 6724
rect 6420 6672 6426 6724
rect 8202 6672 8208 6724
rect 8260 6712 8266 6724
rect 10704 6712 10732 6752
rect 8260 6684 10732 6712
rect 12406 6712 12434 6752
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 13906 6780 13912 6792
rect 13403 6752 13912 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6780 14703 6783
rect 14826 6780 14832 6792
rect 14691 6752 14832 6780
rect 14691 6749 14703 6752
rect 14645 6743 14703 6749
rect 14826 6740 14832 6752
rect 14884 6740 14890 6792
rect 15194 6780 15200 6792
rect 14936 6752 15200 6780
rect 14936 6712 14964 6752
rect 15194 6740 15200 6752
rect 15252 6740 15258 6792
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 15657 6783 15715 6789
rect 15657 6780 15669 6783
rect 15344 6752 15669 6780
rect 15344 6740 15350 6752
rect 15657 6749 15669 6752
rect 15703 6749 15715 6783
rect 15657 6743 15715 6749
rect 18138 6740 18144 6792
rect 18196 6780 18202 6792
rect 18248 6789 18276 6820
rect 19242 6808 19248 6820
rect 19300 6848 19306 6860
rect 19300 6820 20116 6848
rect 19300 6808 19306 6820
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 18196 6752 18245 6780
rect 18196 6740 18202 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 19058 6780 19064 6792
rect 18840 6752 19064 6780
rect 18840 6740 18846 6752
rect 19058 6740 19064 6752
rect 19116 6740 19122 6792
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 19886 6740 19892 6792
rect 19944 6740 19950 6792
rect 20088 6789 20116 6820
rect 20073 6783 20131 6789
rect 20073 6749 20085 6783
rect 20119 6749 20131 6783
rect 20073 6743 20131 6749
rect 12406 6684 14964 6712
rect 15013 6715 15071 6721
rect 8260 6672 8266 6684
rect 15013 6681 15025 6715
rect 15059 6712 15071 6715
rect 15102 6712 15108 6724
rect 15059 6684 15108 6712
rect 15059 6681 15071 6684
rect 15013 6675 15071 6681
rect 15102 6672 15108 6684
rect 15160 6672 15166 6724
rect 15473 6715 15531 6721
rect 15473 6681 15485 6715
rect 15519 6681 15531 6715
rect 15473 6675 15531 6681
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 2961 6647 3019 6653
rect 2961 6644 2973 6647
rect 2188 6616 2973 6644
rect 2188 6604 2194 6616
rect 2961 6613 2973 6616
rect 3007 6613 3019 6647
rect 2961 6607 3019 6613
rect 5905 6647 5963 6653
rect 5905 6613 5917 6647
rect 5951 6644 5963 6647
rect 6914 6644 6920 6656
rect 5951 6616 6920 6644
rect 5951 6613 5963 6616
rect 5905 6607 5963 6613
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 7650 6604 7656 6656
rect 7708 6604 7714 6656
rect 12986 6604 12992 6656
rect 13044 6604 13050 6656
rect 13449 6647 13507 6653
rect 13449 6613 13461 6647
rect 13495 6644 13507 6647
rect 14369 6647 14427 6653
rect 14369 6644 14381 6647
rect 13495 6616 14381 6644
rect 13495 6613 13507 6616
rect 13449 6607 13507 6613
rect 14369 6613 14381 6616
rect 14415 6613 14427 6647
rect 14369 6607 14427 6613
rect 15194 6604 15200 6656
rect 15252 6644 15258 6656
rect 15488 6644 15516 6675
rect 17034 6672 17040 6724
rect 17092 6712 17098 6724
rect 18049 6715 18107 6721
rect 18049 6712 18061 6715
rect 17092 6684 18061 6712
rect 17092 6672 17098 6684
rect 18049 6681 18061 6684
rect 18095 6681 18107 6715
rect 18049 6675 18107 6681
rect 15252 6616 15516 6644
rect 15252 6604 15258 6616
rect 19058 6604 19064 6656
rect 19116 6644 19122 6656
rect 19429 6647 19487 6653
rect 19429 6644 19441 6647
rect 19116 6616 19441 6644
rect 19116 6604 19122 6616
rect 19429 6613 19441 6616
rect 19475 6613 19487 6647
rect 19429 6607 19487 6613
rect 1104 6554 21043 6576
rect 1104 6502 5894 6554
rect 5946 6502 5958 6554
rect 6010 6502 6022 6554
rect 6074 6502 6086 6554
rect 6138 6502 6150 6554
rect 6202 6502 10839 6554
rect 10891 6502 10903 6554
rect 10955 6502 10967 6554
rect 11019 6502 11031 6554
rect 11083 6502 11095 6554
rect 11147 6502 15784 6554
rect 15836 6502 15848 6554
rect 15900 6502 15912 6554
rect 15964 6502 15976 6554
rect 16028 6502 16040 6554
rect 16092 6502 20729 6554
rect 20781 6502 20793 6554
rect 20845 6502 20857 6554
rect 20909 6502 20921 6554
rect 20973 6502 20985 6554
rect 21037 6502 21043 6554
rect 1104 6480 21043 6502
rect 9214 6440 9220 6452
rect 4724 6412 9220 6440
rect 2952 6375 3010 6381
rect 2952 6341 2964 6375
rect 2998 6372 3010 6375
rect 4724 6372 4752 6412
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 11149 6443 11207 6449
rect 9355 6412 9996 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 2998 6344 4752 6372
rect 4792 6375 4850 6381
rect 2998 6341 3010 6344
rect 2952 6335 3010 6341
rect 4792 6341 4804 6375
rect 4838 6372 4850 6375
rect 5442 6372 5448 6384
rect 4838 6344 5448 6372
rect 4838 6341 4850 6344
rect 4792 6335 4850 6341
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 8202 6381 8208 6384
rect 8196 6372 8208 6381
rect 8163 6344 8208 6372
rect 8196 6335 8208 6344
rect 8202 6332 8208 6335
rect 8260 6332 8266 6384
rect 2682 6264 2688 6316
rect 2740 6264 2746 6316
rect 7834 6264 7840 6316
rect 7892 6304 7898 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7892 6276 7941 6304
rect 7892 6264 7898 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 9766 6264 9772 6316
rect 9824 6264 9830 6316
rect 9968 6304 9996 6412
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 13170 6440 13176 6452
rect 11195 6412 13176 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 13633 6443 13691 6449
rect 13633 6409 13645 6443
rect 13679 6440 13691 6443
rect 13814 6440 13820 6452
rect 13679 6412 13820 6440
rect 13679 6409 13691 6412
rect 13633 6403 13691 6409
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 15194 6440 15200 6452
rect 14860 6412 15200 6440
rect 10036 6375 10094 6381
rect 10036 6341 10048 6375
rect 10082 6372 10094 6375
rect 11882 6372 11888 6384
rect 10082 6344 11888 6372
rect 10082 6341 10094 6344
rect 10036 6335 10094 6341
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 14090 6372 14096 6384
rect 11992 6344 14096 6372
rect 11992 6304 12020 6344
rect 14090 6332 14096 6344
rect 14148 6332 14154 6384
rect 9968 6276 12020 6304
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 13541 6307 13599 6313
rect 13541 6304 13553 6307
rect 13228 6276 13553 6304
rect 13228 6264 13234 6276
rect 13541 6273 13553 6276
rect 13587 6304 13599 6307
rect 14860 6304 14888 6412
rect 15194 6400 15200 6412
rect 15252 6400 15258 6452
rect 15286 6400 15292 6452
rect 15344 6400 15350 6452
rect 18690 6400 18696 6452
rect 18748 6400 18754 6452
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 19797 6443 19855 6449
rect 19797 6440 19809 6443
rect 19300 6412 19809 6440
rect 19300 6400 19306 6412
rect 19797 6409 19809 6412
rect 19843 6409 19855 6443
rect 19797 6403 19855 6409
rect 15105 6375 15163 6381
rect 15105 6341 15117 6375
rect 15151 6341 15163 6375
rect 15105 6335 15163 6341
rect 13587 6276 14888 6304
rect 13587 6273 13599 6276
rect 13541 6267 13599 6273
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 4525 6239 4583 6245
rect 4525 6236 4537 6239
rect 4304 6208 4537 6236
rect 4304 6196 4310 6208
rect 4525 6205 4537 6208
rect 4571 6205 4583 6239
rect 4525 6199 4583 6205
rect 13722 6196 13728 6248
rect 13780 6196 13786 6248
rect 15120 6236 15148 6335
rect 15212 6304 15240 6400
rect 18046 6332 18052 6384
rect 18104 6372 18110 6384
rect 18104 6344 19932 6372
rect 18104 6332 18110 6344
rect 15381 6307 15439 6313
rect 15381 6304 15393 6307
rect 15212 6276 15393 6304
rect 15381 6273 15393 6276
rect 15427 6273 15439 6307
rect 15381 6267 15439 6273
rect 16942 6264 16948 6316
rect 17000 6264 17006 6316
rect 17034 6264 17040 6316
rect 17092 6264 17098 6316
rect 18693 6307 18751 6313
rect 18693 6273 18705 6307
rect 18739 6304 18751 6307
rect 18782 6304 18788 6316
rect 18739 6276 18788 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 18874 6264 18880 6316
rect 18932 6264 18938 6316
rect 19058 6264 19064 6316
rect 19116 6264 19122 6316
rect 19904 6313 19932 6344
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 19889 6307 19947 6313
rect 19889 6273 19901 6307
rect 19935 6273 19947 6307
rect 19889 6267 19947 6273
rect 17402 6236 17408 6248
rect 15028 6208 17408 6236
rect 6454 6168 6460 6180
rect 5460 6140 6460 6168
rect 4065 6103 4123 6109
rect 4065 6069 4077 6103
rect 4111 6100 4123 6103
rect 5460 6100 5488 6140
rect 6454 6128 6460 6140
rect 6512 6128 6518 6180
rect 15028 6168 15056 6208
rect 17402 6196 17408 6208
rect 17460 6236 17466 6248
rect 17770 6236 17776 6248
rect 17460 6208 17776 6236
rect 17460 6196 17466 6208
rect 17770 6196 17776 6208
rect 17828 6236 17834 6248
rect 19720 6236 19748 6267
rect 17828 6208 19748 6236
rect 17828 6196 17834 6208
rect 12360 6140 15056 6168
rect 4111 6072 5488 6100
rect 4111 6069 4123 6072
rect 4065 6063 4123 6069
rect 5902 6060 5908 6112
rect 5960 6060 5966 6112
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 12360 6100 12388 6140
rect 15102 6128 15108 6180
rect 15160 6128 15166 6180
rect 9640 6072 12388 6100
rect 9640 6060 9646 6072
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 13173 6103 13231 6109
rect 13173 6100 13185 6103
rect 12860 6072 13185 6100
rect 12860 6060 12866 6072
rect 13173 6069 13185 6072
rect 13219 6069 13231 6103
rect 13173 6063 13231 6069
rect 17221 6103 17279 6109
rect 17221 6069 17233 6103
rect 17267 6100 17279 6103
rect 17402 6100 17408 6112
rect 17267 6072 17408 6100
rect 17267 6069 17279 6072
rect 17221 6063 17279 6069
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 1104 6010 20884 6032
rect 1104 5958 3422 6010
rect 3474 5958 3486 6010
rect 3538 5958 3550 6010
rect 3602 5958 3614 6010
rect 3666 5958 3678 6010
rect 3730 5958 8367 6010
rect 8419 5958 8431 6010
rect 8483 5958 8495 6010
rect 8547 5958 8559 6010
rect 8611 5958 8623 6010
rect 8675 5958 13312 6010
rect 13364 5958 13376 6010
rect 13428 5958 13440 6010
rect 13492 5958 13504 6010
rect 13556 5958 13568 6010
rect 13620 5958 18257 6010
rect 18309 5958 18321 6010
rect 18373 5958 18385 6010
rect 18437 5958 18449 6010
rect 18501 5958 18513 6010
rect 18565 5958 20884 6010
rect 1104 5936 20884 5958
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 9582 5896 9588 5908
rect 5684 5868 9588 5896
rect 5684 5856 5690 5868
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 16393 5899 16451 5905
rect 16393 5896 16405 5899
rect 9692 5868 16405 5896
rect 1578 5652 1584 5704
rect 1636 5692 1642 5704
rect 4246 5692 4252 5704
rect 1636 5664 4252 5692
rect 1636 5652 1642 5664
rect 4246 5652 4252 5664
rect 4304 5652 4310 5704
rect 4522 5652 4528 5704
rect 4580 5652 4586 5704
rect 7098 5652 7104 5704
rect 7156 5652 7162 5704
rect 7368 5695 7426 5701
rect 7368 5661 7380 5695
rect 7414 5692 7426 5695
rect 9692 5692 9720 5868
rect 16393 5865 16405 5868
rect 16439 5865 16451 5899
rect 16393 5859 16451 5865
rect 11149 5831 11207 5837
rect 11149 5797 11161 5831
rect 11195 5828 11207 5831
rect 13906 5828 13912 5840
rect 11195 5800 13912 5828
rect 11195 5797 11207 5800
rect 11149 5791 11207 5797
rect 13906 5788 13912 5800
rect 13964 5788 13970 5840
rect 15562 5788 15568 5840
rect 15620 5828 15626 5840
rect 18782 5828 18788 5840
rect 15620 5800 18788 5828
rect 15620 5788 15626 5800
rect 18782 5788 18788 5800
rect 18840 5788 18846 5840
rect 13173 5763 13231 5769
rect 13173 5729 13185 5763
rect 13219 5760 13231 5763
rect 13630 5760 13636 5772
rect 13219 5732 13636 5760
rect 13219 5729 13231 5732
rect 13173 5723 13231 5729
rect 13630 5720 13636 5732
rect 13688 5760 13694 5772
rect 15580 5760 15608 5788
rect 13688 5732 15608 5760
rect 17037 5763 17095 5769
rect 13688 5720 13694 5732
rect 17037 5729 17049 5763
rect 17083 5760 17095 5763
rect 17402 5760 17408 5772
rect 17083 5732 17408 5760
rect 17083 5729 17095 5732
rect 17037 5723 17095 5729
rect 17402 5720 17408 5732
rect 17460 5720 17466 5772
rect 7414 5664 9720 5692
rect 7414 5661 7426 5664
rect 7368 5655 7426 5661
rect 9766 5652 9772 5704
rect 9824 5652 9830 5704
rect 10036 5695 10094 5701
rect 10036 5661 10048 5695
rect 10082 5692 10094 5695
rect 12986 5692 12992 5704
rect 10082 5664 12992 5692
rect 10082 5661 10094 5664
rect 10036 5655 10094 5661
rect 12986 5652 12992 5664
rect 13044 5652 13050 5704
rect 17310 5652 17316 5704
rect 17368 5692 17374 5704
rect 17589 5695 17647 5701
rect 17589 5692 17601 5695
rect 17368 5664 17601 5692
rect 17368 5652 17374 5664
rect 17589 5661 17601 5664
rect 17635 5661 17647 5695
rect 17589 5655 17647 5661
rect 17770 5652 17776 5704
rect 17828 5652 17834 5704
rect 16666 5624 16672 5636
rect 8496 5596 16672 5624
rect 8496 5565 8524 5596
rect 16666 5584 16672 5596
rect 16724 5624 16730 5636
rect 16761 5627 16819 5633
rect 16761 5624 16773 5627
rect 16724 5596 16773 5624
rect 16724 5584 16730 5596
rect 16761 5593 16773 5596
rect 16807 5593 16819 5627
rect 16761 5587 16819 5593
rect 8481 5559 8539 5565
rect 8481 5525 8493 5559
rect 8527 5525 8539 5559
rect 8481 5519 8539 5525
rect 11330 5516 11336 5568
rect 11388 5556 11394 5568
rect 12529 5559 12587 5565
rect 12529 5556 12541 5559
rect 11388 5528 12541 5556
rect 11388 5516 11394 5528
rect 12529 5525 12541 5528
rect 12575 5525 12587 5559
rect 12529 5519 12587 5525
rect 12894 5516 12900 5568
rect 12952 5516 12958 5568
rect 12986 5516 12992 5568
rect 13044 5516 13050 5568
rect 16853 5559 16911 5565
rect 16853 5525 16865 5559
rect 16899 5556 16911 5559
rect 17681 5559 17739 5565
rect 17681 5556 17693 5559
rect 16899 5528 17693 5556
rect 16899 5525 16911 5528
rect 16853 5519 16911 5525
rect 17681 5525 17693 5528
rect 17727 5525 17739 5559
rect 17681 5519 17739 5525
rect 1104 5466 21043 5488
rect 1104 5414 5894 5466
rect 5946 5414 5958 5466
rect 6010 5414 6022 5466
rect 6074 5414 6086 5466
rect 6138 5414 6150 5466
rect 6202 5414 10839 5466
rect 10891 5414 10903 5466
rect 10955 5414 10967 5466
rect 11019 5414 11031 5466
rect 11083 5414 11095 5466
rect 11147 5414 15784 5466
rect 15836 5414 15848 5466
rect 15900 5414 15912 5466
rect 15964 5414 15976 5466
rect 16028 5414 16040 5466
rect 16092 5414 20729 5466
rect 20781 5414 20793 5466
rect 20845 5414 20857 5466
rect 20909 5414 20921 5466
rect 20973 5414 20985 5466
rect 21037 5414 21043 5466
rect 1104 5392 21043 5414
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6914 5352 6920 5364
rect 6043 5324 6920 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 14829 5355 14887 5361
rect 14829 5352 14841 5355
rect 7024 5324 14841 5352
rect 1578 5176 1584 5228
rect 1636 5176 1642 5228
rect 1854 5225 1860 5228
rect 1848 5179 1860 5225
rect 1854 5176 1860 5179
rect 1912 5176 1918 5228
rect 4884 5219 4942 5225
rect 7024 5222 7052 5324
rect 14829 5321 14841 5324
rect 14875 5321 14887 5355
rect 14829 5315 14887 5321
rect 10036 5287 10094 5293
rect 10036 5253 10048 5287
rect 10082 5284 10094 5287
rect 11330 5284 11336 5296
rect 10082 5256 11336 5284
rect 10082 5253 10094 5256
rect 10036 5247 10094 5253
rect 11330 5244 11336 5256
rect 11388 5244 11394 5296
rect 12526 5244 12532 5296
rect 12584 5284 12590 5296
rect 12584 5256 13124 5284
rect 12584 5244 12590 5256
rect 4884 5185 4896 5219
rect 4930 5216 4942 5219
rect 6932 5216 7052 5222
rect 4930 5194 7052 5216
rect 4930 5188 6960 5194
rect 4930 5185 4942 5188
rect 4884 5179 4942 5185
rect 7098 5176 7104 5228
rect 7156 5176 7162 5228
rect 7368 5219 7426 5225
rect 7368 5185 7380 5219
rect 7414 5216 7426 5219
rect 12802 5216 12808 5228
rect 7414 5188 12808 5216
rect 7414 5185 7426 5188
rect 7368 5179 7426 5185
rect 12802 5176 12808 5188
rect 12860 5176 12866 5228
rect 13096 5225 13124 5256
rect 13630 5244 13636 5296
rect 13688 5244 13694 5296
rect 15933 5287 15991 5293
rect 15933 5253 15945 5287
rect 15979 5284 15991 5287
rect 16298 5284 16304 5296
rect 15979 5256 16304 5284
rect 15979 5253 15991 5256
rect 15933 5247 15991 5253
rect 16298 5244 16304 5256
rect 16356 5244 16362 5296
rect 17034 5244 17040 5296
rect 17092 5284 17098 5296
rect 17681 5287 17739 5293
rect 17681 5284 17693 5287
rect 17092 5256 17693 5284
rect 17092 5244 17098 5256
rect 17681 5253 17693 5256
rect 17727 5253 17739 5287
rect 17681 5247 17739 5253
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 14182 5176 14188 5228
rect 14240 5176 14246 5228
rect 14274 5176 14280 5228
rect 14332 5216 14338 5228
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 14332 5188 14381 5216
rect 14332 5176 14338 5188
rect 14369 5185 14381 5188
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 4617 5151 4675 5157
rect 4617 5148 4629 5151
rect 4304 5120 4629 5148
rect 4304 5108 4310 5120
rect 4617 5117 4629 5120
rect 4663 5117 4675 5151
rect 4617 5111 4675 5117
rect 9766 5108 9772 5160
rect 9824 5108 9830 5160
rect 11149 5083 11207 5089
rect 8404 5052 9812 5080
rect 2958 4972 2964 5024
rect 3016 4972 3022 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 8404 5012 8432 5052
rect 6972 4984 8432 5012
rect 8481 5015 8539 5021
rect 6972 4972 6978 4984
rect 8481 4981 8493 5015
rect 8527 5012 8539 5015
rect 9674 5012 9680 5024
rect 8527 4984 9680 5012
rect 8527 4981 8539 4984
rect 8481 4975 8539 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 9784 5012 9812 5052
rect 11149 5049 11161 5083
rect 11195 5080 11207 5083
rect 12986 5080 12992 5092
rect 11195 5052 12992 5080
rect 11195 5049 11207 5052
rect 11149 5043 11207 5049
rect 12986 5040 12992 5052
rect 13044 5040 13050 5092
rect 14384 5080 14412 5179
rect 14458 5176 14464 5228
rect 14516 5176 14522 5228
rect 14550 5176 14556 5228
rect 14608 5176 14614 5228
rect 15286 5176 15292 5228
rect 15344 5176 15350 5228
rect 15473 5219 15531 5225
rect 15473 5185 15485 5219
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 15565 5219 15623 5225
rect 15565 5185 15577 5219
rect 15611 5185 15623 5219
rect 15565 5179 15623 5185
rect 15488 5080 15516 5179
rect 14384 5052 15516 5080
rect 12894 5012 12900 5024
rect 9784 4984 12900 5012
rect 12894 4972 12900 4984
rect 12952 5012 12958 5024
rect 14366 5012 14372 5024
rect 12952 4984 14372 5012
rect 12952 4972 12958 4984
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 14458 4972 14464 5024
rect 14516 5012 14522 5024
rect 15580 5012 15608 5179
rect 15654 5176 15660 5228
rect 15712 5176 15718 5228
rect 17402 5176 17408 5228
rect 17460 5176 17466 5228
rect 17310 5108 17316 5160
rect 17368 5108 17374 5160
rect 17770 5108 17776 5160
rect 17828 5108 17834 5160
rect 14516 4984 15608 5012
rect 14516 4972 14522 4984
rect 17126 4972 17132 5024
rect 17184 4972 17190 5024
rect 1104 4922 20884 4944
rect 1104 4870 3422 4922
rect 3474 4870 3486 4922
rect 3538 4870 3550 4922
rect 3602 4870 3614 4922
rect 3666 4870 3678 4922
rect 3730 4870 8367 4922
rect 8419 4870 8431 4922
rect 8483 4870 8495 4922
rect 8547 4870 8559 4922
rect 8611 4870 8623 4922
rect 8675 4870 13312 4922
rect 13364 4870 13376 4922
rect 13428 4870 13440 4922
rect 13492 4870 13504 4922
rect 13556 4870 13568 4922
rect 13620 4870 18257 4922
rect 18309 4870 18321 4922
rect 18373 4870 18385 4922
rect 18437 4870 18449 4922
rect 18501 4870 18513 4922
rect 18565 4870 20884 4922
rect 1104 4848 20884 4870
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 13170 4808 13176 4820
rect 9732 4780 13176 4808
rect 9732 4768 9738 4780
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 14369 4811 14427 4817
rect 14369 4777 14381 4811
rect 14415 4808 14427 4811
rect 15286 4808 15292 4820
rect 14415 4780 15292 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 16666 4768 16672 4820
rect 16724 4808 16730 4820
rect 16942 4808 16948 4820
rect 16724 4780 16948 4808
rect 16724 4768 16730 4780
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 17310 4768 17316 4820
rect 17368 4808 17374 4820
rect 17681 4811 17739 4817
rect 17681 4808 17693 4811
rect 17368 4780 17693 4808
rect 17368 4768 17374 4780
rect 17681 4777 17693 4780
rect 17727 4777 17739 4811
rect 17681 4771 17739 4777
rect 17770 4768 17776 4820
rect 17828 4808 17834 4820
rect 18325 4811 18383 4817
rect 18325 4808 18337 4811
rect 17828 4780 18337 4808
rect 17828 4768 17834 4780
rect 18325 4777 18337 4780
rect 18371 4777 18383 4811
rect 18325 4771 18383 4777
rect 11701 4743 11759 4749
rect 11701 4709 11713 4743
rect 11747 4740 11759 4743
rect 11747 4712 12434 4740
rect 11747 4709 11759 4712
rect 11701 4703 11759 4709
rect 12406 4672 12434 4712
rect 14550 4700 14556 4752
rect 14608 4740 14614 4752
rect 15105 4743 15163 4749
rect 15105 4740 15117 4743
rect 14608 4712 15117 4740
rect 14608 4700 14614 4712
rect 15105 4709 15117 4712
rect 15151 4740 15163 4743
rect 15654 4740 15660 4752
rect 15151 4712 15660 4740
rect 15151 4709 15163 4712
rect 15105 4703 15163 4709
rect 15654 4700 15660 4712
rect 15712 4700 15718 4752
rect 17218 4740 17224 4752
rect 16592 4712 17224 4740
rect 16592 4672 16620 4712
rect 17218 4700 17224 4712
rect 17276 4700 17282 4752
rect 12406 4644 16620 4672
rect 9766 4564 9772 4616
rect 9824 4604 9830 4616
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 9824 4576 10333 4604
rect 9824 4564 9830 4576
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13044 4576 14289 4604
rect 13044 4564 13050 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 14550 4564 14556 4616
rect 14608 4604 14614 4616
rect 16592 4613 16620 4644
rect 16776 4644 17632 4672
rect 16776 4616 16804 4644
rect 15197 4607 15255 4613
rect 15197 4604 15209 4607
rect 14608 4576 15209 4604
rect 14608 4564 14614 4576
rect 15197 4573 15209 4576
rect 15243 4573 15255 4607
rect 15197 4567 15255 4573
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4573 16635 4607
rect 16577 4567 16635 4573
rect 16758 4564 16764 4616
rect 16816 4564 16822 4616
rect 17034 4564 17040 4616
rect 17092 4604 17098 4616
rect 17604 4613 17632 4644
rect 17129 4607 17187 4613
rect 17129 4604 17141 4607
rect 17092 4576 17141 4604
rect 17092 4564 17098 4576
rect 17129 4573 17141 4576
rect 17175 4573 17187 4607
rect 17129 4567 17187 4573
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 18104 4576 18245 4604
rect 18104 4564 18110 4576
rect 18233 4573 18245 4576
rect 18279 4604 18291 4607
rect 18598 4604 18604 4616
rect 18279 4576 18604 4604
rect 18279 4573 18291 4576
rect 18233 4567 18291 4573
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 10588 4539 10646 4545
rect 10588 4505 10600 4539
rect 10634 4536 10646 4539
rect 16666 4536 16672 4548
rect 10634 4508 16672 4536
rect 10634 4505 10646 4508
rect 10588 4499 10646 4505
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 16574 4428 16580 4480
rect 16632 4468 16638 4480
rect 16945 4471 17003 4477
rect 16945 4468 16957 4471
rect 16632 4440 16957 4468
rect 16632 4428 16638 4440
rect 16945 4437 16957 4440
rect 16991 4437 17003 4471
rect 16945 4431 17003 4437
rect 1104 4378 21043 4400
rect 1104 4326 5894 4378
rect 5946 4326 5958 4378
rect 6010 4326 6022 4378
rect 6074 4326 6086 4378
rect 6138 4326 6150 4378
rect 6202 4326 10839 4378
rect 10891 4326 10903 4378
rect 10955 4326 10967 4378
rect 11019 4326 11031 4378
rect 11083 4326 11095 4378
rect 11147 4326 15784 4378
rect 15836 4326 15848 4378
rect 15900 4326 15912 4378
rect 15964 4326 15976 4378
rect 16028 4326 16040 4378
rect 16092 4326 20729 4378
rect 20781 4326 20793 4378
rect 20845 4326 20857 4378
rect 20909 4326 20921 4378
rect 20973 4326 20985 4378
rect 21037 4326 21043 4378
rect 1104 4304 21043 4326
rect 1854 4224 1860 4276
rect 1912 4224 1918 4276
rect 2958 4196 2964 4208
rect 2792 4168 2964 4196
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4128 1823 4131
rect 1854 4128 1860 4140
rect 1811 4100 1860 4128
rect 1811 4097 1823 4100
rect 1765 4091 1823 4097
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4128 2007 4131
rect 2792 4128 2820 4168
rect 2958 4156 2964 4168
rect 3016 4156 3022 4208
rect 1995 4100 2820 4128
rect 3044 4131 3102 4137
rect 1995 4097 2007 4100
rect 1949 4091 2007 4097
rect 3044 4097 3056 4131
rect 3090 4128 3102 4131
rect 4062 4128 4068 4140
rect 3090 4100 4068 4128
rect 3090 4097 3102 4100
rect 3044 4091 3102 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4246 4088 4252 4140
rect 4304 4128 4310 4140
rect 4617 4131 4675 4137
rect 4617 4128 4629 4131
rect 4304 4100 4629 4128
rect 4304 4088 4310 4100
rect 4617 4097 4629 4100
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 4884 4131 4942 4137
rect 4884 4097 4896 4131
rect 4930 4128 4942 4131
rect 4930 4100 6914 4128
rect 4930 4097 4942 4100
rect 4884 4091 4942 4097
rect 1578 4020 1584 4072
rect 1636 4060 1642 4072
rect 2777 4063 2835 4069
rect 2777 4060 2789 4063
rect 1636 4032 2789 4060
rect 1636 4020 1642 4032
rect 2777 4029 2789 4032
rect 2823 4029 2835 4063
rect 2777 4023 2835 4029
rect 4154 3884 4160 3936
rect 4212 3884 4218 3936
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 6546 3924 6552 3936
rect 6043 3896 6552 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 6886 3924 6914 4100
rect 7098 4088 7104 4140
rect 7156 4088 7162 4140
rect 7368 4131 7426 4137
rect 7368 4097 7380 4131
rect 7414 4128 7426 4131
rect 9858 4128 9864 4140
rect 7414 4100 9864 4128
rect 7414 4097 7426 4100
rect 7368 4091 7426 4097
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 10036 4131 10094 4137
rect 10036 4097 10048 4131
rect 10082 4128 10094 4131
rect 10082 4100 12434 4128
rect 10082 4097 10094 4100
rect 10036 4091 10094 4097
rect 9766 4020 9772 4072
rect 9824 4020 9830 4072
rect 12406 4060 12434 4100
rect 13906 4088 13912 4140
rect 13964 4088 13970 4140
rect 14090 4088 14096 4140
rect 14148 4088 14154 4140
rect 14366 4088 14372 4140
rect 14424 4088 14430 4140
rect 14458 4088 14464 4140
rect 14516 4088 14522 4140
rect 14642 4088 14648 4140
rect 14700 4088 14706 4140
rect 17126 4060 17132 4072
rect 12406 4032 17132 4060
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 11149 3995 11207 4001
rect 11149 3961 11161 3995
rect 11195 3992 11207 3995
rect 16758 3992 16764 4004
rect 11195 3964 16764 3992
rect 11195 3961 11207 3964
rect 11149 3955 11207 3961
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 7282 3924 7288 3936
rect 6886 3896 7288 3924
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3924 8539 3927
rect 8754 3924 8760 3936
rect 8527 3896 8760 3924
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 1104 3834 20884 3856
rect 1104 3782 3422 3834
rect 3474 3782 3486 3834
rect 3538 3782 3550 3834
rect 3602 3782 3614 3834
rect 3666 3782 3678 3834
rect 3730 3782 8367 3834
rect 8419 3782 8431 3834
rect 8483 3782 8495 3834
rect 8547 3782 8559 3834
rect 8611 3782 8623 3834
rect 8675 3782 13312 3834
rect 13364 3782 13376 3834
rect 13428 3782 13440 3834
rect 13492 3782 13504 3834
rect 13556 3782 13568 3834
rect 13620 3782 18257 3834
rect 18309 3782 18321 3834
rect 18373 3782 18385 3834
rect 18437 3782 18449 3834
rect 18501 3782 18513 3834
rect 18565 3782 20884 3834
rect 1104 3760 20884 3782
rect 4062 3680 4068 3732
rect 4120 3680 4126 3732
rect 8205 3723 8263 3729
rect 8205 3689 8217 3723
rect 8251 3720 8263 3723
rect 12342 3720 12348 3732
rect 8251 3692 12348 3720
rect 8251 3689 8263 3692
rect 8205 3683 8263 3689
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 12452 3692 14228 3720
rect 3234 3612 3240 3664
rect 3292 3652 3298 3664
rect 6362 3652 6368 3664
rect 3292 3624 6368 3652
rect 3292 3612 3298 3624
rect 6362 3612 6368 3624
rect 6420 3612 6426 3664
rect 12452 3661 12480 3692
rect 12437 3655 12495 3661
rect 12437 3621 12449 3655
rect 12483 3621 12495 3655
rect 14200 3652 14228 3692
rect 14274 3680 14280 3732
rect 14332 3680 14338 3732
rect 16666 3680 16672 3732
rect 16724 3680 16730 3732
rect 17129 3723 17187 3729
rect 17129 3689 17141 3723
rect 17175 3720 17187 3723
rect 17402 3720 17408 3732
rect 17175 3692 17408 3720
rect 17175 3689 17187 3692
rect 17129 3683 17187 3689
rect 17402 3680 17408 3692
rect 17460 3720 17466 3732
rect 17773 3723 17831 3729
rect 17773 3720 17785 3723
rect 17460 3692 17785 3720
rect 17460 3680 17466 3692
rect 17773 3689 17785 3692
rect 17819 3689 17831 3723
rect 17773 3683 17831 3689
rect 17034 3652 17040 3664
rect 12437 3615 12495 3621
rect 12912 3624 13124 3652
rect 14200 3624 17040 3652
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 1765 3587 1823 3593
rect 1765 3584 1777 3587
rect 1636 3556 1777 3584
rect 1636 3544 1642 3556
rect 1765 3553 1777 3556
rect 1811 3553 1823 3587
rect 1765 3547 1823 3553
rect 4157 3587 4215 3593
rect 4157 3553 4169 3587
rect 4203 3584 4215 3587
rect 5626 3584 5632 3596
rect 4203 3556 5632 3584
rect 4203 3553 4215 3556
rect 4157 3547 4215 3553
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 12912 3584 12940 3624
rect 12400 3556 12940 3584
rect 12400 3544 12406 3556
rect 12986 3544 12992 3596
rect 13044 3544 13050 3596
rect 1854 3476 1860 3528
rect 1912 3516 1918 3528
rect 1912 3488 4016 3516
rect 1912 3476 1918 3488
rect 2032 3451 2090 3457
rect 2032 3417 2044 3451
rect 2078 3448 2090 3451
rect 2406 3448 2412 3460
rect 2078 3420 2412 3448
rect 2078 3417 2090 3420
rect 2032 3411 2090 3417
rect 2406 3408 2412 3420
rect 2464 3408 2470 3460
rect 3988 3457 4016 3488
rect 4246 3476 4252 3528
rect 4304 3476 4310 3528
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 6914 3516 6920 3528
rect 6871 3488 6920 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 6914 3476 6920 3488
rect 6972 3516 6978 3528
rect 9122 3516 9128 3528
rect 6972 3488 9128 3516
rect 6972 3476 6978 3488
rect 9122 3476 9128 3488
rect 9180 3516 9186 3528
rect 9766 3516 9772 3528
rect 9180 3488 9772 3516
rect 9180 3476 9186 3488
rect 9766 3476 9772 3488
rect 9824 3516 9830 3528
rect 11057 3519 11115 3525
rect 11057 3516 11069 3519
rect 9824 3488 11069 3516
rect 9824 3476 9830 3488
rect 11057 3485 11069 3488
rect 11103 3485 11115 3519
rect 13096 3516 13124 3624
rect 17034 3612 17040 3624
rect 17092 3652 17098 3664
rect 17678 3652 17684 3664
rect 17092 3624 17684 3652
rect 17092 3612 17098 3624
rect 17678 3612 17684 3624
rect 17736 3612 17742 3664
rect 13357 3587 13415 3593
rect 13357 3553 13369 3587
rect 13403 3584 13415 3587
rect 13906 3584 13912 3596
rect 13403 3556 13912 3584
rect 13403 3553 13415 3556
rect 13357 3547 13415 3553
rect 13906 3544 13912 3556
rect 13964 3584 13970 3596
rect 13964 3556 14780 3584
rect 13964 3544 13970 3556
rect 14752 3528 14780 3556
rect 14826 3544 14832 3596
rect 14884 3544 14890 3596
rect 16868 3556 18092 3584
rect 13161 3519 13219 3525
rect 13161 3516 13173 3519
rect 13096 3488 13173 3516
rect 11057 3479 11115 3485
rect 13161 3485 13173 3488
rect 13207 3485 13219 3519
rect 13161 3479 13219 3485
rect 14134 3488 14320 3516
rect 3973 3451 4031 3457
rect 3973 3417 3985 3451
rect 4019 3448 4031 3451
rect 4522 3448 4528 3460
rect 4019 3420 4528 3448
rect 4019 3417 4031 3420
rect 3973 3411 4031 3417
rect 4522 3408 4528 3420
rect 4580 3408 4586 3460
rect 7092 3451 7150 3457
rect 7092 3417 7104 3451
rect 7138 3448 7150 3451
rect 9392 3451 9450 3457
rect 7138 3420 9352 3448
rect 7138 3417 7150 3420
rect 7092 3411 7150 3417
rect 3142 3340 3148 3392
rect 3200 3340 3206 3392
rect 9324 3380 9352 3420
rect 9392 3417 9404 3451
rect 9438 3448 9450 3451
rect 11324 3451 11382 3457
rect 9438 3420 11284 3448
rect 9438 3417 9450 3420
rect 9392 3411 9450 3417
rect 10134 3380 10140 3392
rect 9324 3352 10140 3380
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 10502 3340 10508 3392
rect 10560 3340 10566 3392
rect 11256 3380 11284 3420
rect 11324 3417 11336 3451
rect 11370 3448 11382 3451
rect 14134 3448 14162 3488
rect 11370 3420 14162 3448
rect 14292 3448 14320 3488
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 14424 3488 14473 3516
rect 14424 3476 14430 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3516 14611 3519
rect 14642 3516 14648 3528
rect 14599 3488 14648 3516
rect 14599 3485 14611 3488
rect 14553 3479 14611 3485
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 14792 3488 14933 3516
rect 14792 3476 14798 3488
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 14921 3479 14979 3485
rect 15378 3476 15384 3528
rect 15436 3476 15442 3528
rect 15562 3476 15568 3528
rect 15620 3476 15626 3528
rect 16868 3525 16896 3556
rect 18064 3528 18092 3556
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 16942 3476 16948 3528
rect 17000 3476 17006 3528
rect 17218 3476 17224 3528
rect 17276 3476 17282 3528
rect 17678 3476 17684 3528
rect 17736 3476 17742 3528
rect 17954 3476 17960 3528
rect 18012 3476 18018 3528
rect 18046 3476 18052 3528
rect 18104 3476 18110 3528
rect 18233 3451 18291 3457
rect 18233 3448 18245 3451
rect 14292 3420 18245 3448
rect 11370 3417 11382 3420
rect 11324 3411 11382 3417
rect 18233 3417 18245 3420
rect 18279 3417 18291 3451
rect 18233 3411 18291 3417
rect 13262 3380 13268 3392
rect 11256 3352 13268 3380
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 14550 3340 14556 3392
rect 14608 3380 14614 3392
rect 14645 3383 14703 3389
rect 14645 3380 14657 3383
rect 14608 3352 14657 3380
rect 14608 3340 14614 3352
rect 14645 3349 14657 3352
rect 14691 3349 14703 3383
rect 14645 3343 14703 3349
rect 15470 3340 15476 3392
rect 15528 3340 15534 3392
rect 1104 3290 21043 3312
rect 1104 3238 5894 3290
rect 5946 3238 5958 3290
rect 6010 3238 6022 3290
rect 6074 3238 6086 3290
rect 6138 3238 6150 3290
rect 6202 3238 10839 3290
rect 10891 3238 10903 3290
rect 10955 3238 10967 3290
rect 11019 3238 11031 3290
rect 11083 3238 11095 3290
rect 11147 3238 15784 3290
rect 15836 3238 15848 3290
rect 15900 3238 15912 3290
rect 15964 3238 15976 3290
rect 16028 3238 16040 3290
rect 16092 3238 20729 3290
rect 20781 3238 20793 3290
rect 20845 3238 20857 3290
rect 20909 3238 20921 3290
rect 20973 3238 20985 3290
rect 21037 3238 21043 3290
rect 1104 3216 21043 3238
rect 7009 3179 7067 3185
rect 4356 3148 6914 3176
rect 1578 3068 1584 3120
rect 1636 3108 1642 3120
rect 4356 3117 4384 3148
rect 2593 3111 2651 3117
rect 2593 3108 2605 3111
rect 1636 3080 2605 3108
rect 1636 3068 1642 3080
rect 2593 3077 2605 3080
rect 2639 3077 2651 3111
rect 2593 3071 2651 3077
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3077 4399 3111
rect 4341 3071 4399 3077
rect 5350 3068 5356 3120
rect 5408 3108 5414 3120
rect 5629 3111 5687 3117
rect 5629 3108 5641 3111
rect 5408 3080 5641 3108
rect 5408 3068 5414 3080
rect 5629 3077 5641 3080
rect 5675 3077 5687 3111
rect 6886 3108 6914 3148
rect 7009 3145 7021 3179
rect 7055 3176 7067 3179
rect 7282 3176 7288 3188
rect 7055 3148 7288 3176
rect 7055 3145 7067 3148
rect 7009 3139 7067 3145
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 9122 3136 9128 3188
rect 9180 3136 9186 3188
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 9916 3148 10057 3176
rect 9916 3136 9922 3148
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 10045 3139 10103 3145
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 12253 3179 12311 3185
rect 12253 3176 12265 3179
rect 10192 3148 12265 3176
rect 10192 3136 10198 3148
rect 12253 3145 12265 3148
rect 12299 3145 12311 3179
rect 12253 3139 12311 3145
rect 7650 3108 7656 3120
rect 6886 3080 7656 3108
rect 5629 3071 5687 3077
rect 7650 3068 7656 3080
rect 7708 3108 7714 3120
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 7708 3080 7849 3108
rect 7708 3068 7714 3080
rect 7837 3077 7849 3080
rect 7883 3077 7895 3111
rect 7837 3071 7895 3077
rect 11054 3068 11060 3120
rect 11112 3108 11118 3120
rect 13541 3111 13599 3117
rect 13541 3108 13553 3111
rect 11112 3080 13553 3108
rect 11112 3068 11118 3080
rect 13541 3077 13553 3080
rect 13587 3077 13599 3111
rect 15470 3108 15476 3120
rect 13541 3071 13599 3077
rect 13740 3080 15476 3108
rect 5442 3000 5448 3052
rect 5500 3000 5506 3052
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 6546 3040 6552 3052
rect 5583 3012 6552 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 6822 3000 6828 3052
rect 6880 3000 6886 3052
rect 9950 3000 9956 3052
rect 10008 3040 10014 3052
rect 10229 3043 10287 3049
rect 10229 3040 10241 3043
rect 10008 3012 10241 3040
rect 10008 3000 10014 3012
rect 10229 3009 10241 3012
rect 10275 3009 10287 3043
rect 10229 3003 10287 3009
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3040 12311 3043
rect 12434 3040 12440 3052
rect 12299 3012 12440 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 12434 3000 12440 3012
rect 12492 3000 12498 3052
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3040 12587 3043
rect 13630 3040 13636 3052
rect 12575 3012 13636 3040
rect 12575 3009 12587 3012
rect 12529 3003 12587 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 13740 3049 13768 3080
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3040 14703 3043
rect 14734 3040 14740 3052
rect 14691 3012 14740 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 14826 3000 14832 3052
rect 14884 3000 14890 3052
rect 15654 3000 15660 3052
rect 15712 3000 15718 3052
rect 15930 3000 15936 3052
rect 15988 3000 15994 3052
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 5258 2932 5264 2984
rect 5316 2932 5322 2984
rect 5997 2975 6055 2981
rect 5997 2941 6009 2975
rect 6043 2972 6055 2975
rect 6730 2972 6736 2984
rect 6043 2944 6736 2972
rect 6043 2941 6055 2944
rect 5997 2935 6055 2941
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 10505 2975 10563 2981
rect 10505 2972 10517 2975
rect 8812 2944 10517 2972
rect 8812 2932 8818 2944
rect 10505 2941 10517 2944
rect 10551 2941 10563 2975
rect 10505 2935 10563 2941
rect 5626 2864 5632 2916
rect 5684 2904 5690 2916
rect 6641 2907 6699 2913
rect 6641 2904 6653 2907
rect 5684 2876 6653 2904
rect 5684 2864 5690 2876
rect 6641 2873 6653 2876
rect 6687 2873 6699 2907
rect 6641 2867 6699 2873
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 10413 2839 10471 2845
rect 10413 2836 10425 2839
rect 9732 2808 10425 2836
rect 9732 2796 9738 2808
rect 10413 2805 10425 2808
rect 10459 2805 10471 2839
rect 10520 2836 10548 2935
rect 13998 2932 14004 2984
rect 14056 2932 14062 2984
rect 14550 2932 14556 2984
rect 14608 2972 14614 2984
rect 15838 2972 15844 2984
rect 14608 2944 15844 2972
rect 14608 2932 14614 2944
rect 15838 2932 15844 2944
rect 15896 2972 15902 2984
rect 16132 2972 16160 3003
rect 16942 3000 16948 3052
rect 17000 3040 17006 3052
rect 17129 3043 17187 3049
rect 17129 3040 17141 3043
rect 17000 3012 17141 3040
rect 17000 3000 17006 3012
rect 17129 3009 17141 3012
rect 17175 3009 17187 3043
rect 17129 3003 17187 3009
rect 15896 2944 16160 2972
rect 15896 2932 15902 2944
rect 17218 2932 17224 2984
rect 17276 2932 17282 2984
rect 17497 2975 17555 2981
rect 17497 2941 17509 2975
rect 17543 2972 17555 2975
rect 17954 2972 17960 2984
rect 17543 2944 17960 2972
rect 17543 2941 17555 2944
rect 17497 2935 17555 2941
rect 17954 2932 17960 2944
rect 18012 2932 18018 2984
rect 12345 2907 12403 2913
rect 12345 2873 12357 2907
rect 12391 2904 12403 2907
rect 13909 2907 13967 2913
rect 13909 2904 13921 2907
rect 12391 2876 13921 2904
rect 12391 2873 12403 2876
rect 12345 2867 12403 2873
rect 13909 2873 13921 2876
rect 13955 2904 13967 2907
rect 14461 2907 14519 2913
rect 14461 2904 14473 2907
rect 13955 2876 14473 2904
rect 13955 2873 13967 2876
rect 13909 2867 13967 2873
rect 14461 2873 14473 2876
rect 14507 2873 14519 2907
rect 14461 2867 14519 2873
rect 12618 2836 12624 2848
rect 10520 2808 12624 2836
rect 10413 2799 10471 2805
rect 12618 2796 12624 2808
rect 12676 2836 12682 2848
rect 12986 2836 12992 2848
rect 12676 2808 12992 2836
rect 12676 2796 12682 2808
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 13320 2808 15485 2836
rect 13320 2796 13326 2808
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 1104 2746 20884 2768
rect 1104 2694 3422 2746
rect 3474 2694 3486 2746
rect 3538 2694 3550 2746
rect 3602 2694 3614 2746
rect 3666 2694 3678 2746
rect 3730 2694 8367 2746
rect 8419 2694 8431 2746
rect 8483 2694 8495 2746
rect 8547 2694 8559 2746
rect 8611 2694 8623 2746
rect 8675 2694 13312 2746
rect 13364 2694 13376 2746
rect 13428 2694 13440 2746
rect 13492 2694 13504 2746
rect 13556 2694 13568 2746
rect 13620 2694 18257 2746
rect 18309 2694 18321 2746
rect 18373 2694 18385 2746
rect 18437 2694 18449 2746
rect 18501 2694 18513 2746
rect 18565 2694 20884 2746
rect 1104 2672 20884 2694
rect 2406 2592 2412 2644
rect 2464 2592 2470 2644
rect 4246 2592 4252 2644
rect 4304 2632 4310 2644
rect 4341 2635 4399 2641
rect 4341 2632 4353 2635
rect 4304 2604 4353 2632
rect 4304 2592 4310 2604
rect 4341 2601 4353 2604
rect 4387 2601 4399 2635
rect 4341 2595 4399 2601
rect 5353 2635 5411 2641
rect 5353 2601 5365 2635
rect 5399 2632 5411 2635
rect 5442 2632 5448 2644
rect 5399 2604 5448 2632
rect 5399 2601 5411 2604
rect 5353 2595 5411 2601
rect 1673 2567 1731 2573
rect 1673 2533 1685 2567
rect 1719 2533 1731 2567
rect 5368 2564 5396 2595
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 5537 2635 5595 2641
rect 5537 2601 5549 2635
rect 5583 2632 5595 2635
rect 5626 2632 5632 2644
rect 5583 2604 5632 2632
rect 5583 2601 5595 2604
rect 5537 2595 5595 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6733 2635 6791 2641
rect 6733 2601 6745 2635
rect 6779 2632 6791 2635
rect 6822 2632 6828 2644
rect 6779 2604 6828 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 9950 2632 9956 2644
rect 8619 2604 9956 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 12434 2592 12440 2644
rect 12492 2592 12498 2644
rect 14826 2592 14832 2644
rect 14884 2592 14890 2644
rect 15565 2635 15623 2641
rect 15565 2601 15577 2635
rect 15611 2632 15623 2635
rect 15654 2632 15660 2644
rect 15611 2604 15660 2632
rect 15611 2601 15623 2604
rect 15565 2595 15623 2601
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 1673 2527 1731 2533
rect 4356 2536 5396 2564
rect 11149 2567 11207 2573
rect 1688 2496 1716 2527
rect 2777 2499 2835 2505
rect 1688 2468 2636 2496
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 1854 2428 1860 2440
rect 1719 2400 1860 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 2608 2437 2636 2468
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 2823 2468 3188 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2397 2651 2431
rect 2593 2391 2651 2397
rect 1964 2360 1992 2391
rect 2792 2360 2820 2459
rect 3160 2440 3188 2468
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 2958 2428 2964 2440
rect 2915 2400 2964 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 1964 2332 2820 2360
rect 1857 2295 1915 2301
rect 1857 2261 1869 2295
rect 1903 2292 1915 2295
rect 2884 2292 2912 2391
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 3142 2388 3148 2440
rect 3200 2428 3206 2440
rect 4065 2431 4123 2437
rect 4065 2428 4077 2431
rect 3200 2400 4077 2428
rect 3200 2388 3206 2400
rect 4065 2397 4077 2400
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 4080 2360 4108 2391
rect 4154 2388 4160 2440
rect 4212 2428 4218 2440
rect 4356 2437 4384 2536
rect 11149 2533 11161 2567
rect 11195 2564 11207 2567
rect 13998 2564 14004 2576
rect 11195 2536 14004 2564
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 13998 2524 14004 2536
rect 14056 2524 14062 2576
rect 9674 2496 9680 2508
rect 8312 2468 9680 2496
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 4212 2400 4353 2428
rect 4212 2388 4218 2400
rect 4341 2397 4353 2400
rect 4387 2397 4399 2431
rect 4341 2391 4399 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 4580 2400 6561 2428
rect 4580 2388 4586 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 4080 2332 4292 2360
rect 4154 2292 4160 2304
rect 1903 2264 4160 2292
rect 1903 2261 1915 2264
rect 1857 2255 1915 2261
rect 4154 2252 4160 2264
rect 4212 2252 4218 2304
rect 4264 2292 4292 2332
rect 4430 2320 4436 2372
rect 4488 2360 4494 2372
rect 5169 2363 5227 2369
rect 5169 2360 5181 2363
rect 4488 2332 5181 2360
rect 4488 2320 4494 2332
rect 5169 2329 5181 2332
rect 5215 2360 5227 2363
rect 5258 2360 5264 2372
rect 5215 2332 5264 2360
rect 5215 2329 5227 2332
rect 5169 2323 5227 2329
rect 5258 2320 5264 2332
rect 5316 2320 5322 2372
rect 5350 2320 5356 2372
rect 5408 2369 5414 2372
rect 5408 2363 5427 2369
rect 5415 2329 5427 2363
rect 6564 2360 6592 2391
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 8312 2437 8340 2468
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 9766 2456 9772 2508
rect 9824 2456 9830 2508
rect 14090 2496 14096 2508
rect 12728 2468 14096 2496
rect 8297 2431 8355 2437
rect 8297 2428 8309 2431
rect 6788 2400 8309 2428
rect 6788 2388 6794 2400
rect 8297 2397 8309 2400
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8754 2428 8760 2440
rect 8435 2400 8760 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 8573 2363 8631 2369
rect 8573 2360 8585 2363
rect 6564 2332 8585 2360
rect 5408 2323 5427 2329
rect 8573 2329 8585 2332
rect 8619 2329 8631 2363
rect 9692 2360 9720 2456
rect 10036 2431 10094 2437
rect 10036 2397 10048 2431
rect 10082 2428 10094 2431
rect 11054 2428 11060 2440
rect 10082 2400 11060 2428
rect 10082 2397 10094 2400
rect 10036 2391 10094 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 12437 2431 12495 2437
rect 12437 2428 12449 2431
rect 12400 2400 12449 2428
rect 12400 2388 12406 2400
rect 12437 2397 12449 2400
rect 12483 2397 12495 2431
rect 12437 2391 12495 2397
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 12728 2437 12756 2468
rect 14090 2456 14096 2468
rect 14148 2496 14154 2508
rect 14844 2496 14872 2592
rect 14148 2468 14872 2496
rect 14148 2456 14154 2468
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2397 12771 2431
rect 12713 2391 12771 2397
rect 12728 2360 12756 2391
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15620 2400 15761 2428
rect 15620 2388 15626 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 15930 2388 15936 2440
rect 15988 2428 15994 2440
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 15988 2400 16037 2428
rect 15988 2388 15994 2400
rect 16025 2397 16037 2400
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 9692 2332 12756 2360
rect 8573 2323 8631 2329
rect 5408 2320 5414 2323
rect 13998 2320 14004 2372
rect 14056 2360 14062 2372
rect 14642 2360 14648 2372
rect 14056 2332 14648 2360
rect 14056 2320 14062 2332
rect 14642 2320 14648 2332
rect 14700 2320 14706 2372
rect 14734 2320 14740 2372
rect 14792 2360 14798 2372
rect 14845 2363 14903 2369
rect 14845 2360 14857 2363
rect 14792 2332 14857 2360
rect 14792 2320 14798 2332
rect 14845 2329 14857 2332
rect 14891 2329 14903 2363
rect 15378 2360 15384 2372
rect 14845 2323 14903 2329
rect 15028 2332 15384 2360
rect 5368 2292 5396 2320
rect 15028 2301 15056 2332
rect 15378 2320 15384 2332
rect 15436 2360 15442 2372
rect 16040 2360 16068 2391
rect 15436 2332 16068 2360
rect 15436 2320 15442 2332
rect 4264 2264 5396 2292
rect 15013 2295 15071 2301
rect 15013 2261 15025 2295
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 15838 2252 15844 2304
rect 15896 2292 15902 2304
rect 15933 2295 15991 2301
rect 15933 2292 15945 2295
rect 15896 2264 15945 2292
rect 15896 2252 15902 2264
rect 15933 2261 15945 2264
rect 15979 2261 15991 2295
rect 15933 2255 15991 2261
rect 1104 2202 21043 2224
rect 1104 2150 5894 2202
rect 5946 2150 5958 2202
rect 6010 2150 6022 2202
rect 6074 2150 6086 2202
rect 6138 2150 6150 2202
rect 6202 2150 10839 2202
rect 10891 2150 10903 2202
rect 10955 2150 10967 2202
rect 11019 2150 11031 2202
rect 11083 2150 11095 2202
rect 11147 2150 15784 2202
rect 15836 2150 15848 2202
rect 15900 2150 15912 2202
rect 15964 2150 15976 2202
rect 16028 2150 16040 2202
rect 16092 2150 20729 2202
rect 20781 2150 20793 2202
rect 20845 2150 20857 2202
rect 20909 2150 20921 2202
rect 20973 2150 20985 2202
rect 21037 2150 21043 2202
rect 1104 2128 21043 2150
<< via1 >>
rect 5894 19558 5946 19610
rect 5958 19558 6010 19610
rect 6022 19558 6074 19610
rect 6086 19558 6138 19610
rect 6150 19558 6202 19610
rect 10839 19558 10891 19610
rect 10903 19558 10955 19610
rect 10967 19558 11019 19610
rect 11031 19558 11083 19610
rect 11095 19558 11147 19610
rect 15784 19558 15836 19610
rect 15848 19558 15900 19610
rect 15912 19558 15964 19610
rect 15976 19558 16028 19610
rect 16040 19558 16092 19610
rect 20729 19558 20781 19610
rect 20793 19558 20845 19610
rect 20857 19558 20909 19610
rect 20921 19558 20973 19610
rect 20985 19558 21037 19610
rect 3422 19014 3474 19066
rect 3486 19014 3538 19066
rect 3550 19014 3602 19066
rect 3614 19014 3666 19066
rect 3678 19014 3730 19066
rect 8367 19014 8419 19066
rect 8431 19014 8483 19066
rect 8495 19014 8547 19066
rect 8559 19014 8611 19066
rect 8623 19014 8675 19066
rect 13312 19014 13364 19066
rect 13376 19014 13428 19066
rect 13440 19014 13492 19066
rect 13504 19014 13556 19066
rect 13568 19014 13620 19066
rect 18257 19014 18309 19066
rect 18321 19014 18373 19066
rect 18385 19014 18437 19066
rect 18449 19014 18501 19066
rect 18513 19014 18565 19066
rect 2504 18708 2556 18760
rect 940 18640 992 18692
rect 5894 18470 5946 18522
rect 5958 18470 6010 18522
rect 6022 18470 6074 18522
rect 6086 18470 6138 18522
rect 6150 18470 6202 18522
rect 10839 18470 10891 18522
rect 10903 18470 10955 18522
rect 10967 18470 11019 18522
rect 11031 18470 11083 18522
rect 11095 18470 11147 18522
rect 15784 18470 15836 18522
rect 15848 18470 15900 18522
rect 15912 18470 15964 18522
rect 15976 18470 16028 18522
rect 16040 18470 16092 18522
rect 20729 18470 20781 18522
rect 20793 18470 20845 18522
rect 20857 18470 20909 18522
rect 20921 18470 20973 18522
rect 20985 18470 21037 18522
rect 3422 17926 3474 17978
rect 3486 17926 3538 17978
rect 3550 17926 3602 17978
rect 3614 17926 3666 17978
rect 3678 17926 3730 17978
rect 8367 17926 8419 17978
rect 8431 17926 8483 17978
rect 8495 17926 8547 17978
rect 8559 17926 8611 17978
rect 8623 17926 8675 17978
rect 13312 17926 13364 17978
rect 13376 17926 13428 17978
rect 13440 17926 13492 17978
rect 13504 17926 13556 17978
rect 13568 17926 13620 17978
rect 18257 17926 18309 17978
rect 18321 17926 18373 17978
rect 18385 17926 18437 17978
rect 18449 17926 18501 17978
rect 18513 17926 18565 17978
rect 5894 17382 5946 17434
rect 5958 17382 6010 17434
rect 6022 17382 6074 17434
rect 6086 17382 6138 17434
rect 6150 17382 6202 17434
rect 10839 17382 10891 17434
rect 10903 17382 10955 17434
rect 10967 17382 11019 17434
rect 11031 17382 11083 17434
rect 11095 17382 11147 17434
rect 15784 17382 15836 17434
rect 15848 17382 15900 17434
rect 15912 17382 15964 17434
rect 15976 17382 16028 17434
rect 16040 17382 16092 17434
rect 20729 17382 20781 17434
rect 20793 17382 20845 17434
rect 20857 17382 20909 17434
rect 20921 17382 20973 17434
rect 20985 17382 21037 17434
rect 3056 17144 3108 17196
rect 4068 17144 4120 17196
rect 6000 17144 6052 17196
rect 8116 17144 8168 17196
rect 3332 17008 3384 17060
rect 7748 17076 7800 17128
rect 4068 17008 4120 17060
rect 3148 16940 3200 16992
rect 5448 16983 5500 16992
rect 5448 16949 5457 16983
rect 5457 16949 5491 16983
rect 5491 16949 5500 16983
rect 5448 16940 5500 16949
rect 7288 16940 7340 16992
rect 3422 16838 3474 16890
rect 3486 16838 3538 16890
rect 3550 16838 3602 16890
rect 3614 16838 3666 16890
rect 3678 16838 3730 16890
rect 8367 16838 8419 16890
rect 8431 16838 8483 16890
rect 8495 16838 8547 16890
rect 8559 16838 8611 16890
rect 8623 16838 8675 16890
rect 13312 16838 13364 16890
rect 13376 16838 13428 16890
rect 13440 16838 13492 16890
rect 13504 16838 13556 16890
rect 13568 16838 13620 16890
rect 18257 16838 18309 16890
rect 18321 16838 18373 16890
rect 18385 16838 18437 16890
rect 18449 16838 18501 16890
rect 18513 16838 18565 16890
rect 5816 16736 5868 16788
rect 4068 16668 4120 16720
rect 3148 16575 3200 16584
rect 3148 16541 3157 16575
rect 3157 16541 3191 16575
rect 3191 16541 3200 16575
rect 3148 16532 3200 16541
rect 3240 16575 3292 16584
rect 3240 16541 3249 16575
rect 3249 16541 3283 16575
rect 3283 16541 3292 16575
rect 3240 16532 3292 16541
rect 4068 16532 4120 16584
rect 6000 16668 6052 16720
rect 7564 16668 7616 16720
rect 5448 16600 5500 16652
rect 5724 16643 5776 16652
rect 5724 16609 5733 16643
rect 5733 16609 5767 16643
rect 5767 16609 5776 16643
rect 5724 16600 5776 16609
rect 5816 16575 5868 16584
rect 5816 16541 5825 16575
rect 5825 16541 5859 16575
rect 5859 16541 5868 16575
rect 5816 16532 5868 16541
rect 6000 16532 6052 16584
rect 4344 16464 4396 16516
rect 3148 16439 3200 16448
rect 3148 16405 3157 16439
rect 3157 16405 3191 16439
rect 3191 16405 3200 16439
rect 3148 16396 3200 16405
rect 4804 16439 4856 16448
rect 4804 16405 4813 16439
rect 4813 16405 4847 16439
rect 4847 16405 4856 16439
rect 4804 16396 4856 16405
rect 5264 16396 5316 16448
rect 7196 16464 7248 16516
rect 7748 16532 7800 16584
rect 11336 16532 11388 16584
rect 7380 16464 7432 16516
rect 7472 16396 7524 16448
rect 8116 16464 8168 16516
rect 11612 16439 11664 16448
rect 11612 16405 11621 16439
rect 11621 16405 11655 16439
rect 11655 16405 11664 16439
rect 11612 16396 11664 16405
rect 13084 16396 13136 16448
rect 5894 16294 5946 16346
rect 5958 16294 6010 16346
rect 6022 16294 6074 16346
rect 6086 16294 6138 16346
rect 6150 16294 6202 16346
rect 10839 16294 10891 16346
rect 10903 16294 10955 16346
rect 10967 16294 11019 16346
rect 11031 16294 11083 16346
rect 11095 16294 11147 16346
rect 15784 16294 15836 16346
rect 15848 16294 15900 16346
rect 15912 16294 15964 16346
rect 15976 16294 16028 16346
rect 16040 16294 16092 16346
rect 20729 16294 20781 16346
rect 20793 16294 20845 16346
rect 20857 16294 20909 16346
rect 20921 16294 20973 16346
rect 20985 16294 21037 16346
rect 8024 16192 8076 16244
rect 3240 16124 3292 16176
rect 3332 16167 3384 16176
rect 3332 16133 3341 16167
rect 3341 16133 3375 16167
rect 3375 16133 3384 16167
rect 3332 16124 3384 16133
rect 12716 16124 12768 16176
rect 5448 16099 5500 16108
rect 5448 16065 5457 16099
rect 5457 16065 5491 16099
rect 5491 16065 5500 16099
rect 5448 16056 5500 16065
rect 7288 16099 7340 16108
rect 7288 16065 7297 16099
rect 7297 16065 7331 16099
rect 7331 16065 7340 16099
rect 7288 16056 7340 16065
rect 7472 16099 7524 16108
rect 7472 16065 7481 16099
rect 7481 16065 7515 16099
rect 7515 16065 7524 16099
rect 7472 16056 7524 16065
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 8944 16056 8996 16108
rect 4804 15988 4856 16040
rect 5632 15988 5684 16040
rect 5816 15988 5868 16040
rect 6828 15988 6880 16040
rect 11612 16056 11664 16108
rect 12440 16056 12492 16108
rect 10416 15988 10468 16040
rect 11704 15988 11756 16040
rect 11888 16031 11940 16040
rect 11888 15997 11897 16031
rect 11897 15997 11931 16031
rect 11931 15997 11940 16031
rect 11888 15988 11940 15997
rect 13084 16099 13136 16108
rect 13084 16065 13093 16099
rect 13093 16065 13127 16099
rect 13127 16065 13136 16099
rect 13084 16056 13136 16065
rect 14464 16124 14516 16176
rect 13176 15988 13228 16040
rect 14372 16056 14424 16108
rect 13728 15988 13780 16040
rect 14648 16099 14700 16108
rect 14648 16065 14658 16099
rect 14658 16065 14692 16099
rect 14692 16065 14700 16099
rect 14648 16056 14700 16065
rect 14832 16099 14884 16108
rect 14832 16065 14841 16099
rect 14841 16065 14875 16099
rect 14875 16065 14884 16099
rect 14832 16056 14884 16065
rect 15016 16099 15068 16108
rect 15016 16065 15030 16099
rect 15030 16065 15064 16099
rect 15064 16065 15068 16099
rect 15016 16056 15068 16065
rect 15108 15988 15160 16040
rect 11612 15920 11664 15972
rect 15660 15920 15712 15972
rect 3240 15852 3292 15904
rect 6736 15852 6788 15904
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 3422 15750 3474 15802
rect 3486 15750 3538 15802
rect 3550 15750 3602 15802
rect 3614 15750 3666 15802
rect 3678 15750 3730 15802
rect 8367 15750 8419 15802
rect 8431 15750 8483 15802
rect 8495 15750 8547 15802
rect 8559 15750 8611 15802
rect 8623 15750 8675 15802
rect 13312 15750 13364 15802
rect 13376 15750 13428 15802
rect 13440 15750 13492 15802
rect 13504 15750 13556 15802
rect 13568 15750 13620 15802
rect 18257 15750 18309 15802
rect 18321 15750 18373 15802
rect 18385 15750 18437 15802
rect 18449 15750 18501 15802
rect 18513 15750 18565 15802
rect 3976 15648 4028 15700
rect 5632 15691 5684 15700
rect 5632 15657 5641 15691
rect 5641 15657 5675 15691
rect 5675 15657 5684 15691
rect 5632 15648 5684 15657
rect 4068 15580 4120 15632
rect 5724 15580 5776 15632
rect 6828 15691 6880 15700
rect 6828 15657 6837 15691
rect 6837 15657 6871 15691
rect 6871 15657 6880 15691
rect 6828 15648 6880 15657
rect 7380 15691 7432 15700
rect 7380 15657 7389 15691
rect 7389 15657 7423 15691
rect 7423 15657 7432 15691
rect 7380 15648 7432 15657
rect 11244 15648 11296 15700
rect 7104 15580 7156 15632
rect 3332 15512 3384 15564
rect 4344 15512 4396 15564
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 3240 15487 3292 15496
rect 3240 15453 3249 15487
rect 3249 15453 3283 15487
rect 3283 15453 3292 15487
rect 3240 15444 3292 15453
rect 3976 15444 4028 15496
rect 4712 15444 4764 15496
rect 6920 15555 6972 15564
rect 6920 15521 6929 15555
rect 6929 15521 6963 15555
rect 6963 15521 6972 15555
rect 6920 15512 6972 15521
rect 3700 15376 3752 15428
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 10324 15555 10376 15564
rect 10324 15521 10333 15555
rect 10333 15521 10367 15555
rect 10367 15521 10376 15555
rect 10324 15512 10376 15521
rect 6368 15376 6420 15428
rect 8116 15376 8168 15428
rect 10232 15444 10284 15496
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 11152 15580 11204 15632
rect 11796 15580 11848 15632
rect 12440 15580 12492 15632
rect 13176 15580 13228 15632
rect 15016 15648 15068 15700
rect 15108 15648 15160 15700
rect 18144 15648 18196 15700
rect 11060 15444 11112 15496
rect 11152 15376 11204 15428
rect 3332 15308 3384 15360
rect 4988 15308 5040 15360
rect 9864 15351 9916 15360
rect 9864 15317 9873 15351
rect 9873 15317 9907 15351
rect 9907 15317 9916 15351
rect 9864 15308 9916 15317
rect 10692 15308 10744 15360
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 11520 15487 11572 15496
rect 11520 15453 11529 15487
rect 11529 15453 11563 15487
rect 11563 15453 11572 15487
rect 11520 15444 11572 15453
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 12900 15444 12952 15496
rect 11888 15376 11940 15428
rect 14648 15444 14700 15496
rect 15016 15444 15068 15496
rect 13820 15376 13872 15428
rect 12992 15308 13044 15360
rect 16764 15623 16816 15632
rect 16764 15589 16773 15623
rect 16773 15589 16807 15623
rect 16807 15589 16816 15623
rect 16764 15580 16816 15589
rect 15292 15487 15344 15496
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 18880 15512 18932 15564
rect 15660 15487 15712 15496
rect 15660 15453 15669 15487
rect 15669 15453 15703 15487
rect 15703 15453 15712 15487
rect 15660 15444 15712 15453
rect 16488 15444 16540 15496
rect 17408 15444 17460 15496
rect 15660 15308 15712 15360
rect 17868 15308 17920 15360
rect 5894 15206 5946 15258
rect 5958 15206 6010 15258
rect 6022 15206 6074 15258
rect 6086 15206 6138 15258
rect 6150 15206 6202 15258
rect 10839 15206 10891 15258
rect 10903 15206 10955 15258
rect 10967 15206 11019 15258
rect 11031 15206 11083 15258
rect 11095 15206 11147 15258
rect 15784 15206 15836 15258
rect 15848 15206 15900 15258
rect 15912 15206 15964 15258
rect 15976 15206 16028 15258
rect 16040 15206 16092 15258
rect 20729 15206 20781 15258
rect 20793 15206 20845 15258
rect 20857 15206 20909 15258
rect 20921 15206 20973 15258
rect 20985 15206 21037 15258
rect 3148 15104 3200 15156
rect 2228 15036 2280 15088
rect 3240 15036 3292 15088
rect 3700 15011 3752 15020
rect 3700 14977 3709 15011
rect 3709 14977 3743 15011
rect 3743 14977 3752 15011
rect 3700 14968 3752 14977
rect 3976 15011 4028 15020
rect 3976 14977 3985 15011
rect 3985 14977 4019 15011
rect 4019 14977 4028 15011
rect 3976 14968 4028 14977
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 4712 15011 4764 15020
rect 4712 14977 4721 15011
rect 4721 14977 4755 15011
rect 4755 14977 4764 15011
rect 4712 14968 4764 14977
rect 6828 15104 6880 15156
rect 7748 15104 7800 15156
rect 6368 15036 6420 15088
rect 8024 15079 8076 15088
rect 8024 15045 8033 15079
rect 8033 15045 8067 15079
rect 8067 15045 8076 15079
rect 8024 15036 8076 15045
rect 6644 14968 6696 15020
rect 7840 14968 7892 15020
rect 10232 15104 10284 15156
rect 10324 15104 10376 15156
rect 11428 15104 11480 15156
rect 11520 15104 11572 15156
rect 11796 15104 11848 15156
rect 14832 15104 14884 15156
rect 9128 15036 9180 15088
rect 12808 15036 12860 15088
rect 16856 15104 16908 15156
rect 9864 14968 9916 15020
rect 11796 14968 11848 15020
rect 11888 15011 11940 15020
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 12256 15011 12308 15020
rect 12256 14977 12265 15011
rect 12265 14977 12299 15011
rect 12299 14977 12308 15011
rect 12256 14968 12308 14977
rect 2320 14943 2372 14952
rect 2320 14909 2329 14943
rect 2329 14909 2363 14943
rect 2363 14909 2372 14943
rect 2320 14900 2372 14909
rect 3056 14900 3108 14952
rect 4988 14943 5040 14952
rect 4988 14909 4997 14943
rect 4997 14909 5031 14943
rect 5031 14909 5040 14943
rect 4988 14900 5040 14909
rect 6460 14900 6512 14952
rect 6920 14900 6972 14952
rect 8944 14943 8996 14952
rect 8944 14909 8953 14943
rect 8953 14909 8987 14943
rect 8987 14909 8996 14943
rect 8944 14900 8996 14909
rect 4804 14875 4856 14884
rect 4804 14841 4813 14875
rect 4813 14841 4847 14875
rect 4847 14841 4856 14875
rect 4804 14832 4856 14841
rect 9220 14832 9272 14884
rect 2044 14764 2096 14816
rect 4252 14807 4304 14816
rect 4252 14773 4261 14807
rect 4261 14773 4295 14807
rect 4295 14773 4304 14807
rect 4252 14764 4304 14773
rect 4896 14807 4948 14816
rect 4896 14773 4905 14807
rect 4905 14773 4939 14807
rect 4939 14773 4948 14807
rect 4896 14764 4948 14773
rect 8852 14764 8904 14816
rect 11244 14900 11296 14952
rect 12164 14943 12216 14952
rect 12164 14909 12173 14943
rect 12173 14909 12207 14943
rect 12207 14909 12216 14943
rect 12164 14900 12216 14909
rect 11704 14832 11756 14884
rect 12808 14900 12860 14952
rect 13636 14968 13688 15020
rect 14832 15011 14884 15020
rect 14832 14977 14841 15011
rect 14841 14977 14875 15011
rect 14875 14977 14884 15011
rect 14832 14968 14884 14977
rect 15200 14968 15252 15020
rect 15752 15011 15804 15020
rect 15752 14977 15761 15011
rect 15761 14977 15795 15011
rect 15795 14977 15804 15011
rect 15752 14968 15804 14977
rect 16764 14968 16816 15020
rect 18604 14968 18656 15020
rect 18972 15011 19024 15020
rect 18972 14977 18981 15011
rect 18981 14977 19015 15011
rect 19015 14977 19024 15011
rect 18972 14968 19024 14977
rect 19248 15011 19300 15020
rect 19248 14977 19257 15011
rect 19257 14977 19291 15011
rect 19291 14977 19300 15011
rect 19248 14968 19300 14977
rect 13084 14900 13136 14952
rect 15568 14943 15620 14952
rect 15568 14909 15577 14943
rect 15577 14909 15611 14943
rect 15611 14909 15620 14943
rect 15568 14900 15620 14909
rect 15384 14832 15436 14884
rect 17132 14943 17184 14952
rect 17132 14909 17141 14943
rect 17141 14909 17175 14943
rect 17175 14909 17184 14943
rect 17132 14900 17184 14909
rect 17592 14943 17644 14952
rect 17592 14909 17601 14943
rect 17601 14909 17635 14943
rect 17635 14909 17644 14943
rect 17592 14900 17644 14909
rect 17408 14875 17460 14884
rect 17408 14841 17417 14875
rect 17417 14841 17451 14875
rect 17451 14841 17460 14875
rect 17408 14832 17460 14841
rect 18880 14832 18932 14884
rect 12072 14764 12124 14816
rect 12624 14764 12676 14816
rect 13084 14764 13136 14816
rect 13176 14807 13228 14816
rect 13176 14773 13185 14807
rect 13185 14773 13219 14807
rect 13219 14773 13228 14807
rect 13176 14764 13228 14773
rect 15660 14764 15712 14816
rect 18052 14764 18104 14816
rect 3422 14662 3474 14714
rect 3486 14662 3538 14714
rect 3550 14662 3602 14714
rect 3614 14662 3666 14714
rect 3678 14662 3730 14714
rect 8367 14662 8419 14714
rect 8431 14662 8483 14714
rect 8495 14662 8547 14714
rect 8559 14662 8611 14714
rect 8623 14662 8675 14714
rect 13312 14662 13364 14714
rect 13376 14662 13428 14714
rect 13440 14662 13492 14714
rect 13504 14662 13556 14714
rect 13568 14662 13620 14714
rect 18257 14662 18309 14714
rect 18321 14662 18373 14714
rect 18385 14662 18437 14714
rect 18449 14662 18501 14714
rect 18513 14662 18565 14714
rect 13176 14560 13228 14612
rect 14372 14560 14424 14612
rect 12256 14492 12308 14544
rect 14648 14492 14700 14544
rect 14832 14560 14884 14612
rect 14924 14492 14976 14544
rect 19248 14560 19300 14612
rect 8944 14424 8996 14476
rect 13728 14424 13780 14476
rect 6460 14356 6512 14408
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 9220 14399 9272 14408
rect 9220 14365 9262 14399
rect 9262 14365 9272 14399
rect 9220 14356 9272 14365
rect 9588 14356 9640 14408
rect 11704 14356 11756 14408
rect 11888 14356 11940 14408
rect 12256 14399 12308 14408
rect 12256 14365 12265 14399
rect 12265 14365 12299 14399
rect 12299 14365 12308 14399
rect 12256 14356 12308 14365
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 12900 14356 12952 14408
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 14832 14356 14884 14408
rect 15292 14356 15344 14408
rect 5724 14288 5776 14340
rect 6920 14263 6972 14272
rect 6920 14229 6929 14263
rect 6929 14229 6963 14263
rect 6963 14229 6972 14263
rect 6920 14220 6972 14229
rect 7104 14331 7156 14340
rect 7104 14297 7113 14331
rect 7113 14297 7147 14331
rect 7147 14297 7156 14331
rect 7104 14288 7156 14297
rect 11244 14331 11296 14340
rect 11244 14297 11253 14331
rect 11253 14297 11287 14331
rect 11287 14297 11296 14331
rect 11244 14288 11296 14297
rect 14556 14288 14608 14340
rect 16580 14356 16632 14408
rect 9220 14220 9272 14272
rect 9312 14263 9364 14272
rect 9312 14229 9321 14263
rect 9321 14229 9355 14263
rect 9355 14229 9364 14263
rect 9312 14220 9364 14229
rect 11612 14220 11664 14272
rect 11796 14220 11848 14272
rect 12992 14220 13044 14272
rect 15476 14220 15528 14272
rect 16120 14288 16172 14340
rect 17592 14399 17644 14408
rect 17592 14365 17601 14399
rect 17601 14365 17635 14399
rect 17635 14365 17644 14399
rect 17592 14356 17644 14365
rect 18144 14399 18196 14408
rect 18144 14365 18153 14399
rect 18153 14365 18187 14399
rect 18187 14365 18196 14399
rect 18144 14356 18196 14365
rect 18604 14424 18656 14476
rect 19892 14424 19944 14476
rect 19984 14399 20036 14408
rect 19984 14365 19993 14399
rect 19993 14365 20027 14399
rect 20027 14365 20036 14399
rect 19984 14356 20036 14365
rect 17408 14220 17460 14272
rect 18144 14220 18196 14272
rect 19616 14263 19668 14272
rect 19616 14229 19625 14263
rect 19625 14229 19659 14263
rect 19659 14229 19668 14263
rect 19616 14220 19668 14229
rect 5894 14118 5946 14170
rect 5958 14118 6010 14170
rect 6022 14118 6074 14170
rect 6086 14118 6138 14170
rect 6150 14118 6202 14170
rect 10839 14118 10891 14170
rect 10903 14118 10955 14170
rect 10967 14118 11019 14170
rect 11031 14118 11083 14170
rect 11095 14118 11147 14170
rect 15784 14118 15836 14170
rect 15848 14118 15900 14170
rect 15912 14118 15964 14170
rect 15976 14118 16028 14170
rect 16040 14118 16092 14170
rect 20729 14118 20781 14170
rect 20793 14118 20845 14170
rect 20857 14118 20909 14170
rect 20921 14118 20973 14170
rect 20985 14118 21037 14170
rect 1768 14016 1820 14068
rect 2044 14059 2096 14068
rect 2044 14025 2053 14059
rect 2053 14025 2087 14059
rect 2087 14025 2096 14059
rect 2044 14016 2096 14025
rect 9312 14016 9364 14068
rect 4804 13948 4856 14000
rect 2044 13880 2096 13932
rect 3332 13880 3384 13932
rect 2320 13812 2372 13864
rect 2412 13744 2464 13796
rect 3884 13923 3936 13932
rect 3884 13889 3893 13923
rect 3893 13889 3927 13923
rect 3927 13889 3936 13923
rect 3884 13880 3936 13889
rect 3792 13812 3844 13864
rect 5264 13923 5316 13932
rect 5264 13889 5273 13923
rect 5273 13889 5307 13923
rect 5307 13889 5316 13923
rect 5264 13880 5316 13889
rect 5356 13812 5408 13864
rect 11888 14016 11940 14068
rect 12072 14016 12124 14068
rect 9680 13948 9732 14000
rect 11612 13880 11664 13932
rect 8760 13812 8812 13864
rect 11336 13812 11388 13864
rect 11428 13812 11480 13864
rect 11888 13880 11940 13932
rect 12072 13923 12124 13932
rect 12072 13889 12081 13923
rect 12081 13889 12115 13923
rect 12115 13889 12124 13923
rect 12072 13880 12124 13889
rect 12532 14016 12584 14068
rect 12808 14016 12860 14068
rect 14464 14016 14516 14068
rect 11796 13812 11848 13864
rect 12808 13812 12860 13864
rect 5448 13744 5500 13796
rect 9036 13744 9088 13796
rect 12440 13744 12492 13796
rect 12992 13880 13044 13932
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 13728 13880 13780 13932
rect 14648 14059 14700 14068
rect 14648 14025 14657 14059
rect 14657 14025 14691 14059
rect 14691 14025 14700 14059
rect 14648 14016 14700 14025
rect 15568 14016 15620 14068
rect 14464 13812 14516 13864
rect 13636 13744 13688 13796
rect 3332 13719 3384 13728
rect 3332 13685 3341 13719
rect 3341 13685 3375 13719
rect 3375 13685 3384 13719
rect 3332 13676 3384 13685
rect 11704 13719 11756 13728
rect 11704 13685 11713 13719
rect 11713 13685 11747 13719
rect 11747 13685 11756 13719
rect 11704 13676 11756 13685
rect 12992 13676 13044 13728
rect 16212 13923 16264 13932
rect 16212 13889 16221 13923
rect 16221 13889 16255 13923
rect 16255 13889 16264 13923
rect 16212 13880 16264 13889
rect 16488 13880 16540 13932
rect 17776 13923 17828 13932
rect 17776 13889 17785 13923
rect 17785 13889 17819 13923
rect 17819 13889 17828 13923
rect 17776 13880 17828 13889
rect 18052 13991 18104 14000
rect 18052 13957 18061 13991
rect 18061 13957 18095 13991
rect 18095 13957 18104 13991
rect 18052 13948 18104 13957
rect 18144 13991 18196 14000
rect 18144 13957 18153 13991
rect 18153 13957 18187 13991
rect 18187 13957 18196 13991
rect 18144 13948 18196 13957
rect 19892 13880 19944 13932
rect 17684 13855 17736 13864
rect 17684 13821 17693 13855
rect 17693 13821 17727 13855
rect 17727 13821 17736 13855
rect 17684 13812 17736 13821
rect 16856 13744 16908 13796
rect 17592 13744 17644 13796
rect 16672 13676 16724 13728
rect 17500 13719 17552 13728
rect 17500 13685 17509 13719
rect 17509 13685 17543 13719
rect 17543 13685 17552 13719
rect 17500 13676 17552 13685
rect 3422 13574 3474 13626
rect 3486 13574 3538 13626
rect 3550 13574 3602 13626
rect 3614 13574 3666 13626
rect 3678 13574 3730 13626
rect 8367 13574 8419 13626
rect 8431 13574 8483 13626
rect 8495 13574 8547 13626
rect 8559 13574 8611 13626
rect 8623 13574 8675 13626
rect 13312 13574 13364 13626
rect 13376 13574 13428 13626
rect 13440 13574 13492 13626
rect 13504 13574 13556 13626
rect 13568 13574 13620 13626
rect 18257 13574 18309 13626
rect 18321 13574 18373 13626
rect 18385 13574 18437 13626
rect 18449 13574 18501 13626
rect 18513 13574 18565 13626
rect 3884 13472 3936 13524
rect 13084 13472 13136 13524
rect 16396 13472 16448 13524
rect 16488 13515 16540 13524
rect 16488 13481 16497 13515
rect 16497 13481 16531 13515
rect 16531 13481 16540 13515
rect 16488 13472 16540 13481
rect 17684 13515 17736 13524
rect 17684 13481 17693 13515
rect 17693 13481 17727 13515
rect 17727 13481 17736 13515
rect 17684 13472 17736 13481
rect 19892 13515 19944 13524
rect 19892 13481 19901 13515
rect 19901 13481 19935 13515
rect 19935 13481 19944 13515
rect 19892 13472 19944 13481
rect 2412 13379 2464 13388
rect 2412 13345 2421 13379
rect 2421 13345 2455 13379
rect 2455 13345 2464 13379
rect 2412 13336 2464 13345
rect 4896 13336 4948 13388
rect 5448 13379 5500 13388
rect 5448 13345 5457 13379
rect 5457 13345 5491 13379
rect 5491 13345 5500 13379
rect 5448 13336 5500 13345
rect 2320 13200 2372 13252
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4160 13268 4212 13277
rect 6920 13336 6972 13388
rect 9680 13447 9732 13456
rect 9680 13413 9689 13447
rect 9689 13413 9723 13447
rect 9723 13413 9732 13447
rect 9680 13404 9732 13413
rect 12164 13404 12216 13456
rect 13176 13404 13228 13456
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 7380 13336 7432 13388
rect 8944 13336 8996 13388
rect 8024 13268 8076 13320
rect 8300 13268 8352 13320
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 11428 13268 11480 13320
rect 11612 13379 11664 13388
rect 11612 13345 11621 13379
rect 11621 13345 11655 13379
rect 11655 13345 11664 13379
rect 18880 13404 18932 13456
rect 11612 13336 11664 13345
rect 11796 13268 11848 13320
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 12992 13268 13044 13277
rect 13636 13268 13688 13320
rect 17500 13336 17552 13388
rect 15476 13268 15528 13320
rect 16304 13311 16356 13320
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 16580 13311 16632 13320
rect 16580 13277 16589 13311
rect 16589 13277 16623 13311
rect 16623 13277 16632 13311
rect 16580 13268 16632 13277
rect 17040 13268 17092 13320
rect 18144 13379 18196 13388
rect 18144 13345 18153 13379
rect 18153 13345 18187 13379
rect 18187 13345 18196 13379
rect 18144 13336 18196 13345
rect 17684 13268 17736 13320
rect 18052 13311 18104 13320
rect 18052 13277 18061 13311
rect 18061 13277 18095 13311
rect 18095 13277 18104 13311
rect 18052 13268 18104 13277
rect 19708 13268 19760 13320
rect 1676 13132 1728 13184
rect 2228 13175 2280 13184
rect 2228 13141 2237 13175
rect 2237 13141 2271 13175
rect 2271 13141 2280 13175
rect 2228 13132 2280 13141
rect 3148 13132 3200 13184
rect 6920 13243 6972 13252
rect 6920 13209 6955 13243
rect 6955 13209 6972 13243
rect 6920 13200 6972 13209
rect 11520 13200 11572 13252
rect 12256 13200 12308 13252
rect 5080 13132 5132 13184
rect 5816 13132 5868 13184
rect 6276 13132 6328 13184
rect 6736 13132 6788 13184
rect 11336 13175 11388 13184
rect 11336 13141 11345 13175
rect 11345 13141 11379 13175
rect 11379 13141 11388 13175
rect 11336 13132 11388 13141
rect 12900 13132 12952 13184
rect 14188 13132 14240 13184
rect 15292 13243 15344 13252
rect 15292 13209 15301 13243
rect 15301 13209 15335 13243
rect 15335 13209 15344 13243
rect 15292 13200 15344 13209
rect 15660 13132 15712 13184
rect 15936 13132 15988 13184
rect 19616 13200 19668 13252
rect 5894 13030 5946 13082
rect 5958 13030 6010 13082
rect 6022 13030 6074 13082
rect 6086 13030 6138 13082
rect 6150 13030 6202 13082
rect 10839 13030 10891 13082
rect 10903 13030 10955 13082
rect 10967 13030 11019 13082
rect 11031 13030 11083 13082
rect 11095 13030 11147 13082
rect 15784 13030 15836 13082
rect 15848 13030 15900 13082
rect 15912 13030 15964 13082
rect 15976 13030 16028 13082
rect 16040 13030 16092 13082
rect 20729 13030 20781 13082
rect 20793 13030 20845 13082
rect 20857 13030 20909 13082
rect 20921 13030 20973 13082
rect 20985 13030 21037 13082
rect 3148 12928 3200 12980
rect 5080 12971 5132 12980
rect 5080 12937 5089 12971
rect 5089 12937 5123 12971
rect 5123 12937 5132 12971
rect 5080 12928 5132 12937
rect 8760 12928 8812 12980
rect 2228 12860 2280 12912
rect 2780 12860 2832 12912
rect 3976 12860 4028 12912
rect 4804 12860 4856 12912
rect 2044 12792 2096 12844
rect 2688 12835 2740 12844
rect 2688 12801 2697 12835
rect 2697 12801 2731 12835
rect 2731 12801 2740 12835
rect 2688 12792 2740 12801
rect 4160 12792 4212 12844
rect 6276 12792 6328 12844
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 8024 12835 8076 12844
rect 8024 12801 8033 12835
rect 8033 12801 8067 12835
rect 8067 12801 8076 12835
rect 8024 12792 8076 12801
rect 9128 12928 9180 12980
rect 12716 12928 12768 12980
rect 9036 12903 9088 12912
rect 9036 12869 9045 12903
rect 9045 12869 9079 12903
rect 9079 12869 9088 12903
rect 9036 12860 9088 12869
rect 12440 12860 12492 12912
rect 13084 12860 13136 12912
rect 14096 12860 14148 12912
rect 15292 12860 15344 12912
rect 9312 12792 9364 12844
rect 10784 12792 10836 12844
rect 12992 12792 13044 12844
rect 3056 12656 3108 12708
rect 3792 12724 3844 12776
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 7380 12767 7432 12776
rect 7380 12733 7389 12767
rect 7389 12733 7423 12767
rect 7423 12733 7432 12767
rect 7380 12724 7432 12733
rect 8300 12724 8352 12776
rect 9128 12767 9180 12776
rect 9128 12733 9137 12767
rect 9137 12733 9171 12767
rect 9171 12733 9180 12767
rect 9128 12724 9180 12733
rect 11336 12656 11388 12708
rect 12808 12724 12860 12776
rect 15108 12724 15160 12776
rect 16304 12928 16356 12980
rect 17684 12928 17736 12980
rect 18696 12928 18748 12980
rect 19248 12928 19300 12980
rect 16396 12860 16448 12912
rect 17040 12903 17092 12912
rect 17040 12869 17051 12903
rect 17051 12869 17092 12903
rect 17040 12860 17092 12869
rect 17132 12860 17184 12912
rect 18052 12860 18104 12912
rect 17316 12792 17368 12844
rect 17868 12792 17920 12844
rect 18604 12792 18656 12844
rect 19248 12835 19300 12844
rect 19248 12801 19257 12835
rect 19257 12801 19291 12835
rect 19291 12801 19300 12835
rect 19248 12792 19300 12801
rect 19708 12792 19760 12844
rect 19340 12724 19392 12776
rect 4620 12631 4672 12640
rect 4620 12597 4629 12631
rect 4629 12597 4663 12631
rect 4663 12597 4672 12631
rect 4620 12588 4672 12597
rect 7932 12588 7984 12640
rect 8116 12588 8168 12640
rect 10508 12588 10560 12640
rect 12532 12588 12584 12640
rect 12808 12588 12860 12640
rect 15292 12656 15344 12708
rect 15752 12656 15804 12708
rect 18972 12656 19024 12708
rect 13636 12631 13688 12640
rect 13636 12597 13645 12631
rect 13645 12597 13679 12631
rect 13679 12597 13688 12631
rect 13636 12588 13688 12597
rect 17040 12631 17092 12640
rect 17040 12597 17049 12631
rect 17049 12597 17083 12631
rect 17083 12597 17092 12631
rect 17040 12588 17092 12597
rect 20076 12631 20128 12640
rect 20076 12597 20085 12631
rect 20085 12597 20119 12631
rect 20119 12597 20128 12631
rect 20076 12588 20128 12597
rect 3422 12486 3474 12538
rect 3486 12486 3538 12538
rect 3550 12486 3602 12538
rect 3614 12486 3666 12538
rect 3678 12486 3730 12538
rect 8367 12486 8419 12538
rect 8431 12486 8483 12538
rect 8495 12486 8547 12538
rect 8559 12486 8611 12538
rect 8623 12486 8675 12538
rect 13312 12486 13364 12538
rect 13376 12486 13428 12538
rect 13440 12486 13492 12538
rect 13504 12486 13556 12538
rect 13568 12486 13620 12538
rect 18257 12486 18309 12538
rect 18321 12486 18373 12538
rect 18385 12486 18437 12538
rect 18449 12486 18501 12538
rect 18513 12486 18565 12538
rect 6736 12427 6788 12436
rect 6736 12393 6745 12427
rect 6745 12393 6779 12427
rect 6779 12393 6788 12427
rect 6736 12384 6788 12393
rect 7104 12384 7156 12436
rect 7840 12384 7892 12436
rect 9128 12384 9180 12436
rect 11244 12384 11296 12436
rect 12532 12384 12584 12436
rect 13636 12384 13688 12436
rect 14372 12384 14424 12436
rect 15016 12384 15068 12436
rect 15752 12384 15804 12436
rect 17316 12384 17368 12436
rect 17776 12384 17828 12436
rect 2320 12316 2372 12368
rect 4252 12248 4304 12300
rect 12716 12316 12768 12368
rect 11520 12248 11572 12300
rect 14740 12291 14792 12300
rect 14740 12257 14749 12291
rect 14749 12257 14783 12291
rect 14783 12257 14792 12291
rect 14740 12248 14792 12257
rect 16580 12248 16632 12300
rect 3056 12180 3108 12232
rect 4068 12180 4120 12232
rect 6736 12223 6788 12232
rect 6736 12189 6745 12223
rect 6745 12189 6779 12223
rect 6779 12189 6788 12223
rect 6736 12180 6788 12189
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 10416 12180 10468 12232
rect 11336 12223 11388 12232
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11336 12180 11388 12189
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 13176 12180 13228 12232
rect 14096 12180 14148 12232
rect 14280 12180 14332 12232
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 14556 12223 14608 12232
rect 14556 12189 14566 12223
rect 14566 12189 14600 12223
rect 14600 12189 14608 12223
rect 14556 12180 14608 12189
rect 2136 12112 2188 12164
rect 2412 12112 2464 12164
rect 4528 12112 4580 12164
rect 10784 12112 10836 12164
rect 14648 12112 14700 12164
rect 15292 12223 15344 12232
rect 15292 12189 15301 12223
rect 15301 12189 15335 12223
rect 15335 12189 15344 12223
rect 15292 12180 15344 12189
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15476 12180 15528 12189
rect 17316 12180 17368 12232
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 18696 12248 18748 12300
rect 19984 12316 20036 12368
rect 18236 12180 18288 12232
rect 18604 12180 18656 12232
rect 19064 12180 19116 12232
rect 20076 12223 20128 12232
rect 20076 12189 20085 12223
rect 20085 12189 20119 12223
rect 20119 12189 20128 12223
rect 20076 12180 20128 12189
rect 4436 12044 4488 12096
rect 4804 12044 4856 12096
rect 7288 12044 7340 12096
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 13176 12044 13228 12096
rect 14004 12044 14056 12096
rect 15200 12044 15252 12096
rect 16488 12044 16540 12096
rect 16580 12044 16632 12096
rect 19340 12112 19392 12164
rect 5894 11942 5946 11994
rect 5958 11942 6010 11994
rect 6022 11942 6074 11994
rect 6086 11942 6138 11994
rect 6150 11942 6202 11994
rect 10839 11942 10891 11994
rect 10903 11942 10955 11994
rect 10967 11942 11019 11994
rect 11031 11942 11083 11994
rect 11095 11942 11147 11994
rect 15784 11942 15836 11994
rect 15848 11942 15900 11994
rect 15912 11942 15964 11994
rect 15976 11942 16028 11994
rect 16040 11942 16092 11994
rect 20729 11942 20781 11994
rect 20793 11942 20845 11994
rect 20857 11942 20909 11994
rect 20921 11942 20973 11994
rect 20985 11942 21037 11994
rect 3332 11840 3384 11892
rect 4436 11883 4488 11892
rect 4436 11849 4445 11883
rect 4445 11849 4479 11883
rect 4479 11849 4488 11883
rect 4436 11840 4488 11849
rect 7196 11840 7248 11892
rect 3056 11772 3108 11824
rect 4896 11772 4948 11824
rect 2964 11704 3016 11756
rect 3884 11704 3936 11756
rect 2136 11636 2188 11688
rect 3056 11679 3108 11688
rect 3056 11645 3065 11679
rect 3065 11645 3099 11679
rect 3099 11645 3108 11679
rect 3056 11636 3108 11645
rect 1952 11568 2004 11620
rect 2688 11568 2740 11620
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 4988 11704 5040 11756
rect 5356 11815 5408 11824
rect 5356 11781 5365 11815
rect 5365 11781 5399 11815
rect 5399 11781 5408 11815
rect 5356 11772 5408 11781
rect 5816 11704 5868 11756
rect 6736 11636 6788 11688
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 11244 11840 11296 11892
rect 11796 11883 11848 11892
rect 11796 11849 11805 11883
rect 11805 11849 11839 11883
rect 11839 11849 11848 11883
rect 11796 11840 11848 11849
rect 13820 11840 13872 11892
rect 16028 11840 16080 11892
rect 9496 11772 9548 11824
rect 11704 11772 11756 11824
rect 12072 11815 12124 11824
rect 12072 11781 12081 11815
rect 12081 11781 12115 11815
rect 12115 11781 12124 11815
rect 12072 11772 12124 11781
rect 2136 11543 2188 11552
rect 2136 11509 2145 11543
rect 2145 11509 2179 11543
rect 2179 11509 2188 11543
rect 2136 11500 2188 11509
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 2872 11543 2924 11552
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 3976 11543 4028 11552
rect 3976 11509 3985 11543
rect 3985 11509 4019 11543
rect 4019 11509 4028 11543
rect 3976 11500 4028 11509
rect 4712 11500 4764 11552
rect 7012 11500 7064 11552
rect 8208 11704 8260 11756
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 9588 11704 9640 11756
rect 10324 11704 10376 11756
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 10600 11747 10652 11756
rect 10600 11713 10609 11747
rect 10609 11713 10643 11747
rect 10643 11713 10652 11747
rect 10600 11704 10652 11713
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 11612 11704 11664 11756
rect 11336 11636 11388 11688
rect 11796 11636 11848 11688
rect 13176 11747 13228 11756
rect 13176 11713 13185 11747
rect 13185 11713 13219 11747
rect 13219 11713 13228 11747
rect 13176 11704 13228 11713
rect 11888 11568 11940 11620
rect 12716 11636 12768 11688
rect 14740 11704 14792 11756
rect 15016 11747 15068 11756
rect 15016 11713 15025 11747
rect 15025 11713 15059 11747
rect 15059 11713 15068 11747
rect 15016 11704 15068 11713
rect 15936 11815 15988 11824
rect 15936 11781 15945 11815
rect 15945 11781 15979 11815
rect 15979 11781 15988 11815
rect 15936 11772 15988 11781
rect 16488 11772 16540 11824
rect 15292 11704 15344 11756
rect 14832 11636 14884 11688
rect 16028 11747 16080 11756
rect 16028 11713 16037 11747
rect 16037 11713 16071 11747
rect 16071 11713 16080 11747
rect 16028 11704 16080 11713
rect 16120 11747 16172 11756
rect 16120 11713 16134 11747
rect 16134 11713 16168 11747
rect 16168 11713 16172 11747
rect 16120 11704 16172 11713
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 18144 11772 18196 11824
rect 18972 11840 19024 11892
rect 19616 11840 19668 11892
rect 19524 11772 19576 11824
rect 17960 11747 18012 11756
rect 17960 11713 17969 11747
rect 17969 11713 18003 11747
rect 18003 11713 18012 11747
rect 17960 11704 18012 11713
rect 18788 11704 18840 11756
rect 15476 11568 15528 11620
rect 16028 11568 16080 11620
rect 18052 11636 18104 11688
rect 18880 11636 18932 11688
rect 17960 11568 18012 11620
rect 8944 11500 8996 11552
rect 10048 11500 10100 11552
rect 15200 11543 15252 11552
rect 15200 11509 15209 11543
rect 15209 11509 15243 11543
rect 15243 11509 15252 11543
rect 15200 11500 15252 11509
rect 15292 11500 15344 11552
rect 16120 11500 16172 11552
rect 16212 11500 16264 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 18604 11500 18656 11552
rect 20076 11568 20128 11620
rect 19340 11543 19392 11552
rect 19340 11509 19349 11543
rect 19349 11509 19383 11543
rect 19383 11509 19392 11543
rect 19340 11500 19392 11509
rect 3422 11398 3474 11450
rect 3486 11398 3538 11450
rect 3550 11398 3602 11450
rect 3614 11398 3666 11450
rect 3678 11398 3730 11450
rect 8367 11398 8419 11450
rect 8431 11398 8483 11450
rect 8495 11398 8547 11450
rect 8559 11398 8611 11450
rect 8623 11398 8675 11450
rect 13312 11398 13364 11450
rect 13376 11398 13428 11450
rect 13440 11398 13492 11450
rect 13504 11398 13556 11450
rect 13568 11398 13620 11450
rect 18257 11398 18309 11450
rect 18321 11398 18373 11450
rect 18385 11398 18437 11450
rect 18449 11398 18501 11450
rect 18513 11398 18565 11450
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 2504 11339 2556 11348
rect 2504 11305 2513 11339
rect 2513 11305 2547 11339
rect 2547 11305 2556 11339
rect 2504 11296 2556 11305
rect 4988 11339 5040 11348
rect 4988 11305 4997 11339
rect 4997 11305 5031 11339
rect 5031 11305 5040 11339
rect 4988 11296 5040 11305
rect 5172 11296 5224 11348
rect 4896 11228 4948 11280
rect 8760 11296 8812 11348
rect 11428 11339 11480 11348
rect 11428 11305 11437 11339
rect 11437 11305 11471 11339
rect 11471 11305 11480 11339
rect 11428 11296 11480 11305
rect 14464 11296 14516 11348
rect 16856 11296 16908 11348
rect 18144 11296 18196 11348
rect 18696 11339 18748 11348
rect 18696 11305 18724 11339
rect 18724 11305 18748 11339
rect 18696 11296 18748 11305
rect 3056 11160 3108 11212
rect 4068 11160 4120 11212
rect 2596 11092 2648 11144
rect 2964 11092 3016 11144
rect 4528 11092 4580 11144
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 5632 11092 5684 11144
rect 7012 11203 7064 11212
rect 7012 11169 7021 11203
rect 7021 11169 7055 11203
rect 7055 11169 7064 11203
rect 7012 11160 7064 11169
rect 14372 11228 14424 11280
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 14096 11160 14148 11212
rect 8944 11092 8996 11144
rect 940 11024 992 11076
rect 6920 11067 6972 11076
rect 6920 11033 6929 11067
rect 6929 11033 6963 11067
rect 6963 11033 6972 11067
rect 6920 11024 6972 11033
rect 8208 11024 8260 11076
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 11704 11135 11756 11144
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 11704 11092 11756 11101
rect 11796 11135 11848 11144
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 11796 11092 11848 11101
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 6552 10999 6604 11008
rect 6552 10965 6561 10999
rect 6561 10965 6595 10999
rect 6595 10965 6604 10999
rect 6552 10956 6604 10965
rect 8116 10956 8168 11008
rect 10324 11024 10376 11076
rect 10416 11024 10468 11076
rect 12716 11024 12768 11076
rect 13084 11024 13136 11076
rect 14556 11092 14608 11144
rect 16580 11228 16632 11280
rect 14832 11024 14884 11076
rect 17960 11092 18012 11144
rect 18788 11160 18840 11212
rect 18880 11160 18932 11212
rect 18696 11092 18748 11144
rect 18880 11067 18932 11076
rect 18880 11033 18889 11067
rect 18889 11033 18923 11067
rect 18923 11033 18932 11067
rect 18880 11024 18932 11033
rect 16948 10956 17000 11008
rect 5894 10854 5946 10906
rect 5958 10854 6010 10906
rect 6022 10854 6074 10906
rect 6086 10854 6138 10906
rect 6150 10854 6202 10906
rect 10839 10854 10891 10906
rect 10903 10854 10955 10906
rect 10967 10854 11019 10906
rect 11031 10854 11083 10906
rect 11095 10854 11147 10906
rect 15784 10854 15836 10906
rect 15848 10854 15900 10906
rect 15912 10854 15964 10906
rect 15976 10854 16028 10906
rect 16040 10854 16092 10906
rect 20729 10854 20781 10906
rect 20793 10854 20845 10906
rect 20857 10854 20909 10906
rect 20921 10854 20973 10906
rect 20985 10854 21037 10906
rect 2964 10752 3016 10804
rect 12440 10752 12492 10804
rect 18880 10752 18932 10804
rect 2136 10684 2188 10736
rect 11704 10684 11756 10736
rect 2228 10616 2280 10668
rect 12716 10616 12768 10668
rect 14832 10684 14884 10736
rect 14924 10684 14976 10736
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 15200 10616 15252 10668
rect 15844 10616 15896 10668
rect 16212 10659 16264 10668
rect 16212 10625 16221 10659
rect 16221 10625 16255 10659
rect 16255 10625 16264 10659
rect 16212 10616 16264 10625
rect 18972 10684 19024 10736
rect 10600 10480 10652 10532
rect 12440 10480 12492 10532
rect 1860 10412 1912 10464
rect 9588 10412 9640 10464
rect 13912 10591 13964 10600
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 17040 10548 17092 10600
rect 18604 10659 18656 10668
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 18696 10616 18748 10668
rect 19524 10616 19576 10668
rect 20076 10659 20128 10668
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 14280 10480 14332 10532
rect 16028 10480 16080 10532
rect 16948 10480 17000 10532
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 12992 10412 13044 10421
rect 3422 10310 3474 10362
rect 3486 10310 3538 10362
rect 3550 10310 3602 10362
rect 3614 10310 3666 10362
rect 3678 10310 3730 10362
rect 8367 10310 8419 10362
rect 8431 10310 8483 10362
rect 8495 10310 8547 10362
rect 8559 10310 8611 10362
rect 8623 10310 8675 10362
rect 13312 10310 13364 10362
rect 13376 10310 13428 10362
rect 13440 10310 13492 10362
rect 13504 10310 13556 10362
rect 13568 10310 13620 10362
rect 18257 10310 18309 10362
rect 18321 10310 18373 10362
rect 18385 10310 18437 10362
rect 18449 10310 18501 10362
rect 18513 10310 18565 10362
rect 2964 10251 3016 10260
rect 2964 10217 2973 10251
rect 2973 10217 3007 10251
rect 3007 10217 3016 10251
rect 2964 10208 3016 10217
rect 9496 10208 9548 10260
rect 11704 10251 11756 10260
rect 11704 10217 11713 10251
rect 11713 10217 11747 10251
rect 11747 10217 11756 10251
rect 11704 10208 11756 10217
rect 13912 10208 13964 10260
rect 14740 10208 14792 10260
rect 15844 10251 15896 10260
rect 15844 10217 15853 10251
rect 15853 10217 15887 10251
rect 15887 10217 15896 10251
rect 15844 10208 15896 10217
rect 16028 10251 16080 10260
rect 16028 10217 16037 10251
rect 16037 10217 16071 10251
rect 16071 10217 16080 10251
rect 16028 10208 16080 10217
rect 16672 10208 16724 10260
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 1860 10047 1912 10056
rect 1860 10013 1894 10047
rect 1894 10013 1912 10047
rect 1860 10004 1912 10013
rect 7840 10004 7892 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 8116 9936 8168 9988
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 14740 10047 14792 10056
rect 14740 10013 14749 10047
rect 14749 10013 14783 10047
rect 14783 10013 14792 10047
rect 14740 10004 14792 10013
rect 12992 9936 13044 9988
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 18144 10047 18196 10056
rect 18144 10013 18153 10047
rect 18153 10013 18187 10047
rect 18187 10013 18196 10047
rect 18144 10004 18196 10013
rect 19064 10072 19116 10124
rect 18880 10047 18932 10056
rect 18880 10013 18889 10047
rect 18889 10013 18923 10047
rect 18923 10013 18932 10047
rect 18880 10004 18932 10013
rect 16396 9936 16448 9988
rect 16580 9936 16632 9988
rect 14740 9868 14792 9920
rect 5894 9766 5946 9818
rect 5958 9766 6010 9818
rect 6022 9766 6074 9818
rect 6086 9766 6138 9818
rect 6150 9766 6202 9818
rect 10839 9766 10891 9818
rect 10903 9766 10955 9818
rect 10967 9766 11019 9818
rect 11031 9766 11083 9818
rect 11095 9766 11147 9818
rect 15784 9766 15836 9818
rect 15848 9766 15900 9818
rect 15912 9766 15964 9818
rect 15976 9766 16028 9818
rect 16040 9766 16092 9818
rect 20729 9766 20781 9818
rect 20793 9766 20845 9818
rect 20857 9766 20909 9818
rect 20921 9766 20973 9818
rect 20985 9766 21037 9818
rect 3976 9596 4028 9648
rect 4620 9596 4672 9648
rect 7840 9528 7892 9580
rect 10324 9596 10376 9648
rect 15108 9596 15160 9648
rect 16764 9596 16816 9648
rect 10048 9571 10100 9580
rect 10048 9537 10082 9571
rect 10082 9537 10100 9571
rect 10048 9528 10100 9537
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 1584 9460 1636 9512
rect 4436 9460 4488 9512
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 8852 9460 8904 9512
rect 3884 9392 3936 9444
rect 14740 9392 14792 9444
rect 16120 9528 16172 9580
rect 18144 9528 18196 9580
rect 18972 9571 19024 9580
rect 18972 9537 18981 9571
rect 18981 9537 19015 9571
rect 19015 9537 19024 9571
rect 18972 9528 19024 9537
rect 20076 9528 20128 9580
rect 19340 9392 19392 9444
rect 4804 9324 4856 9376
rect 13176 9324 13228 9376
rect 15200 9324 15252 9376
rect 16672 9324 16724 9376
rect 3422 9222 3474 9274
rect 3486 9222 3538 9274
rect 3550 9222 3602 9274
rect 3614 9222 3666 9274
rect 3678 9222 3730 9274
rect 8367 9222 8419 9274
rect 8431 9222 8483 9274
rect 8495 9222 8547 9274
rect 8559 9222 8611 9274
rect 8623 9222 8675 9274
rect 13312 9222 13364 9274
rect 13376 9222 13428 9274
rect 13440 9222 13492 9274
rect 13504 9222 13556 9274
rect 13568 9222 13620 9274
rect 18257 9222 18309 9274
rect 18321 9222 18373 9274
rect 18385 9222 18437 9274
rect 18449 9222 18501 9274
rect 18513 9222 18565 9274
rect 3056 9120 3108 9172
rect 5816 9163 5868 9172
rect 5816 9129 5825 9163
rect 5825 9129 5859 9163
rect 5859 9129 5868 9163
rect 5816 9120 5868 9129
rect 8024 9120 8076 9172
rect 1584 8984 1636 9036
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 2872 8916 2924 8968
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 4712 8959 4764 8968
rect 4712 8925 4746 8959
rect 4746 8925 4764 8959
rect 4712 8916 4764 8925
rect 11796 9120 11848 9172
rect 14096 9120 14148 9172
rect 18144 9120 18196 9172
rect 18788 9163 18840 9172
rect 18788 9129 18797 9163
rect 18797 9129 18831 9163
rect 18831 9129 18840 9163
rect 18788 9120 18840 9129
rect 14188 9052 14240 9104
rect 13084 8984 13136 9036
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 13176 8916 13228 8968
rect 14924 8984 14976 9036
rect 14740 8916 14792 8968
rect 16304 8959 16356 8968
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 16672 8916 16724 8968
rect 17040 9027 17092 9036
rect 17040 8993 17049 9027
rect 17049 8993 17083 9027
rect 17083 8993 17092 9027
rect 17040 8984 17092 8993
rect 17868 8984 17920 9036
rect 18880 9052 18932 9104
rect 16948 8916 17000 8968
rect 13820 8848 13872 8900
rect 14464 8891 14516 8900
rect 14464 8857 14473 8891
rect 14473 8857 14507 8891
rect 14507 8857 14516 8891
rect 14464 8848 14516 8857
rect 15660 8848 15712 8900
rect 18144 8848 18196 8900
rect 13912 8780 13964 8832
rect 16304 8780 16356 8832
rect 18052 8780 18104 8832
rect 18420 8780 18472 8832
rect 5894 8678 5946 8730
rect 5958 8678 6010 8730
rect 6022 8678 6074 8730
rect 6086 8678 6138 8730
rect 6150 8678 6202 8730
rect 10839 8678 10891 8730
rect 10903 8678 10955 8730
rect 10967 8678 11019 8730
rect 11031 8678 11083 8730
rect 11095 8678 11147 8730
rect 15784 8678 15836 8730
rect 15848 8678 15900 8730
rect 15912 8678 15964 8730
rect 15976 8678 16028 8730
rect 16040 8678 16092 8730
rect 20729 8678 20781 8730
rect 20793 8678 20845 8730
rect 20857 8678 20909 8730
rect 20921 8678 20973 8730
rect 20985 8678 21037 8730
rect 11888 8576 11940 8628
rect 17040 8576 17092 8628
rect 18880 8576 18932 8628
rect 10324 8508 10376 8560
rect 13912 8551 13964 8560
rect 13912 8517 13921 8551
rect 13921 8517 13955 8551
rect 13955 8517 13964 8551
rect 13912 8508 13964 8517
rect 14004 8551 14056 8560
rect 14004 8517 14013 8551
rect 14013 8517 14047 8551
rect 14047 8517 14056 8551
rect 14004 8508 14056 8517
rect 11520 8440 11572 8492
rect 13820 8483 13872 8492
rect 13820 8449 13829 8483
rect 13829 8449 13863 8483
rect 13863 8449 13872 8483
rect 13820 8440 13872 8449
rect 14096 8483 14148 8492
rect 14096 8449 14131 8483
rect 14131 8449 14148 8483
rect 14096 8440 14148 8449
rect 14740 8483 14792 8492
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 14740 8440 14792 8449
rect 14924 8483 14976 8492
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 15108 8440 15160 8492
rect 16580 8440 16632 8492
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 18144 8483 18196 8492
rect 18144 8449 18153 8483
rect 18153 8449 18187 8483
rect 18187 8449 18196 8483
rect 18144 8440 18196 8449
rect 18236 8483 18288 8492
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 18512 8483 18564 8492
rect 18512 8449 18521 8483
rect 18521 8449 18555 8483
rect 18555 8449 18564 8483
rect 18512 8440 18564 8449
rect 18696 8372 18748 8424
rect 16948 8304 17000 8356
rect 13636 8279 13688 8288
rect 13636 8245 13645 8279
rect 13645 8245 13679 8279
rect 13679 8245 13688 8279
rect 13636 8236 13688 8245
rect 14832 8279 14884 8288
rect 14832 8245 14841 8279
rect 14841 8245 14875 8279
rect 14875 8245 14884 8279
rect 14832 8236 14884 8245
rect 3422 8134 3474 8186
rect 3486 8134 3538 8186
rect 3550 8134 3602 8186
rect 3614 8134 3666 8186
rect 3678 8134 3730 8186
rect 8367 8134 8419 8186
rect 8431 8134 8483 8186
rect 8495 8134 8547 8186
rect 8559 8134 8611 8186
rect 8623 8134 8675 8186
rect 13312 8134 13364 8186
rect 13376 8134 13428 8186
rect 13440 8134 13492 8186
rect 13504 8134 13556 8186
rect 13568 8134 13620 8186
rect 18257 8134 18309 8186
rect 18321 8134 18373 8186
rect 18385 8134 18437 8186
rect 18449 8134 18501 8186
rect 18513 8134 18565 8186
rect 2780 8032 2832 8084
rect 6460 8032 6512 8084
rect 8208 8075 8260 8084
rect 8208 8041 8217 8075
rect 8217 8041 8251 8075
rect 8251 8041 8260 8075
rect 8208 8032 8260 8041
rect 15660 8032 15712 8084
rect 16672 7964 16724 8016
rect 1584 7939 1636 7948
rect 1584 7905 1593 7939
rect 1593 7905 1627 7939
rect 1627 7905 1636 7939
rect 1584 7896 1636 7905
rect 2688 7896 2740 7948
rect 4436 7896 4488 7948
rect 13728 7896 13780 7948
rect 17040 7896 17092 7948
rect 17408 7896 17460 7948
rect 1676 7828 1728 7880
rect 7840 7828 7892 7880
rect 10324 7828 10376 7880
rect 10508 7828 10560 7880
rect 13636 7828 13688 7880
rect 7104 7803 7156 7812
rect 7104 7769 7138 7803
rect 7138 7769 7156 7803
rect 7104 7760 7156 7769
rect 15568 7828 15620 7880
rect 16764 7828 16816 7880
rect 17132 7828 17184 7880
rect 18052 7896 18104 7948
rect 18696 7939 18748 7948
rect 18696 7905 18705 7939
rect 18705 7905 18739 7939
rect 18739 7905 18748 7939
rect 18696 7896 18748 7905
rect 18144 7828 18196 7880
rect 18420 7871 18472 7880
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 18604 7871 18656 7880
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 15108 7760 15160 7812
rect 11888 7692 11940 7744
rect 13176 7692 13228 7744
rect 15200 7692 15252 7744
rect 16856 7692 16908 7744
rect 18880 7735 18932 7744
rect 18880 7701 18889 7735
rect 18889 7701 18923 7735
rect 18923 7701 18932 7735
rect 18880 7692 18932 7701
rect 5894 7590 5946 7642
rect 5958 7590 6010 7642
rect 6022 7590 6074 7642
rect 6086 7590 6138 7642
rect 6150 7590 6202 7642
rect 10839 7590 10891 7642
rect 10903 7590 10955 7642
rect 10967 7590 11019 7642
rect 11031 7590 11083 7642
rect 11095 7590 11147 7642
rect 15784 7590 15836 7642
rect 15848 7590 15900 7642
rect 15912 7590 15964 7642
rect 15976 7590 16028 7642
rect 16040 7590 16092 7642
rect 20729 7590 20781 7642
rect 20793 7590 20845 7642
rect 20857 7590 20909 7642
rect 20921 7590 20973 7642
rect 20985 7590 21037 7642
rect 16764 7488 16816 7540
rect 16856 7531 16908 7540
rect 16856 7497 16865 7531
rect 16865 7497 16899 7531
rect 16899 7497 16908 7531
rect 16856 7488 16908 7497
rect 1584 7420 1636 7472
rect 2688 7420 2740 7472
rect 10324 7420 10376 7472
rect 14464 7420 14516 7472
rect 7656 7352 7708 7404
rect 14832 7352 14884 7404
rect 17868 7463 17920 7472
rect 17868 7429 17877 7463
rect 17877 7429 17911 7463
rect 17911 7429 17920 7463
rect 17868 7420 17920 7429
rect 13176 7284 13228 7336
rect 15292 7284 15344 7336
rect 15936 7327 15988 7336
rect 15936 7293 15945 7327
rect 15945 7293 15979 7327
rect 15979 7293 15988 7327
rect 15936 7284 15988 7293
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 19064 7488 19116 7540
rect 18420 7420 18472 7472
rect 18604 7352 18656 7404
rect 13912 7216 13964 7268
rect 13820 7191 13872 7200
rect 13820 7157 13829 7191
rect 13829 7157 13863 7191
rect 13863 7157 13872 7191
rect 13820 7148 13872 7157
rect 14004 7148 14056 7200
rect 14280 7148 14332 7200
rect 15108 7148 15160 7200
rect 18144 7191 18196 7200
rect 18144 7157 18153 7191
rect 18153 7157 18187 7191
rect 18187 7157 18196 7191
rect 18144 7148 18196 7157
rect 18604 7148 18656 7200
rect 19892 7148 19944 7200
rect 3422 7046 3474 7098
rect 3486 7046 3538 7098
rect 3550 7046 3602 7098
rect 3614 7046 3666 7098
rect 3678 7046 3730 7098
rect 8367 7046 8419 7098
rect 8431 7046 8483 7098
rect 8495 7046 8547 7098
rect 8559 7046 8611 7098
rect 8623 7046 8675 7098
rect 13312 7046 13364 7098
rect 13376 7046 13428 7098
rect 13440 7046 13492 7098
rect 13504 7046 13556 7098
rect 13568 7046 13620 7098
rect 18257 7046 18309 7098
rect 18321 7046 18373 7098
rect 18385 7046 18437 7098
rect 18449 7046 18501 7098
rect 18513 7046 18565 7098
rect 4436 6808 4488 6860
rect 14464 6876 14516 6928
rect 13728 6808 13780 6860
rect 15936 6944 15988 6996
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 1860 6783 1912 6792
rect 1860 6749 1894 6783
rect 1894 6749 1912 6783
rect 1860 6740 1912 6749
rect 6552 6740 6604 6792
rect 9772 6740 9824 6792
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 10600 6783 10652 6792
rect 10600 6749 10634 6783
rect 10634 6749 10652 6783
rect 10600 6740 10652 6749
rect 6368 6715 6420 6724
rect 6368 6681 6377 6715
rect 6377 6681 6411 6715
rect 6411 6681 6420 6715
rect 6368 6672 6420 6681
rect 8208 6672 8260 6724
rect 13912 6740 13964 6792
rect 14832 6740 14884 6792
rect 15200 6740 15252 6792
rect 15292 6740 15344 6792
rect 18144 6740 18196 6792
rect 19248 6808 19300 6860
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 19064 6740 19116 6792
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 19892 6783 19944 6792
rect 19892 6749 19901 6783
rect 19901 6749 19935 6783
rect 19935 6749 19944 6783
rect 19892 6740 19944 6749
rect 15108 6672 15160 6724
rect 2136 6604 2188 6656
rect 6920 6604 6972 6656
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 7656 6604 7708 6613
rect 12992 6647 13044 6656
rect 12992 6613 13001 6647
rect 13001 6613 13035 6647
rect 13035 6613 13044 6647
rect 12992 6604 13044 6613
rect 15200 6604 15252 6656
rect 17040 6672 17092 6724
rect 19064 6604 19116 6656
rect 5894 6502 5946 6554
rect 5958 6502 6010 6554
rect 6022 6502 6074 6554
rect 6086 6502 6138 6554
rect 6150 6502 6202 6554
rect 10839 6502 10891 6554
rect 10903 6502 10955 6554
rect 10967 6502 11019 6554
rect 11031 6502 11083 6554
rect 11095 6502 11147 6554
rect 15784 6502 15836 6554
rect 15848 6502 15900 6554
rect 15912 6502 15964 6554
rect 15976 6502 16028 6554
rect 16040 6502 16092 6554
rect 20729 6502 20781 6554
rect 20793 6502 20845 6554
rect 20857 6502 20909 6554
rect 20921 6502 20973 6554
rect 20985 6502 21037 6554
rect 9220 6400 9272 6452
rect 5448 6332 5500 6384
rect 8208 6375 8260 6384
rect 8208 6341 8242 6375
rect 8242 6341 8260 6375
rect 8208 6332 8260 6341
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 7840 6264 7892 6316
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 13176 6400 13228 6452
rect 13820 6400 13872 6452
rect 11888 6332 11940 6384
rect 14096 6332 14148 6384
rect 13176 6264 13228 6316
rect 15200 6400 15252 6452
rect 15292 6443 15344 6452
rect 15292 6409 15301 6443
rect 15301 6409 15335 6443
rect 15335 6409 15344 6443
rect 15292 6400 15344 6409
rect 18696 6443 18748 6452
rect 18696 6409 18705 6443
rect 18705 6409 18739 6443
rect 18739 6409 18748 6443
rect 18696 6400 18748 6409
rect 19248 6400 19300 6452
rect 4252 6196 4304 6248
rect 13728 6239 13780 6248
rect 13728 6205 13737 6239
rect 13737 6205 13771 6239
rect 13771 6205 13780 6239
rect 13728 6196 13780 6205
rect 18052 6332 18104 6384
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 18788 6264 18840 6316
rect 18880 6307 18932 6316
rect 18880 6273 18889 6307
rect 18889 6273 18923 6307
rect 18923 6273 18932 6307
rect 18880 6264 18932 6273
rect 19064 6307 19116 6316
rect 19064 6273 19073 6307
rect 19073 6273 19107 6307
rect 19107 6273 19116 6307
rect 19064 6264 19116 6273
rect 6460 6128 6512 6180
rect 17408 6196 17460 6248
rect 17776 6196 17828 6248
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 9588 6060 9640 6112
rect 15108 6171 15160 6180
rect 15108 6137 15117 6171
rect 15117 6137 15151 6171
rect 15151 6137 15160 6171
rect 15108 6128 15160 6137
rect 12808 6060 12860 6112
rect 17408 6060 17460 6112
rect 3422 5958 3474 6010
rect 3486 5958 3538 6010
rect 3550 5958 3602 6010
rect 3614 5958 3666 6010
rect 3678 5958 3730 6010
rect 8367 5958 8419 6010
rect 8431 5958 8483 6010
rect 8495 5958 8547 6010
rect 8559 5958 8611 6010
rect 8623 5958 8675 6010
rect 13312 5958 13364 6010
rect 13376 5958 13428 6010
rect 13440 5958 13492 6010
rect 13504 5958 13556 6010
rect 13568 5958 13620 6010
rect 18257 5958 18309 6010
rect 18321 5958 18373 6010
rect 18385 5958 18437 6010
rect 18449 5958 18501 6010
rect 18513 5958 18565 6010
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 9588 5856 9640 5908
rect 1584 5652 1636 5704
rect 4252 5695 4304 5704
rect 4252 5661 4261 5695
rect 4261 5661 4295 5695
rect 4295 5661 4304 5695
rect 4252 5652 4304 5661
rect 4528 5695 4580 5704
rect 4528 5661 4537 5695
rect 4537 5661 4571 5695
rect 4571 5661 4580 5695
rect 4528 5652 4580 5661
rect 7104 5695 7156 5704
rect 7104 5661 7113 5695
rect 7113 5661 7147 5695
rect 7147 5661 7156 5695
rect 7104 5652 7156 5661
rect 13912 5788 13964 5840
rect 15568 5788 15620 5840
rect 18788 5788 18840 5840
rect 13636 5720 13688 5772
rect 17408 5720 17460 5772
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 12992 5652 13044 5704
rect 17316 5652 17368 5704
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 16672 5584 16724 5636
rect 11336 5516 11388 5568
rect 12900 5559 12952 5568
rect 12900 5525 12909 5559
rect 12909 5525 12943 5559
rect 12943 5525 12952 5559
rect 12900 5516 12952 5525
rect 12992 5559 13044 5568
rect 12992 5525 13001 5559
rect 13001 5525 13035 5559
rect 13035 5525 13044 5559
rect 12992 5516 13044 5525
rect 5894 5414 5946 5466
rect 5958 5414 6010 5466
rect 6022 5414 6074 5466
rect 6086 5414 6138 5466
rect 6150 5414 6202 5466
rect 10839 5414 10891 5466
rect 10903 5414 10955 5466
rect 10967 5414 11019 5466
rect 11031 5414 11083 5466
rect 11095 5414 11147 5466
rect 15784 5414 15836 5466
rect 15848 5414 15900 5466
rect 15912 5414 15964 5466
rect 15976 5414 16028 5466
rect 16040 5414 16092 5466
rect 20729 5414 20781 5466
rect 20793 5414 20845 5466
rect 20857 5414 20909 5466
rect 20921 5414 20973 5466
rect 20985 5414 21037 5466
rect 6920 5312 6972 5364
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 1860 5219 1912 5228
rect 1860 5185 1894 5219
rect 1894 5185 1912 5219
rect 1860 5176 1912 5185
rect 11336 5244 11388 5296
rect 12532 5244 12584 5296
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 12808 5176 12860 5228
rect 13636 5287 13688 5296
rect 13636 5253 13645 5287
rect 13645 5253 13679 5287
rect 13679 5253 13688 5287
rect 13636 5244 13688 5253
rect 16304 5244 16356 5296
rect 17040 5244 17092 5296
rect 14188 5219 14240 5228
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 14280 5176 14332 5228
rect 4252 5108 4304 5160
rect 9772 5151 9824 5160
rect 9772 5117 9781 5151
rect 9781 5117 9815 5151
rect 9815 5117 9824 5151
rect 9772 5108 9824 5117
rect 2964 5015 3016 5024
rect 2964 4981 2973 5015
rect 2973 4981 3007 5015
rect 3007 4981 3016 5015
rect 2964 4972 3016 4981
rect 6920 4972 6972 5024
rect 9680 4972 9732 5024
rect 12992 5040 13044 5092
rect 14464 5219 14516 5228
rect 14464 5185 14473 5219
rect 14473 5185 14507 5219
rect 14507 5185 14516 5219
rect 14464 5176 14516 5185
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 15292 5219 15344 5228
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 15292 5176 15344 5185
rect 12900 4972 12952 5024
rect 14372 4972 14424 5024
rect 14464 4972 14516 5024
rect 15660 5219 15712 5228
rect 15660 5185 15670 5219
rect 15670 5185 15704 5219
rect 15704 5185 15712 5219
rect 15660 5176 15712 5185
rect 17408 5219 17460 5228
rect 17408 5185 17417 5219
rect 17417 5185 17451 5219
rect 17451 5185 17460 5219
rect 17408 5176 17460 5185
rect 17316 5151 17368 5160
rect 17316 5117 17325 5151
rect 17325 5117 17359 5151
rect 17359 5117 17368 5151
rect 17316 5108 17368 5117
rect 17776 5151 17828 5160
rect 17776 5117 17785 5151
rect 17785 5117 17819 5151
rect 17819 5117 17828 5151
rect 17776 5108 17828 5117
rect 17132 5015 17184 5024
rect 17132 4981 17141 5015
rect 17141 4981 17175 5015
rect 17175 4981 17184 5015
rect 17132 4972 17184 4981
rect 3422 4870 3474 4922
rect 3486 4870 3538 4922
rect 3550 4870 3602 4922
rect 3614 4870 3666 4922
rect 3678 4870 3730 4922
rect 8367 4870 8419 4922
rect 8431 4870 8483 4922
rect 8495 4870 8547 4922
rect 8559 4870 8611 4922
rect 8623 4870 8675 4922
rect 13312 4870 13364 4922
rect 13376 4870 13428 4922
rect 13440 4870 13492 4922
rect 13504 4870 13556 4922
rect 13568 4870 13620 4922
rect 18257 4870 18309 4922
rect 18321 4870 18373 4922
rect 18385 4870 18437 4922
rect 18449 4870 18501 4922
rect 18513 4870 18565 4922
rect 9680 4768 9732 4820
rect 13176 4768 13228 4820
rect 15292 4768 15344 4820
rect 16672 4811 16724 4820
rect 16672 4777 16681 4811
rect 16681 4777 16715 4811
rect 16715 4777 16724 4811
rect 16672 4768 16724 4777
rect 16948 4768 17000 4820
rect 17316 4768 17368 4820
rect 17776 4768 17828 4820
rect 14556 4700 14608 4752
rect 15660 4700 15712 4752
rect 17224 4700 17276 4752
rect 9772 4564 9824 4616
rect 12992 4564 13044 4616
rect 14556 4564 14608 4616
rect 16764 4607 16816 4616
rect 16764 4573 16773 4607
rect 16773 4573 16807 4607
rect 16807 4573 16816 4607
rect 16764 4564 16816 4573
rect 17040 4564 17092 4616
rect 18052 4564 18104 4616
rect 18604 4564 18656 4616
rect 16672 4496 16724 4548
rect 16580 4428 16632 4480
rect 5894 4326 5946 4378
rect 5958 4326 6010 4378
rect 6022 4326 6074 4378
rect 6086 4326 6138 4378
rect 6150 4326 6202 4378
rect 10839 4326 10891 4378
rect 10903 4326 10955 4378
rect 10967 4326 11019 4378
rect 11031 4326 11083 4378
rect 11095 4326 11147 4378
rect 15784 4326 15836 4378
rect 15848 4326 15900 4378
rect 15912 4326 15964 4378
rect 15976 4326 16028 4378
rect 16040 4326 16092 4378
rect 20729 4326 20781 4378
rect 20793 4326 20845 4378
rect 20857 4326 20909 4378
rect 20921 4326 20973 4378
rect 20985 4326 21037 4378
rect 1860 4267 1912 4276
rect 1860 4233 1869 4267
rect 1869 4233 1903 4267
rect 1903 4233 1912 4267
rect 1860 4224 1912 4233
rect 1860 4088 1912 4140
rect 2964 4156 3016 4208
rect 4068 4088 4120 4140
rect 4252 4088 4304 4140
rect 1584 4020 1636 4072
rect 4160 3927 4212 3936
rect 4160 3893 4169 3927
rect 4169 3893 4203 3927
rect 4203 3893 4212 3927
rect 4160 3884 4212 3893
rect 6552 3884 6604 3936
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 9864 4088 9916 4140
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 14096 4131 14148 4140
rect 14096 4097 14105 4131
rect 14105 4097 14139 4131
rect 14139 4097 14148 4131
rect 14096 4088 14148 4097
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 14464 4131 14516 4140
rect 14464 4097 14473 4131
rect 14473 4097 14507 4131
rect 14507 4097 14516 4131
rect 14464 4088 14516 4097
rect 14648 4131 14700 4140
rect 14648 4097 14657 4131
rect 14657 4097 14691 4131
rect 14691 4097 14700 4131
rect 14648 4088 14700 4097
rect 17132 4020 17184 4072
rect 16764 3952 16816 4004
rect 7288 3884 7340 3936
rect 8760 3884 8812 3936
rect 3422 3782 3474 3834
rect 3486 3782 3538 3834
rect 3550 3782 3602 3834
rect 3614 3782 3666 3834
rect 3678 3782 3730 3834
rect 8367 3782 8419 3834
rect 8431 3782 8483 3834
rect 8495 3782 8547 3834
rect 8559 3782 8611 3834
rect 8623 3782 8675 3834
rect 13312 3782 13364 3834
rect 13376 3782 13428 3834
rect 13440 3782 13492 3834
rect 13504 3782 13556 3834
rect 13568 3782 13620 3834
rect 18257 3782 18309 3834
rect 18321 3782 18373 3834
rect 18385 3782 18437 3834
rect 18449 3782 18501 3834
rect 18513 3782 18565 3834
rect 4068 3723 4120 3732
rect 4068 3689 4077 3723
rect 4077 3689 4111 3723
rect 4111 3689 4120 3723
rect 4068 3680 4120 3689
rect 12348 3680 12400 3732
rect 3240 3612 3292 3664
rect 6368 3612 6420 3664
rect 14280 3723 14332 3732
rect 14280 3689 14289 3723
rect 14289 3689 14323 3723
rect 14323 3689 14332 3723
rect 14280 3680 14332 3689
rect 16672 3723 16724 3732
rect 16672 3689 16681 3723
rect 16681 3689 16715 3723
rect 16715 3689 16724 3723
rect 16672 3680 16724 3689
rect 17408 3680 17460 3732
rect 1584 3544 1636 3596
rect 5632 3544 5684 3596
rect 12348 3544 12400 3596
rect 12992 3587 13044 3596
rect 12992 3553 13001 3587
rect 13001 3553 13035 3587
rect 13035 3553 13044 3587
rect 12992 3544 13044 3553
rect 1860 3476 1912 3528
rect 2412 3408 2464 3460
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4252 3476 4304 3485
rect 6920 3476 6972 3528
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 9772 3476 9824 3528
rect 17040 3612 17092 3664
rect 17684 3612 17736 3664
rect 13912 3544 13964 3596
rect 14832 3587 14884 3596
rect 14832 3553 14841 3587
rect 14841 3553 14875 3587
rect 14875 3553 14884 3587
rect 14832 3544 14884 3553
rect 4528 3408 4580 3460
rect 3148 3383 3200 3392
rect 3148 3349 3157 3383
rect 3157 3349 3191 3383
rect 3191 3349 3200 3383
rect 3148 3340 3200 3349
rect 10140 3340 10192 3392
rect 10508 3383 10560 3392
rect 10508 3349 10517 3383
rect 10517 3349 10551 3383
rect 10551 3349 10560 3383
rect 10508 3340 10560 3349
rect 14372 3476 14424 3528
rect 14648 3476 14700 3528
rect 14740 3476 14792 3528
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 15568 3519 15620 3528
rect 15568 3485 15577 3519
rect 15577 3485 15611 3519
rect 15611 3485 15620 3519
rect 15568 3476 15620 3485
rect 16948 3519 17000 3528
rect 16948 3485 16957 3519
rect 16957 3485 16991 3519
rect 16991 3485 17000 3519
rect 16948 3476 17000 3485
rect 17224 3519 17276 3528
rect 17224 3485 17233 3519
rect 17233 3485 17267 3519
rect 17267 3485 17276 3519
rect 17224 3476 17276 3485
rect 17684 3519 17736 3528
rect 17684 3485 17693 3519
rect 17693 3485 17727 3519
rect 17727 3485 17736 3519
rect 17684 3476 17736 3485
rect 17960 3519 18012 3528
rect 17960 3485 17969 3519
rect 17969 3485 18003 3519
rect 18003 3485 18012 3519
rect 17960 3476 18012 3485
rect 18052 3519 18104 3528
rect 18052 3485 18061 3519
rect 18061 3485 18095 3519
rect 18095 3485 18104 3519
rect 18052 3476 18104 3485
rect 13268 3340 13320 3392
rect 14556 3340 14608 3392
rect 15476 3383 15528 3392
rect 15476 3349 15485 3383
rect 15485 3349 15519 3383
rect 15519 3349 15528 3383
rect 15476 3340 15528 3349
rect 5894 3238 5946 3290
rect 5958 3238 6010 3290
rect 6022 3238 6074 3290
rect 6086 3238 6138 3290
rect 6150 3238 6202 3290
rect 10839 3238 10891 3290
rect 10903 3238 10955 3290
rect 10967 3238 11019 3290
rect 11031 3238 11083 3290
rect 11095 3238 11147 3290
rect 15784 3238 15836 3290
rect 15848 3238 15900 3290
rect 15912 3238 15964 3290
rect 15976 3238 16028 3290
rect 16040 3238 16092 3290
rect 20729 3238 20781 3290
rect 20793 3238 20845 3290
rect 20857 3238 20909 3290
rect 20921 3238 20973 3290
rect 20985 3238 21037 3290
rect 1584 3068 1636 3120
rect 5356 3068 5408 3120
rect 7288 3136 7340 3188
rect 9128 3179 9180 3188
rect 9128 3145 9137 3179
rect 9137 3145 9171 3179
rect 9171 3145 9180 3179
rect 9128 3136 9180 3145
rect 9864 3136 9916 3188
rect 10140 3136 10192 3188
rect 7656 3068 7708 3120
rect 11060 3068 11112 3120
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 9956 3000 10008 3052
rect 12440 3000 12492 3052
rect 13636 3000 13688 3052
rect 15476 3068 15528 3120
rect 14740 3000 14792 3052
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 15660 3043 15712 3052
rect 15660 3009 15669 3043
rect 15669 3009 15703 3043
rect 15703 3009 15712 3043
rect 15660 3000 15712 3009
rect 15936 3043 15988 3052
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 5264 2975 5316 2984
rect 5264 2941 5273 2975
rect 5273 2941 5307 2975
rect 5307 2941 5316 2975
rect 5264 2932 5316 2941
rect 6736 2932 6788 2984
rect 8760 2932 8812 2984
rect 5632 2864 5684 2916
rect 9680 2796 9732 2848
rect 14004 2975 14056 2984
rect 14004 2941 14013 2975
rect 14013 2941 14047 2975
rect 14047 2941 14056 2975
rect 14004 2932 14056 2941
rect 14556 2932 14608 2984
rect 15844 2932 15896 2984
rect 16948 3000 17000 3052
rect 17224 2975 17276 2984
rect 17224 2941 17233 2975
rect 17233 2941 17267 2975
rect 17267 2941 17276 2975
rect 17224 2932 17276 2941
rect 17960 2932 18012 2984
rect 12624 2796 12676 2848
rect 12992 2796 13044 2848
rect 13268 2796 13320 2848
rect 3422 2694 3474 2746
rect 3486 2694 3538 2746
rect 3550 2694 3602 2746
rect 3614 2694 3666 2746
rect 3678 2694 3730 2746
rect 8367 2694 8419 2746
rect 8431 2694 8483 2746
rect 8495 2694 8547 2746
rect 8559 2694 8611 2746
rect 8623 2694 8675 2746
rect 13312 2694 13364 2746
rect 13376 2694 13428 2746
rect 13440 2694 13492 2746
rect 13504 2694 13556 2746
rect 13568 2694 13620 2746
rect 18257 2694 18309 2746
rect 18321 2694 18373 2746
rect 18385 2694 18437 2746
rect 18449 2694 18501 2746
rect 18513 2694 18565 2746
rect 2412 2635 2464 2644
rect 2412 2601 2421 2635
rect 2421 2601 2455 2635
rect 2455 2601 2464 2635
rect 2412 2592 2464 2601
rect 4252 2592 4304 2644
rect 5448 2592 5500 2644
rect 5632 2592 5684 2644
rect 6828 2592 6880 2644
rect 9956 2592 10008 2644
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 14832 2635 14884 2644
rect 14832 2601 14841 2635
rect 14841 2601 14875 2635
rect 14875 2601 14884 2635
rect 14832 2592 14884 2601
rect 15660 2592 15712 2644
rect 1860 2388 1912 2440
rect 2964 2388 3016 2440
rect 3148 2388 3200 2440
rect 4160 2388 4212 2440
rect 14004 2524 14056 2576
rect 4528 2388 4580 2440
rect 4160 2295 4212 2304
rect 4160 2261 4169 2295
rect 4169 2261 4203 2295
rect 4203 2261 4212 2295
rect 4160 2252 4212 2261
rect 4436 2320 4488 2372
rect 5264 2320 5316 2372
rect 5356 2363 5408 2372
rect 5356 2329 5381 2363
rect 5381 2329 5408 2363
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 9680 2456 9732 2508
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 6736 2388 6788 2397
rect 8760 2388 8812 2440
rect 5356 2320 5408 2329
rect 11060 2388 11112 2440
rect 12348 2388 12400 2440
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 14096 2456 14148 2508
rect 15568 2388 15620 2440
rect 15936 2388 15988 2440
rect 14004 2320 14056 2372
rect 14648 2363 14700 2372
rect 14648 2329 14657 2363
rect 14657 2329 14691 2363
rect 14691 2329 14700 2363
rect 14648 2320 14700 2329
rect 14740 2320 14792 2372
rect 15384 2320 15436 2372
rect 15844 2252 15896 2304
rect 5894 2150 5946 2202
rect 5958 2150 6010 2202
rect 6022 2150 6074 2202
rect 6086 2150 6138 2202
rect 6150 2150 6202 2202
rect 10839 2150 10891 2202
rect 10903 2150 10955 2202
rect 10967 2150 11019 2202
rect 11031 2150 11083 2202
rect 11095 2150 11147 2202
rect 15784 2150 15836 2202
rect 15848 2150 15900 2202
rect 15912 2150 15964 2202
rect 15976 2150 16028 2202
rect 16040 2150 16092 2202
rect 20729 2150 20781 2202
rect 20793 2150 20845 2202
rect 20857 2150 20909 2202
rect 20921 2150 20973 2202
rect 20985 2150 21037 2202
<< metal2 >>
rect 5894 19612 6202 19621
rect 5894 19610 5900 19612
rect 5956 19610 5980 19612
rect 6036 19610 6060 19612
rect 6116 19610 6140 19612
rect 6196 19610 6202 19612
rect 5956 19558 5958 19610
rect 6138 19558 6140 19610
rect 5894 19556 5900 19558
rect 5956 19556 5980 19558
rect 6036 19556 6060 19558
rect 6116 19556 6140 19558
rect 6196 19556 6202 19558
rect 5894 19547 6202 19556
rect 10839 19612 11147 19621
rect 10839 19610 10845 19612
rect 10901 19610 10925 19612
rect 10981 19610 11005 19612
rect 11061 19610 11085 19612
rect 11141 19610 11147 19612
rect 10901 19558 10903 19610
rect 11083 19558 11085 19610
rect 10839 19556 10845 19558
rect 10901 19556 10925 19558
rect 10981 19556 11005 19558
rect 11061 19556 11085 19558
rect 11141 19556 11147 19558
rect 10839 19547 11147 19556
rect 15784 19612 16092 19621
rect 15784 19610 15790 19612
rect 15846 19610 15870 19612
rect 15926 19610 15950 19612
rect 16006 19610 16030 19612
rect 16086 19610 16092 19612
rect 15846 19558 15848 19610
rect 16028 19558 16030 19610
rect 15784 19556 15790 19558
rect 15846 19556 15870 19558
rect 15926 19556 15950 19558
rect 16006 19556 16030 19558
rect 16086 19556 16092 19558
rect 15784 19547 16092 19556
rect 20729 19612 21037 19621
rect 20729 19610 20735 19612
rect 20791 19610 20815 19612
rect 20871 19610 20895 19612
rect 20951 19610 20975 19612
rect 21031 19610 21037 19612
rect 20791 19558 20793 19610
rect 20973 19558 20975 19610
rect 20729 19556 20735 19558
rect 20791 19556 20815 19558
rect 20871 19556 20895 19558
rect 20951 19556 20975 19558
rect 21031 19556 21037 19558
rect 20729 19547 21037 19556
rect 3422 19068 3730 19077
rect 3422 19066 3428 19068
rect 3484 19066 3508 19068
rect 3564 19066 3588 19068
rect 3644 19066 3668 19068
rect 3724 19066 3730 19068
rect 3484 19014 3486 19066
rect 3666 19014 3668 19066
rect 3422 19012 3428 19014
rect 3484 19012 3508 19014
rect 3564 19012 3588 19014
rect 3644 19012 3668 19014
rect 3724 19012 3730 19014
rect 3422 19003 3730 19012
rect 8367 19068 8675 19077
rect 8367 19066 8373 19068
rect 8429 19066 8453 19068
rect 8509 19066 8533 19068
rect 8589 19066 8613 19068
rect 8669 19066 8675 19068
rect 8429 19014 8431 19066
rect 8611 19014 8613 19066
rect 8367 19012 8373 19014
rect 8429 19012 8453 19014
rect 8509 19012 8533 19014
rect 8589 19012 8613 19014
rect 8669 19012 8675 19014
rect 8367 19003 8675 19012
rect 13312 19068 13620 19077
rect 13312 19066 13318 19068
rect 13374 19066 13398 19068
rect 13454 19066 13478 19068
rect 13534 19066 13558 19068
rect 13614 19066 13620 19068
rect 13374 19014 13376 19066
rect 13556 19014 13558 19066
rect 13312 19012 13318 19014
rect 13374 19012 13398 19014
rect 13454 19012 13478 19014
rect 13534 19012 13558 19014
rect 13614 19012 13620 19014
rect 13312 19003 13620 19012
rect 18257 19068 18565 19077
rect 18257 19066 18263 19068
rect 18319 19066 18343 19068
rect 18399 19066 18423 19068
rect 18479 19066 18503 19068
rect 18559 19066 18565 19068
rect 18319 19014 18321 19066
rect 18501 19014 18503 19066
rect 18257 19012 18263 19014
rect 18319 19012 18343 19014
rect 18399 19012 18423 19014
rect 18479 19012 18503 19014
rect 18559 19012 18565 19014
rect 18257 19003 18565 19012
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 940 18692 992 18698
rect 940 18634 992 18640
rect 952 18329 980 18634
rect 938 18320 994 18329
rect 938 18255 994 18264
rect 2228 15088 2280 15094
rect 2228 15030 2280 15036
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 2056 14074 2084 14758
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 940 11076 992 11082
rect 940 11018 992 11024
rect 952 10985 980 11018
rect 938 10976 994 10985
rect 938 10911 994 10920
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9518 1624 9998
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 9042 1624 9454
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1596 7954 1624 8978
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1596 7478 1624 7890
rect 1688 7886 1716 13126
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1780 6914 1808 14010
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 2056 12850 2084 13874
rect 2240 13190 2268 15030
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2332 13870 2360 14894
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2332 13258 2360 13806
rect 2412 13796 2464 13802
rect 2412 13738 2464 13744
rect 2424 13394 2452 13738
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12918 2268 13126
rect 2228 12912 2280 12918
rect 2228 12854 2280 12860
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1952 11620 2004 11626
rect 1952 11562 2004 11568
rect 1964 11354 1992 11562
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 1872 10062 1900 10406
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 2056 6914 2084 12786
rect 2332 12374 2360 13194
rect 2320 12368 2372 12374
rect 2320 12310 2372 12316
rect 2136 12164 2188 12170
rect 2136 12106 2188 12112
rect 2148 11694 2176 12106
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2228 11552 2280 11558
rect 2332 11540 2360 12310
rect 2424 12170 2452 13330
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2280 11512 2360 11540
rect 2228 11494 2280 11500
rect 2148 10742 2176 11494
rect 2136 10736 2188 10742
rect 2136 10678 2188 10684
rect 2240 10674 2268 11494
rect 2516 11354 2544 18702
rect 5894 18524 6202 18533
rect 5894 18522 5900 18524
rect 5956 18522 5980 18524
rect 6036 18522 6060 18524
rect 6116 18522 6140 18524
rect 6196 18522 6202 18524
rect 5956 18470 5958 18522
rect 6138 18470 6140 18522
rect 5894 18468 5900 18470
rect 5956 18468 5980 18470
rect 6036 18468 6060 18470
rect 6116 18468 6140 18470
rect 6196 18468 6202 18470
rect 5894 18459 6202 18468
rect 10839 18524 11147 18533
rect 10839 18522 10845 18524
rect 10901 18522 10925 18524
rect 10981 18522 11005 18524
rect 11061 18522 11085 18524
rect 11141 18522 11147 18524
rect 10901 18470 10903 18522
rect 11083 18470 11085 18522
rect 10839 18468 10845 18470
rect 10901 18468 10925 18470
rect 10981 18468 11005 18470
rect 11061 18468 11085 18470
rect 11141 18468 11147 18470
rect 10839 18459 11147 18468
rect 15784 18524 16092 18533
rect 15784 18522 15790 18524
rect 15846 18522 15870 18524
rect 15926 18522 15950 18524
rect 16006 18522 16030 18524
rect 16086 18522 16092 18524
rect 15846 18470 15848 18522
rect 16028 18470 16030 18522
rect 15784 18468 15790 18470
rect 15846 18468 15870 18470
rect 15926 18468 15950 18470
rect 16006 18468 16030 18470
rect 16086 18468 16092 18470
rect 15784 18459 16092 18468
rect 20729 18524 21037 18533
rect 20729 18522 20735 18524
rect 20791 18522 20815 18524
rect 20871 18522 20895 18524
rect 20951 18522 20975 18524
rect 21031 18522 21037 18524
rect 20791 18470 20793 18522
rect 20973 18470 20975 18522
rect 20729 18468 20735 18470
rect 20791 18468 20815 18470
rect 20871 18468 20895 18470
rect 20951 18468 20975 18470
rect 21031 18468 21037 18470
rect 20729 18459 21037 18468
rect 3422 17980 3730 17989
rect 3422 17978 3428 17980
rect 3484 17978 3508 17980
rect 3564 17978 3588 17980
rect 3644 17978 3668 17980
rect 3724 17978 3730 17980
rect 3484 17926 3486 17978
rect 3666 17926 3668 17978
rect 3422 17924 3428 17926
rect 3484 17924 3508 17926
rect 3564 17924 3588 17926
rect 3644 17924 3668 17926
rect 3724 17924 3730 17926
rect 3422 17915 3730 17924
rect 8367 17980 8675 17989
rect 8367 17978 8373 17980
rect 8429 17978 8453 17980
rect 8509 17978 8533 17980
rect 8589 17978 8613 17980
rect 8669 17978 8675 17980
rect 8429 17926 8431 17978
rect 8611 17926 8613 17978
rect 8367 17924 8373 17926
rect 8429 17924 8453 17926
rect 8509 17924 8533 17926
rect 8589 17924 8613 17926
rect 8669 17924 8675 17926
rect 8367 17915 8675 17924
rect 13312 17980 13620 17989
rect 13312 17978 13318 17980
rect 13374 17978 13398 17980
rect 13454 17978 13478 17980
rect 13534 17978 13558 17980
rect 13614 17978 13620 17980
rect 13374 17926 13376 17978
rect 13556 17926 13558 17978
rect 13312 17924 13318 17926
rect 13374 17924 13398 17926
rect 13454 17924 13478 17926
rect 13534 17924 13558 17926
rect 13614 17924 13620 17926
rect 13312 17915 13620 17924
rect 18257 17980 18565 17989
rect 18257 17978 18263 17980
rect 18319 17978 18343 17980
rect 18399 17978 18423 17980
rect 18479 17978 18503 17980
rect 18559 17978 18565 17980
rect 18319 17926 18321 17978
rect 18501 17926 18503 17978
rect 18257 17924 18263 17926
rect 18319 17924 18343 17926
rect 18399 17924 18423 17926
rect 18479 17924 18503 17926
rect 18559 17924 18565 17926
rect 18257 17915 18565 17924
rect 5894 17436 6202 17445
rect 5894 17434 5900 17436
rect 5956 17434 5980 17436
rect 6036 17434 6060 17436
rect 6116 17434 6140 17436
rect 6196 17434 6202 17436
rect 5956 17382 5958 17434
rect 6138 17382 6140 17434
rect 5894 17380 5900 17382
rect 5956 17380 5980 17382
rect 6036 17380 6060 17382
rect 6116 17380 6140 17382
rect 6196 17380 6202 17382
rect 5894 17371 6202 17380
rect 10839 17436 11147 17445
rect 10839 17434 10845 17436
rect 10901 17434 10925 17436
rect 10981 17434 11005 17436
rect 11061 17434 11085 17436
rect 11141 17434 11147 17436
rect 10901 17382 10903 17434
rect 11083 17382 11085 17434
rect 10839 17380 10845 17382
rect 10901 17380 10925 17382
rect 10981 17380 11005 17382
rect 11061 17380 11085 17382
rect 11141 17380 11147 17382
rect 10839 17371 11147 17380
rect 15784 17436 16092 17445
rect 15784 17434 15790 17436
rect 15846 17434 15870 17436
rect 15926 17434 15950 17436
rect 16006 17434 16030 17436
rect 16086 17434 16092 17436
rect 15846 17382 15848 17434
rect 16028 17382 16030 17434
rect 15784 17380 15790 17382
rect 15846 17380 15870 17382
rect 15926 17380 15950 17382
rect 16006 17380 16030 17382
rect 16086 17380 16092 17382
rect 15784 17371 16092 17380
rect 20729 17436 21037 17445
rect 20729 17434 20735 17436
rect 20791 17434 20815 17436
rect 20871 17434 20895 17436
rect 20951 17434 20975 17436
rect 21031 17434 21037 17436
rect 20791 17382 20793 17434
rect 20973 17382 20975 17434
rect 20729 17380 20735 17382
rect 20791 17380 20815 17382
rect 20871 17380 20895 17382
rect 20951 17380 20975 17382
rect 21031 17380 21037 17382
rect 20729 17371 21037 17380
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 3068 15502 3096 17138
rect 4080 17066 4108 17138
rect 3332 17060 3384 17066
rect 3332 17002 3384 17008
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 3160 16590 3188 16934
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 3068 14958 3096 15438
rect 3160 15162 3188 16390
rect 3252 16182 3280 16526
rect 3344 16182 3372 17002
rect 3422 16892 3730 16901
rect 3422 16890 3428 16892
rect 3484 16890 3508 16892
rect 3564 16890 3588 16892
rect 3644 16890 3668 16892
rect 3724 16890 3730 16892
rect 3484 16838 3486 16890
rect 3666 16838 3668 16890
rect 3422 16836 3428 16838
rect 3484 16836 3508 16838
rect 3564 16836 3588 16838
rect 3644 16836 3668 16838
rect 3724 16836 3730 16838
rect 3422 16827 3730 16836
rect 4080 16726 4108 17002
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 5460 16658 5488 16934
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 3240 16176 3292 16182
rect 3240 16118 3292 16124
rect 3332 16176 3384 16182
rect 3332 16118 3384 16124
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3252 15502 3280 15846
rect 3344 15570 3372 16118
rect 3422 15804 3730 15813
rect 3422 15802 3428 15804
rect 3484 15802 3508 15804
rect 3564 15802 3588 15804
rect 3644 15802 3668 15804
rect 3724 15802 3730 15804
rect 3484 15750 3486 15802
rect 3666 15750 3668 15802
rect 3422 15748 3428 15750
rect 3484 15748 3508 15750
rect 3564 15748 3588 15750
rect 3644 15748 3668 15750
rect 3724 15748 3730 15750
rect 3422 15739 3730 15748
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3988 15502 4016 15642
rect 4080 15638 4108 16526
rect 4344 16516 4396 16522
rect 4344 16458 4396 16464
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3252 15094 3280 15438
rect 3700 15428 3752 15434
rect 3700 15370 3752 15376
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 3344 13938 3372 15302
rect 3712 15026 3740 15370
rect 3988 15026 4016 15438
rect 4080 15026 4108 15574
rect 4356 15570 4384 16458
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 4816 16046 4844 16390
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4816 15586 4844 15982
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4724 15558 4844 15586
rect 4724 15502 4752 15558
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4724 15026 4752 15438
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 5000 14958 5028 15302
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 3422 14716 3730 14725
rect 3422 14714 3428 14716
rect 3484 14714 3508 14716
rect 3564 14714 3588 14716
rect 3644 14714 3668 14716
rect 3724 14714 3730 14716
rect 3484 14662 3486 14714
rect 3666 14662 3668 14714
rect 3422 14660 3428 14662
rect 3484 14660 3508 14662
rect 3564 14660 3588 14662
rect 3644 14660 3668 14662
rect 3724 14660 3730 14662
rect 3422 14651 3730 14660
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12986 3188 13126
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2700 11626 2728 12786
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 1780 6886 1900 6914
rect 2056 6886 2176 6914
rect 1872 6798 1900 6886
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1596 5710 1624 6734
rect 2148 6662 2176 6886
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2608 6225 2636 11086
rect 2792 8090 2820 12854
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 3068 12238 3096 12650
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3068 11830 3096 12174
rect 3344 11898 3372 13670
rect 3422 13628 3730 13637
rect 3422 13626 3428 13628
rect 3484 13626 3508 13628
rect 3564 13626 3588 13628
rect 3644 13626 3668 13628
rect 3724 13626 3730 13628
rect 3484 13574 3486 13626
rect 3666 13574 3668 13626
rect 3422 13572 3428 13574
rect 3484 13572 3508 13574
rect 3564 13572 3588 13574
rect 3644 13572 3668 13574
rect 3724 13572 3730 13574
rect 3422 13563 3730 13572
rect 3804 12782 3832 13806
rect 3896 13530 3924 13874
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 3988 12918 4016 13262
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 4172 12850 4200 13262
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3422 12540 3730 12549
rect 3422 12538 3428 12540
rect 3484 12538 3508 12540
rect 3564 12538 3588 12540
rect 3644 12538 3668 12540
rect 3724 12538 3730 12540
rect 3484 12486 3486 12538
rect 3666 12486 3668 12538
rect 3422 12484 3428 12486
rect 3484 12484 3508 12486
rect 3564 12484 3588 12486
rect 3644 12484 3668 12486
rect 3724 12484 3730 12486
rect 3422 12475 3730 12484
rect 4264 12306 4292 14758
rect 4816 14006 4844 14826
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4908 13394 4936 14758
rect 5276 13938 5304 16390
rect 5460 16114 5488 16594
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5644 15706 5672 15982
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5736 15638 5764 16594
rect 5828 16590 5856 16730
rect 6012 16726 6040 17138
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6012 16590 6040 16662
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 6000 16584 6052 16590
rect 7300 16538 7328 16934
rect 7564 16720 7616 16726
rect 7564 16662 7616 16668
rect 6000 16526 6052 16532
rect 5828 16046 5856 16526
rect 7208 16522 7328 16538
rect 7196 16516 7328 16522
rect 7248 16510 7328 16516
rect 7196 16458 7248 16464
rect 5894 16348 6202 16357
rect 5894 16346 5900 16348
rect 5956 16346 5980 16348
rect 6036 16346 6060 16348
rect 6116 16346 6140 16348
rect 6196 16346 6202 16348
rect 5956 16294 5958 16346
rect 6138 16294 6140 16346
rect 5894 16292 5900 16294
rect 5956 16292 5980 16294
rect 6036 16292 6060 16294
rect 6116 16292 6140 16294
rect 6196 16292 6202 16294
rect 5894 16283 6202 16292
rect 7300 16114 7328 16510
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 5724 15632 5776 15638
rect 5724 15574 5776 15580
rect 5736 14346 5764 15574
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 5894 15260 6202 15269
rect 5894 15258 5900 15260
rect 5956 15258 5980 15260
rect 6036 15258 6060 15260
rect 6116 15258 6140 15260
rect 6196 15258 6202 15260
rect 5956 15206 5958 15258
rect 6138 15206 6140 15258
rect 5894 15204 5900 15206
rect 5956 15204 5980 15206
rect 6036 15204 6060 15206
rect 6116 15204 6140 15206
rect 6196 15204 6202 15206
rect 5894 15195 6202 15204
rect 6380 15094 6408 15370
rect 6368 15088 6420 15094
rect 6368 15030 6420 15036
rect 5724 14340 5776 14346
rect 5724 14282 5776 14288
rect 5894 14172 6202 14181
rect 5894 14170 5900 14172
rect 5956 14170 5980 14172
rect 6036 14170 6060 14172
rect 6116 14170 6140 14172
rect 6196 14170 6202 14172
rect 5956 14118 5958 14170
rect 6138 14118 6140 14170
rect 5894 14116 5900 14118
rect 5956 14116 5980 14118
rect 6036 14116 6060 14118
rect 6116 14116 6140 14118
rect 6196 14116 6202 14118
rect 5894 14107 6202 14116
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5092 12986 5120 13126
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2884 8974 2912 11494
rect 2976 11150 3004 11698
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 3068 11218 3096 11630
rect 3422 11452 3730 11461
rect 3422 11450 3428 11452
rect 3484 11450 3508 11452
rect 3564 11450 3588 11452
rect 3644 11450 3668 11452
rect 3724 11450 3730 11452
rect 3484 11398 3486 11450
rect 3666 11398 3668 11450
rect 3422 11396 3428 11398
rect 3484 11396 3508 11398
rect 3564 11396 3588 11398
rect 3644 11396 3668 11398
rect 3724 11396 3730 11398
rect 3422 11387 3730 11396
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2976 10810 3004 11086
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2976 10266 3004 10746
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 3068 9178 3096 11154
rect 3422 10364 3730 10373
rect 3422 10362 3428 10364
rect 3484 10362 3508 10364
rect 3564 10362 3588 10364
rect 3644 10362 3668 10364
rect 3724 10362 3730 10364
rect 3484 10310 3486 10362
rect 3666 10310 3668 10362
rect 3422 10308 3428 10310
rect 3484 10308 3508 10310
rect 3564 10308 3588 10310
rect 3644 10308 3668 10310
rect 3724 10308 3730 10310
rect 3422 10299 3730 10308
rect 3896 9450 3924 11698
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3988 9654 4016 11494
rect 4080 11218 4108 12174
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4448 11898 4476 12038
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4540 11694 4568 12106
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4540 11150 4568 11630
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4632 9654 4660 12582
rect 4816 12102 4844 12854
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3422 9276 3730 9285
rect 3422 9274 3428 9276
rect 3484 9274 3508 9276
rect 3564 9274 3588 9276
rect 3644 9274 3668 9276
rect 3724 9274 3730 9276
rect 3484 9222 3486 9274
rect 3666 9222 3668 9274
rect 3422 9220 3428 9222
rect 3484 9220 3508 9222
rect 3564 9220 3588 9222
rect 3644 9220 3668 9222
rect 3724 9220 3730 9222
rect 3422 9211 3730 9220
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 4448 8974 4476 9454
rect 4724 8974 4752 11494
rect 4816 9382 4844 12038
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 4908 11286 4936 11766
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5000 11354 5028 11698
rect 5184 11354 5212 12718
rect 5368 11830 5396 13806
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 13394 5488 13738
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5828 11762 5856 13126
rect 5894 13084 6202 13093
rect 5894 13082 5900 13084
rect 5956 13082 5980 13084
rect 6036 13082 6060 13084
rect 6116 13082 6140 13084
rect 6196 13082 6202 13084
rect 5956 13030 5958 13082
rect 6138 13030 6140 13082
rect 5894 13028 5900 13030
rect 5956 13028 5980 13030
rect 6036 13028 6060 13030
rect 6116 13028 6140 13030
rect 6196 13028 6202 13030
rect 5894 13019 6202 13028
rect 6288 12850 6316 13126
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 5894 11996 6202 12005
rect 5894 11994 5900 11996
rect 5956 11994 5980 11996
rect 6036 11994 6060 11996
rect 6116 11994 6140 11996
rect 6196 11994 6202 11996
rect 5956 11942 5958 11994
rect 6138 11942 6140 11994
rect 5894 11940 5900 11942
rect 5956 11940 5980 11942
rect 6036 11940 6060 11942
rect 6116 11940 6140 11942
rect 6196 11940 6202 11942
rect 5894 11931 6202 11940
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 3422 8188 3730 8197
rect 3422 8186 3428 8188
rect 3484 8186 3508 8188
rect 3564 8186 3588 8188
rect 3644 8186 3668 8188
rect 3724 8186 3730 8188
rect 3484 8134 3486 8186
rect 3666 8134 3668 8186
rect 3422 8132 3428 8134
rect 3484 8132 3508 8134
rect 3564 8132 3588 8134
rect 3644 8132 3668 8134
rect 3724 8132 3730 8134
rect 3422 8123 3730 8132
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 4448 7954 4476 8910
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 2700 7478 2728 7890
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2700 6322 2728 7414
rect 3422 7100 3730 7109
rect 3422 7098 3428 7100
rect 3484 7098 3508 7100
rect 3564 7098 3588 7100
rect 3644 7098 3668 7100
rect 3724 7098 3730 7100
rect 3484 7046 3486 7098
rect 3666 7046 3668 7098
rect 3422 7044 3428 7046
rect 3484 7044 3508 7046
rect 3564 7044 3588 7046
rect 3644 7044 3668 7046
rect 3724 7044 3730 7046
rect 3422 7035 3730 7044
rect 4448 6866 4476 7890
rect 4908 6914 4936 11222
rect 5184 11150 5212 11290
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 4540 6886 4936 6914
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 4252 6248 4304 6254
rect 2594 6216 2650 6225
rect 4252 6190 4304 6196
rect 2594 6151 2650 6160
rect 3422 6012 3730 6021
rect 3422 6010 3428 6012
rect 3484 6010 3508 6012
rect 3564 6010 3588 6012
rect 3644 6010 3668 6012
rect 3724 6010 3730 6012
rect 3484 5958 3486 6010
rect 3666 5958 3668 6010
rect 3422 5956 3428 5958
rect 3484 5956 3508 5958
rect 3564 5956 3588 5958
rect 3644 5956 3668 5958
rect 3724 5956 3730 5958
rect 3422 5947 3730 5956
rect 4264 5710 4292 6190
rect 4540 5710 4568 6886
rect 5448 6384 5500 6390
rect 5446 6352 5448 6361
rect 5500 6352 5502 6361
rect 5446 6287 5502 6296
rect 5644 5914 5672 11086
rect 5828 9178 5856 11698
rect 5894 10908 6202 10917
rect 5894 10906 5900 10908
rect 5956 10906 5980 10908
rect 6036 10906 6060 10908
rect 6116 10906 6140 10908
rect 6196 10906 6202 10908
rect 5956 10854 5958 10906
rect 6138 10854 6140 10906
rect 5894 10852 5900 10854
rect 5956 10852 5980 10854
rect 6036 10852 6060 10854
rect 6116 10852 6140 10854
rect 6196 10852 6202 10854
rect 5894 10843 6202 10852
rect 5894 9820 6202 9829
rect 5894 9818 5900 9820
rect 5956 9818 5980 9820
rect 6036 9818 6060 9820
rect 6116 9818 6140 9820
rect 6196 9818 6202 9820
rect 5956 9766 5958 9818
rect 6138 9766 6140 9818
rect 5894 9764 5900 9766
rect 5956 9764 5980 9766
rect 6036 9764 6060 9766
rect 6116 9764 6140 9766
rect 6196 9764 6202 9766
rect 5894 9755 6202 9764
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5894 8732 6202 8741
rect 5894 8730 5900 8732
rect 5956 8730 5980 8732
rect 6036 8730 6060 8732
rect 6116 8730 6140 8732
rect 6196 8730 6202 8732
rect 5956 8678 5958 8730
rect 6138 8678 6140 8730
rect 5894 8676 5900 8678
rect 5956 8676 5980 8678
rect 6036 8676 6060 8678
rect 6116 8676 6140 8678
rect 6196 8676 6202 8678
rect 5894 8667 6202 8676
rect 5894 7644 6202 7653
rect 5894 7642 5900 7644
rect 5956 7642 5980 7644
rect 6036 7642 6060 7644
rect 6116 7642 6140 7644
rect 6196 7642 6202 7644
rect 5956 7590 5958 7642
rect 6138 7590 6140 7642
rect 5894 7588 5900 7590
rect 5956 7588 5980 7590
rect 6036 7588 6060 7590
rect 6116 7588 6140 7590
rect 6196 7588 6202 7590
rect 5894 7579 6202 7588
rect 6380 6914 6408 15030
rect 6656 15026 6684 15438
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6472 14414 6500 14894
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6472 8090 6500 14350
rect 6748 13326 6776 15846
rect 6840 15706 6868 15982
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6748 12442 6776 13126
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6748 11694 6776 12174
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6380 6886 6500 6914
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 5894 6556 6202 6565
rect 5894 6554 5900 6556
rect 5956 6554 5980 6556
rect 6036 6554 6060 6556
rect 6116 6554 6140 6556
rect 6196 6554 6202 6556
rect 5956 6502 5958 6554
rect 6138 6502 6140 6554
rect 5894 6500 5900 6502
rect 5956 6500 5980 6502
rect 6036 6500 6060 6502
rect 6116 6500 6140 6502
rect 6196 6500 6202 6502
rect 5894 6491 6202 6500
rect 5906 6216 5962 6225
rect 5906 6151 5962 6160
rect 5920 6118 5948 6151
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 1596 5234 1624 5646
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1596 4078 1624 5170
rect 1872 4282 1900 5170
rect 4264 5166 4292 5646
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 2976 4214 3004 4966
rect 3422 4924 3730 4933
rect 3422 4922 3428 4924
rect 3484 4922 3508 4924
rect 3564 4922 3588 4924
rect 3644 4922 3668 4924
rect 3724 4922 3730 4924
rect 3484 4870 3486 4922
rect 3666 4870 3668 4922
rect 3422 4868 3428 4870
rect 3484 4868 3508 4870
rect 3564 4868 3588 4870
rect 3644 4868 3668 4870
rect 3724 4868 3730 4870
rect 3422 4859 3730 4868
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1596 3602 1624 4014
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1596 3126 1624 3538
rect 1872 3534 1900 4082
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1584 3120 1636 3126
rect 1584 3062 1636 3068
rect 1872 2446 1900 3470
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2424 2650 2452 3402
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 2976 2446 3004 4150
rect 4264 4146 4292 5102
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 3422 3836 3730 3845
rect 3422 3834 3428 3836
rect 3484 3834 3508 3836
rect 3564 3834 3588 3836
rect 3644 3834 3668 3836
rect 3724 3834 3730 3836
rect 3484 3782 3486 3834
rect 3666 3782 3668 3834
rect 3422 3780 3428 3782
rect 3484 3780 3508 3782
rect 3564 3780 3588 3782
rect 3644 3780 3668 3782
rect 3724 3780 3730 3782
rect 3422 3771 3730 3780
rect 4080 3738 4108 4082
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 3240 3664 3292 3670
rect 3238 3632 3240 3641
rect 3292 3632 3294 3641
rect 3238 3567 3294 3576
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3160 2446 3188 3334
rect 3422 2748 3730 2757
rect 3422 2746 3428 2748
rect 3484 2746 3508 2748
rect 3564 2746 3588 2748
rect 3644 2746 3668 2748
rect 3724 2746 3730 2748
rect 3484 2694 3486 2746
rect 3666 2694 3668 2746
rect 3422 2692 3428 2694
rect 3484 2692 3508 2694
rect 3564 2692 3588 2694
rect 3644 2692 3668 2694
rect 3724 2692 3730 2694
rect 3422 2683 3730 2692
rect 4172 2446 4200 3878
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4264 2650 4292 3470
rect 4540 3466 4568 5646
rect 5894 5468 6202 5477
rect 5894 5466 5900 5468
rect 5956 5466 5980 5468
rect 6036 5466 6060 5468
rect 6116 5466 6140 5468
rect 6196 5466 6202 5468
rect 5956 5414 5958 5466
rect 6138 5414 6140 5466
rect 5894 5412 5900 5414
rect 5956 5412 5980 5414
rect 6036 5412 6060 5414
rect 6116 5412 6140 5414
rect 6196 5412 6202 5414
rect 5894 5403 6202 5412
rect 5894 4380 6202 4389
rect 5894 4378 5900 4380
rect 5956 4378 5980 4380
rect 6036 4378 6060 4380
rect 6116 4378 6140 4380
rect 6196 4378 6202 4380
rect 5956 4326 5958 4378
rect 6138 4326 6140 4378
rect 5894 4324 5900 4326
rect 5956 4324 5980 4326
rect 6036 4324 6060 4326
rect 6116 4324 6140 4326
rect 6196 4324 6202 4326
rect 5894 4315 6202 4324
rect 6380 3670 6408 6666
rect 6472 6186 6500 6886
rect 6564 6798 6592 10950
rect 6840 9518 6868 15098
rect 6932 14958 6960 15506
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 7116 14346 7144 15574
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6932 13394 6960 14214
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6932 12238 6960 13194
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6932 11082 6960 12174
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 7024 11218 7052 11494
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6932 6662 6960 11018
rect 7116 7818 7144 12378
rect 7208 11898 7236 15846
rect 7392 15706 7420 16458
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7484 16114 7512 16390
rect 7576 16114 7604 16662
rect 7760 16590 7788 17070
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7760 15162 7788 16526
rect 8128 16522 8156 17138
rect 8367 16892 8675 16901
rect 8367 16890 8373 16892
rect 8429 16890 8453 16892
rect 8509 16890 8533 16892
rect 8589 16890 8613 16892
rect 8669 16890 8675 16892
rect 8429 16838 8431 16890
rect 8611 16838 8613 16890
rect 8367 16836 8373 16838
rect 8429 16836 8453 16838
rect 8509 16836 8533 16838
rect 8589 16836 8613 16838
rect 8669 16836 8675 16838
rect 8367 16827 8675 16836
rect 13312 16892 13620 16901
rect 13312 16890 13318 16892
rect 13374 16890 13398 16892
rect 13454 16890 13478 16892
rect 13534 16890 13558 16892
rect 13614 16890 13620 16892
rect 13374 16838 13376 16890
rect 13556 16838 13558 16890
rect 13312 16836 13318 16838
rect 13374 16836 13398 16838
rect 13454 16836 13478 16838
rect 13534 16836 13558 16838
rect 13614 16836 13620 16838
rect 13312 16827 13620 16836
rect 18257 16892 18565 16901
rect 18257 16890 18263 16892
rect 18319 16890 18343 16892
rect 18399 16890 18423 16892
rect 18479 16890 18503 16892
rect 18559 16890 18565 16892
rect 18319 16838 18321 16890
rect 18501 16838 18503 16890
rect 18257 16836 18263 16838
rect 18319 16836 18343 16838
rect 18399 16836 18423 16838
rect 18479 16836 18503 16838
rect 18559 16836 18565 16838
rect 18257 16827 18565 16836
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 8024 16244 8076 16250
rect 8024 16186 8076 16192
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 8036 15094 8064 16186
rect 8128 15434 8156 16458
rect 10839 16348 11147 16357
rect 10839 16346 10845 16348
rect 10901 16346 10925 16348
rect 10981 16346 11005 16348
rect 11061 16346 11085 16348
rect 11141 16346 11147 16348
rect 10901 16294 10903 16346
rect 11083 16294 11085 16346
rect 10839 16292 10845 16294
rect 10901 16292 10925 16294
rect 10981 16292 11005 16294
rect 11061 16292 11085 16294
rect 11141 16292 11147 16294
rect 10839 16283 11147 16292
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8367 15804 8675 15813
rect 8367 15802 8373 15804
rect 8429 15802 8453 15804
rect 8509 15802 8533 15804
rect 8589 15802 8613 15804
rect 8669 15802 8675 15804
rect 8429 15750 8431 15802
rect 8611 15750 8613 15802
rect 8367 15748 8373 15750
rect 8429 15748 8453 15750
rect 8509 15748 8533 15750
rect 8589 15748 8613 15750
rect 8669 15748 8675 15750
rect 8367 15739 8675 15748
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8024 15088 8076 15094
rect 7944 15048 8024 15076
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7300 12102 7328 12786
rect 7392 12782 7420 13330
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7392 11694 7420 12718
rect 7852 12442 7880 14962
rect 7944 12646 7972 15048
rect 8024 15030 8076 15036
rect 8128 14414 8156 15370
rect 8956 14958 8984 16050
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8367 14716 8675 14725
rect 8367 14714 8373 14716
rect 8429 14714 8453 14716
rect 8509 14714 8533 14716
rect 8589 14714 8613 14716
rect 8669 14714 8675 14716
rect 8429 14662 8431 14714
rect 8611 14662 8613 14714
rect 8367 14660 8373 14662
rect 8429 14660 8453 14662
rect 8509 14660 8533 14662
rect 8589 14660 8613 14662
rect 8669 14660 8675 14662
rect 8367 14651 8675 14660
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8036 12850 8064 13262
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 8128 12730 8156 14350
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8367 13628 8675 13637
rect 8367 13626 8373 13628
rect 8429 13626 8453 13628
rect 8509 13626 8533 13628
rect 8589 13626 8613 13628
rect 8669 13626 8675 13628
rect 8429 13574 8431 13626
rect 8611 13574 8613 13626
rect 8367 13572 8373 13574
rect 8429 13572 8453 13574
rect 8509 13572 8533 13574
rect 8589 13572 8613 13574
rect 8669 13572 8675 13574
rect 8367 13563 8675 13572
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8312 12782 8340 13262
rect 8772 12986 8800 13806
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8036 12702 8156 12730
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7852 9586 7880 9998
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7852 9042 7880 9522
rect 8036 9178 8064 12702
rect 8116 12640 8168 12646
rect 8312 12594 8340 12718
rect 8116 12582 8168 12588
rect 8128 11014 8156 12582
rect 8220 12566 8340 12594
rect 8220 11762 8248 12566
rect 8367 12540 8675 12549
rect 8367 12538 8373 12540
rect 8429 12538 8453 12540
rect 8509 12538 8533 12540
rect 8589 12538 8613 12540
rect 8669 12538 8675 12540
rect 8429 12486 8431 12538
rect 8611 12486 8613 12538
rect 8367 12484 8373 12486
rect 8429 12484 8453 12486
rect 8509 12484 8533 12486
rect 8589 12484 8613 12486
rect 8669 12484 8675 12486
rect 8367 12475 8675 12484
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8220 11082 8248 11698
rect 8367 11452 8675 11461
rect 8367 11450 8373 11452
rect 8429 11450 8453 11452
rect 8509 11450 8533 11452
rect 8589 11450 8613 11452
rect 8669 11450 8675 11452
rect 8429 11398 8431 11450
rect 8611 11398 8613 11450
rect 8367 11396 8373 11398
rect 8429 11396 8453 11398
rect 8509 11396 8533 11398
rect 8589 11396 8613 11398
rect 8669 11396 8675 11398
rect 8367 11387 8675 11396
rect 8772 11354 8800 11698
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 9994 8156 10950
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7852 7886 7880 8978
rect 8220 8090 8248 11018
rect 8367 10364 8675 10373
rect 8367 10362 8373 10364
rect 8429 10362 8453 10364
rect 8509 10362 8533 10364
rect 8589 10362 8613 10364
rect 8669 10362 8675 10364
rect 8429 10310 8431 10362
rect 8611 10310 8613 10362
rect 8367 10308 8373 10310
rect 8429 10308 8453 10310
rect 8509 10308 8533 10310
rect 8589 10308 8613 10310
rect 8669 10308 8675 10310
rect 8367 10299 8675 10308
rect 8864 9518 8892 14758
rect 8956 14482 8984 14894
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 8944 13388 8996 13394
rect 8944 13330 8996 13336
rect 8956 11558 8984 13330
rect 9048 12918 9076 13738
rect 9140 12986 9168 15030
rect 9876 15026 9904 15302
rect 10244 15162 10272 15438
rect 10336 15162 10364 15506
rect 10428 15502 10456 15982
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11152 15632 11204 15638
rect 11072 15592 11152 15620
rect 11072 15502 11100 15592
rect 11152 15574 11204 15580
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 11060 15496 11112 15502
rect 11256 15450 11284 15642
rect 11348 15502 11376 16526
rect 11612 16448 11664 16454
rect 11612 16390 11664 16396
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 11624 16114 11652 16390
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11612 15972 11664 15978
rect 11612 15914 11664 15920
rect 11624 15502 11652 15914
rect 11336 15496 11388 15502
rect 11060 15438 11112 15444
rect 11164 15434 11284 15450
rect 11152 15428 11284 15434
rect 11204 15422 11284 15428
rect 11152 15370 11204 15376
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9220 14884 9272 14890
rect 9220 14826 9272 14832
rect 9232 14414 9260 14826
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9140 12442 9168 12718
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8956 11150 8984 11494
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8367 9276 8675 9285
rect 8367 9274 8373 9276
rect 8429 9274 8453 9276
rect 8509 9274 8533 9276
rect 8589 9274 8613 9276
rect 8669 9274 8675 9276
rect 8429 9222 8431 9274
rect 8611 9222 8613 9274
rect 8367 9220 8373 9222
rect 8429 9220 8453 9222
rect 8509 9220 8533 9222
rect 8589 9220 8613 9222
rect 8669 9220 8675 9222
rect 8367 9211 8675 9220
rect 8367 8188 8675 8197
rect 8367 8186 8373 8188
rect 8429 8186 8453 8188
rect 8509 8186 8533 8188
rect 8589 8186 8613 8188
rect 8669 8186 8675 8188
rect 8429 8134 8431 8186
rect 8611 8134 8613 8186
rect 8367 8132 8373 8134
rect 8429 8132 8453 8134
rect 8509 8132 8533 8134
rect 8589 8132 8613 8134
rect 8669 8132 8675 8134
rect 8367 8123 8675 8132
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7668 6662 7696 7346
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6932 5030 6960 5306
rect 7116 5234 7144 5646
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 7116 4146 7144 5170
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 4528 3460 4580 3466
rect 4528 3402 4580 3408
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4540 2446 4568 3402
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5276 2378 5304 2926
rect 5368 2378 5396 3062
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5460 2650 5488 2994
rect 5644 2922 5672 3538
rect 5894 3292 6202 3301
rect 5894 3290 5900 3292
rect 5956 3290 5980 3292
rect 6036 3290 6060 3292
rect 6116 3290 6140 3292
rect 6196 3290 6202 3292
rect 5956 3238 5958 3290
rect 6138 3238 6140 3290
rect 5894 3236 5900 3238
rect 5956 3236 5980 3238
rect 6036 3236 6060 3238
rect 6116 3236 6140 3238
rect 6196 3236 6202 3238
rect 5894 3227 6202 3236
rect 6564 3058 6592 3878
rect 6920 3528 6972 3534
rect 7116 3516 7144 4082
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 6972 3488 7144 3516
rect 6920 3470 6972 3476
rect 7300 3194 7328 3878
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7668 3126 7696 6598
rect 7852 6322 7880 7822
rect 8367 7100 8675 7109
rect 8367 7098 8373 7100
rect 8429 7098 8453 7100
rect 8509 7098 8533 7100
rect 8589 7098 8613 7100
rect 8669 7098 8675 7100
rect 8429 7046 8431 7098
rect 8611 7046 8613 7098
rect 8367 7044 8373 7046
rect 8429 7044 8453 7046
rect 8509 7044 8533 7046
rect 8589 7044 8613 7046
rect 8669 7044 8675 7046
rect 8367 7035 8675 7044
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8220 6390 8248 6666
rect 9232 6458 9260 14214
rect 9324 14074 9352 14214
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9324 12850 9352 13262
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9508 11150 9536 11766
rect 9600 11762 9628 14350
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 9692 13462 9720 13942
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9508 10266 9536 11086
rect 9600 10470 9628 11698
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 10060 9586 10088 11494
rect 10336 11082 10364 11698
rect 10428 11082 10456 12174
rect 10520 11762 10548 12582
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11762 10640 12038
rect 10704 11762 10732 15302
rect 10839 15260 11147 15269
rect 10839 15258 10845 15260
rect 10901 15258 10925 15260
rect 10981 15258 11005 15260
rect 11061 15258 11085 15260
rect 11141 15258 11147 15260
rect 10901 15206 10903 15258
rect 11083 15206 11085 15258
rect 10839 15204 10845 15206
rect 10901 15204 10925 15206
rect 10981 15204 11005 15206
rect 11061 15204 11085 15206
rect 11141 15204 11147 15206
rect 10839 15195 11147 15204
rect 11256 14958 11284 15422
rect 11334 15464 11336 15473
rect 11520 15496 11572 15502
rect 11388 15464 11390 15473
rect 11520 15438 11572 15444
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11334 15399 11390 15408
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 10839 14172 11147 14181
rect 10839 14170 10845 14172
rect 10901 14170 10925 14172
rect 10981 14170 11005 14172
rect 11061 14170 11085 14172
rect 11141 14170 11147 14172
rect 10901 14118 10903 14170
rect 11083 14118 11085 14170
rect 10839 14116 10845 14118
rect 10901 14116 10925 14118
rect 10981 14116 11005 14118
rect 11061 14116 11085 14118
rect 11141 14116 11147 14118
rect 10839 14107 11147 14116
rect 10839 13084 11147 13093
rect 10839 13082 10845 13084
rect 10901 13082 10925 13084
rect 10981 13082 11005 13084
rect 11061 13082 11085 13084
rect 11141 13082 11147 13084
rect 10901 13030 10903 13082
rect 11083 13030 11085 13082
rect 10839 13028 10845 13030
rect 10901 13028 10925 13030
rect 10981 13028 11005 13030
rect 11061 13028 11085 13030
rect 11141 13028 11147 13030
rect 10839 13019 11147 13028
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10796 12170 10824 12786
rect 11256 12442 11284 14282
rect 11348 13870 11376 15399
rect 11532 15162 11560 15438
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 11440 13870 11468 15098
rect 11716 14890 11744 15982
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11808 15162 11836 15574
rect 11900 15434 11928 15982
rect 12452 15638 12480 16050
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 11888 15428 11940 15434
rect 11888 15370 11940 15376
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11900 15026 11928 15370
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 12256 15020 12308 15026
rect 12452 15008 12480 15574
rect 12452 14980 12664 15008
rect 12256 14962 12308 14968
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11624 13938 11652 14214
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11624 13394 11652 13874
rect 11716 13734 11744 14350
rect 11808 14278 11836 14962
rect 11900 14414 11928 14962
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 13870 11836 14214
rect 11900 14074 11928 14350
rect 12084 14074 12112 14758
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12084 13938 12112 14010
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11348 12714 11376 13126
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10839 11996 11147 12005
rect 10839 11994 10845 11996
rect 10901 11994 10925 11996
rect 10981 11994 11005 11996
rect 11061 11994 11085 11996
rect 11141 11994 11147 11996
rect 10901 11942 10903 11994
rect 11083 11942 11085 11994
rect 10839 11940 10845 11942
rect 10901 11940 10925 11942
rect 10981 11940 11005 11942
rect 11061 11940 11085 11942
rect 11141 11940 11147 11942
rect 10839 11931 11147 11940
rect 11256 11898 11284 12378
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 11348 11694 11376 12174
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11440 11354 11468 13262
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11532 12306 11560 13194
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10336 9654 10364 9998
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10336 8974 10364 9590
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10336 8566 10364 8910
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10336 7886 10364 8502
rect 10324 7880 10376 7886
rect 10428 7868 10456 11018
rect 10839 10908 11147 10917
rect 10839 10906 10845 10908
rect 10901 10906 10925 10908
rect 10981 10906 11005 10908
rect 11061 10906 11085 10908
rect 11141 10906 11147 10908
rect 10901 10854 10903 10906
rect 11083 10854 11085 10906
rect 10839 10852 10845 10854
rect 10901 10852 10925 10854
rect 10981 10852 11005 10854
rect 11061 10852 11085 10854
rect 11141 10852 11147 10854
rect 10839 10843 11147 10852
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10508 7880 10560 7886
rect 10428 7840 10508 7868
rect 10324 7822 10376 7828
rect 10508 7822 10560 7828
rect 10336 7478 10364 7822
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 10336 6798 10364 7414
rect 10612 6798 10640 10474
rect 10839 9820 11147 9829
rect 10839 9818 10845 9820
rect 10901 9818 10925 9820
rect 10981 9818 11005 9820
rect 11061 9818 11085 9820
rect 11141 9818 11147 9820
rect 10901 9766 10903 9818
rect 11083 9766 11085 9818
rect 10839 9764 10845 9766
rect 10901 9764 10925 9766
rect 10981 9764 11005 9766
rect 11061 9764 11085 9766
rect 11141 9764 11147 9766
rect 10839 9755 11147 9764
rect 10839 8732 11147 8741
rect 10839 8730 10845 8732
rect 10901 8730 10925 8732
rect 10981 8730 11005 8732
rect 11061 8730 11085 8732
rect 11141 8730 11147 8732
rect 10901 8678 10903 8730
rect 11083 8678 11085 8730
rect 10839 8676 10845 8678
rect 10901 8676 10925 8678
rect 10981 8676 11005 8678
rect 11061 8676 11085 8678
rect 11141 8676 11147 8678
rect 10839 8667 11147 8676
rect 11532 8498 11560 12242
rect 11808 11898 11836 13262
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11624 11218 11652 11698
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11716 11150 11744 11766
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11808 11150 11836 11630
rect 11900 11626 11928 13874
rect 12176 13462 12204 14894
rect 12268 14550 12296 14962
rect 12636 14822 12664 14980
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12256 14408 12308 14414
rect 12440 14408 12492 14414
rect 12256 14350 12308 14356
rect 12438 14376 12440 14385
rect 12492 14376 12494 14385
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 12268 13258 12296 14350
rect 12438 14311 12494 14320
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12452 12918 12480 13738
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12544 12646 12572 14010
rect 12728 12986 12756 16118
rect 13096 16114 13124 16390
rect 15784 16348 16092 16357
rect 15784 16346 15790 16348
rect 15846 16346 15870 16348
rect 15926 16346 15950 16348
rect 16006 16346 16030 16348
rect 16086 16346 16092 16348
rect 15846 16294 15848 16346
rect 16028 16294 16030 16346
rect 15784 16292 15790 16294
rect 15846 16292 15870 16294
rect 15926 16292 15950 16294
rect 16006 16292 16030 16294
rect 16086 16292 16092 16294
rect 15784 16283 16092 16292
rect 20729 16348 21037 16357
rect 20729 16346 20735 16348
rect 20791 16346 20815 16348
rect 20871 16346 20895 16348
rect 20951 16346 20975 16348
rect 21031 16346 21037 16348
rect 20791 16294 20793 16346
rect 20973 16294 20975 16346
rect 20729 16292 20735 16294
rect 20791 16292 20815 16294
rect 20871 16292 20895 16294
rect 20951 16292 20975 16294
rect 21031 16292 21037 16294
rect 20729 16283 21037 16292
rect 14464 16176 14516 16182
rect 14464 16118 14516 16124
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15094 12848 15846
rect 12898 15600 12954 15609
rect 12898 15535 12954 15544
rect 12912 15502 12940 15535
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12820 14074 12848 14894
rect 12912 14414 12940 15438
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12084 11830 12112 12174
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11900 11150 11928 11562
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11716 10742 11744 11086
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11716 10266 11744 10678
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11808 9178 11836 11086
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11900 8634 11928 11086
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12452 10538 12480 10746
rect 12440 10532 12492 10538
rect 12440 10474 12492 10480
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 10839 7644 11147 7653
rect 10839 7642 10845 7644
rect 10901 7642 10925 7644
rect 10981 7642 11005 7644
rect 11061 7642 11085 7644
rect 11141 7642 11147 7644
rect 10901 7590 10903 7642
rect 11083 7590 11085 7642
rect 10839 7588 10845 7590
rect 10901 7588 10925 7590
rect 10981 7588 11005 7590
rect 11061 7588 11085 7590
rect 11141 7588 11147 7590
rect 10839 7579 11147 7588
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 9784 6322 9812 6734
rect 10839 6556 11147 6565
rect 10839 6554 10845 6556
rect 10901 6554 10925 6556
rect 10981 6554 11005 6556
rect 11061 6554 11085 6556
rect 11141 6554 11147 6556
rect 10901 6502 10903 6554
rect 11083 6502 11085 6554
rect 10839 6500 10845 6502
rect 10901 6500 10925 6502
rect 10981 6500 11005 6502
rect 11061 6500 11085 6502
rect 11141 6500 11147 6502
rect 10839 6491 11147 6500
rect 11900 6390 11928 7686
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 8367 6012 8675 6021
rect 8367 6010 8373 6012
rect 8429 6010 8453 6012
rect 8509 6010 8533 6012
rect 8589 6010 8613 6012
rect 8669 6010 8675 6012
rect 8429 5958 8431 6010
rect 8611 5958 8613 6010
rect 8367 5956 8373 5958
rect 8429 5956 8453 5958
rect 8509 5956 8533 5958
rect 8589 5956 8613 5958
rect 8669 5956 8675 5958
rect 8367 5947 8675 5956
rect 9600 5914 9628 6054
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9784 5166 9812 5646
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 10839 5468 11147 5477
rect 10839 5466 10845 5468
rect 10901 5466 10925 5468
rect 10981 5466 11005 5468
rect 11061 5466 11085 5468
rect 11141 5466 11147 5468
rect 10901 5414 10903 5466
rect 11083 5414 11085 5466
rect 10839 5412 10845 5414
rect 10901 5412 10925 5414
rect 10981 5412 11005 5414
rect 11061 5412 11085 5414
rect 11141 5412 11147 5414
rect 10839 5403 11147 5412
rect 11348 5302 11376 5510
rect 12544 5302 12572 12378
rect 12728 12374 12756 12922
rect 12820 12782 12848 13806
rect 12912 13190 12940 14350
rect 13004 14278 13032 15302
rect 13096 14958 13124 16050
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13188 15638 13216 15982
rect 13312 15804 13620 15813
rect 13312 15802 13318 15804
rect 13374 15802 13398 15804
rect 13454 15802 13478 15804
rect 13534 15802 13558 15804
rect 13614 15802 13620 15804
rect 13374 15750 13376 15802
rect 13556 15750 13558 15802
rect 13312 15748 13318 15750
rect 13374 15748 13398 15750
rect 13454 15748 13478 15750
rect 13534 15748 13558 15750
rect 13614 15748 13620 15750
rect 13312 15739 13620 15748
rect 13176 15632 13228 15638
rect 13176 15574 13228 15580
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 13188 14822 13216 15574
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 13004 13938 13032 14214
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 13004 13326 13032 13670
rect 13096 13530 13124 14758
rect 13188 14618 13216 14758
rect 13312 14716 13620 14725
rect 13312 14714 13318 14716
rect 13374 14714 13398 14716
rect 13454 14714 13478 14716
rect 13534 14714 13558 14716
rect 13614 14714 13620 14716
rect 13374 14662 13376 14714
rect 13556 14662 13558 14714
rect 13312 14660 13318 14662
rect 13374 14660 13398 14662
rect 13454 14660 13478 14662
rect 13534 14660 13558 14662
rect 13614 14660 13620 14662
rect 13312 14651 13620 14660
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13360 14408 13412 14414
rect 13358 14376 13360 14385
rect 13412 14376 13414 14385
rect 13358 14311 13414 14320
rect 13372 13938 13400 14311
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13648 13802 13676 14962
rect 13740 14482 13768 15982
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13832 14929 13860 15370
rect 13818 14920 13874 14929
rect 13818 14855 13874 14864
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13312 13628 13620 13637
rect 13312 13626 13318 13628
rect 13374 13626 13398 13628
rect 13454 13626 13478 13628
rect 13534 13626 13558 13628
rect 13614 13626 13620 13628
rect 13374 13574 13376 13626
rect 13556 13574 13558 13626
rect 13312 13572 13318 13574
rect 13374 13572 13398 13574
rect 13454 13572 13478 13574
rect 13534 13572 13558 13574
rect 13614 13572 13620 13574
rect 13312 13563 13620 13572
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 13004 12850 13032 13262
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12728 11082 12756 11630
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12728 10674 12756 11018
rect 12820 10962 12848 12582
rect 13096 11082 13124 12854
rect 13188 12238 13216 13398
rect 13648 13326 13676 13738
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13312 12540 13620 12549
rect 13312 12538 13318 12540
rect 13374 12538 13398 12540
rect 13454 12538 13478 12540
rect 13534 12538 13558 12540
rect 13614 12538 13620 12540
rect 13374 12486 13376 12538
rect 13556 12486 13558 12538
rect 13312 12484 13318 12486
rect 13374 12484 13398 12486
rect 13454 12484 13478 12486
rect 13534 12484 13558 12486
rect 13614 12484 13620 12486
rect 13312 12475 13620 12484
rect 13648 12442 13676 12582
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11762 13216 12038
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13312 11452 13620 11461
rect 13312 11450 13318 11452
rect 13374 11450 13398 11452
rect 13454 11450 13478 11452
rect 13534 11450 13558 11452
rect 13614 11450 13620 11452
rect 13374 11398 13376 11450
rect 13556 11398 13558 11450
rect 13312 11396 13318 11398
rect 13374 11396 13398 11398
rect 13454 11396 13478 11398
rect 13534 11396 13558 11398
rect 13614 11396 13620 11398
rect 13312 11387 13620 11396
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 12820 10934 13032 10962
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 13004 10470 13032 10934
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 9994 13032 10406
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 13096 9042 13124 11018
rect 13312 10364 13620 10373
rect 13312 10362 13318 10364
rect 13374 10362 13398 10364
rect 13454 10362 13478 10364
rect 13534 10362 13558 10364
rect 13614 10362 13620 10364
rect 13374 10310 13376 10362
rect 13556 10310 13558 10362
rect 13312 10308 13318 10310
rect 13374 10308 13398 10310
rect 13454 10308 13478 10310
rect 13534 10308 13558 10310
rect 13614 10308 13620 10310
rect 13312 10299 13620 10308
rect 13740 10169 13768 13874
rect 13832 11898 13860 14855
rect 14384 14618 14412 16050
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 14108 12238 14136 12854
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 14016 10674 14044 12038
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13924 10266 13952 10542
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13542 10160 13598 10169
rect 13542 10095 13598 10104
rect 13726 10160 13782 10169
rect 13726 10095 13782 10104
rect 13556 10062 13584 10095
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13188 8974 13216 9318
rect 13312 9276 13620 9285
rect 13312 9274 13318 9276
rect 13374 9274 13398 9276
rect 13454 9274 13478 9276
rect 13534 9274 13558 9276
rect 13614 9274 13620 9276
rect 13374 9222 13376 9274
rect 13556 9222 13558 9274
rect 13312 9220 13318 9222
rect 13374 9220 13398 9222
rect 13454 9220 13478 9222
rect 13534 9220 13558 9222
rect 13614 9220 13620 9222
rect 13312 9211 13620 9220
rect 14108 9178 14136 11154
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14200 9110 14228 13126
rect 14292 12434 14320 14350
rect 14476 14074 14504 16118
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 14660 15502 14688 16050
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14844 15162 14872 16050
rect 15028 15706 15056 16050
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15120 15706 15148 15982
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14844 14618 14872 14962
rect 15028 14906 15056 15438
rect 15212 15026 15240 15846
rect 15672 15502 15700 15914
rect 18257 15804 18565 15813
rect 18257 15802 18263 15804
rect 18319 15802 18343 15804
rect 18399 15802 18423 15804
rect 18479 15802 18503 15804
rect 18559 15802 18565 15804
rect 18319 15750 18321 15802
rect 18501 15750 18503 15802
rect 18257 15748 18263 15750
rect 18319 15748 18343 15750
rect 18399 15748 18423 15750
rect 18479 15748 18503 15750
rect 18559 15748 18565 15750
rect 18257 15739 18565 15748
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 16764 15632 16816 15638
rect 16762 15600 16764 15609
rect 16816 15600 16818 15609
rect 16762 15535 16818 15544
rect 15292 15496 15344 15502
rect 15290 15464 15292 15473
rect 15660 15496 15712 15502
rect 15344 15464 15346 15473
rect 15660 15438 15712 15444
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 15290 15399 15346 15408
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15028 14878 15240 14906
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14648 14544 14700 14550
rect 14648 14486 14700 14492
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14372 12436 14424 12442
rect 14292 12406 14372 12434
rect 14372 12378 14424 12384
rect 14476 12238 14504 13806
rect 14568 12238 14596 14282
rect 14660 14074 14688 14486
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14292 10538 14320 12174
rect 14476 11354 14504 12174
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14292 10062 14320 10474
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13832 8498 13860 8842
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13924 8566 13952 8774
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13312 8188 13620 8197
rect 13312 8186 13318 8188
rect 13374 8186 13398 8188
rect 13454 8186 13478 8188
rect 13534 8186 13558 8188
rect 13614 8186 13620 8188
rect 13374 8134 13376 8186
rect 13556 8134 13558 8186
rect 13312 8132 13318 8134
rect 13374 8132 13398 8134
rect 13454 8132 13478 8134
rect 13534 8132 13558 8134
rect 13614 8132 13620 8134
rect 13312 8123 13620 8132
rect 13648 7886 13676 8230
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13188 7342 13216 7686
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12820 5234 12848 6054
rect 13004 5710 13032 6598
rect 13188 6458 13216 7278
rect 13312 7100 13620 7109
rect 13312 7098 13318 7100
rect 13374 7098 13398 7100
rect 13454 7098 13478 7100
rect 13534 7098 13558 7100
rect 13614 7098 13620 7100
rect 13374 7046 13376 7098
rect 13556 7046 13558 7098
rect 13312 7044 13318 7046
rect 13374 7044 13398 7046
rect 13454 7044 13478 7046
rect 13534 7044 13558 7046
rect 13614 7044 13620 7046
rect 13312 7035 13620 7044
rect 13740 6866 13768 7890
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 8367 4924 8675 4933
rect 8367 4922 8373 4924
rect 8429 4922 8453 4924
rect 8509 4922 8533 4924
rect 8589 4922 8613 4924
rect 8669 4922 8675 4924
rect 8429 4870 8431 4922
rect 8611 4870 8613 4922
rect 8367 4868 8373 4870
rect 8429 4868 8453 4870
rect 8509 4868 8533 4870
rect 8589 4868 8613 4870
rect 8669 4868 8675 4870
rect 8367 4859 8675 4868
rect 9692 4826 9720 4966
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9784 4622 9812 5102
rect 12912 5030 12940 5510
rect 13004 5098 13032 5510
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 13004 4622 13032 5034
rect 13188 4826 13216 6258
rect 13740 6254 13768 6802
rect 13832 6458 13860 7142
rect 13924 6798 13952 7210
rect 14016 7206 14044 8502
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14108 7154 14136 8434
rect 14280 7200 14332 7206
rect 14108 7148 14280 7154
rect 14108 7142 14332 7148
rect 14108 7126 14320 7142
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13312 6012 13620 6021
rect 13312 6010 13318 6012
rect 13374 6010 13398 6012
rect 13454 6010 13478 6012
rect 13534 6010 13558 6012
rect 13614 6010 13620 6012
rect 13374 5958 13376 6010
rect 13556 5958 13558 6010
rect 13312 5956 13318 5958
rect 13374 5956 13398 5958
rect 13454 5956 13478 5958
rect 13534 5956 13558 5958
rect 13614 5956 13620 5958
rect 13312 5947 13620 5956
rect 13924 5846 13952 6734
rect 14108 6390 14136 7126
rect 14384 7018 14412 11222
rect 14568 11150 14596 12174
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14660 10044 14688 12106
rect 14752 11762 14780 12242
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14752 10266 14780 11698
rect 14844 11694 14872 14350
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14844 10742 14872 11018
rect 14936 10742 14964 14486
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15028 11762 15056 12378
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14740 10056 14792 10062
rect 14660 10016 14740 10044
rect 14740 9998 14792 10004
rect 14752 9926 14780 9998
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14752 9450 14780 9862
rect 15120 9654 15148 12718
rect 15212 12102 15240 14878
rect 15304 14414 15332 15399
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15672 15008 15700 15302
rect 15784 15260 16092 15269
rect 15784 15258 15790 15260
rect 15846 15258 15870 15260
rect 15926 15258 15950 15260
rect 16006 15258 16030 15260
rect 16086 15258 16092 15260
rect 15846 15206 15848 15258
rect 16028 15206 16030 15258
rect 15784 15204 15790 15206
rect 15846 15204 15870 15206
rect 15926 15204 15950 15206
rect 16006 15204 16030 15206
rect 16086 15204 16092 15206
rect 15784 15195 16092 15204
rect 15752 15020 15804 15026
rect 15672 14980 15752 15008
rect 15752 14962 15804 14968
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15292 13252 15344 13258
rect 15396 13240 15424 14826
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 13326 15516 14214
rect 15580 14074 15608 14894
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15672 13682 15700 14758
rect 16120 14340 16172 14346
rect 16120 14282 16172 14288
rect 15784 14172 16092 14181
rect 15784 14170 15790 14172
rect 15846 14170 15870 14172
rect 15926 14170 15950 14172
rect 16006 14170 16030 14172
rect 16086 14170 16092 14172
rect 15846 14118 15848 14170
rect 16028 14118 16030 14170
rect 15784 14116 15790 14118
rect 15846 14116 15870 14118
rect 15926 14116 15950 14118
rect 16006 14116 16030 14118
rect 16086 14116 16092 14118
rect 15784 14107 16092 14116
rect 15580 13654 15700 13682
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15344 13212 15424 13240
rect 15292 13194 15344 13200
rect 15304 12918 15332 13194
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15304 12238 15332 12650
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15304 11558 15332 11698
rect 15488 11626 15516 12174
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15212 10674 15240 11494
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15108 9648 15160 9654
rect 15108 9590 15160 9596
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14476 7478 14504 8842
rect 14752 8498 14780 8910
rect 14936 8498 14964 8978
rect 15120 8498 15148 9590
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15212 9382 15240 9522
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14200 6990 14412 7018
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13648 5302 13676 5714
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13312 4924 13620 4933
rect 13312 4922 13318 4924
rect 13374 4922 13398 4924
rect 13454 4922 13478 4924
rect 13534 4922 13558 4924
rect 13614 4922 13620 4924
rect 13374 4870 13376 4922
rect 13556 4870 13558 4922
rect 13312 4868 13318 4870
rect 13374 4868 13398 4870
rect 13454 4868 13478 4870
rect 13534 4868 13558 4870
rect 13614 4868 13620 4870
rect 13312 4859 13620 4868
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 9784 4078 9812 4558
rect 10839 4380 11147 4389
rect 10839 4378 10845 4380
rect 10901 4378 10925 4380
rect 10981 4378 11005 4380
rect 11061 4378 11085 4380
rect 11141 4378 11147 4380
rect 10901 4326 10903 4378
rect 11083 4326 11085 4378
rect 10839 4324 10845 4326
rect 10901 4324 10925 4326
rect 10981 4324 11005 4326
rect 11061 4324 11085 4326
rect 11141 4324 11147 4326
rect 10839 4315 11147 4324
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8367 3836 8675 3845
rect 8367 3834 8373 3836
rect 8429 3834 8453 3836
rect 8509 3834 8533 3836
rect 8589 3834 8613 3836
rect 8669 3834 8675 3836
rect 8429 3782 8431 3834
rect 8611 3782 8613 3834
rect 8367 3780 8373 3782
rect 8429 3780 8453 3782
rect 8509 3780 8533 3782
rect 8589 3780 8613 3782
rect 8669 3780 8675 3782
rect 8367 3771 8675 3780
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5644 2650 5672 2858
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 6748 2446 6776 2926
rect 6840 2650 6868 2994
rect 8772 2990 8800 3878
rect 9784 3534 9812 4014
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9140 3194 9168 3470
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8367 2748 8675 2757
rect 8367 2746 8373 2748
rect 8429 2746 8453 2748
rect 8509 2746 8533 2748
rect 8589 2746 8613 2748
rect 8669 2746 8675 2748
rect 8429 2694 8431 2746
rect 8611 2694 8613 2746
rect 8367 2692 8373 2694
rect 8429 2692 8453 2694
rect 8509 2692 8533 2694
rect 8589 2692 8613 2694
rect 8669 2692 8675 2694
rect 8367 2683 8675 2692
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 8772 2446 8800 2926
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9692 2514 9720 2790
rect 9784 2514 9812 3470
rect 9876 3194 9904 4082
rect 13312 3836 13620 3845
rect 13312 3834 13318 3836
rect 13374 3834 13398 3836
rect 13454 3834 13478 3836
rect 13534 3834 13558 3836
rect 13614 3834 13620 3836
rect 13374 3782 13376 3834
rect 13556 3782 13558 3834
rect 13312 3780 13318 3782
rect 13374 3780 13398 3782
rect 13454 3780 13478 3782
rect 13534 3780 13558 3782
rect 13614 3780 13620 3782
rect 13312 3771 13620 3780
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12360 3602 12388 3674
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 10506 3496 10562 3505
rect 10506 3431 10562 3440
rect 10520 3398 10548 3431
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10152 3194 10180 3334
rect 10839 3292 11147 3301
rect 10839 3290 10845 3292
rect 10901 3290 10925 3292
rect 10981 3290 11005 3292
rect 11061 3290 11085 3292
rect 11141 3290 11147 3292
rect 10901 3238 10903 3290
rect 11083 3238 11085 3290
rect 10839 3236 10845 3238
rect 10901 3236 10925 3238
rect 10981 3236 11005 3238
rect 11061 3236 11085 3238
rect 11141 3236 11147 3238
rect 10839 3227 11147 3236
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 9968 2650 9996 2994
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 11072 2446 11100 3062
rect 12360 2446 12388 3538
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12452 2650 12480 2994
rect 13004 2854 13032 3538
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13280 2854 13308 3334
rect 13648 3058 13676 5238
rect 14200 5234 14228 6990
rect 14476 6934 14504 7414
rect 14844 7410 14872 8230
rect 15580 7886 15608 13654
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15936 13184 15988 13190
rect 16132 13172 16160 14282
rect 16500 13938 16528 15438
rect 16776 15026 16804 15535
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16212 13932 16264 13938
rect 16488 13932 16540 13938
rect 16264 13892 16344 13920
rect 16212 13874 16264 13880
rect 16316 13326 16344 13892
rect 16488 13874 16540 13880
rect 16500 13530 16528 13874
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 15988 13144 16160 13172
rect 15936 13126 15988 13132
rect 15672 11812 15700 13126
rect 15784 13084 16092 13093
rect 15784 13082 15790 13084
rect 15846 13082 15870 13084
rect 15926 13082 15950 13084
rect 16006 13082 16030 13084
rect 16086 13082 16092 13084
rect 15846 13030 15848 13082
rect 16028 13030 16030 13082
rect 15784 13028 15790 13030
rect 15846 13028 15870 13030
rect 15926 13028 15950 13030
rect 16006 13028 16030 13030
rect 16086 13028 16092 13030
rect 15784 13019 16092 13028
rect 16316 12986 16344 13262
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16408 12918 16436 13466
rect 16592 13326 16620 14350
rect 16868 13802 16896 15098
rect 17132 14952 17184 14958
rect 17130 14920 17132 14929
rect 17184 14920 17186 14929
rect 17420 14890 17448 15438
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17130 14855 17186 14864
rect 17408 14884 17460 14890
rect 16856 13796 16908 13802
rect 16856 13738 16908 13744
rect 16672 13728 16724 13734
rect 16672 13670 16724 13676
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15764 12442 15792 12650
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15784 11996 16092 12005
rect 15784 11994 15790 11996
rect 15846 11994 15870 11996
rect 15926 11994 15950 11996
rect 16006 11994 16030 11996
rect 16086 11994 16092 11996
rect 15846 11942 15848 11994
rect 16028 11942 16030 11994
rect 15784 11940 15790 11942
rect 15846 11940 15870 11942
rect 15926 11940 15950 11942
rect 16006 11940 16030 11942
rect 16086 11940 16092 11942
rect 15784 11931 16092 11940
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 15936 11824 15988 11830
rect 15672 11784 15936 11812
rect 15936 11766 15988 11772
rect 16040 11762 16068 11834
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16040 11626 16068 11698
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 16040 11098 16068 11562
rect 16132 11558 16160 11698
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16040 11070 16160 11098
rect 15784 10908 16092 10917
rect 15784 10906 15790 10908
rect 15846 10906 15870 10908
rect 15926 10906 15950 10908
rect 16006 10906 16030 10908
rect 16086 10906 16092 10908
rect 15846 10854 15848 10906
rect 16028 10854 16030 10906
rect 15784 10852 15790 10854
rect 15846 10852 15870 10854
rect 15926 10852 15950 10854
rect 16006 10852 16030 10854
rect 16086 10852 16092 10854
rect 15784 10843 16092 10852
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15856 10266 15884 10610
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 16040 10266 16068 10474
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15856 10169 15884 10202
rect 15842 10160 15898 10169
rect 15842 10095 15898 10104
rect 15784 9820 16092 9829
rect 15784 9818 15790 9820
rect 15846 9818 15870 9820
rect 15926 9818 15950 9820
rect 16006 9818 16030 9820
rect 16086 9818 16092 9820
rect 15846 9766 15848 9818
rect 16028 9766 16030 9818
rect 15784 9764 15790 9766
rect 15846 9764 15870 9766
rect 15926 9764 15950 9766
rect 16006 9764 16030 9766
rect 16086 9764 16092 9766
rect 15784 9755 16092 9764
rect 16132 9586 16160 11070
rect 16224 10674 16252 11494
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16408 9994 16436 12854
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16592 12102 16620 12242
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16500 11830 16528 12038
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 16592 11286 16620 12038
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16592 9994 16620 11222
rect 16684 10266 16712 13670
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17052 12918 17080 13262
rect 17144 12918 17172 14855
rect 17408 14826 17460 14832
rect 17420 14278 17448 14826
rect 17604 14414 17632 14894
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17776 13932 17828 13938
rect 17776 13874 17828 13880
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17512 13394 17540 13670
rect 17604 13410 17632 13738
rect 17696 13530 17724 13806
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17500 13388 17552 13394
rect 17604 13382 17724 13410
rect 17500 13330 17552 13336
rect 17696 13326 17724 13382
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17696 12986 17724 13262
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16868 11354 16896 11698
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16960 11014 16988 11494
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16960 10538 16988 10950
rect 17052 10606 17080 12582
rect 17328 12442 17356 12786
rect 17788 12442 17816 13874
rect 17880 12850 17908 15302
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 18064 14006 18092 14758
rect 18156 14414 18184 15642
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18257 14716 18565 14725
rect 18257 14714 18263 14716
rect 18319 14714 18343 14716
rect 18399 14714 18423 14716
rect 18479 14714 18503 14716
rect 18559 14714 18565 14716
rect 18319 14662 18321 14714
rect 18501 14662 18503 14714
rect 18257 14660 18263 14662
rect 18319 14660 18343 14662
rect 18399 14660 18423 14662
rect 18479 14660 18503 14662
rect 18559 14660 18565 14662
rect 18257 14651 18565 14660
rect 18616 14482 18644 14962
rect 18892 14890 18920 15506
rect 20729 15260 21037 15269
rect 20729 15258 20735 15260
rect 20791 15258 20815 15260
rect 20871 15258 20895 15260
rect 20951 15258 20975 15260
rect 21031 15258 21037 15260
rect 20791 15206 20793 15258
rect 20973 15206 20975 15258
rect 20729 15204 20735 15206
rect 20791 15204 20815 15206
rect 20871 15204 20895 15206
rect 20951 15204 20975 15206
rect 21031 15204 21037 15206
rect 20729 15195 21037 15204
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18604 14476 18656 14482
rect 18656 14436 18736 14464
rect 18604 14418 18656 14424
rect 18144 14408 18196 14414
rect 18196 14356 18276 14362
rect 18144 14350 18276 14356
rect 18156 14334 18276 14350
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18156 14006 18184 14214
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18248 13818 18276 14334
rect 18156 13790 18276 13818
rect 18156 13394 18184 13790
rect 18257 13628 18565 13637
rect 18257 13626 18263 13628
rect 18319 13626 18343 13628
rect 18399 13626 18423 13628
rect 18479 13626 18503 13628
rect 18559 13626 18565 13628
rect 18319 13574 18321 13626
rect 18501 13574 18503 13626
rect 18257 13572 18263 13574
rect 18319 13572 18343 13574
rect 18399 13572 18423 13574
rect 18479 13572 18503 13574
rect 18559 13572 18565 13574
rect 18257 13563 18565 13572
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18064 12918 18092 13262
rect 18708 12986 18736 14436
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17328 12238 17356 12378
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17972 11762 18000 12174
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 18064 11694 18092 12854
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18257 12540 18565 12549
rect 18257 12538 18263 12540
rect 18319 12538 18343 12540
rect 18399 12538 18423 12540
rect 18479 12538 18503 12540
rect 18559 12538 18565 12540
rect 18319 12486 18321 12538
rect 18501 12486 18503 12538
rect 18257 12484 18263 12486
rect 18319 12484 18343 12486
rect 18399 12484 18423 12486
rect 18479 12484 18503 12486
rect 18559 12484 18565 12486
rect 18257 12475 18565 12484
rect 18616 12238 18644 12786
rect 18708 12306 18736 12922
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18236 12232 18288 12238
rect 18156 12192 18236 12220
rect 18156 11830 18184 12192
rect 18236 12174 18288 12180
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18144 11824 18196 11830
rect 18144 11766 18196 11772
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 17972 11150 18000 11562
rect 18156 11354 18184 11766
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18257 11452 18565 11461
rect 18257 11450 18263 11452
rect 18319 11450 18343 11452
rect 18399 11450 18423 11452
rect 18479 11450 18503 11452
rect 18559 11450 18565 11452
rect 18319 11398 18321 11450
rect 18501 11398 18503 11450
rect 18257 11396 18263 11398
rect 18319 11396 18343 11398
rect 18399 11396 18423 11398
rect 18479 11396 18503 11398
rect 18559 11396 18565 11398
rect 18257 11387 18565 11396
rect 18616 11370 18644 11494
rect 18616 11354 18736 11370
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18616 11348 18748 11354
rect 18616 11342 18696 11348
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 18616 10674 18644 11342
rect 18696 11290 18748 11296
rect 18800 11218 18828 11698
rect 18892 11694 18920 13398
rect 18984 12714 19012 14962
rect 19260 14618 19288 14962
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19628 13258 19656 14214
rect 19904 13938 19932 14418
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 19904 13530 19932 13874
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19616 13252 19668 13258
rect 19616 13194 19668 13200
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19260 12850 19288 12922
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 18972 12708 19024 12714
rect 18972 12650 19024 12656
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18892 11218 18920 11630
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18708 10674 18736 11086
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 18257 10364 18565 10373
rect 18257 10362 18263 10364
rect 18319 10362 18343 10364
rect 18399 10362 18423 10364
rect 18479 10362 18503 10364
rect 18559 10362 18565 10364
rect 18319 10310 18321 10362
rect 18501 10310 18503 10362
rect 18257 10308 18263 10310
rect 18319 10308 18343 10310
rect 18399 10308 18423 10310
rect 18479 10308 18503 10310
rect 18559 10308 18565 10310
rect 18257 10299 18565 10308
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 16776 9654 16804 9998
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 18156 9586 18184 9998
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16684 8974 16712 9318
rect 18156 9178 18184 9522
rect 18257 9276 18565 9285
rect 18257 9274 18263 9276
rect 18319 9274 18343 9276
rect 18399 9274 18423 9276
rect 18479 9274 18503 9276
rect 18559 9274 18565 9276
rect 18319 9222 18321 9274
rect 18501 9222 18503 9274
rect 18257 9220 18263 9222
rect 18319 9220 18343 9222
rect 18399 9220 18423 9222
rect 18479 9220 18503 9222
rect 18559 9220 18565 9222
rect 18257 9211 18565 9220
rect 18800 9178 18828 11154
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 18892 10810 18920 11018
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18984 10742 19012 11834
rect 18972 10736 19024 10742
rect 18972 10678 19024 10684
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18892 9110 18920 9998
rect 18984 9586 19012 10678
rect 19076 10130 19104 12174
rect 19352 12170 19380 12718
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19352 11558 19380 12106
rect 19628 11898 19656 13194
rect 19720 12850 19748 13262
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19524 11824 19576 11830
rect 19720 11778 19748 12786
rect 19996 12374 20024 14350
rect 20729 14172 21037 14181
rect 20729 14170 20735 14172
rect 20791 14170 20815 14172
rect 20871 14170 20895 14172
rect 20951 14170 20975 14172
rect 21031 14170 21037 14172
rect 20791 14118 20793 14170
rect 20973 14118 20975 14170
rect 20729 14116 20735 14118
rect 20791 14116 20815 14118
rect 20871 14116 20895 14118
rect 20951 14116 20975 14118
rect 21031 14116 21037 14118
rect 20729 14107 21037 14116
rect 20729 13084 21037 13093
rect 20729 13082 20735 13084
rect 20791 13082 20815 13084
rect 20871 13082 20895 13084
rect 20951 13082 20975 13084
rect 21031 13082 21037 13084
rect 20791 13030 20793 13082
rect 20973 13030 20975 13082
rect 20729 13028 20735 13030
rect 20791 13028 20815 13030
rect 20871 13028 20895 13030
rect 20951 13028 20975 13030
rect 21031 13028 21037 13030
rect 20729 13019 21037 13028
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 19984 12368 20036 12374
rect 19984 12310 20036 12316
rect 20088 12238 20116 12582
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20729 11996 21037 12005
rect 20729 11994 20735 11996
rect 20791 11994 20815 11996
rect 20871 11994 20895 11996
rect 20951 11994 20975 11996
rect 21031 11994 21037 11996
rect 20791 11942 20793 11994
rect 20973 11942 20975 11994
rect 20729 11940 20735 11942
rect 20791 11940 20815 11942
rect 20871 11940 20895 11942
rect 20951 11940 20975 11942
rect 21031 11940 21037 11942
rect 20729 11931 21037 11940
rect 19576 11772 19748 11778
rect 19524 11766 19748 11772
rect 19536 11750 19748 11766
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18880 9104 18932 9110
rect 18880 9046 18932 9052
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15672 8090 15700 8842
rect 16316 8838 16344 8910
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 15784 8732 16092 8741
rect 15784 8730 15790 8732
rect 15846 8730 15870 8732
rect 15926 8730 15950 8732
rect 16006 8730 16030 8732
rect 16086 8730 16092 8732
rect 15846 8678 15848 8730
rect 16028 8678 16030 8730
rect 15784 8676 15790 8678
rect 15846 8676 15870 8678
rect 15926 8676 15950 8678
rect 16006 8676 16030 8678
rect 16086 8676 16092 8678
rect 15784 8667 16092 8676
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14464 6928 14516 6934
rect 14464 6870 14516 6876
rect 14844 6798 14872 7346
rect 15120 7206 15148 7754
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15212 6798 15240 7686
rect 15784 7644 16092 7653
rect 15784 7642 15790 7644
rect 15846 7642 15870 7644
rect 15926 7642 15950 7644
rect 16006 7642 16030 7644
rect 16086 7642 16092 7644
rect 15846 7590 15848 7642
rect 16028 7590 16030 7642
rect 15784 7588 15790 7590
rect 15846 7588 15870 7590
rect 15926 7588 15950 7590
rect 16006 7588 16030 7590
rect 16086 7588 16092 7590
rect 15784 7579 16092 7588
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15304 6798 15332 7278
rect 15948 7002 15976 7278
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 15120 6186 15148 6666
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15212 6458 15240 6598
rect 15304 6458 15332 6734
rect 15784 6556 16092 6565
rect 15784 6554 15790 6556
rect 15846 6554 15870 6556
rect 15926 6554 15950 6556
rect 16006 6554 16030 6556
rect 16086 6554 16092 6556
rect 15846 6502 15848 6554
rect 16028 6502 16030 6554
rect 15784 6500 15790 6502
rect 15846 6500 15870 6502
rect 15926 6500 15950 6502
rect 16006 6500 16030 6502
rect 16086 6500 16092 6502
rect 15784 6491 16092 6500
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 13924 3602 13952 4082
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12636 2446 12664 2790
rect 13312 2748 13620 2757
rect 13312 2746 13318 2748
rect 13374 2746 13398 2748
rect 13454 2746 13478 2748
rect 13534 2746 13558 2748
rect 13614 2746 13620 2748
rect 13374 2694 13376 2746
rect 13556 2694 13558 2746
rect 13312 2692 13318 2694
rect 13374 2692 13398 2694
rect 13454 2692 13478 2694
rect 13534 2692 13558 2694
rect 13614 2692 13620 2694
rect 13312 2683 13620 2692
rect 14016 2582 14044 2926
rect 14004 2576 14056 2582
rect 14004 2518 14056 2524
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 14016 2378 14044 2518
rect 14108 2514 14136 4082
rect 14292 3738 14320 5170
rect 14476 5030 14504 5170
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14384 4146 14412 4966
rect 14476 4146 14504 4966
rect 14568 4758 14596 5170
rect 15304 4826 15332 5170
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14384 3534 14412 4082
rect 14372 3528 14424 3534
rect 14568 3505 14596 4558
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14660 3534 14688 4082
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14648 3528 14700 3534
rect 14372 3470 14424 3476
rect 14554 3496 14610 3505
rect 14648 3470 14700 3476
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14554 3431 14610 3440
rect 14568 3398 14596 3431
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14568 2990 14596 3334
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 14660 2378 14688 3470
rect 14752 3058 14780 3470
rect 14844 3058 14872 3538
rect 15580 3534 15608 5782
rect 15784 5468 16092 5477
rect 15784 5466 15790 5468
rect 15846 5466 15870 5468
rect 15926 5466 15950 5468
rect 16006 5466 16030 5468
rect 16086 5466 16092 5468
rect 15846 5414 15848 5466
rect 16028 5414 16030 5466
rect 15784 5412 15790 5414
rect 15846 5412 15870 5414
rect 15926 5412 15950 5414
rect 16006 5412 16030 5414
rect 16086 5412 16092 5414
rect 15784 5403 16092 5412
rect 16316 5302 16344 8774
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16304 5296 16356 5302
rect 16304 5238 16356 5244
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15672 4758 15700 5170
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 16592 4486 16620 8434
rect 16684 8022 16712 8910
rect 16960 8362 16988 8910
rect 17052 8634 17080 8978
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16776 7546 16804 7822
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16868 7546 16896 7686
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16960 6322 16988 8298
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 17052 6730 17080 7890
rect 17144 7886 17172 8434
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17420 7410 17448 7890
rect 17880 7478 17908 8978
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 7954 18092 8774
rect 18156 8498 18184 8842
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18432 8498 18460 8774
rect 18892 8634 18920 9046
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18248 8378 18276 8434
rect 18156 8350 18276 8378
rect 18524 8378 18552 8434
rect 18696 8424 18748 8430
rect 18524 8350 18644 8378
rect 18696 8366 18748 8372
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17040 6724 17092 6730
rect 17040 6666 17092 6672
rect 17052 6322 17080 6666
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17420 6254 17448 7346
rect 18064 6390 18092 7890
rect 18156 7886 18184 8350
rect 18257 8188 18565 8197
rect 18257 8186 18263 8188
rect 18319 8186 18343 8188
rect 18399 8186 18423 8188
rect 18479 8186 18503 8188
rect 18559 8186 18565 8188
rect 18319 8134 18321 8186
rect 18501 8134 18503 8186
rect 18257 8132 18263 8134
rect 18319 8132 18343 8134
rect 18399 8132 18423 8134
rect 18479 8132 18503 8134
rect 18559 8132 18565 8134
rect 18257 8123 18565 8132
rect 18616 7886 18644 8350
rect 18708 7954 18736 8366
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18432 7478 18460 7822
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18616 7410 18644 7822
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18156 6798 18184 7142
rect 18257 7100 18565 7109
rect 18257 7098 18263 7100
rect 18319 7098 18343 7100
rect 18399 7098 18423 7100
rect 18479 7098 18503 7100
rect 18559 7098 18565 7100
rect 18319 7046 18321 7098
rect 18501 7046 18503 7098
rect 18257 7044 18263 7046
rect 18319 7044 18343 7046
rect 18399 7044 18423 7046
rect 18479 7044 18503 7046
rect 18559 7044 18565 7046
rect 18257 7035 18565 7044
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17420 5778 17448 6054
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16684 4826 16712 5578
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 15784 4380 16092 4389
rect 15784 4378 15790 4380
rect 15846 4378 15870 4380
rect 15926 4378 15950 4380
rect 16006 4378 16030 4380
rect 16086 4378 16092 4380
rect 15846 4326 15848 4378
rect 16028 4326 16030 4378
rect 15784 4324 15790 4326
rect 15846 4324 15870 4326
rect 15926 4324 15950 4326
rect 16006 4324 16030 4326
rect 16086 4324 16092 4326
rect 15784 4315 16092 4324
rect 16684 3738 16712 4490
rect 16776 4010 16804 4558
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16960 3534 16988 4762
rect 17052 4622 17080 5238
rect 17328 5166 17356 5646
rect 17420 5234 17448 5714
rect 17788 5710 17816 6190
rect 18257 6012 18565 6021
rect 18257 6010 18263 6012
rect 18319 6010 18343 6012
rect 18399 6010 18423 6012
rect 18479 6010 18503 6012
rect 18559 6010 18565 6012
rect 18319 5958 18321 6010
rect 18501 5958 18503 6010
rect 18257 5956 18263 5958
rect 18319 5956 18343 5958
rect 18399 5956 18423 5958
rect 18479 5956 18503 5958
rect 18559 5956 18565 5958
rect 18257 5947 18565 5956
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 17052 3670 17080 4558
rect 17144 4078 17172 4966
rect 17328 4826 17356 5102
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17224 4752 17276 4758
rect 17224 4694 17276 4700
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 17236 3534 17264 4694
rect 17420 3738 17448 5170
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17788 4826 17816 5102
rect 18257 4924 18565 4933
rect 18257 4922 18263 4924
rect 18319 4922 18343 4924
rect 18399 4922 18423 4924
rect 18479 4922 18503 4924
rect 18559 4922 18565 4924
rect 18319 4870 18321 4922
rect 18501 4870 18503 4922
rect 18257 4868 18263 4870
rect 18319 4868 18343 4870
rect 18399 4868 18423 4870
rect 18479 4868 18503 4870
rect 18559 4868 18565 4870
rect 18257 4859 18565 4868
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 18616 4622 18644 7142
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18708 6361 18736 6394
rect 18694 6352 18750 6361
rect 18800 6322 18828 6734
rect 18892 6322 18920 7686
rect 19076 7546 19104 10066
rect 19352 9450 19380 11494
rect 19536 10674 19564 11750
rect 20076 11620 20128 11626
rect 20076 11562 20128 11568
rect 20088 10674 20116 11562
rect 20729 10908 21037 10917
rect 20729 10906 20735 10908
rect 20791 10906 20815 10908
rect 20871 10906 20895 10908
rect 20951 10906 20975 10908
rect 21031 10906 21037 10908
rect 20791 10854 20793 10906
rect 20973 10854 20975 10906
rect 20729 10852 20735 10854
rect 20791 10852 20815 10854
rect 20871 10852 20895 10854
rect 20951 10852 20975 10854
rect 21031 10852 21037 10854
rect 20729 10843 21037 10852
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20088 9586 20116 10610
rect 20729 9820 21037 9829
rect 20729 9818 20735 9820
rect 20791 9818 20815 9820
rect 20871 9818 20895 9820
rect 20951 9818 20975 9820
rect 21031 9818 21037 9820
rect 20791 9766 20793 9818
rect 20973 9766 20975 9818
rect 20729 9764 20735 9766
rect 20791 9764 20815 9766
rect 20871 9764 20895 9766
rect 20951 9764 20975 9766
rect 21031 9764 21037 9766
rect 20729 9755 21037 9764
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 20729 8732 21037 8741
rect 20729 8730 20735 8732
rect 20791 8730 20815 8732
rect 20871 8730 20895 8732
rect 20951 8730 20975 8732
rect 21031 8730 21037 8732
rect 20791 8678 20793 8730
rect 20973 8678 20975 8730
rect 20729 8676 20735 8678
rect 20791 8676 20815 8678
rect 20871 8676 20895 8678
rect 20951 8676 20975 8678
rect 21031 8676 21037 8678
rect 20729 8667 21037 8676
rect 20729 7644 21037 7653
rect 20729 7642 20735 7644
rect 20791 7642 20815 7644
rect 20871 7642 20895 7644
rect 20951 7642 20975 7644
rect 21031 7642 21037 7644
rect 20791 7590 20793 7642
rect 20973 7590 20975 7642
rect 20729 7588 20735 7590
rect 20791 7588 20815 7590
rect 20871 7588 20895 7590
rect 20951 7588 20975 7590
rect 21031 7588 21037 7590
rect 20729 7579 21037 7588
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19076 6798 19104 7482
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 19076 6322 19104 6598
rect 19260 6458 19288 6802
rect 19904 6798 19932 7142
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 18694 6287 18750 6296
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 18800 5846 18828 6258
rect 19628 6225 19656 6734
rect 20729 6556 21037 6565
rect 20729 6554 20735 6556
rect 20791 6554 20815 6556
rect 20871 6554 20895 6556
rect 20951 6554 20975 6556
rect 21031 6554 21037 6556
rect 20791 6502 20793 6554
rect 20973 6502 20975 6554
rect 20729 6500 20735 6502
rect 20791 6500 20815 6502
rect 20871 6500 20895 6502
rect 20951 6500 20975 6502
rect 21031 6500 21037 6502
rect 20729 6491 21037 6500
rect 19614 6216 19670 6225
rect 19614 6151 19670 6160
rect 18788 5840 18840 5846
rect 18788 5782 18840 5788
rect 20729 5468 21037 5477
rect 20729 5466 20735 5468
rect 20791 5466 20815 5468
rect 20871 5466 20895 5468
rect 20951 5466 20975 5468
rect 21031 5466 21037 5468
rect 20791 5414 20793 5466
rect 20973 5414 20975 5466
rect 20729 5412 20735 5414
rect 20791 5412 20815 5414
rect 20871 5412 20895 5414
rect 20951 5412 20975 5414
rect 21031 5412 21037 5414
rect 20729 5403 21037 5412
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 17696 3534 17724 3606
rect 18064 3534 18092 4558
rect 20729 4380 21037 4389
rect 20729 4378 20735 4380
rect 20791 4378 20815 4380
rect 20871 4378 20895 4380
rect 20951 4378 20975 4380
rect 21031 4378 21037 4380
rect 20791 4326 20793 4378
rect 20973 4326 20975 4378
rect 20729 4324 20735 4326
rect 20791 4324 20815 4326
rect 20871 4324 20895 4326
rect 20951 4324 20975 4326
rect 21031 4324 21037 4326
rect 20729 4315 21037 4324
rect 18257 3836 18565 3845
rect 18257 3834 18263 3836
rect 18319 3834 18343 3836
rect 18399 3834 18423 3836
rect 18479 3834 18503 3836
rect 18559 3834 18565 3836
rect 18319 3782 18321 3834
rect 18501 3782 18503 3834
rect 18257 3780 18263 3782
rect 18319 3780 18343 3782
rect 18399 3780 18423 3782
rect 18479 3780 18503 3782
rect 18559 3780 18565 3782
rect 18257 3771 18565 3780
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14752 2378 14780 2994
rect 14844 2650 14872 2994
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 15396 2378 15424 3470
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15488 3126 15516 3334
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 15580 2446 15608 3470
rect 15784 3292 16092 3301
rect 15784 3290 15790 3292
rect 15846 3290 15870 3292
rect 15926 3290 15950 3292
rect 16006 3290 16030 3292
rect 16086 3290 16092 3292
rect 15846 3238 15848 3290
rect 16028 3238 16030 3290
rect 15784 3236 15790 3238
rect 15846 3236 15870 3238
rect 15926 3236 15950 3238
rect 16006 3236 16030 3238
rect 16086 3236 16092 3238
rect 15784 3227 16092 3236
rect 16960 3058 16988 3470
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 15672 2650 15700 2994
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 5356 2372 5408 2378
rect 5356 2314 5408 2320
rect 14004 2372 14056 2378
rect 14004 2314 14056 2320
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 14740 2372 14792 2378
rect 14740 2314 14792 2320
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 4160 2304 4212 2310
rect 4448 2258 4476 2314
rect 15856 2310 15884 2926
rect 15948 2446 15976 2994
rect 17236 2990 17264 3470
rect 17972 2990 18000 3470
rect 20729 3292 21037 3301
rect 20729 3290 20735 3292
rect 20791 3290 20815 3292
rect 20871 3290 20895 3292
rect 20951 3290 20975 3292
rect 21031 3290 21037 3292
rect 20791 3238 20793 3290
rect 20973 3238 20975 3290
rect 20729 3236 20735 3238
rect 20791 3236 20815 3238
rect 20871 3236 20895 3238
rect 20951 3236 20975 3238
rect 21031 3236 21037 3238
rect 20729 3227 21037 3236
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 18257 2748 18565 2757
rect 18257 2746 18263 2748
rect 18319 2746 18343 2748
rect 18399 2746 18423 2748
rect 18479 2746 18503 2748
rect 18559 2746 18565 2748
rect 18319 2694 18321 2746
rect 18501 2694 18503 2746
rect 18257 2692 18263 2694
rect 18319 2692 18343 2694
rect 18399 2692 18423 2694
rect 18479 2692 18503 2694
rect 18559 2692 18565 2694
rect 18257 2683 18565 2692
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 4212 2252 4476 2258
rect 4160 2246 4476 2252
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 4172 2230 4476 2246
rect 5894 2204 6202 2213
rect 5894 2202 5900 2204
rect 5956 2202 5980 2204
rect 6036 2202 6060 2204
rect 6116 2202 6140 2204
rect 6196 2202 6202 2204
rect 5956 2150 5958 2202
rect 6138 2150 6140 2202
rect 5894 2148 5900 2150
rect 5956 2148 5980 2150
rect 6036 2148 6060 2150
rect 6116 2148 6140 2150
rect 6196 2148 6202 2150
rect 5894 2139 6202 2148
rect 10839 2204 11147 2213
rect 10839 2202 10845 2204
rect 10901 2202 10925 2204
rect 10981 2202 11005 2204
rect 11061 2202 11085 2204
rect 11141 2202 11147 2204
rect 10901 2150 10903 2202
rect 11083 2150 11085 2202
rect 10839 2148 10845 2150
rect 10901 2148 10925 2150
rect 10981 2148 11005 2150
rect 11061 2148 11085 2150
rect 11141 2148 11147 2150
rect 10839 2139 11147 2148
rect 15784 2204 16092 2213
rect 15784 2202 15790 2204
rect 15846 2202 15870 2204
rect 15926 2202 15950 2204
rect 16006 2202 16030 2204
rect 16086 2202 16092 2204
rect 15846 2150 15848 2202
rect 16028 2150 16030 2202
rect 15784 2148 15790 2150
rect 15846 2148 15870 2150
rect 15926 2148 15950 2150
rect 16006 2148 16030 2150
rect 16086 2148 16092 2150
rect 15784 2139 16092 2148
rect 20729 2204 21037 2213
rect 20729 2202 20735 2204
rect 20791 2202 20815 2204
rect 20871 2202 20895 2204
rect 20951 2202 20975 2204
rect 21031 2202 21037 2204
rect 20791 2150 20793 2202
rect 20973 2150 20975 2202
rect 20729 2148 20735 2150
rect 20791 2148 20815 2150
rect 20871 2148 20895 2150
rect 20951 2148 20975 2150
rect 21031 2148 21037 2150
rect 20729 2139 21037 2148
<< via2 >>
rect 5900 19610 5956 19612
rect 5980 19610 6036 19612
rect 6060 19610 6116 19612
rect 6140 19610 6196 19612
rect 5900 19558 5946 19610
rect 5946 19558 5956 19610
rect 5980 19558 6010 19610
rect 6010 19558 6022 19610
rect 6022 19558 6036 19610
rect 6060 19558 6074 19610
rect 6074 19558 6086 19610
rect 6086 19558 6116 19610
rect 6140 19558 6150 19610
rect 6150 19558 6196 19610
rect 5900 19556 5956 19558
rect 5980 19556 6036 19558
rect 6060 19556 6116 19558
rect 6140 19556 6196 19558
rect 10845 19610 10901 19612
rect 10925 19610 10981 19612
rect 11005 19610 11061 19612
rect 11085 19610 11141 19612
rect 10845 19558 10891 19610
rect 10891 19558 10901 19610
rect 10925 19558 10955 19610
rect 10955 19558 10967 19610
rect 10967 19558 10981 19610
rect 11005 19558 11019 19610
rect 11019 19558 11031 19610
rect 11031 19558 11061 19610
rect 11085 19558 11095 19610
rect 11095 19558 11141 19610
rect 10845 19556 10901 19558
rect 10925 19556 10981 19558
rect 11005 19556 11061 19558
rect 11085 19556 11141 19558
rect 15790 19610 15846 19612
rect 15870 19610 15926 19612
rect 15950 19610 16006 19612
rect 16030 19610 16086 19612
rect 15790 19558 15836 19610
rect 15836 19558 15846 19610
rect 15870 19558 15900 19610
rect 15900 19558 15912 19610
rect 15912 19558 15926 19610
rect 15950 19558 15964 19610
rect 15964 19558 15976 19610
rect 15976 19558 16006 19610
rect 16030 19558 16040 19610
rect 16040 19558 16086 19610
rect 15790 19556 15846 19558
rect 15870 19556 15926 19558
rect 15950 19556 16006 19558
rect 16030 19556 16086 19558
rect 20735 19610 20791 19612
rect 20815 19610 20871 19612
rect 20895 19610 20951 19612
rect 20975 19610 21031 19612
rect 20735 19558 20781 19610
rect 20781 19558 20791 19610
rect 20815 19558 20845 19610
rect 20845 19558 20857 19610
rect 20857 19558 20871 19610
rect 20895 19558 20909 19610
rect 20909 19558 20921 19610
rect 20921 19558 20951 19610
rect 20975 19558 20985 19610
rect 20985 19558 21031 19610
rect 20735 19556 20791 19558
rect 20815 19556 20871 19558
rect 20895 19556 20951 19558
rect 20975 19556 21031 19558
rect 3428 19066 3484 19068
rect 3508 19066 3564 19068
rect 3588 19066 3644 19068
rect 3668 19066 3724 19068
rect 3428 19014 3474 19066
rect 3474 19014 3484 19066
rect 3508 19014 3538 19066
rect 3538 19014 3550 19066
rect 3550 19014 3564 19066
rect 3588 19014 3602 19066
rect 3602 19014 3614 19066
rect 3614 19014 3644 19066
rect 3668 19014 3678 19066
rect 3678 19014 3724 19066
rect 3428 19012 3484 19014
rect 3508 19012 3564 19014
rect 3588 19012 3644 19014
rect 3668 19012 3724 19014
rect 8373 19066 8429 19068
rect 8453 19066 8509 19068
rect 8533 19066 8589 19068
rect 8613 19066 8669 19068
rect 8373 19014 8419 19066
rect 8419 19014 8429 19066
rect 8453 19014 8483 19066
rect 8483 19014 8495 19066
rect 8495 19014 8509 19066
rect 8533 19014 8547 19066
rect 8547 19014 8559 19066
rect 8559 19014 8589 19066
rect 8613 19014 8623 19066
rect 8623 19014 8669 19066
rect 8373 19012 8429 19014
rect 8453 19012 8509 19014
rect 8533 19012 8589 19014
rect 8613 19012 8669 19014
rect 13318 19066 13374 19068
rect 13398 19066 13454 19068
rect 13478 19066 13534 19068
rect 13558 19066 13614 19068
rect 13318 19014 13364 19066
rect 13364 19014 13374 19066
rect 13398 19014 13428 19066
rect 13428 19014 13440 19066
rect 13440 19014 13454 19066
rect 13478 19014 13492 19066
rect 13492 19014 13504 19066
rect 13504 19014 13534 19066
rect 13558 19014 13568 19066
rect 13568 19014 13614 19066
rect 13318 19012 13374 19014
rect 13398 19012 13454 19014
rect 13478 19012 13534 19014
rect 13558 19012 13614 19014
rect 18263 19066 18319 19068
rect 18343 19066 18399 19068
rect 18423 19066 18479 19068
rect 18503 19066 18559 19068
rect 18263 19014 18309 19066
rect 18309 19014 18319 19066
rect 18343 19014 18373 19066
rect 18373 19014 18385 19066
rect 18385 19014 18399 19066
rect 18423 19014 18437 19066
rect 18437 19014 18449 19066
rect 18449 19014 18479 19066
rect 18503 19014 18513 19066
rect 18513 19014 18559 19066
rect 18263 19012 18319 19014
rect 18343 19012 18399 19014
rect 18423 19012 18479 19014
rect 18503 19012 18559 19014
rect 938 18264 994 18320
rect 938 10920 994 10976
rect 5900 18522 5956 18524
rect 5980 18522 6036 18524
rect 6060 18522 6116 18524
rect 6140 18522 6196 18524
rect 5900 18470 5946 18522
rect 5946 18470 5956 18522
rect 5980 18470 6010 18522
rect 6010 18470 6022 18522
rect 6022 18470 6036 18522
rect 6060 18470 6074 18522
rect 6074 18470 6086 18522
rect 6086 18470 6116 18522
rect 6140 18470 6150 18522
rect 6150 18470 6196 18522
rect 5900 18468 5956 18470
rect 5980 18468 6036 18470
rect 6060 18468 6116 18470
rect 6140 18468 6196 18470
rect 10845 18522 10901 18524
rect 10925 18522 10981 18524
rect 11005 18522 11061 18524
rect 11085 18522 11141 18524
rect 10845 18470 10891 18522
rect 10891 18470 10901 18522
rect 10925 18470 10955 18522
rect 10955 18470 10967 18522
rect 10967 18470 10981 18522
rect 11005 18470 11019 18522
rect 11019 18470 11031 18522
rect 11031 18470 11061 18522
rect 11085 18470 11095 18522
rect 11095 18470 11141 18522
rect 10845 18468 10901 18470
rect 10925 18468 10981 18470
rect 11005 18468 11061 18470
rect 11085 18468 11141 18470
rect 15790 18522 15846 18524
rect 15870 18522 15926 18524
rect 15950 18522 16006 18524
rect 16030 18522 16086 18524
rect 15790 18470 15836 18522
rect 15836 18470 15846 18522
rect 15870 18470 15900 18522
rect 15900 18470 15912 18522
rect 15912 18470 15926 18522
rect 15950 18470 15964 18522
rect 15964 18470 15976 18522
rect 15976 18470 16006 18522
rect 16030 18470 16040 18522
rect 16040 18470 16086 18522
rect 15790 18468 15846 18470
rect 15870 18468 15926 18470
rect 15950 18468 16006 18470
rect 16030 18468 16086 18470
rect 20735 18522 20791 18524
rect 20815 18522 20871 18524
rect 20895 18522 20951 18524
rect 20975 18522 21031 18524
rect 20735 18470 20781 18522
rect 20781 18470 20791 18522
rect 20815 18470 20845 18522
rect 20845 18470 20857 18522
rect 20857 18470 20871 18522
rect 20895 18470 20909 18522
rect 20909 18470 20921 18522
rect 20921 18470 20951 18522
rect 20975 18470 20985 18522
rect 20985 18470 21031 18522
rect 20735 18468 20791 18470
rect 20815 18468 20871 18470
rect 20895 18468 20951 18470
rect 20975 18468 21031 18470
rect 3428 17978 3484 17980
rect 3508 17978 3564 17980
rect 3588 17978 3644 17980
rect 3668 17978 3724 17980
rect 3428 17926 3474 17978
rect 3474 17926 3484 17978
rect 3508 17926 3538 17978
rect 3538 17926 3550 17978
rect 3550 17926 3564 17978
rect 3588 17926 3602 17978
rect 3602 17926 3614 17978
rect 3614 17926 3644 17978
rect 3668 17926 3678 17978
rect 3678 17926 3724 17978
rect 3428 17924 3484 17926
rect 3508 17924 3564 17926
rect 3588 17924 3644 17926
rect 3668 17924 3724 17926
rect 8373 17978 8429 17980
rect 8453 17978 8509 17980
rect 8533 17978 8589 17980
rect 8613 17978 8669 17980
rect 8373 17926 8419 17978
rect 8419 17926 8429 17978
rect 8453 17926 8483 17978
rect 8483 17926 8495 17978
rect 8495 17926 8509 17978
rect 8533 17926 8547 17978
rect 8547 17926 8559 17978
rect 8559 17926 8589 17978
rect 8613 17926 8623 17978
rect 8623 17926 8669 17978
rect 8373 17924 8429 17926
rect 8453 17924 8509 17926
rect 8533 17924 8589 17926
rect 8613 17924 8669 17926
rect 13318 17978 13374 17980
rect 13398 17978 13454 17980
rect 13478 17978 13534 17980
rect 13558 17978 13614 17980
rect 13318 17926 13364 17978
rect 13364 17926 13374 17978
rect 13398 17926 13428 17978
rect 13428 17926 13440 17978
rect 13440 17926 13454 17978
rect 13478 17926 13492 17978
rect 13492 17926 13504 17978
rect 13504 17926 13534 17978
rect 13558 17926 13568 17978
rect 13568 17926 13614 17978
rect 13318 17924 13374 17926
rect 13398 17924 13454 17926
rect 13478 17924 13534 17926
rect 13558 17924 13614 17926
rect 18263 17978 18319 17980
rect 18343 17978 18399 17980
rect 18423 17978 18479 17980
rect 18503 17978 18559 17980
rect 18263 17926 18309 17978
rect 18309 17926 18319 17978
rect 18343 17926 18373 17978
rect 18373 17926 18385 17978
rect 18385 17926 18399 17978
rect 18423 17926 18437 17978
rect 18437 17926 18449 17978
rect 18449 17926 18479 17978
rect 18503 17926 18513 17978
rect 18513 17926 18559 17978
rect 18263 17924 18319 17926
rect 18343 17924 18399 17926
rect 18423 17924 18479 17926
rect 18503 17924 18559 17926
rect 5900 17434 5956 17436
rect 5980 17434 6036 17436
rect 6060 17434 6116 17436
rect 6140 17434 6196 17436
rect 5900 17382 5946 17434
rect 5946 17382 5956 17434
rect 5980 17382 6010 17434
rect 6010 17382 6022 17434
rect 6022 17382 6036 17434
rect 6060 17382 6074 17434
rect 6074 17382 6086 17434
rect 6086 17382 6116 17434
rect 6140 17382 6150 17434
rect 6150 17382 6196 17434
rect 5900 17380 5956 17382
rect 5980 17380 6036 17382
rect 6060 17380 6116 17382
rect 6140 17380 6196 17382
rect 10845 17434 10901 17436
rect 10925 17434 10981 17436
rect 11005 17434 11061 17436
rect 11085 17434 11141 17436
rect 10845 17382 10891 17434
rect 10891 17382 10901 17434
rect 10925 17382 10955 17434
rect 10955 17382 10967 17434
rect 10967 17382 10981 17434
rect 11005 17382 11019 17434
rect 11019 17382 11031 17434
rect 11031 17382 11061 17434
rect 11085 17382 11095 17434
rect 11095 17382 11141 17434
rect 10845 17380 10901 17382
rect 10925 17380 10981 17382
rect 11005 17380 11061 17382
rect 11085 17380 11141 17382
rect 15790 17434 15846 17436
rect 15870 17434 15926 17436
rect 15950 17434 16006 17436
rect 16030 17434 16086 17436
rect 15790 17382 15836 17434
rect 15836 17382 15846 17434
rect 15870 17382 15900 17434
rect 15900 17382 15912 17434
rect 15912 17382 15926 17434
rect 15950 17382 15964 17434
rect 15964 17382 15976 17434
rect 15976 17382 16006 17434
rect 16030 17382 16040 17434
rect 16040 17382 16086 17434
rect 15790 17380 15846 17382
rect 15870 17380 15926 17382
rect 15950 17380 16006 17382
rect 16030 17380 16086 17382
rect 20735 17434 20791 17436
rect 20815 17434 20871 17436
rect 20895 17434 20951 17436
rect 20975 17434 21031 17436
rect 20735 17382 20781 17434
rect 20781 17382 20791 17434
rect 20815 17382 20845 17434
rect 20845 17382 20857 17434
rect 20857 17382 20871 17434
rect 20895 17382 20909 17434
rect 20909 17382 20921 17434
rect 20921 17382 20951 17434
rect 20975 17382 20985 17434
rect 20985 17382 21031 17434
rect 20735 17380 20791 17382
rect 20815 17380 20871 17382
rect 20895 17380 20951 17382
rect 20975 17380 21031 17382
rect 3428 16890 3484 16892
rect 3508 16890 3564 16892
rect 3588 16890 3644 16892
rect 3668 16890 3724 16892
rect 3428 16838 3474 16890
rect 3474 16838 3484 16890
rect 3508 16838 3538 16890
rect 3538 16838 3550 16890
rect 3550 16838 3564 16890
rect 3588 16838 3602 16890
rect 3602 16838 3614 16890
rect 3614 16838 3644 16890
rect 3668 16838 3678 16890
rect 3678 16838 3724 16890
rect 3428 16836 3484 16838
rect 3508 16836 3564 16838
rect 3588 16836 3644 16838
rect 3668 16836 3724 16838
rect 3428 15802 3484 15804
rect 3508 15802 3564 15804
rect 3588 15802 3644 15804
rect 3668 15802 3724 15804
rect 3428 15750 3474 15802
rect 3474 15750 3484 15802
rect 3508 15750 3538 15802
rect 3538 15750 3550 15802
rect 3550 15750 3564 15802
rect 3588 15750 3602 15802
rect 3602 15750 3614 15802
rect 3614 15750 3644 15802
rect 3668 15750 3678 15802
rect 3678 15750 3724 15802
rect 3428 15748 3484 15750
rect 3508 15748 3564 15750
rect 3588 15748 3644 15750
rect 3668 15748 3724 15750
rect 3428 14714 3484 14716
rect 3508 14714 3564 14716
rect 3588 14714 3644 14716
rect 3668 14714 3724 14716
rect 3428 14662 3474 14714
rect 3474 14662 3484 14714
rect 3508 14662 3538 14714
rect 3538 14662 3550 14714
rect 3550 14662 3564 14714
rect 3588 14662 3602 14714
rect 3602 14662 3614 14714
rect 3614 14662 3644 14714
rect 3668 14662 3678 14714
rect 3678 14662 3724 14714
rect 3428 14660 3484 14662
rect 3508 14660 3564 14662
rect 3588 14660 3644 14662
rect 3668 14660 3724 14662
rect 3428 13626 3484 13628
rect 3508 13626 3564 13628
rect 3588 13626 3644 13628
rect 3668 13626 3724 13628
rect 3428 13574 3474 13626
rect 3474 13574 3484 13626
rect 3508 13574 3538 13626
rect 3538 13574 3550 13626
rect 3550 13574 3564 13626
rect 3588 13574 3602 13626
rect 3602 13574 3614 13626
rect 3614 13574 3644 13626
rect 3668 13574 3678 13626
rect 3678 13574 3724 13626
rect 3428 13572 3484 13574
rect 3508 13572 3564 13574
rect 3588 13572 3644 13574
rect 3668 13572 3724 13574
rect 3428 12538 3484 12540
rect 3508 12538 3564 12540
rect 3588 12538 3644 12540
rect 3668 12538 3724 12540
rect 3428 12486 3474 12538
rect 3474 12486 3484 12538
rect 3508 12486 3538 12538
rect 3538 12486 3550 12538
rect 3550 12486 3564 12538
rect 3588 12486 3602 12538
rect 3602 12486 3614 12538
rect 3614 12486 3644 12538
rect 3668 12486 3678 12538
rect 3678 12486 3724 12538
rect 3428 12484 3484 12486
rect 3508 12484 3564 12486
rect 3588 12484 3644 12486
rect 3668 12484 3724 12486
rect 5900 16346 5956 16348
rect 5980 16346 6036 16348
rect 6060 16346 6116 16348
rect 6140 16346 6196 16348
rect 5900 16294 5946 16346
rect 5946 16294 5956 16346
rect 5980 16294 6010 16346
rect 6010 16294 6022 16346
rect 6022 16294 6036 16346
rect 6060 16294 6074 16346
rect 6074 16294 6086 16346
rect 6086 16294 6116 16346
rect 6140 16294 6150 16346
rect 6150 16294 6196 16346
rect 5900 16292 5956 16294
rect 5980 16292 6036 16294
rect 6060 16292 6116 16294
rect 6140 16292 6196 16294
rect 5900 15258 5956 15260
rect 5980 15258 6036 15260
rect 6060 15258 6116 15260
rect 6140 15258 6196 15260
rect 5900 15206 5946 15258
rect 5946 15206 5956 15258
rect 5980 15206 6010 15258
rect 6010 15206 6022 15258
rect 6022 15206 6036 15258
rect 6060 15206 6074 15258
rect 6074 15206 6086 15258
rect 6086 15206 6116 15258
rect 6140 15206 6150 15258
rect 6150 15206 6196 15258
rect 5900 15204 5956 15206
rect 5980 15204 6036 15206
rect 6060 15204 6116 15206
rect 6140 15204 6196 15206
rect 5900 14170 5956 14172
rect 5980 14170 6036 14172
rect 6060 14170 6116 14172
rect 6140 14170 6196 14172
rect 5900 14118 5946 14170
rect 5946 14118 5956 14170
rect 5980 14118 6010 14170
rect 6010 14118 6022 14170
rect 6022 14118 6036 14170
rect 6060 14118 6074 14170
rect 6074 14118 6086 14170
rect 6086 14118 6116 14170
rect 6140 14118 6150 14170
rect 6150 14118 6196 14170
rect 5900 14116 5956 14118
rect 5980 14116 6036 14118
rect 6060 14116 6116 14118
rect 6140 14116 6196 14118
rect 3428 11450 3484 11452
rect 3508 11450 3564 11452
rect 3588 11450 3644 11452
rect 3668 11450 3724 11452
rect 3428 11398 3474 11450
rect 3474 11398 3484 11450
rect 3508 11398 3538 11450
rect 3538 11398 3550 11450
rect 3550 11398 3564 11450
rect 3588 11398 3602 11450
rect 3602 11398 3614 11450
rect 3614 11398 3644 11450
rect 3668 11398 3678 11450
rect 3678 11398 3724 11450
rect 3428 11396 3484 11398
rect 3508 11396 3564 11398
rect 3588 11396 3644 11398
rect 3668 11396 3724 11398
rect 3428 10362 3484 10364
rect 3508 10362 3564 10364
rect 3588 10362 3644 10364
rect 3668 10362 3724 10364
rect 3428 10310 3474 10362
rect 3474 10310 3484 10362
rect 3508 10310 3538 10362
rect 3538 10310 3550 10362
rect 3550 10310 3564 10362
rect 3588 10310 3602 10362
rect 3602 10310 3614 10362
rect 3614 10310 3644 10362
rect 3668 10310 3678 10362
rect 3678 10310 3724 10362
rect 3428 10308 3484 10310
rect 3508 10308 3564 10310
rect 3588 10308 3644 10310
rect 3668 10308 3724 10310
rect 3428 9274 3484 9276
rect 3508 9274 3564 9276
rect 3588 9274 3644 9276
rect 3668 9274 3724 9276
rect 3428 9222 3474 9274
rect 3474 9222 3484 9274
rect 3508 9222 3538 9274
rect 3538 9222 3550 9274
rect 3550 9222 3564 9274
rect 3588 9222 3602 9274
rect 3602 9222 3614 9274
rect 3614 9222 3644 9274
rect 3668 9222 3678 9274
rect 3678 9222 3724 9274
rect 3428 9220 3484 9222
rect 3508 9220 3564 9222
rect 3588 9220 3644 9222
rect 3668 9220 3724 9222
rect 5900 13082 5956 13084
rect 5980 13082 6036 13084
rect 6060 13082 6116 13084
rect 6140 13082 6196 13084
rect 5900 13030 5946 13082
rect 5946 13030 5956 13082
rect 5980 13030 6010 13082
rect 6010 13030 6022 13082
rect 6022 13030 6036 13082
rect 6060 13030 6074 13082
rect 6074 13030 6086 13082
rect 6086 13030 6116 13082
rect 6140 13030 6150 13082
rect 6150 13030 6196 13082
rect 5900 13028 5956 13030
rect 5980 13028 6036 13030
rect 6060 13028 6116 13030
rect 6140 13028 6196 13030
rect 5900 11994 5956 11996
rect 5980 11994 6036 11996
rect 6060 11994 6116 11996
rect 6140 11994 6196 11996
rect 5900 11942 5946 11994
rect 5946 11942 5956 11994
rect 5980 11942 6010 11994
rect 6010 11942 6022 11994
rect 6022 11942 6036 11994
rect 6060 11942 6074 11994
rect 6074 11942 6086 11994
rect 6086 11942 6116 11994
rect 6140 11942 6150 11994
rect 6150 11942 6196 11994
rect 5900 11940 5956 11942
rect 5980 11940 6036 11942
rect 6060 11940 6116 11942
rect 6140 11940 6196 11942
rect 3428 8186 3484 8188
rect 3508 8186 3564 8188
rect 3588 8186 3644 8188
rect 3668 8186 3724 8188
rect 3428 8134 3474 8186
rect 3474 8134 3484 8186
rect 3508 8134 3538 8186
rect 3538 8134 3550 8186
rect 3550 8134 3564 8186
rect 3588 8134 3602 8186
rect 3602 8134 3614 8186
rect 3614 8134 3644 8186
rect 3668 8134 3678 8186
rect 3678 8134 3724 8186
rect 3428 8132 3484 8134
rect 3508 8132 3564 8134
rect 3588 8132 3644 8134
rect 3668 8132 3724 8134
rect 3428 7098 3484 7100
rect 3508 7098 3564 7100
rect 3588 7098 3644 7100
rect 3668 7098 3724 7100
rect 3428 7046 3474 7098
rect 3474 7046 3484 7098
rect 3508 7046 3538 7098
rect 3538 7046 3550 7098
rect 3550 7046 3564 7098
rect 3588 7046 3602 7098
rect 3602 7046 3614 7098
rect 3614 7046 3644 7098
rect 3668 7046 3678 7098
rect 3678 7046 3724 7098
rect 3428 7044 3484 7046
rect 3508 7044 3564 7046
rect 3588 7044 3644 7046
rect 3668 7044 3724 7046
rect 2594 6160 2650 6216
rect 3428 6010 3484 6012
rect 3508 6010 3564 6012
rect 3588 6010 3644 6012
rect 3668 6010 3724 6012
rect 3428 5958 3474 6010
rect 3474 5958 3484 6010
rect 3508 5958 3538 6010
rect 3538 5958 3550 6010
rect 3550 5958 3564 6010
rect 3588 5958 3602 6010
rect 3602 5958 3614 6010
rect 3614 5958 3644 6010
rect 3668 5958 3678 6010
rect 3678 5958 3724 6010
rect 3428 5956 3484 5958
rect 3508 5956 3564 5958
rect 3588 5956 3644 5958
rect 3668 5956 3724 5958
rect 5446 6332 5448 6352
rect 5448 6332 5500 6352
rect 5500 6332 5502 6352
rect 5446 6296 5502 6332
rect 5900 10906 5956 10908
rect 5980 10906 6036 10908
rect 6060 10906 6116 10908
rect 6140 10906 6196 10908
rect 5900 10854 5946 10906
rect 5946 10854 5956 10906
rect 5980 10854 6010 10906
rect 6010 10854 6022 10906
rect 6022 10854 6036 10906
rect 6060 10854 6074 10906
rect 6074 10854 6086 10906
rect 6086 10854 6116 10906
rect 6140 10854 6150 10906
rect 6150 10854 6196 10906
rect 5900 10852 5956 10854
rect 5980 10852 6036 10854
rect 6060 10852 6116 10854
rect 6140 10852 6196 10854
rect 5900 9818 5956 9820
rect 5980 9818 6036 9820
rect 6060 9818 6116 9820
rect 6140 9818 6196 9820
rect 5900 9766 5946 9818
rect 5946 9766 5956 9818
rect 5980 9766 6010 9818
rect 6010 9766 6022 9818
rect 6022 9766 6036 9818
rect 6060 9766 6074 9818
rect 6074 9766 6086 9818
rect 6086 9766 6116 9818
rect 6140 9766 6150 9818
rect 6150 9766 6196 9818
rect 5900 9764 5956 9766
rect 5980 9764 6036 9766
rect 6060 9764 6116 9766
rect 6140 9764 6196 9766
rect 5900 8730 5956 8732
rect 5980 8730 6036 8732
rect 6060 8730 6116 8732
rect 6140 8730 6196 8732
rect 5900 8678 5946 8730
rect 5946 8678 5956 8730
rect 5980 8678 6010 8730
rect 6010 8678 6022 8730
rect 6022 8678 6036 8730
rect 6060 8678 6074 8730
rect 6074 8678 6086 8730
rect 6086 8678 6116 8730
rect 6140 8678 6150 8730
rect 6150 8678 6196 8730
rect 5900 8676 5956 8678
rect 5980 8676 6036 8678
rect 6060 8676 6116 8678
rect 6140 8676 6196 8678
rect 5900 7642 5956 7644
rect 5980 7642 6036 7644
rect 6060 7642 6116 7644
rect 6140 7642 6196 7644
rect 5900 7590 5946 7642
rect 5946 7590 5956 7642
rect 5980 7590 6010 7642
rect 6010 7590 6022 7642
rect 6022 7590 6036 7642
rect 6060 7590 6074 7642
rect 6074 7590 6086 7642
rect 6086 7590 6116 7642
rect 6140 7590 6150 7642
rect 6150 7590 6196 7642
rect 5900 7588 5956 7590
rect 5980 7588 6036 7590
rect 6060 7588 6116 7590
rect 6140 7588 6196 7590
rect 5900 6554 5956 6556
rect 5980 6554 6036 6556
rect 6060 6554 6116 6556
rect 6140 6554 6196 6556
rect 5900 6502 5946 6554
rect 5946 6502 5956 6554
rect 5980 6502 6010 6554
rect 6010 6502 6022 6554
rect 6022 6502 6036 6554
rect 6060 6502 6074 6554
rect 6074 6502 6086 6554
rect 6086 6502 6116 6554
rect 6140 6502 6150 6554
rect 6150 6502 6196 6554
rect 5900 6500 5956 6502
rect 5980 6500 6036 6502
rect 6060 6500 6116 6502
rect 6140 6500 6196 6502
rect 5906 6160 5962 6216
rect 3428 4922 3484 4924
rect 3508 4922 3564 4924
rect 3588 4922 3644 4924
rect 3668 4922 3724 4924
rect 3428 4870 3474 4922
rect 3474 4870 3484 4922
rect 3508 4870 3538 4922
rect 3538 4870 3550 4922
rect 3550 4870 3564 4922
rect 3588 4870 3602 4922
rect 3602 4870 3614 4922
rect 3614 4870 3644 4922
rect 3668 4870 3678 4922
rect 3678 4870 3724 4922
rect 3428 4868 3484 4870
rect 3508 4868 3564 4870
rect 3588 4868 3644 4870
rect 3668 4868 3724 4870
rect 3428 3834 3484 3836
rect 3508 3834 3564 3836
rect 3588 3834 3644 3836
rect 3668 3834 3724 3836
rect 3428 3782 3474 3834
rect 3474 3782 3484 3834
rect 3508 3782 3538 3834
rect 3538 3782 3550 3834
rect 3550 3782 3564 3834
rect 3588 3782 3602 3834
rect 3602 3782 3614 3834
rect 3614 3782 3644 3834
rect 3668 3782 3678 3834
rect 3678 3782 3724 3834
rect 3428 3780 3484 3782
rect 3508 3780 3564 3782
rect 3588 3780 3644 3782
rect 3668 3780 3724 3782
rect 3238 3612 3240 3632
rect 3240 3612 3292 3632
rect 3292 3612 3294 3632
rect 3238 3576 3294 3612
rect 3428 2746 3484 2748
rect 3508 2746 3564 2748
rect 3588 2746 3644 2748
rect 3668 2746 3724 2748
rect 3428 2694 3474 2746
rect 3474 2694 3484 2746
rect 3508 2694 3538 2746
rect 3538 2694 3550 2746
rect 3550 2694 3564 2746
rect 3588 2694 3602 2746
rect 3602 2694 3614 2746
rect 3614 2694 3644 2746
rect 3668 2694 3678 2746
rect 3678 2694 3724 2746
rect 3428 2692 3484 2694
rect 3508 2692 3564 2694
rect 3588 2692 3644 2694
rect 3668 2692 3724 2694
rect 5900 5466 5956 5468
rect 5980 5466 6036 5468
rect 6060 5466 6116 5468
rect 6140 5466 6196 5468
rect 5900 5414 5946 5466
rect 5946 5414 5956 5466
rect 5980 5414 6010 5466
rect 6010 5414 6022 5466
rect 6022 5414 6036 5466
rect 6060 5414 6074 5466
rect 6074 5414 6086 5466
rect 6086 5414 6116 5466
rect 6140 5414 6150 5466
rect 6150 5414 6196 5466
rect 5900 5412 5956 5414
rect 5980 5412 6036 5414
rect 6060 5412 6116 5414
rect 6140 5412 6196 5414
rect 5900 4378 5956 4380
rect 5980 4378 6036 4380
rect 6060 4378 6116 4380
rect 6140 4378 6196 4380
rect 5900 4326 5946 4378
rect 5946 4326 5956 4378
rect 5980 4326 6010 4378
rect 6010 4326 6022 4378
rect 6022 4326 6036 4378
rect 6060 4326 6074 4378
rect 6074 4326 6086 4378
rect 6086 4326 6116 4378
rect 6140 4326 6150 4378
rect 6150 4326 6196 4378
rect 5900 4324 5956 4326
rect 5980 4324 6036 4326
rect 6060 4324 6116 4326
rect 6140 4324 6196 4326
rect 8373 16890 8429 16892
rect 8453 16890 8509 16892
rect 8533 16890 8589 16892
rect 8613 16890 8669 16892
rect 8373 16838 8419 16890
rect 8419 16838 8429 16890
rect 8453 16838 8483 16890
rect 8483 16838 8495 16890
rect 8495 16838 8509 16890
rect 8533 16838 8547 16890
rect 8547 16838 8559 16890
rect 8559 16838 8589 16890
rect 8613 16838 8623 16890
rect 8623 16838 8669 16890
rect 8373 16836 8429 16838
rect 8453 16836 8509 16838
rect 8533 16836 8589 16838
rect 8613 16836 8669 16838
rect 13318 16890 13374 16892
rect 13398 16890 13454 16892
rect 13478 16890 13534 16892
rect 13558 16890 13614 16892
rect 13318 16838 13364 16890
rect 13364 16838 13374 16890
rect 13398 16838 13428 16890
rect 13428 16838 13440 16890
rect 13440 16838 13454 16890
rect 13478 16838 13492 16890
rect 13492 16838 13504 16890
rect 13504 16838 13534 16890
rect 13558 16838 13568 16890
rect 13568 16838 13614 16890
rect 13318 16836 13374 16838
rect 13398 16836 13454 16838
rect 13478 16836 13534 16838
rect 13558 16836 13614 16838
rect 18263 16890 18319 16892
rect 18343 16890 18399 16892
rect 18423 16890 18479 16892
rect 18503 16890 18559 16892
rect 18263 16838 18309 16890
rect 18309 16838 18319 16890
rect 18343 16838 18373 16890
rect 18373 16838 18385 16890
rect 18385 16838 18399 16890
rect 18423 16838 18437 16890
rect 18437 16838 18449 16890
rect 18449 16838 18479 16890
rect 18503 16838 18513 16890
rect 18513 16838 18559 16890
rect 18263 16836 18319 16838
rect 18343 16836 18399 16838
rect 18423 16836 18479 16838
rect 18503 16836 18559 16838
rect 10845 16346 10901 16348
rect 10925 16346 10981 16348
rect 11005 16346 11061 16348
rect 11085 16346 11141 16348
rect 10845 16294 10891 16346
rect 10891 16294 10901 16346
rect 10925 16294 10955 16346
rect 10955 16294 10967 16346
rect 10967 16294 10981 16346
rect 11005 16294 11019 16346
rect 11019 16294 11031 16346
rect 11031 16294 11061 16346
rect 11085 16294 11095 16346
rect 11095 16294 11141 16346
rect 10845 16292 10901 16294
rect 10925 16292 10981 16294
rect 11005 16292 11061 16294
rect 11085 16292 11141 16294
rect 8373 15802 8429 15804
rect 8453 15802 8509 15804
rect 8533 15802 8589 15804
rect 8613 15802 8669 15804
rect 8373 15750 8419 15802
rect 8419 15750 8429 15802
rect 8453 15750 8483 15802
rect 8483 15750 8495 15802
rect 8495 15750 8509 15802
rect 8533 15750 8547 15802
rect 8547 15750 8559 15802
rect 8559 15750 8589 15802
rect 8613 15750 8623 15802
rect 8623 15750 8669 15802
rect 8373 15748 8429 15750
rect 8453 15748 8509 15750
rect 8533 15748 8589 15750
rect 8613 15748 8669 15750
rect 8373 14714 8429 14716
rect 8453 14714 8509 14716
rect 8533 14714 8589 14716
rect 8613 14714 8669 14716
rect 8373 14662 8419 14714
rect 8419 14662 8429 14714
rect 8453 14662 8483 14714
rect 8483 14662 8495 14714
rect 8495 14662 8509 14714
rect 8533 14662 8547 14714
rect 8547 14662 8559 14714
rect 8559 14662 8589 14714
rect 8613 14662 8623 14714
rect 8623 14662 8669 14714
rect 8373 14660 8429 14662
rect 8453 14660 8509 14662
rect 8533 14660 8589 14662
rect 8613 14660 8669 14662
rect 8373 13626 8429 13628
rect 8453 13626 8509 13628
rect 8533 13626 8589 13628
rect 8613 13626 8669 13628
rect 8373 13574 8419 13626
rect 8419 13574 8429 13626
rect 8453 13574 8483 13626
rect 8483 13574 8495 13626
rect 8495 13574 8509 13626
rect 8533 13574 8547 13626
rect 8547 13574 8559 13626
rect 8559 13574 8589 13626
rect 8613 13574 8623 13626
rect 8623 13574 8669 13626
rect 8373 13572 8429 13574
rect 8453 13572 8509 13574
rect 8533 13572 8589 13574
rect 8613 13572 8669 13574
rect 8373 12538 8429 12540
rect 8453 12538 8509 12540
rect 8533 12538 8589 12540
rect 8613 12538 8669 12540
rect 8373 12486 8419 12538
rect 8419 12486 8429 12538
rect 8453 12486 8483 12538
rect 8483 12486 8495 12538
rect 8495 12486 8509 12538
rect 8533 12486 8547 12538
rect 8547 12486 8559 12538
rect 8559 12486 8589 12538
rect 8613 12486 8623 12538
rect 8623 12486 8669 12538
rect 8373 12484 8429 12486
rect 8453 12484 8509 12486
rect 8533 12484 8589 12486
rect 8613 12484 8669 12486
rect 8373 11450 8429 11452
rect 8453 11450 8509 11452
rect 8533 11450 8589 11452
rect 8613 11450 8669 11452
rect 8373 11398 8419 11450
rect 8419 11398 8429 11450
rect 8453 11398 8483 11450
rect 8483 11398 8495 11450
rect 8495 11398 8509 11450
rect 8533 11398 8547 11450
rect 8547 11398 8559 11450
rect 8559 11398 8589 11450
rect 8613 11398 8623 11450
rect 8623 11398 8669 11450
rect 8373 11396 8429 11398
rect 8453 11396 8509 11398
rect 8533 11396 8589 11398
rect 8613 11396 8669 11398
rect 8373 10362 8429 10364
rect 8453 10362 8509 10364
rect 8533 10362 8589 10364
rect 8613 10362 8669 10364
rect 8373 10310 8419 10362
rect 8419 10310 8429 10362
rect 8453 10310 8483 10362
rect 8483 10310 8495 10362
rect 8495 10310 8509 10362
rect 8533 10310 8547 10362
rect 8547 10310 8559 10362
rect 8559 10310 8589 10362
rect 8613 10310 8623 10362
rect 8623 10310 8669 10362
rect 8373 10308 8429 10310
rect 8453 10308 8509 10310
rect 8533 10308 8589 10310
rect 8613 10308 8669 10310
rect 8373 9274 8429 9276
rect 8453 9274 8509 9276
rect 8533 9274 8589 9276
rect 8613 9274 8669 9276
rect 8373 9222 8419 9274
rect 8419 9222 8429 9274
rect 8453 9222 8483 9274
rect 8483 9222 8495 9274
rect 8495 9222 8509 9274
rect 8533 9222 8547 9274
rect 8547 9222 8559 9274
rect 8559 9222 8589 9274
rect 8613 9222 8623 9274
rect 8623 9222 8669 9274
rect 8373 9220 8429 9222
rect 8453 9220 8509 9222
rect 8533 9220 8589 9222
rect 8613 9220 8669 9222
rect 8373 8186 8429 8188
rect 8453 8186 8509 8188
rect 8533 8186 8589 8188
rect 8613 8186 8669 8188
rect 8373 8134 8419 8186
rect 8419 8134 8429 8186
rect 8453 8134 8483 8186
rect 8483 8134 8495 8186
rect 8495 8134 8509 8186
rect 8533 8134 8547 8186
rect 8547 8134 8559 8186
rect 8559 8134 8589 8186
rect 8613 8134 8623 8186
rect 8623 8134 8669 8186
rect 8373 8132 8429 8134
rect 8453 8132 8509 8134
rect 8533 8132 8589 8134
rect 8613 8132 8669 8134
rect 5900 3290 5956 3292
rect 5980 3290 6036 3292
rect 6060 3290 6116 3292
rect 6140 3290 6196 3292
rect 5900 3238 5946 3290
rect 5946 3238 5956 3290
rect 5980 3238 6010 3290
rect 6010 3238 6022 3290
rect 6022 3238 6036 3290
rect 6060 3238 6074 3290
rect 6074 3238 6086 3290
rect 6086 3238 6116 3290
rect 6140 3238 6150 3290
rect 6150 3238 6196 3290
rect 5900 3236 5956 3238
rect 5980 3236 6036 3238
rect 6060 3236 6116 3238
rect 6140 3236 6196 3238
rect 8373 7098 8429 7100
rect 8453 7098 8509 7100
rect 8533 7098 8589 7100
rect 8613 7098 8669 7100
rect 8373 7046 8419 7098
rect 8419 7046 8429 7098
rect 8453 7046 8483 7098
rect 8483 7046 8495 7098
rect 8495 7046 8509 7098
rect 8533 7046 8547 7098
rect 8547 7046 8559 7098
rect 8559 7046 8589 7098
rect 8613 7046 8623 7098
rect 8623 7046 8669 7098
rect 8373 7044 8429 7046
rect 8453 7044 8509 7046
rect 8533 7044 8589 7046
rect 8613 7044 8669 7046
rect 10845 15258 10901 15260
rect 10925 15258 10981 15260
rect 11005 15258 11061 15260
rect 11085 15258 11141 15260
rect 10845 15206 10891 15258
rect 10891 15206 10901 15258
rect 10925 15206 10955 15258
rect 10955 15206 10967 15258
rect 10967 15206 10981 15258
rect 11005 15206 11019 15258
rect 11019 15206 11031 15258
rect 11031 15206 11061 15258
rect 11085 15206 11095 15258
rect 11095 15206 11141 15258
rect 10845 15204 10901 15206
rect 10925 15204 10981 15206
rect 11005 15204 11061 15206
rect 11085 15204 11141 15206
rect 11334 15444 11336 15464
rect 11336 15444 11388 15464
rect 11388 15444 11390 15464
rect 11334 15408 11390 15444
rect 10845 14170 10901 14172
rect 10925 14170 10981 14172
rect 11005 14170 11061 14172
rect 11085 14170 11141 14172
rect 10845 14118 10891 14170
rect 10891 14118 10901 14170
rect 10925 14118 10955 14170
rect 10955 14118 10967 14170
rect 10967 14118 10981 14170
rect 11005 14118 11019 14170
rect 11019 14118 11031 14170
rect 11031 14118 11061 14170
rect 11085 14118 11095 14170
rect 11095 14118 11141 14170
rect 10845 14116 10901 14118
rect 10925 14116 10981 14118
rect 11005 14116 11061 14118
rect 11085 14116 11141 14118
rect 10845 13082 10901 13084
rect 10925 13082 10981 13084
rect 11005 13082 11061 13084
rect 11085 13082 11141 13084
rect 10845 13030 10891 13082
rect 10891 13030 10901 13082
rect 10925 13030 10955 13082
rect 10955 13030 10967 13082
rect 10967 13030 10981 13082
rect 11005 13030 11019 13082
rect 11019 13030 11031 13082
rect 11031 13030 11061 13082
rect 11085 13030 11095 13082
rect 11095 13030 11141 13082
rect 10845 13028 10901 13030
rect 10925 13028 10981 13030
rect 11005 13028 11061 13030
rect 11085 13028 11141 13030
rect 10845 11994 10901 11996
rect 10925 11994 10981 11996
rect 11005 11994 11061 11996
rect 11085 11994 11141 11996
rect 10845 11942 10891 11994
rect 10891 11942 10901 11994
rect 10925 11942 10955 11994
rect 10955 11942 10967 11994
rect 10967 11942 10981 11994
rect 11005 11942 11019 11994
rect 11019 11942 11031 11994
rect 11031 11942 11061 11994
rect 11085 11942 11095 11994
rect 11095 11942 11141 11994
rect 10845 11940 10901 11942
rect 10925 11940 10981 11942
rect 11005 11940 11061 11942
rect 11085 11940 11141 11942
rect 10845 10906 10901 10908
rect 10925 10906 10981 10908
rect 11005 10906 11061 10908
rect 11085 10906 11141 10908
rect 10845 10854 10891 10906
rect 10891 10854 10901 10906
rect 10925 10854 10955 10906
rect 10955 10854 10967 10906
rect 10967 10854 10981 10906
rect 11005 10854 11019 10906
rect 11019 10854 11031 10906
rect 11031 10854 11061 10906
rect 11085 10854 11095 10906
rect 11095 10854 11141 10906
rect 10845 10852 10901 10854
rect 10925 10852 10981 10854
rect 11005 10852 11061 10854
rect 11085 10852 11141 10854
rect 10845 9818 10901 9820
rect 10925 9818 10981 9820
rect 11005 9818 11061 9820
rect 11085 9818 11141 9820
rect 10845 9766 10891 9818
rect 10891 9766 10901 9818
rect 10925 9766 10955 9818
rect 10955 9766 10967 9818
rect 10967 9766 10981 9818
rect 11005 9766 11019 9818
rect 11019 9766 11031 9818
rect 11031 9766 11061 9818
rect 11085 9766 11095 9818
rect 11095 9766 11141 9818
rect 10845 9764 10901 9766
rect 10925 9764 10981 9766
rect 11005 9764 11061 9766
rect 11085 9764 11141 9766
rect 10845 8730 10901 8732
rect 10925 8730 10981 8732
rect 11005 8730 11061 8732
rect 11085 8730 11141 8732
rect 10845 8678 10891 8730
rect 10891 8678 10901 8730
rect 10925 8678 10955 8730
rect 10955 8678 10967 8730
rect 10967 8678 10981 8730
rect 11005 8678 11019 8730
rect 11019 8678 11031 8730
rect 11031 8678 11061 8730
rect 11085 8678 11095 8730
rect 11095 8678 11141 8730
rect 10845 8676 10901 8678
rect 10925 8676 10981 8678
rect 11005 8676 11061 8678
rect 11085 8676 11141 8678
rect 12438 14356 12440 14376
rect 12440 14356 12492 14376
rect 12492 14356 12494 14376
rect 12438 14320 12494 14356
rect 15790 16346 15846 16348
rect 15870 16346 15926 16348
rect 15950 16346 16006 16348
rect 16030 16346 16086 16348
rect 15790 16294 15836 16346
rect 15836 16294 15846 16346
rect 15870 16294 15900 16346
rect 15900 16294 15912 16346
rect 15912 16294 15926 16346
rect 15950 16294 15964 16346
rect 15964 16294 15976 16346
rect 15976 16294 16006 16346
rect 16030 16294 16040 16346
rect 16040 16294 16086 16346
rect 15790 16292 15846 16294
rect 15870 16292 15926 16294
rect 15950 16292 16006 16294
rect 16030 16292 16086 16294
rect 20735 16346 20791 16348
rect 20815 16346 20871 16348
rect 20895 16346 20951 16348
rect 20975 16346 21031 16348
rect 20735 16294 20781 16346
rect 20781 16294 20791 16346
rect 20815 16294 20845 16346
rect 20845 16294 20857 16346
rect 20857 16294 20871 16346
rect 20895 16294 20909 16346
rect 20909 16294 20921 16346
rect 20921 16294 20951 16346
rect 20975 16294 20985 16346
rect 20985 16294 21031 16346
rect 20735 16292 20791 16294
rect 20815 16292 20871 16294
rect 20895 16292 20951 16294
rect 20975 16292 21031 16294
rect 12898 15544 12954 15600
rect 10845 7642 10901 7644
rect 10925 7642 10981 7644
rect 11005 7642 11061 7644
rect 11085 7642 11141 7644
rect 10845 7590 10891 7642
rect 10891 7590 10901 7642
rect 10925 7590 10955 7642
rect 10955 7590 10967 7642
rect 10967 7590 10981 7642
rect 11005 7590 11019 7642
rect 11019 7590 11031 7642
rect 11031 7590 11061 7642
rect 11085 7590 11095 7642
rect 11095 7590 11141 7642
rect 10845 7588 10901 7590
rect 10925 7588 10981 7590
rect 11005 7588 11061 7590
rect 11085 7588 11141 7590
rect 10845 6554 10901 6556
rect 10925 6554 10981 6556
rect 11005 6554 11061 6556
rect 11085 6554 11141 6556
rect 10845 6502 10891 6554
rect 10891 6502 10901 6554
rect 10925 6502 10955 6554
rect 10955 6502 10967 6554
rect 10967 6502 10981 6554
rect 11005 6502 11019 6554
rect 11019 6502 11031 6554
rect 11031 6502 11061 6554
rect 11085 6502 11095 6554
rect 11095 6502 11141 6554
rect 10845 6500 10901 6502
rect 10925 6500 10981 6502
rect 11005 6500 11061 6502
rect 11085 6500 11141 6502
rect 8373 6010 8429 6012
rect 8453 6010 8509 6012
rect 8533 6010 8589 6012
rect 8613 6010 8669 6012
rect 8373 5958 8419 6010
rect 8419 5958 8429 6010
rect 8453 5958 8483 6010
rect 8483 5958 8495 6010
rect 8495 5958 8509 6010
rect 8533 5958 8547 6010
rect 8547 5958 8559 6010
rect 8559 5958 8589 6010
rect 8613 5958 8623 6010
rect 8623 5958 8669 6010
rect 8373 5956 8429 5958
rect 8453 5956 8509 5958
rect 8533 5956 8589 5958
rect 8613 5956 8669 5958
rect 10845 5466 10901 5468
rect 10925 5466 10981 5468
rect 11005 5466 11061 5468
rect 11085 5466 11141 5468
rect 10845 5414 10891 5466
rect 10891 5414 10901 5466
rect 10925 5414 10955 5466
rect 10955 5414 10967 5466
rect 10967 5414 10981 5466
rect 11005 5414 11019 5466
rect 11019 5414 11031 5466
rect 11031 5414 11061 5466
rect 11085 5414 11095 5466
rect 11095 5414 11141 5466
rect 10845 5412 10901 5414
rect 10925 5412 10981 5414
rect 11005 5412 11061 5414
rect 11085 5412 11141 5414
rect 13318 15802 13374 15804
rect 13398 15802 13454 15804
rect 13478 15802 13534 15804
rect 13558 15802 13614 15804
rect 13318 15750 13364 15802
rect 13364 15750 13374 15802
rect 13398 15750 13428 15802
rect 13428 15750 13440 15802
rect 13440 15750 13454 15802
rect 13478 15750 13492 15802
rect 13492 15750 13504 15802
rect 13504 15750 13534 15802
rect 13558 15750 13568 15802
rect 13568 15750 13614 15802
rect 13318 15748 13374 15750
rect 13398 15748 13454 15750
rect 13478 15748 13534 15750
rect 13558 15748 13614 15750
rect 13318 14714 13374 14716
rect 13398 14714 13454 14716
rect 13478 14714 13534 14716
rect 13558 14714 13614 14716
rect 13318 14662 13364 14714
rect 13364 14662 13374 14714
rect 13398 14662 13428 14714
rect 13428 14662 13440 14714
rect 13440 14662 13454 14714
rect 13478 14662 13492 14714
rect 13492 14662 13504 14714
rect 13504 14662 13534 14714
rect 13558 14662 13568 14714
rect 13568 14662 13614 14714
rect 13318 14660 13374 14662
rect 13398 14660 13454 14662
rect 13478 14660 13534 14662
rect 13558 14660 13614 14662
rect 13358 14356 13360 14376
rect 13360 14356 13412 14376
rect 13412 14356 13414 14376
rect 13358 14320 13414 14356
rect 13818 14864 13874 14920
rect 13318 13626 13374 13628
rect 13398 13626 13454 13628
rect 13478 13626 13534 13628
rect 13558 13626 13614 13628
rect 13318 13574 13364 13626
rect 13364 13574 13374 13626
rect 13398 13574 13428 13626
rect 13428 13574 13440 13626
rect 13440 13574 13454 13626
rect 13478 13574 13492 13626
rect 13492 13574 13504 13626
rect 13504 13574 13534 13626
rect 13558 13574 13568 13626
rect 13568 13574 13614 13626
rect 13318 13572 13374 13574
rect 13398 13572 13454 13574
rect 13478 13572 13534 13574
rect 13558 13572 13614 13574
rect 13318 12538 13374 12540
rect 13398 12538 13454 12540
rect 13478 12538 13534 12540
rect 13558 12538 13614 12540
rect 13318 12486 13364 12538
rect 13364 12486 13374 12538
rect 13398 12486 13428 12538
rect 13428 12486 13440 12538
rect 13440 12486 13454 12538
rect 13478 12486 13492 12538
rect 13492 12486 13504 12538
rect 13504 12486 13534 12538
rect 13558 12486 13568 12538
rect 13568 12486 13614 12538
rect 13318 12484 13374 12486
rect 13398 12484 13454 12486
rect 13478 12484 13534 12486
rect 13558 12484 13614 12486
rect 13318 11450 13374 11452
rect 13398 11450 13454 11452
rect 13478 11450 13534 11452
rect 13558 11450 13614 11452
rect 13318 11398 13364 11450
rect 13364 11398 13374 11450
rect 13398 11398 13428 11450
rect 13428 11398 13440 11450
rect 13440 11398 13454 11450
rect 13478 11398 13492 11450
rect 13492 11398 13504 11450
rect 13504 11398 13534 11450
rect 13558 11398 13568 11450
rect 13568 11398 13614 11450
rect 13318 11396 13374 11398
rect 13398 11396 13454 11398
rect 13478 11396 13534 11398
rect 13558 11396 13614 11398
rect 13318 10362 13374 10364
rect 13398 10362 13454 10364
rect 13478 10362 13534 10364
rect 13558 10362 13614 10364
rect 13318 10310 13364 10362
rect 13364 10310 13374 10362
rect 13398 10310 13428 10362
rect 13428 10310 13440 10362
rect 13440 10310 13454 10362
rect 13478 10310 13492 10362
rect 13492 10310 13504 10362
rect 13504 10310 13534 10362
rect 13558 10310 13568 10362
rect 13568 10310 13614 10362
rect 13318 10308 13374 10310
rect 13398 10308 13454 10310
rect 13478 10308 13534 10310
rect 13558 10308 13614 10310
rect 13542 10104 13598 10160
rect 13726 10104 13782 10160
rect 13318 9274 13374 9276
rect 13398 9274 13454 9276
rect 13478 9274 13534 9276
rect 13558 9274 13614 9276
rect 13318 9222 13364 9274
rect 13364 9222 13374 9274
rect 13398 9222 13428 9274
rect 13428 9222 13440 9274
rect 13440 9222 13454 9274
rect 13478 9222 13492 9274
rect 13492 9222 13504 9274
rect 13504 9222 13534 9274
rect 13558 9222 13568 9274
rect 13568 9222 13614 9274
rect 13318 9220 13374 9222
rect 13398 9220 13454 9222
rect 13478 9220 13534 9222
rect 13558 9220 13614 9222
rect 18263 15802 18319 15804
rect 18343 15802 18399 15804
rect 18423 15802 18479 15804
rect 18503 15802 18559 15804
rect 18263 15750 18309 15802
rect 18309 15750 18319 15802
rect 18343 15750 18373 15802
rect 18373 15750 18385 15802
rect 18385 15750 18399 15802
rect 18423 15750 18437 15802
rect 18437 15750 18449 15802
rect 18449 15750 18479 15802
rect 18503 15750 18513 15802
rect 18513 15750 18559 15802
rect 18263 15748 18319 15750
rect 18343 15748 18399 15750
rect 18423 15748 18479 15750
rect 18503 15748 18559 15750
rect 16762 15580 16764 15600
rect 16764 15580 16816 15600
rect 16816 15580 16818 15600
rect 16762 15544 16818 15580
rect 15290 15444 15292 15464
rect 15292 15444 15344 15464
rect 15344 15444 15346 15464
rect 15290 15408 15346 15444
rect 13318 8186 13374 8188
rect 13398 8186 13454 8188
rect 13478 8186 13534 8188
rect 13558 8186 13614 8188
rect 13318 8134 13364 8186
rect 13364 8134 13374 8186
rect 13398 8134 13428 8186
rect 13428 8134 13440 8186
rect 13440 8134 13454 8186
rect 13478 8134 13492 8186
rect 13492 8134 13504 8186
rect 13504 8134 13534 8186
rect 13558 8134 13568 8186
rect 13568 8134 13614 8186
rect 13318 8132 13374 8134
rect 13398 8132 13454 8134
rect 13478 8132 13534 8134
rect 13558 8132 13614 8134
rect 13318 7098 13374 7100
rect 13398 7098 13454 7100
rect 13478 7098 13534 7100
rect 13558 7098 13614 7100
rect 13318 7046 13364 7098
rect 13364 7046 13374 7098
rect 13398 7046 13428 7098
rect 13428 7046 13440 7098
rect 13440 7046 13454 7098
rect 13478 7046 13492 7098
rect 13492 7046 13504 7098
rect 13504 7046 13534 7098
rect 13558 7046 13568 7098
rect 13568 7046 13614 7098
rect 13318 7044 13374 7046
rect 13398 7044 13454 7046
rect 13478 7044 13534 7046
rect 13558 7044 13614 7046
rect 8373 4922 8429 4924
rect 8453 4922 8509 4924
rect 8533 4922 8589 4924
rect 8613 4922 8669 4924
rect 8373 4870 8419 4922
rect 8419 4870 8429 4922
rect 8453 4870 8483 4922
rect 8483 4870 8495 4922
rect 8495 4870 8509 4922
rect 8533 4870 8547 4922
rect 8547 4870 8559 4922
rect 8559 4870 8589 4922
rect 8613 4870 8623 4922
rect 8623 4870 8669 4922
rect 8373 4868 8429 4870
rect 8453 4868 8509 4870
rect 8533 4868 8589 4870
rect 8613 4868 8669 4870
rect 13318 6010 13374 6012
rect 13398 6010 13454 6012
rect 13478 6010 13534 6012
rect 13558 6010 13614 6012
rect 13318 5958 13364 6010
rect 13364 5958 13374 6010
rect 13398 5958 13428 6010
rect 13428 5958 13440 6010
rect 13440 5958 13454 6010
rect 13478 5958 13492 6010
rect 13492 5958 13504 6010
rect 13504 5958 13534 6010
rect 13558 5958 13568 6010
rect 13568 5958 13614 6010
rect 13318 5956 13374 5958
rect 13398 5956 13454 5958
rect 13478 5956 13534 5958
rect 13558 5956 13614 5958
rect 15790 15258 15846 15260
rect 15870 15258 15926 15260
rect 15950 15258 16006 15260
rect 16030 15258 16086 15260
rect 15790 15206 15836 15258
rect 15836 15206 15846 15258
rect 15870 15206 15900 15258
rect 15900 15206 15912 15258
rect 15912 15206 15926 15258
rect 15950 15206 15964 15258
rect 15964 15206 15976 15258
rect 15976 15206 16006 15258
rect 16030 15206 16040 15258
rect 16040 15206 16086 15258
rect 15790 15204 15846 15206
rect 15870 15204 15926 15206
rect 15950 15204 16006 15206
rect 16030 15204 16086 15206
rect 15790 14170 15846 14172
rect 15870 14170 15926 14172
rect 15950 14170 16006 14172
rect 16030 14170 16086 14172
rect 15790 14118 15836 14170
rect 15836 14118 15846 14170
rect 15870 14118 15900 14170
rect 15900 14118 15912 14170
rect 15912 14118 15926 14170
rect 15950 14118 15964 14170
rect 15964 14118 15976 14170
rect 15976 14118 16006 14170
rect 16030 14118 16040 14170
rect 16040 14118 16086 14170
rect 15790 14116 15846 14118
rect 15870 14116 15926 14118
rect 15950 14116 16006 14118
rect 16030 14116 16086 14118
rect 13318 4922 13374 4924
rect 13398 4922 13454 4924
rect 13478 4922 13534 4924
rect 13558 4922 13614 4924
rect 13318 4870 13364 4922
rect 13364 4870 13374 4922
rect 13398 4870 13428 4922
rect 13428 4870 13440 4922
rect 13440 4870 13454 4922
rect 13478 4870 13492 4922
rect 13492 4870 13504 4922
rect 13504 4870 13534 4922
rect 13558 4870 13568 4922
rect 13568 4870 13614 4922
rect 13318 4868 13374 4870
rect 13398 4868 13454 4870
rect 13478 4868 13534 4870
rect 13558 4868 13614 4870
rect 10845 4378 10901 4380
rect 10925 4378 10981 4380
rect 11005 4378 11061 4380
rect 11085 4378 11141 4380
rect 10845 4326 10891 4378
rect 10891 4326 10901 4378
rect 10925 4326 10955 4378
rect 10955 4326 10967 4378
rect 10967 4326 10981 4378
rect 11005 4326 11019 4378
rect 11019 4326 11031 4378
rect 11031 4326 11061 4378
rect 11085 4326 11095 4378
rect 11095 4326 11141 4378
rect 10845 4324 10901 4326
rect 10925 4324 10981 4326
rect 11005 4324 11061 4326
rect 11085 4324 11141 4326
rect 8373 3834 8429 3836
rect 8453 3834 8509 3836
rect 8533 3834 8589 3836
rect 8613 3834 8669 3836
rect 8373 3782 8419 3834
rect 8419 3782 8429 3834
rect 8453 3782 8483 3834
rect 8483 3782 8495 3834
rect 8495 3782 8509 3834
rect 8533 3782 8547 3834
rect 8547 3782 8559 3834
rect 8559 3782 8589 3834
rect 8613 3782 8623 3834
rect 8623 3782 8669 3834
rect 8373 3780 8429 3782
rect 8453 3780 8509 3782
rect 8533 3780 8589 3782
rect 8613 3780 8669 3782
rect 8373 2746 8429 2748
rect 8453 2746 8509 2748
rect 8533 2746 8589 2748
rect 8613 2746 8669 2748
rect 8373 2694 8419 2746
rect 8419 2694 8429 2746
rect 8453 2694 8483 2746
rect 8483 2694 8495 2746
rect 8495 2694 8509 2746
rect 8533 2694 8547 2746
rect 8547 2694 8559 2746
rect 8559 2694 8589 2746
rect 8613 2694 8623 2746
rect 8623 2694 8669 2746
rect 8373 2692 8429 2694
rect 8453 2692 8509 2694
rect 8533 2692 8589 2694
rect 8613 2692 8669 2694
rect 13318 3834 13374 3836
rect 13398 3834 13454 3836
rect 13478 3834 13534 3836
rect 13558 3834 13614 3836
rect 13318 3782 13364 3834
rect 13364 3782 13374 3834
rect 13398 3782 13428 3834
rect 13428 3782 13440 3834
rect 13440 3782 13454 3834
rect 13478 3782 13492 3834
rect 13492 3782 13504 3834
rect 13504 3782 13534 3834
rect 13558 3782 13568 3834
rect 13568 3782 13614 3834
rect 13318 3780 13374 3782
rect 13398 3780 13454 3782
rect 13478 3780 13534 3782
rect 13558 3780 13614 3782
rect 10506 3440 10562 3496
rect 10845 3290 10901 3292
rect 10925 3290 10981 3292
rect 11005 3290 11061 3292
rect 11085 3290 11141 3292
rect 10845 3238 10891 3290
rect 10891 3238 10901 3290
rect 10925 3238 10955 3290
rect 10955 3238 10967 3290
rect 10967 3238 10981 3290
rect 11005 3238 11019 3290
rect 11019 3238 11031 3290
rect 11031 3238 11061 3290
rect 11085 3238 11095 3290
rect 11095 3238 11141 3290
rect 10845 3236 10901 3238
rect 10925 3236 10981 3238
rect 11005 3236 11061 3238
rect 11085 3236 11141 3238
rect 15790 13082 15846 13084
rect 15870 13082 15926 13084
rect 15950 13082 16006 13084
rect 16030 13082 16086 13084
rect 15790 13030 15836 13082
rect 15836 13030 15846 13082
rect 15870 13030 15900 13082
rect 15900 13030 15912 13082
rect 15912 13030 15926 13082
rect 15950 13030 15964 13082
rect 15964 13030 15976 13082
rect 15976 13030 16006 13082
rect 16030 13030 16040 13082
rect 16040 13030 16086 13082
rect 15790 13028 15846 13030
rect 15870 13028 15926 13030
rect 15950 13028 16006 13030
rect 16030 13028 16086 13030
rect 17130 14900 17132 14920
rect 17132 14900 17184 14920
rect 17184 14900 17186 14920
rect 17130 14864 17186 14900
rect 15790 11994 15846 11996
rect 15870 11994 15926 11996
rect 15950 11994 16006 11996
rect 16030 11994 16086 11996
rect 15790 11942 15836 11994
rect 15836 11942 15846 11994
rect 15870 11942 15900 11994
rect 15900 11942 15912 11994
rect 15912 11942 15926 11994
rect 15950 11942 15964 11994
rect 15964 11942 15976 11994
rect 15976 11942 16006 11994
rect 16030 11942 16040 11994
rect 16040 11942 16086 11994
rect 15790 11940 15846 11942
rect 15870 11940 15926 11942
rect 15950 11940 16006 11942
rect 16030 11940 16086 11942
rect 15790 10906 15846 10908
rect 15870 10906 15926 10908
rect 15950 10906 16006 10908
rect 16030 10906 16086 10908
rect 15790 10854 15836 10906
rect 15836 10854 15846 10906
rect 15870 10854 15900 10906
rect 15900 10854 15912 10906
rect 15912 10854 15926 10906
rect 15950 10854 15964 10906
rect 15964 10854 15976 10906
rect 15976 10854 16006 10906
rect 16030 10854 16040 10906
rect 16040 10854 16086 10906
rect 15790 10852 15846 10854
rect 15870 10852 15926 10854
rect 15950 10852 16006 10854
rect 16030 10852 16086 10854
rect 15842 10104 15898 10160
rect 15790 9818 15846 9820
rect 15870 9818 15926 9820
rect 15950 9818 16006 9820
rect 16030 9818 16086 9820
rect 15790 9766 15836 9818
rect 15836 9766 15846 9818
rect 15870 9766 15900 9818
rect 15900 9766 15912 9818
rect 15912 9766 15926 9818
rect 15950 9766 15964 9818
rect 15964 9766 15976 9818
rect 15976 9766 16006 9818
rect 16030 9766 16040 9818
rect 16040 9766 16086 9818
rect 15790 9764 15846 9766
rect 15870 9764 15926 9766
rect 15950 9764 16006 9766
rect 16030 9764 16086 9766
rect 18263 14714 18319 14716
rect 18343 14714 18399 14716
rect 18423 14714 18479 14716
rect 18503 14714 18559 14716
rect 18263 14662 18309 14714
rect 18309 14662 18319 14714
rect 18343 14662 18373 14714
rect 18373 14662 18385 14714
rect 18385 14662 18399 14714
rect 18423 14662 18437 14714
rect 18437 14662 18449 14714
rect 18449 14662 18479 14714
rect 18503 14662 18513 14714
rect 18513 14662 18559 14714
rect 18263 14660 18319 14662
rect 18343 14660 18399 14662
rect 18423 14660 18479 14662
rect 18503 14660 18559 14662
rect 20735 15258 20791 15260
rect 20815 15258 20871 15260
rect 20895 15258 20951 15260
rect 20975 15258 21031 15260
rect 20735 15206 20781 15258
rect 20781 15206 20791 15258
rect 20815 15206 20845 15258
rect 20845 15206 20857 15258
rect 20857 15206 20871 15258
rect 20895 15206 20909 15258
rect 20909 15206 20921 15258
rect 20921 15206 20951 15258
rect 20975 15206 20985 15258
rect 20985 15206 21031 15258
rect 20735 15204 20791 15206
rect 20815 15204 20871 15206
rect 20895 15204 20951 15206
rect 20975 15204 21031 15206
rect 18263 13626 18319 13628
rect 18343 13626 18399 13628
rect 18423 13626 18479 13628
rect 18503 13626 18559 13628
rect 18263 13574 18309 13626
rect 18309 13574 18319 13626
rect 18343 13574 18373 13626
rect 18373 13574 18385 13626
rect 18385 13574 18399 13626
rect 18423 13574 18437 13626
rect 18437 13574 18449 13626
rect 18449 13574 18479 13626
rect 18503 13574 18513 13626
rect 18513 13574 18559 13626
rect 18263 13572 18319 13574
rect 18343 13572 18399 13574
rect 18423 13572 18479 13574
rect 18503 13572 18559 13574
rect 18263 12538 18319 12540
rect 18343 12538 18399 12540
rect 18423 12538 18479 12540
rect 18503 12538 18559 12540
rect 18263 12486 18309 12538
rect 18309 12486 18319 12538
rect 18343 12486 18373 12538
rect 18373 12486 18385 12538
rect 18385 12486 18399 12538
rect 18423 12486 18437 12538
rect 18437 12486 18449 12538
rect 18449 12486 18479 12538
rect 18503 12486 18513 12538
rect 18513 12486 18559 12538
rect 18263 12484 18319 12486
rect 18343 12484 18399 12486
rect 18423 12484 18479 12486
rect 18503 12484 18559 12486
rect 18263 11450 18319 11452
rect 18343 11450 18399 11452
rect 18423 11450 18479 11452
rect 18503 11450 18559 11452
rect 18263 11398 18309 11450
rect 18309 11398 18319 11450
rect 18343 11398 18373 11450
rect 18373 11398 18385 11450
rect 18385 11398 18399 11450
rect 18423 11398 18437 11450
rect 18437 11398 18449 11450
rect 18449 11398 18479 11450
rect 18503 11398 18513 11450
rect 18513 11398 18559 11450
rect 18263 11396 18319 11398
rect 18343 11396 18399 11398
rect 18423 11396 18479 11398
rect 18503 11396 18559 11398
rect 18263 10362 18319 10364
rect 18343 10362 18399 10364
rect 18423 10362 18479 10364
rect 18503 10362 18559 10364
rect 18263 10310 18309 10362
rect 18309 10310 18319 10362
rect 18343 10310 18373 10362
rect 18373 10310 18385 10362
rect 18385 10310 18399 10362
rect 18423 10310 18437 10362
rect 18437 10310 18449 10362
rect 18449 10310 18479 10362
rect 18503 10310 18513 10362
rect 18513 10310 18559 10362
rect 18263 10308 18319 10310
rect 18343 10308 18399 10310
rect 18423 10308 18479 10310
rect 18503 10308 18559 10310
rect 18263 9274 18319 9276
rect 18343 9274 18399 9276
rect 18423 9274 18479 9276
rect 18503 9274 18559 9276
rect 18263 9222 18309 9274
rect 18309 9222 18319 9274
rect 18343 9222 18373 9274
rect 18373 9222 18385 9274
rect 18385 9222 18399 9274
rect 18423 9222 18437 9274
rect 18437 9222 18449 9274
rect 18449 9222 18479 9274
rect 18503 9222 18513 9274
rect 18513 9222 18559 9274
rect 18263 9220 18319 9222
rect 18343 9220 18399 9222
rect 18423 9220 18479 9222
rect 18503 9220 18559 9222
rect 20735 14170 20791 14172
rect 20815 14170 20871 14172
rect 20895 14170 20951 14172
rect 20975 14170 21031 14172
rect 20735 14118 20781 14170
rect 20781 14118 20791 14170
rect 20815 14118 20845 14170
rect 20845 14118 20857 14170
rect 20857 14118 20871 14170
rect 20895 14118 20909 14170
rect 20909 14118 20921 14170
rect 20921 14118 20951 14170
rect 20975 14118 20985 14170
rect 20985 14118 21031 14170
rect 20735 14116 20791 14118
rect 20815 14116 20871 14118
rect 20895 14116 20951 14118
rect 20975 14116 21031 14118
rect 20735 13082 20791 13084
rect 20815 13082 20871 13084
rect 20895 13082 20951 13084
rect 20975 13082 21031 13084
rect 20735 13030 20781 13082
rect 20781 13030 20791 13082
rect 20815 13030 20845 13082
rect 20845 13030 20857 13082
rect 20857 13030 20871 13082
rect 20895 13030 20909 13082
rect 20909 13030 20921 13082
rect 20921 13030 20951 13082
rect 20975 13030 20985 13082
rect 20985 13030 21031 13082
rect 20735 13028 20791 13030
rect 20815 13028 20871 13030
rect 20895 13028 20951 13030
rect 20975 13028 21031 13030
rect 20735 11994 20791 11996
rect 20815 11994 20871 11996
rect 20895 11994 20951 11996
rect 20975 11994 21031 11996
rect 20735 11942 20781 11994
rect 20781 11942 20791 11994
rect 20815 11942 20845 11994
rect 20845 11942 20857 11994
rect 20857 11942 20871 11994
rect 20895 11942 20909 11994
rect 20909 11942 20921 11994
rect 20921 11942 20951 11994
rect 20975 11942 20985 11994
rect 20985 11942 21031 11994
rect 20735 11940 20791 11942
rect 20815 11940 20871 11942
rect 20895 11940 20951 11942
rect 20975 11940 21031 11942
rect 15790 8730 15846 8732
rect 15870 8730 15926 8732
rect 15950 8730 16006 8732
rect 16030 8730 16086 8732
rect 15790 8678 15836 8730
rect 15836 8678 15846 8730
rect 15870 8678 15900 8730
rect 15900 8678 15912 8730
rect 15912 8678 15926 8730
rect 15950 8678 15964 8730
rect 15964 8678 15976 8730
rect 15976 8678 16006 8730
rect 16030 8678 16040 8730
rect 16040 8678 16086 8730
rect 15790 8676 15846 8678
rect 15870 8676 15926 8678
rect 15950 8676 16006 8678
rect 16030 8676 16086 8678
rect 15790 7642 15846 7644
rect 15870 7642 15926 7644
rect 15950 7642 16006 7644
rect 16030 7642 16086 7644
rect 15790 7590 15836 7642
rect 15836 7590 15846 7642
rect 15870 7590 15900 7642
rect 15900 7590 15912 7642
rect 15912 7590 15926 7642
rect 15950 7590 15964 7642
rect 15964 7590 15976 7642
rect 15976 7590 16006 7642
rect 16030 7590 16040 7642
rect 16040 7590 16086 7642
rect 15790 7588 15846 7590
rect 15870 7588 15926 7590
rect 15950 7588 16006 7590
rect 16030 7588 16086 7590
rect 15790 6554 15846 6556
rect 15870 6554 15926 6556
rect 15950 6554 16006 6556
rect 16030 6554 16086 6556
rect 15790 6502 15836 6554
rect 15836 6502 15846 6554
rect 15870 6502 15900 6554
rect 15900 6502 15912 6554
rect 15912 6502 15926 6554
rect 15950 6502 15964 6554
rect 15964 6502 15976 6554
rect 15976 6502 16006 6554
rect 16030 6502 16040 6554
rect 16040 6502 16086 6554
rect 15790 6500 15846 6502
rect 15870 6500 15926 6502
rect 15950 6500 16006 6502
rect 16030 6500 16086 6502
rect 13318 2746 13374 2748
rect 13398 2746 13454 2748
rect 13478 2746 13534 2748
rect 13558 2746 13614 2748
rect 13318 2694 13364 2746
rect 13364 2694 13374 2746
rect 13398 2694 13428 2746
rect 13428 2694 13440 2746
rect 13440 2694 13454 2746
rect 13478 2694 13492 2746
rect 13492 2694 13504 2746
rect 13504 2694 13534 2746
rect 13558 2694 13568 2746
rect 13568 2694 13614 2746
rect 13318 2692 13374 2694
rect 13398 2692 13454 2694
rect 13478 2692 13534 2694
rect 13558 2692 13614 2694
rect 14554 3440 14610 3496
rect 15790 5466 15846 5468
rect 15870 5466 15926 5468
rect 15950 5466 16006 5468
rect 16030 5466 16086 5468
rect 15790 5414 15836 5466
rect 15836 5414 15846 5466
rect 15870 5414 15900 5466
rect 15900 5414 15912 5466
rect 15912 5414 15926 5466
rect 15950 5414 15964 5466
rect 15964 5414 15976 5466
rect 15976 5414 16006 5466
rect 16030 5414 16040 5466
rect 16040 5414 16086 5466
rect 15790 5412 15846 5414
rect 15870 5412 15926 5414
rect 15950 5412 16006 5414
rect 16030 5412 16086 5414
rect 18263 8186 18319 8188
rect 18343 8186 18399 8188
rect 18423 8186 18479 8188
rect 18503 8186 18559 8188
rect 18263 8134 18309 8186
rect 18309 8134 18319 8186
rect 18343 8134 18373 8186
rect 18373 8134 18385 8186
rect 18385 8134 18399 8186
rect 18423 8134 18437 8186
rect 18437 8134 18449 8186
rect 18449 8134 18479 8186
rect 18503 8134 18513 8186
rect 18513 8134 18559 8186
rect 18263 8132 18319 8134
rect 18343 8132 18399 8134
rect 18423 8132 18479 8134
rect 18503 8132 18559 8134
rect 18263 7098 18319 7100
rect 18343 7098 18399 7100
rect 18423 7098 18479 7100
rect 18503 7098 18559 7100
rect 18263 7046 18309 7098
rect 18309 7046 18319 7098
rect 18343 7046 18373 7098
rect 18373 7046 18385 7098
rect 18385 7046 18399 7098
rect 18423 7046 18437 7098
rect 18437 7046 18449 7098
rect 18449 7046 18479 7098
rect 18503 7046 18513 7098
rect 18513 7046 18559 7098
rect 18263 7044 18319 7046
rect 18343 7044 18399 7046
rect 18423 7044 18479 7046
rect 18503 7044 18559 7046
rect 15790 4378 15846 4380
rect 15870 4378 15926 4380
rect 15950 4378 16006 4380
rect 16030 4378 16086 4380
rect 15790 4326 15836 4378
rect 15836 4326 15846 4378
rect 15870 4326 15900 4378
rect 15900 4326 15912 4378
rect 15912 4326 15926 4378
rect 15950 4326 15964 4378
rect 15964 4326 15976 4378
rect 15976 4326 16006 4378
rect 16030 4326 16040 4378
rect 16040 4326 16086 4378
rect 15790 4324 15846 4326
rect 15870 4324 15926 4326
rect 15950 4324 16006 4326
rect 16030 4324 16086 4326
rect 18263 6010 18319 6012
rect 18343 6010 18399 6012
rect 18423 6010 18479 6012
rect 18503 6010 18559 6012
rect 18263 5958 18309 6010
rect 18309 5958 18319 6010
rect 18343 5958 18373 6010
rect 18373 5958 18385 6010
rect 18385 5958 18399 6010
rect 18423 5958 18437 6010
rect 18437 5958 18449 6010
rect 18449 5958 18479 6010
rect 18503 5958 18513 6010
rect 18513 5958 18559 6010
rect 18263 5956 18319 5958
rect 18343 5956 18399 5958
rect 18423 5956 18479 5958
rect 18503 5956 18559 5958
rect 18263 4922 18319 4924
rect 18343 4922 18399 4924
rect 18423 4922 18479 4924
rect 18503 4922 18559 4924
rect 18263 4870 18309 4922
rect 18309 4870 18319 4922
rect 18343 4870 18373 4922
rect 18373 4870 18385 4922
rect 18385 4870 18399 4922
rect 18423 4870 18437 4922
rect 18437 4870 18449 4922
rect 18449 4870 18479 4922
rect 18503 4870 18513 4922
rect 18513 4870 18559 4922
rect 18263 4868 18319 4870
rect 18343 4868 18399 4870
rect 18423 4868 18479 4870
rect 18503 4868 18559 4870
rect 18694 6296 18750 6352
rect 20735 10906 20791 10908
rect 20815 10906 20871 10908
rect 20895 10906 20951 10908
rect 20975 10906 21031 10908
rect 20735 10854 20781 10906
rect 20781 10854 20791 10906
rect 20815 10854 20845 10906
rect 20845 10854 20857 10906
rect 20857 10854 20871 10906
rect 20895 10854 20909 10906
rect 20909 10854 20921 10906
rect 20921 10854 20951 10906
rect 20975 10854 20985 10906
rect 20985 10854 21031 10906
rect 20735 10852 20791 10854
rect 20815 10852 20871 10854
rect 20895 10852 20951 10854
rect 20975 10852 21031 10854
rect 20735 9818 20791 9820
rect 20815 9818 20871 9820
rect 20895 9818 20951 9820
rect 20975 9818 21031 9820
rect 20735 9766 20781 9818
rect 20781 9766 20791 9818
rect 20815 9766 20845 9818
rect 20845 9766 20857 9818
rect 20857 9766 20871 9818
rect 20895 9766 20909 9818
rect 20909 9766 20921 9818
rect 20921 9766 20951 9818
rect 20975 9766 20985 9818
rect 20985 9766 21031 9818
rect 20735 9764 20791 9766
rect 20815 9764 20871 9766
rect 20895 9764 20951 9766
rect 20975 9764 21031 9766
rect 20735 8730 20791 8732
rect 20815 8730 20871 8732
rect 20895 8730 20951 8732
rect 20975 8730 21031 8732
rect 20735 8678 20781 8730
rect 20781 8678 20791 8730
rect 20815 8678 20845 8730
rect 20845 8678 20857 8730
rect 20857 8678 20871 8730
rect 20895 8678 20909 8730
rect 20909 8678 20921 8730
rect 20921 8678 20951 8730
rect 20975 8678 20985 8730
rect 20985 8678 21031 8730
rect 20735 8676 20791 8678
rect 20815 8676 20871 8678
rect 20895 8676 20951 8678
rect 20975 8676 21031 8678
rect 20735 7642 20791 7644
rect 20815 7642 20871 7644
rect 20895 7642 20951 7644
rect 20975 7642 21031 7644
rect 20735 7590 20781 7642
rect 20781 7590 20791 7642
rect 20815 7590 20845 7642
rect 20845 7590 20857 7642
rect 20857 7590 20871 7642
rect 20895 7590 20909 7642
rect 20909 7590 20921 7642
rect 20921 7590 20951 7642
rect 20975 7590 20985 7642
rect 20985 7590 21031 7642
rect 20735 7588 20791 7590
rect 20815 7588 20871 7590
rect 20895 7588 20951 7590
rect 20975 7588 21031 7590
rect 20735 6554 20791 6556
rect 20815 6554 20871 6556
rect 20895 6554 20951 6556
rect 20975 6554 21031 6556
rect 20735 6502 20781 6554
rect 20781 6502 20791 6554
rect 20815 6502 20845 6554
rect 20845 6502 20857 6554
rect 20857 6502 20871 6554
rect 20895 6502 20909 6554
rect 20909 6502 20921 6554
rect 20921 6502 20951 6554
rect 20975 6502 20985 6554
rect 20985 6502 21031 6554
rect 20735 6500 20791 6502
rect 20815 6500 20871 6502
rect 20895 6500 20951 6502
rect 20975 6500 21031 6502
rect 19614 6160 19670 6216
rect 20735 5466 20791 5468
rect 20815 5466 20871 5468
rect 20895 5466 20951 5468
rect 20975 5466 21031 5468
rect 20735 5414 20781 5466
rect 20781 5414 20791 5466
rect 20815 5414 20845 5466
rect 20845 5414 20857 5466
rect 20857 5414 20871 5466
rect 20895 5414 20909 5466
rect 20909 5414 20921 5466
rect 20921 5414 20951 5466
rect 20975 5414 20985 5466
rect 20985 5414 21031 5466
rect 20735 5412 20791 5414
rect 20815 5412 20871 5414
rect 20895 5412 20951 5414
rect 20975 5412 21031 5414
rect 20735 4378 20791 4380
rect 20815 4378 20871 4380
rect 20895 4378 20951 4380
rect 20975 4378 21031 4380
rect 20735 4326 20781 4378
rect 20781 4326 20791 4378
rect 20815 4326 20845 4378
rect 20845 4326 20857 4378
rect 20857 4326 20871 4378
rect 20895 4326 20909 4378
rect 20909 4326 20921 4378
rect 20921 4326 20951 4378
rect 20975 4326 20985 4378
rect 20985 4326 21031 4378
rect 20735 4324 20791 4326
rect 20815 4324 20871 4326
rect 20895 4324 20951 4326
rect 20975 4324 21031 4326
rect 18263 3834 18319 3836
rect 18343 3834 18399 3836
rect 18423 3834 18479 3836
rect 18503 3834 18559 3836
rect 18263 3782 18309 3834
rect 18309 3782 18319 3834
rect 18343 3782 18373 3834
rect 18373 3782 18385 3834
rect 18385 3782 18399 3834
rect 18423 3782 18437 3834
rect 18437 3782 18449 3834
rect 18449 3782 18479 3834
rect 18503 3782 18513 3834
rect 18513 3782 18559 3834
rect 18263 3780 18319 3782
rect 18343 3780 18399 3782
rect 18423 3780 18479 3782
rect 18503 3780 18559 3782
rect 15790 3290 15846 3292
rect 15870 3290 15926 3292
rect 15950 3290 16006 3292
rect 16030 3290 16086 3292
rect 15790 3238 15836 3290
rect 15836 3238 15846 3290
rect 15870 3238 15900 3290
rect 15900 3238 15912 3290
rect 15912 3238 15926 3290
rect 15950 3238 15964 3290
rect 15964 3238 15976 3290
rect 15976 3238 16006 3290
rect 16030 3238 16040 3290
rect 16040 3238 16086 3290
rect 15790 3236 15846 3238
rect 15870 3236 15926 3238
rect 15950 3236 16006 3238
rect 16030 3236 16086 3238
rect 20735 3290 20791 3292
rect 20815 3290 20871 3292
rect 20895 3290 20951 3292
rect 20975 3290 21031 3292
rect 20735 3238 20781 3290
rect 20781 3238 20791 3290
rect 20815 3238 20845 3290
rect 20845 3238 20857 3290
rect 20857 3238 20871 3290
rect 20895 3238 20909 3290
rect 20909 3238 20921 3290
rect 20921 3238 20951 3290
rect 20975 3238 20985 3290
rect 20985 3238 21031 3290
rect 20735 3236 20791 3238
rect 20815 3236 20871 3238
rect 20895 3236 20951 3238
rect 20975 3236 21031 3238
rect 18263 2746 18319 2748
rect 18343 2746 18399 2748
rect 18423 2746 18479 2748
rect 18503 2746 18559 2748
rect 18263 2694 18309 2746
rect 18309 2694 18319 2746
rect 18343 2694 18373 2746
rect 18373 2694 18385 2746
rect 18385 2694 18399 2746
rect 18423 2694 18437 2746
rect 18437 2694 18449 2746
rect 18449 2694 18479 2746
rect 18503 2694 18513 2746
rect 18513 2694 18559 2746
rect 18263 2692 18319 2694
rect 18343 2692 18399 2694
rect 18423 2692 18479 2694
rect 18503 2692 18559 2694
rect 5900 2202 5956 2204
rect 5980 2202 6036 2204
rect 6060 2202 6116 2204
rect 6140 2202 6196 2204
rect 5900 2150 5946 2202
rect 5946 2150 5956 2202
rect 5980 2150 6010 2202
rect 6010 2150 6022 2202
rect 6022 2150 6036 2202
rect 6060 2150 6074 2202
rect 6074 2150 6086 2202
rect 6086 2150 6116 2202
rect 6140 2150 6150 2202
rect 6150 2150 6196 2202
rect 5900 2148 5956 2150
rect 5980 2148 6036 2150
rect 6060 2148 6116 2150
rect 6140 2148 6196 2150
rect 10845 2202 10901 2204
rect 10925 2202 10981 2204
rect 11005 2202 11061 2204
rect 11085 2202 11141 2204
rect 10845 2150 10891 2202
rect 10891 2150 10901 2202
rect 10925 2150 10955 2202
rect 10955 2150 10967 2202
rect 10967 2150 10981 2202
rect 11005 2150 11019 2202
rect 11019 2150 11031 2202
rect 11031 2150 11061 2202
rect 11085 2150 11095 2202
rect 11095 2150 11141 2202
rect 10845 2148 10901 2150
rect 10925 2148 10981 2150
rect 11005 2148 11061 2150
rect 11085 2148 11141 2150
rect 15790 2202 15846 2204
rect 15870 2202 15926 2204
rect 15950 2202 16006 2204
rect 16030 2202 16086 2204
rect 15790 2150 15836 2202
rect 15836 2150 15846 2202
rect 15870 2150 15900 2202
rect 15900 2150 15912 2202
rect 15912 2150 15926 2202
rect 15950 2150 15964 2202
rect 15964 2150 15976 2202
rect 15976 2150 16006 2202
rect 16030 2150 16040 2202
rect 16040 2150 16086 2202
rect 15790 2148 15846 2150
rect 15870 2148 15926 2150
rect 15950 2148 16006 2150
rect 16030 2148 16086 2150
rect 20735 2202 20791 2204
rect 20815 2202 20871 2204
rect 20895 2202 20951 2204
rect 20975 2202 21031 2204
rect 20735 2150 20781 2202
rect 20781 2150 20791 2202
rect 20815 2150 20845 2202
rect 20845 2150 20857 2202
rect 20857 2150 20871 2202
rect 20895 2150 20909 2202
rect 20909 2150 20921 2202
rect 20921 2150 20951 2202
rect 20975 2150 20985 2202
rect 20985 2150 21031 2202
rect 20735 2148 20791 2150
rect 20815 2148 20871 2150
rect 20895 2148 20951 2150
rect 20975 2148 21031 2150
<< metal3 >>
rect 5890 19616 6206 19617
rect 5890 19552 5896 19616
rect 5960 19552 5976 19616
rect 6040 19552 6056 19616
rect 6120 19552 6136 19616
rect 6200 19552 6206 19616
rect 5890 19551 6206 19552
rect 10835 19616 11151 19617
rect 10835 19552 10841 19616
rect 10905 19552 10921 19616
rect 10985 19552 11001 19616
rect 11065 19552 11081 19616
rect 11145 19552 11151 19616
rect 10835 19551 11151 19552
rect 15780 19616 16096 19617
rect 15780 19552 15786 19616
rect 15850 19552 15866 19616
rect 15930 19552 15946 19616
rect 16010 19552 16026 19616
rect 16090 19552 16096 19616
rect 15780 19551 16096 19552
rect 20725 19616 21041 19617
rect 20725 19552 20731 19616
rect 20795 19552 20811 19616
rect 20875 19552 20891 19616
rect 20955 19552 20971 19616
rect 21035 19552 21041 19616
rect 20725 19551 21041 19552
rect 3418 19072 3734 19073
rect 3418 19008 3424 19072
rect 3488 19008 3504 19072
rect 3568 19008 3584 19072
rect 3648 19008 3664 19072
rect 3728 19008 3734 19072
rect 3418 19007 3734 19008
rect 8363 19072 8679 19073
rect 8363 19008 8369 19072
rect 8433 19008 8449 19072
rect 8513 19008 8529 19072
rect 8593 19008 8609 19072
rect 8673 19008 8679 19072
rect 8363 19007 8679 19008
rect 13308 19072 13624 19073
rect 13308 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13554 19072
rect 13618 19008 13624 19072
rect 13308 19007 13624 19008
rect 18253 19072 18569 19073
rect 18253 19008 18259 19072
rect 18323 19008 18339 19072
rect 18403 19008 18419 19072
rect 18483 19008 18499 19072
rect 18563 19008 18569 19072
rect 18253 19007 18569 19008
rect 5890 18528 6206 18529
rect 5890 18464 5896 18528
rect 5960 18464 5976 18528
rect 6040 18464 6056 18528
rect 6120 18464 6136 18528
rect 6200 18464 6206 18528
rect 5890 18463 6206 18464
rect 10835 18528 11151 18529
rect 10835 18464 10841 18528
rect 10905 18464 10921 18528
rect 10985 18464 11001 18528
rect 11065 18464 11081 18528
rect 11145 18464 11151 18528
rect 10835 18463 11151 18464
rect 15780 18528 16096 18529
rect 15780 18464 15786 18528
rect 15850 18464 15866 18528
rect 15930 18464 15946 18528
rect 16010 18464 16026 18528
rect 16090 18464 16096 18528
rect 15780 18463 16096 18464
rect 20725 18528 21041 18529
rect 20725 18464 20731 18528
rect 20795 18464 20811 18528
rect 20875 18464 20891 18528
rect 20955 18464 20971 18528
rect 21035 18464 21041 18528
rect 20725 18463 21041 18464
rect 0 18322 800 18352
rect 933 18322 999 18325
rect 0 18320 999 18322
rect 0 18264 938 18320
rect 994 18264 999 18320
rect 0 18262 999 18264
rect 0 18232 800 18262
rect 933 18259 999 18262
rect 3418 17984 3734 17985
rect 3418 17920 3424 17984
rect 3488 17920 3504 17984
rect 3568 17920 3584 17984
rect 3648 17920 3664 17984
rect 3728 17920 3734 17984
rect 3418 17919 3734 17920
rect 8363 17984 8679 17985
rect 8363 17920 8369 17984
rect 8433 17920 8449 17984
rect 8513 17920 8529 17984
rect 8593 17920 8609 17984
rect 8673 17920 8679 17984
rect 8363 17919 8679 17920
rect 13308 17984 13624 17985
rect 13308 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13554 17984
rect 13618 17920 13624 17984
rect 13308 17919 13624 17920
rect 18253 17984 18569 17985
rect 18253 17920 18259 17984
rect 18323 17920 18339 17984
rect 18403 17920 18419 17984
rect 18483 17920 18499 17984
rect 18563 17920 18569 17984
rect 18253 17919 18569 17920
rect 5890 17440 6206 17441
rect 5890 17376 5896 17440
rect 5960 17376 5976 17440
rect 6040 17376 6056 17440
rect 6120 17376 6136 17440
rect 6200 17376 6206 17440
rect 5890 17375 6206 17376
rect 10835 17440 11151 17441
rect 10835 17376 10841 17440
rect 10905 17376 10921 17440
rect 10985 17376 11001 17440
rect 11065 17376 11081 17440
rect 11145 17376 11151 17440
rect 10835 17375 11151 17376
rect 15780 17440 16096 17441
rect 15780 17376 15786 17440
rect 15850 17376 15866 17440
rect 15930 17376 15946 17440
rect 16010 17376 16026 17440
rect 16090 17376 16096 17440
rect 15780 17375 16096 17376
rect 20725 17440 21041 17441
rect 20725 17376 20731 17440
rect 20795 17376 20811 17440
rect 20875 17376 20891 17440
rect 20955 17376 20971 17440
rect 21035 17376 21041 17440
rect 20725 17375 21041 17376
rect 3418 16896 3734 16897
rect 3418 16832 3424 16896
rect 3488 16832 3504 16896
rect 3568 16832 3584 16896
rect 3648 16832 3664 16896
rect 3728 16832 3734 16896
rect 3418 16831 3734 16832
rect 8363 16896 8679 16897
rect 8363 16832 8369 16896
rect 8433 16832 8449 16896
rect 8513 16832 8529 16896
rect 8593 16832 8609 16896
rect 8673 16832 8679 16896
rect 8363 16831 8679 16832
rect 13308 16896 13624 16897
rect 13308 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13554 16896
rect 13618 16832 13624 16896
rect 13308 16831 13624 16832
rect 18253 16896 18569 16897
rect 18253 16832 18259 16896
rect 18323 16832 18339 16896
rect 18403 16832 18419 16896
rect 18483 16832 18499 16896
rect 18563 16832 18569 16896
rect 18253 16831 18569 16832
rect 5890 16352 6206 16353
rect 5890 16288 5896 16352
rect 5960 16288 5976 16352
rect 6040 16288 6056 16352
rect 6120 16288 6136 16352
rect 6200 16288 6206 16352
rect 5890 16287 6206 16288
rect 10835 16352 11151 16353
rect 10835 16288 10841 16352
rect 10905 16288 10921 16352
rect 10985 16288 11001 16352
rect 11065 16288 11081 16352
rect 11145 16288 11151 16352
rect 10835 16287 11151 16288
rect 15780 16352 16096 16353
rect 15780 16288 15786 16352
rect 15850 16288 15866 16352
rect 15930 16288 15946 16352
rect 16010 16288 16026 16352
rect 16090 16288 16096 16352
rect 15780 16287 16096 16288
rect 20725 16352 21041 16353
rect 20725 16288 20731 16352
rect 20795 16288 20811 16352
rect 20875 16288 20891 16352
rect 20955 16288 20971 16352
rect 21035 16288 21041 16352
rect 20725 16287 21041 16288
rect 3418 15808 3734 15809
rect 3418 15744 3424 15808
rect 3488 15744 3504 15808
rect 3568 15744 3584 15808
rect 3648 15744 3664 15808
rect 3728 15744 3734 15808
rect 3418 15743 3734 15744
rect 8363 15808 8679 15809
rect 8363 15744 8369 15808
rect 8433 15744 8449 15808
rect 8513 15744 8529 15808
rect 8593 15744 8609 15808
rect 8673 15744 8679 15808
rect 8363 15743 8679 15744
rect 13308 15808 13624 15809
rect 13308 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13554 15808
rect 13618 15744 13624 15808
rect 13308 15743 13624 15744
rect 18253 15808 18569 15809
rect 18253 15744 18259 15808
rect 18323 15744 18339 15808
rect 18403 15744 18419 15808
rect 18483 15744 18499 15808
rect 18563 15744 18569 15808
rect 18253 15743 18569 15744
rect 12893 15602 12959 15605
rect 16757 15602 16823 15605
rect 12893 15600 16823 15602
rect 12893 15544 12898 15600
rect 12954 15544 16762 15600
rect 16818 15544 16823 15600
rect 12893 15542 16823 15544
rect 12893 15539 12959 15542
rect 16757 15539 16823 15542
rect 11329 15466 11395 15469
rect 15285 15466 15351 15469
rect 11329 15464 15351 15466
rect 11329 15408 11334 15464
rect 11390 15408 15290 15464
rect 15346 15408 15351 15464
rect 11329 15406 15351 15408
rect 11329 15403 11395 15406
rect 15285 15403 15351 15406
rect 5890 15264 6206 15265
rect 5890 15200 5896 15264
rect 5960 15200 5976 15264
rect 6040 15200 6056 15264
rect 6120 15200 6136 15264
rect 6200 15200 6206 15264
rect 5890 15199 6206 15200
rect 10835 15264 11151 15265
rect 10835 15200 10841 15264
rect 10905 15200 10921 15264
rect 10985 15200 11001 15264
rect 11065 15200 11081 15264
rect 11145 15200 11151 15264
rect 10835 15199 11151 15200
rect 15780 15264 16096 15265
rect 15780 15200 15786 15264
rect 15850 15200 15866 15264
rect 15930 15200 15946 15264
rect 16010 15200 16026 15264
rect 16090 15200 16096 15264
rect 15780 15199 16096 15200
rect 20725 15264 21041 15265
rect 20725 15200 20731 15264
rect 20795 15200 20811 15264
rect 20875 15200 20891 15264
rect 20955 15200 20971 15264
rect 21035 15200 21041 15264
rect 20725 15199 21041 15200
rect 13813 14922 13879 14925
rect 17125 14922 17191 14925
rect 13813 14920 17191 14922
rect 13813 14864 13818 14920
rect 13874 14864 17130 14920
rect 17186 14864 17191 14920
rect 13813 14862 17191 14864
rect 13813 14859 13879 14862
rect 17125 14859 17191 14862
rect 3418 14720 3734 14721
rect 3418 14656 3424 14720
rect 3488 14656 3504 14720
rect 3568 14656 3584 14720
rect 3648 14656 3664 14720
rect 3728 14656 3734 14720
rect 3418 14655 3734 14656
rect 8363 14720 8679 14721
rect 8363 14656 8369 14720
rect 8433 14656 8449 14720
rect 8513 14656 8529 14720
rect 8593 14656 8609 14720
rect 8673 14656 8679 14720
rect 8363 14655 8679 14656
rect 13308 14720 13624 14721
rect 13308 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13554 14720
rect 13618 14656 13624 14720
rect 13308 14655 13624 14656
rect 18253 14720 18569 14721
rect 18253 14656 18259 14720
rect 18323 14656 18339 14720
rect 18403 14656 18419 14720
rect 18483 14656 18499 14720
rect 18563 14656 18569 14720
rect 18253 14655 18569 14656
rect 12433 14378 12499 14381
rect 13353 14378 13419 14381
rect 12433 14376 13419 14378
rect 12433 14320 12438 14376
rect 12494 14320 13358 14376
rect 13414 14320 13419 14376
rect 12433 14318 13419 14320
rect 12433 14315 12499 14318
rect 13353 14315 13419 14318
rect 5890 14176 6206 14177
rect 5890 14112 5896 14176
rect 5960 14112 5976 14176
rect 6040 14112 6056 14176
rect 6120 14112 6136 14176
rect 6200 14112 6206 14176
rect 5890 14111 6206 14112
rect 10835 14176 11151 14177
rect 10835 14112 10841 14176
rect 10905 14112 10921 14176
rect 10985 14112 11001 14176
rect 11065 14112 11081 14176
rect 11145 14112 11151 14176
rect 10835 14111 11151 14112
rect 15780 14176 16096 14177
rect 15780 14112 15786 14176
rect 15850 14112 15866 14176
rect 15930 14112 15946 14176
rect 16010 14112 16026 14176
rect 16090 14112 16096 14176
rect 15780 14111 16096 14112
rect 20725 14176 21041 14177
rect 20725 14112 20731 14176
rect 20795 14112 20811 14176
rect 20875 14112 20891 14176
rect 20955 14112 20971 14176
rect 21035 14112 21041 14176
rect 20725 14111 21041 14112
rect 3418 13632 3734 13633
rect 3418 13568 3424 13632
rect 3488 13568 3504 13632
rect 3568 13568 3584 13632
rect 3648 13568 3664 13632
rect 3728 13568 3734 13632
rect 3418 13567 3734 13568
rect 8363 13632 8679 13633
rect 8363 13568 8369 13632
rect 8433 13568 8449 13632
rect 8513 13568 8529 13632
rect 8593 13568 8609 13632
rect 8673 13568 8679 13632
rect 8363 13567 8679 13568
rect 13308 13632 13624 13633
rect 13308 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13554 13632
rect 13618 13568 13624 13632
rect 13308 13567 13624 13568
rect 18253 13632 18569 13633
rect 18253 13568 18259 13632
rect 18323 13568 18339 13632
rect 18403 13568 18419 13632
rect 18483 13568 18499 13632
rect 18563 13568 18569 13632
rect 18253 13567 18569 13568
rect 5890 13088 6206 13089
rect 5890 13024 5896 13088
rect 5960 13024 5976 13088
rect 6040 13024 6056 13088
rect 6120 13024 6136 13088
rect 6200 13024 6206 13088
rect 5890 13023 6206 13024
rect 10835 13088 11151 13089
rect 10835 13024 10841 13088
rect 10905 13024 10921 13088
rect 10985 13024 11001 13088
rect 11065 13024 11081 13088
rect 11145 13024 11151 13088
rect 10835 13023 11151 13024
rect 15780 13088 16096 13089
rect 15780 13024 15786 13088
rect 15850 13024 15866 13088
rect 15930 13024 15946 13088
rect 16010 13024 16026 13088
rect 16090 13024 16096 13088
rect 15780 13023 16096 13024
rect 20725 13088 21041 13089
rect 20725 13024 20731 13088
rect 20795 13024 20811 13088
rect 20875 13024 20891 13088
rect 20955 13024 20971 13088
rect 21035 13024 21041 13088
rect 20725 13023 21041 13024
rect 3418 12544 3734 12545
rect 3418 12480 3424 12544
rect 3488 12480 3504 12544
rect 3568 12480 3584 12544
rect 3648 12480 3664 12544
rect 3728 12480 3734 12544
rect 3418 12479 3734 12480
rect 8363 12544 8679 12545
rect 8363 12480 8369 12544
rect 8433 12480 8449 12544
rect 8513 12480 8529 12544
rect 8593 12480 8609 12544
rect 8673 12480 8679 12544
rect 8363 12479 8679 12480
rect 13308 12544 13624 12545
rect 13308 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13554 12544
rect 13618 12480 13624 12544
rect 13308 12479 13624 12480
rect 18253 12544 18569 12545
rect 18253 12480 18259 12544
rect 18323 12480 18339 12544
rect 18403 12480 18419 12544
rect 18483 12480 18499 12544
rect 18563 12480 18569 12544
rect 18253 12479 18569 12480
rect 5890 12000 6206 12001
rect 5890 11936 5896 12000
rect 5960 11936 5976 12000
rect 6040 11936 6056 12000
rect 6120 11936 6136 12000
rect 6200 11936 6206 12000
rect 5890 11935 6206 11936
rect 10835 12000 11151 12001
rect 10835 11936 10841 12000
rect 10905 11936 10921 12000
rect 10985 11936 11001 12000
rect 11065 11936 11081 12000
rect 11145 11936 11151 12000
rect 10835 11935 11151 11936
rect 15780 12000 16096 12001
rect 15780 11936 15786 12000
rect 15850 11936 15866 12000
rect 15930 11936 15946 12000
rect 16010 11936 16026 12000
rect 16090 11936 16096 12000
rect 15780 11935 16096 11936
rect 20725 12000 21041 12001
rect 20725 11936 20731 12000
rect 20795 11936 20811 12000
rect 20875 11936 20891 12000
rect 20955 11936 20971 12000
rect 21035 11936 21041 12000
rect 20725 11935 21041 11936
rect 3418 11456 3734 11457
rect 3418 11392 3424 11456
rect 3488 11392 3504 11456
rect 3568 11392 3584 11456
rect 3648 11392 3664 11456
rect 3728 11392 3734 11456
rect 3418 11391 3734 11392
rect 8363 11456 8679 11457
rect 8363 11392 8369 11456
rect 8433 11392 8449 11456
rect 8513 11392 8529 11456
rect 8593 11392 8609 11456
rect 8673 11392 8679 11456
rect 8363 11391 8679 11392
rect 13308 11456 13624 11457
rect 13308 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13554 11456
rect 13618 11392 13624 11456
rect 13308 11391 13624 11392
rect 18253 11456 18569 11457
rect 18253 11392 18259 11456
rect 18323 11392 18339 11456
rect 18403 11392 18419 11456
rect 18483 11392 18499 11456
rect 18563 11392 18569 11456
rect 18253 11391 18569 11392
rect 0 10978 800 11008
rect 933 10978 999 10981
rect 0 10976 999 10978
rect 0 10920 938 10976
rect 994 10920 999 10976
rect 0 10918 999 10920
rect 0 10888 800 10918
rect 933 10915 999 10918
rect 5890 10912 6206 10913
rect 5890 10848 5896 10912
rect 5960 10848 5976 10912
rect 6040 10848 6056 10912
rect 6120 10848 6136 10912
rect 6200 10848 6206 10912
rect 5890 10847 6206 10848
rect 10835 10912 11151 10913
rect 10835 10848 10841 10912
rect 10905 10848 10921 10912
rect 10985 10848 11001 10912
rect 11065 10848 11081 10912
rect 11145 10848 11151 10912
rect 10835 10847 11151 10848
rect 15780 10912 16096 10913
rect 15780 10848 15786 10912
rect 15850 10848 15866 10912
rect 15930 10848 15946 10912
rect 16010 10848 16026 10912
rect 16090 10848 16096 10912
rect 15780 10847 16096 10848
rect 20725 10912 21041 10913
rect 20725 10848 20731 10912
rect 20795 10848 20811 10912
rect 20875 10848 20891 10912
rect 20955 10848 20971 10912
rect 21035 10848 21041 10912
rect 20725 10847 21041 10848
rect 3418 10368 3734 10369
rect 3418 10304 3424 10368
rect 3488 10304 3504 10368
rect 3568 10304 3584 10368
rect 3648 10304 3664 10368
rect 3728 10304 3734 10368
rect 3418 10303 3734 10304
rect 8363 10368 8679 10369
rect 8363 10304 8369 10368
rect 8433 10304 8449 10368
rect 8513 10304 8529 10368
rect 8593 10304 8609 10368
rect 8673 10304 8679 10368
rect 8363 10303 8679 10304
rect 13308 10368 13624 10369
rect 13308 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13554 10368
rect 13618 10304 13624 10368
rect 13308 10303 13624 10304
rect 18253 10368 18569 10369
rect 18253 10304 18259 10368
rect 18323 10304 18339 10368
rect 18403 10304 18419 10368
rect 18483 10304 18499 10368
rect 18563 10304 18569 10368
rect 18253 10303 18569 10304
rect 13537 10162 13603 10165
rect 13721 10162 13787 10165
rect 15837 10162 15903 10165
rect 13537 10160 15903 10162
rect 13537 10104 13542 10160
rect 13598 10104 13726 10160
rect 13782 10104 15842 10160
rect 15898 10104 15903 10160
rect 13537 10102 15903 10104
rect 13537 10099 13603 10102
rect 13721 10099 13787 10102
rect 15837 10099 15903 10102
rect 5890 9824 6206 9825
rect 5890 9760 5896 9824
rect 5960 9760 5976 9824
rect 6040 9760 6056 9824
rect 6120 9760 6136 9824
rect 6200 9760 6206 9824
rect 5890 9759 6206 9760
rect 10835 9824 11151 9825
rect 10835 9760 10841 9824
rect 10905 9760 10921 9824
rect 10985 9760 11001 9824
rect 11065 9760 11081 9824
rect 11145 9760 11151 9824
rect 10835 9759 11151 9760
rect 15780 9824 16096 9825
rect 15780 9760 15786 9824
rect 15850 9760 15866 9824
rect 15930 9760 15946 9824
rect 16010 9760 16026 9824
rect 16090 9760 16096 9824
rect 15780 9759 16096 9760
rect 20725 9824 21041 9825
rect 20725 9760 20731 9824
rect 20795 9760 20811 9824
rect 20875 9760 20891 9824
rect 20955 9760 20971 9824
rect 21035 9760 21041 9824
rect 20725 9759 21041 9760
rect 3418 9280 3734 9281
rect 3418 9216 3424 9280
rect 3488 9216 3504 9280
rect 3568 9216 3584 9280
rect 3648 9216 3664 9280
rect 3728 9216 3734 9280
rect 3418 9215 3734 9216
rect 8363 9280 8679 9281
rect 8363 9216 8369 9280
rect 8433 9216 8449 9280
rect 8513 9216 8529 9280
rect 8593 9216 8609 9280
rect 8673 9216 8679 9280
rect 8363 9215 8679 9216
rect 13308 9280 13624 9281
rect 13308 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13554 9280
rect 13618 9216 13624 9280
rect 13308 9215 13624 9216
rect 18253 9280 18569 9281
rect 18253 9216 18259 9280
rect 18323 9216 18339 9280
rect 18403 9216 18419 9280
rect 18483 9216 18499 9280
rect 18563 9216 18569 9280
rect 18253 9215 18569 9216
rect 5890 8736 6206 8737
rect 5890 8672 5896 8736
rect 5960 8672 5976 8736
rect 6040 8672 6056 8736
rect 6120 8672 6136 8736
rect 6200 8672 6206 8736
rect 5890 8671 6206 8672
rect 10835 8736 11151 8737
rect 10835 8672 10841 8736
rect 10905 8672 10921 8736
rect 10985 8672 11001 8736
rect 11065 8672 11081 8736
rect 11145 8672 11151 8736
rect 10835 8671 11151 8672
rect 15780 8736 16096 8737
rect 15780 8672 15786 8736
rect 15850 8672 15866 8736
rect 15930 8672 15946 8736
rect 16010 8672 16026 8736
rect 16090 8672 16096 8736
rect 15780 8671 16096 8672
rect 20725 8736 21041 8737
rect 20725 8672 20731 8736
rect 20795 8672 20811 8736
rect 20875 8672 20891 8736
rect 20955 8672 20971 8736
rect 21035 8672 21041 8736
rect 20725 8671 21041 8672
rect 3418 8192 3734 8193
rect 3418 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3584 8192
rect 3648 8128 3664 8192
rect 3728 8128 3734 8192
rect 3418 8127 3734 8128
rect 8363 8192 8679 8193
rect 8363 8128 8369 8192
rect 8433 8128 8449 8192
rect 8513 8128 8529 8192
rect 8593 8128 8609 8192
rect 8673 8128 8679 8192
rect 8363 8127 8679 8128
rect 13308 8192 13624 8193
rect 13308 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13554 8192
rect 13618 8128 13624 8192
rect 13308 8127 13624 8128
rect 18253 8192 18569 8193
rect 18253 8128 18259 8192
rect 18323 8128 18339 8192
rect 18403 8128 18419 8192
rect 18483 8128 18499 8192
rect 18563 8128 18569 8192
rect 18253 8127 18569 8128
rect 5890 7648 6206 7649
rect 5890 7584 5896 7648
rect 5960 7584 5976 7648
rect 6040 7584 6056 7648
rect 6120 7584 6136 7648
rect 6200 7584 6206 7648
rect 5890 7583 6206 7584
rect 10835 7648 11151 7649
rect 10835 7584 10841 7648
rect 10905 7584 10921 7648
rect 10985 7584 11001 7648
rect 11065 7584 11081 7648
rect 11145 7584 11151 7648
rect 10835 7583 11151 7584
rect 15780 7648 16096 7649
rect 15780 7584 15786 7648
rect 15850 7584 15866 7648
rect 15930 7584 15946 7648
rect 16010 7584 16026 7648
rect 16090 7584 16096 7648
rect 15780 7583 16096 7584
rect 20725 7648 21041 7649
rect 20725 7584 20731 7648
rect 20795 7584 20811 7648
rect 20875 7584 20891 7648
rect 20955 7584 20971 7648
rect 21035 7584 21041 7648
rect 20725 7583 21041 7584
rect 3418 7104 3734 7105
rect 3418 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3584 7104
rect 3648 7040 3664 7104
rect 3728 7040 3734 7104
rect 3418 7039 3734 7040
rect 8363 7104 8679 7105
rect 8363 7040 8369 7104
rect 8433 7040 8449 7104
rect 8513 7040 8529 7104
rect 8593 7040 8609 7104
rect 8673 7040 8679 7104
rect 8363 7039 8679 7040
rect 13308 7104 13624 7105
rect 13308 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13554 7104
rect 13618 7040 13624 7104
rect 13308 7039 13624 7040
rect 18253 7104 18569 7105
rect 18253 7040 18259 7104
rect 18323 7040 18339 7104
rect 18403 7040 18419 7104
rect 18483 7040 18499 7104
rect 18563 7040 18569 7104
rect 18253 7039 18569 7040
rect 5890 6560 6206 6561
rect 5890 6496 5896 6560
rect 5960 6496 5976 6560
rect 6040 6496 6056 6560
rect 6120 6496 6136 6560
rect 6200 6496 6206 6560
rect 5890 6495 6206 6496
rect 10835 6560 11151 6561
rect 10835 6496 10841 6560
rect 10905 6496 10921 6560
rect 10985 6496 11001 6560
rect 11065 6496 11081 6560
rect 11145 6496 11151 6560
rect 10835 6495 11151 6496
rect 15780 6560 16096 6561
rect 15780 6496 15786 6560
rect 15850 6496 15866 6560
rect 15930 6496 15946 6560
rect 16010 6496 16026 6560
rect 16090 6496 16096 6560
rect 15780 6495 16096 6496
rect 20725 6560 21041 6561
rect 20725 6496 20731 6560
rect 20795 6496 20811 6560
rect 20875 6496 20891 6560
rect 20955 6496 20971 6560
rect 21035 6496 21041 6560
rect 20725 6495 21041 6496
rect 5441 6354 5507 6357
rect 18689 6354 18755 6357
rect 5441 6352 18755 6354
rect 5441 6296 5446 6352
rect 5502 6296 18694 6352
rect 18750 6296 18755 6352
rect 5441 6294 18755 6296
rect 5441 6291 5507 6294
rect 18689 6291 18755 6294
rect 2589 6218 2655 6221
rect 5901 6218 5967 6221
rect 19609 6218 19675 6221
rect 2589 6216 19675 6218
rect 2589 6160 2594 6216
rect 2650 6160 5906 6216
rect 5962 6160 19614 6216
rect 19670 6160 19675 6216
rect 2589 6158 19675 6160
rect 2589 6155 2655 6158
rect 5901 6155 5967 6158
rect 19609 6155 19675 6158
rect 3418 6016 3734 6017
rect 3418 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3584 6016
rect 3648 5952 3664 6016
rect 3728 5952 3734 6016
rect 3418 5951 3734 5952
rect 8363 6016 8679 6017
rect 8363 5952 8369 6016
rect 8433 5952 8449 6016
rect 8513 5952 8529 6016
rect 8593 5952 8609 6016
rect 8673 5952 8679 6016
rect 8363 5951 8679 5952
rect 13308 6016 13624 6017
rect 13308 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13554 6016
rect 13618 5952 13624 6016
rect 13308 5951 13624 5952
rect 18253 6016 18569 6017
rect 18253 5952 18259 6016
rect 18323 5952 18339 6016
rect 18403 5952 18419 6016
rect 18483 5952 18499 6016
rect 18563 5952 18569 6016
rect 18253 5951 18569 5952
rect 5890 5472 6206 5473
rect 5890 5408 5896 5472
rect 5960 5408 5976 5472
rect 6040 5408 6056 5472
rect 6120 5408 6136 5472
rect 6200 5408 6206 5472
rect 5890 5407 6206 5408
rect 10835 5472 11151 5473
rect 10835 5408 10841 5472
rect 10905 5408 10921 5472
rect 10985 5408 11001 5472
rect 11065 5408 11081 5472
rect 11145 5408 11151 5472
rect 10835 5407 11151 5408
rect 15780 5472 16096 5473
rect 15780 5408 15786 5472
rect 15850 5408 15866 5472
rect 15930 5408 15946 5472
rect 16010 5408 16026 5472
rect 16090 5408 16096 5472
rect 15780 5407 16096 5408
rect 20725 5472 21041 5473
rect 20725 5408 20731 5472
rect 20795 5408 20811 5472
rect 20875 5408 20891 5472
rect 20955 5408 20971 5472
rect 21035 5408 21041 5472
rect 20725 5407 21041 5408
rect 3418 4928 3734 4929
rect 3418 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3584 4928
rect 3648 4864 3664 4928
rect 3728 4864 3734 4928
rect 3418 4863 3734 4864
rect 8363 4928 8679 4929
rect 8363 4864 8369 4928
rect 8433 4864 8449 4928
rect 8513 4864 8529 4928
rect 8593 4864 8609 4928
rect 8673 4864 8679 4928
rect 8363 4863 8679 4864
rect 13308 4928 13624 4929
rect 13308 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13554 4928
rect 13618 4864 13624 4928
rect 13308 4863 13624 4864
rect 18253 4928 18569 4929
rect 18253 4864 18259 4928
rect 18323 4864 18339 4928
rect 18403 4864 18419 4928
rect 18483 4864 18499 4928
rect 18563 4864 18569 4928
rect 18253 4863 18569 4864
rect 5890 4384 6206 4385
rect 5890 4320 5896 4384
rect 5960 4320 5976 4384
rect 6040 4320 6056 4384
rect 6120 4320 6136 4384
rect 6200 4320 6206 4384
rect 5890 4319 6206 4320
rect 10835 4384 11151 4385
rect 10835 4320 10841 4384
rect 10905 4320 10921 4384
rect 10985 4320 11001 4384
rect 11065 4320 11081 4384
rect 11145 4320 11151 4384
rect 10835 4319 11151 4320
rect 15780 4384 16096 4385
rect 15780 4320 15786 4384
rect 15850 4320 15866 4384
rect 15930 4320 15946 4384
rect 16010 4320 16026 4384
rect 16090 4320 16096 4384
rect 15780 4319 16096 4320
rect 20725 4384 21041 4385
rect 20725 4320 20731 4384
rect 20795 4320 20811 4384
rect 20875 4320 20891 4384
rect 20955 4320 20971 4384
rect 21035 4320 21041 4384
rect 20725 4319 21041 4320
rect 3418 3840 3734 3841
rect 3418 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3584 3840
rect 3648 3776 3664 3840
rect 3728 3776 3734 3840
rect 3418 3775 3734 3776
rect 8363 3840 8679 3841
rect 8363 3776 8369 3840
rect 8433 3776 8449 3840
rect 8513 3776 8529 3840
rect 8593 3776 8609 3840
rect 8673 3776 8679 3840
rect 8363 3775 8679 3776
rect 13308 3840 13624 3841
rect 13308 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13554 3840
rect 13618 3776 13624 3840
rect 13308 3775 13624 3776
rect 18253 3840 18569 3841
rect 18253 3776 18259 3840
rect 18323 3776 18339 3840
rect 18403 3776 18419 3840
rect 18483 3776 18499 3840
rect 18563 3776 18569 3840
rect 18253 3775 18569 3776
rect 0 3634 800 3664
rect 3233 3634 3299 3637
rect 0 3632 3299 3634
rect 0 3576 3238 3632
rect 3294 3576 3299 3632
rect 0 3574 3299 3576
rect 0 3544 800 3574
rect 3233 3571 3299 3574
rect 10501 3498 10567 3501
rect 14549 3498 14615 3501
rect 10501 3496 14615 3498
rect 10501 3440 10506 3496
rect 10562 3440 14554 3496
rect 14610 3440 14615 3496
rect 10501 3438 14615 3440
rect 10501 3435 10567 3438
rect 14549 3435 14615 3438
rect 5890 3296 6206 3297
rect 5890 3232 5896 3296
rect 5960 3232 5976 3296
rect 6040 3232 6056 3296
rect 6120 3232 6136 3296
rect 6200 3232 6206 3296
rect 5890 3231 6206 3232
rect 10835 3296 11151 3297
rect 10835 3232 10841 3296
rect 10905 3232 10921 3296
rect 10985 3232 11001 3296
rect 11065 3232 11081 3296
rect 11145 3232 11151 3296
rect 10835 3231 11151 3232
rect 15780 3296 16096 3297
rect 15780 3232 15786 3296
rect 15850 3232 15866 3296
rect 15930 3232 15946 3296
rect 16010 3232 16026 3296
rect 16090 3232 16096 3296
rect 15780 3231 16096 3232
rect 20725 3296 21041 3297
rect 20725 3232 20731 3296
rect 20795 3232 20811 3296
rect 20875 3232 20891 3296
rect 20955 3232 20971 3296
rect 21035 3232 21041 3296
rect 20725 3231 21041 3232
rect 3418 2752 3734 2753
rect 3418 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3584 2752
rect 3648 2688 3664 2752
rect 3728 2688 3734 2752
rect 3418 2687 3734 2688
rect 8363 2752 8679 2753
rect 8363 2688 8369 2752
rect 8433 2688 8449 2752
rect 8513 2688 8529 2752
rect 8593 2688 8609 2752
rect 8673 2688 8679 2752
rect 8363 2687 8679 2688
rect 13308 2752 13624 2753
rect 13308 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13554 2752
rect 13618 2688 13624 2752
rect 13308 2687 13624 2688
rect 18253 2752 18569 2753
rect 18253 2688 18259 2752
rect 18323 2688 18339 2752
rect 18403 2688 18419 2752
rect 18483 2688 18499 2752
rect 18563 2688 18569 2752
rect 18253 2687 18569 2688
rect 5890 2208 6206 2209
rect 5890 2144 5896 2208
rect 5960 2144 5976 2208
rect 6040 2144 6056 2208
rect 6120 2144 6136 2208
rect 6200 2144 6206 2208
rect 5890 2143 6206 2144
rect 10835 2208 11151 2209
rect 10835 2144 10841 2208
rect 10905 2144 10921 2208
rect 10985 2144 11001 2208
rect 11065 2144 11081 2208
rect 11145 2144 11151 2208
rect 10835 2143 11151 2144
rect 15780 2208 16096 2209
rect 15780 2144 15786 2208
rect 15850 2144 15866 2208
rect 15930 2144 15946 2208
rect 16010 2144 16026 2208
rect 16090 2144 16096 2208
rect 15780 2143 16096 2144
rect 20725 2208 21041 2209
rect 20725 2144 20731 2208
rect 20795 2144 20811 2208
rect 20875 2144 20891 2208
rect 20955 2144 20971 2208
rect 21035 2144 21041 2208
rect 20725 2143 21041 2144
<< via3 >>
rect 5896 19612 5960 19616
rect 5896 19556 5900 19612
rect 5900 19556 5956 19612
rect 5956 19556 5960 19612
rect 5896 19552 5960 19556
rect 5976 19612 6040 19616
rect 5976 19556 5980 19612
rect 5980 19556 6036 19612
rect 6036 19556 6040 19612
rect 5976 19552 6040 19556
rect 6056 19612 6120 19616
rect 6056 19556 6060 19612
rect 6060 19556 6116 19612
rect 6116 19556 6120 19612
rect 6056 19552 6120 19556
rect 6136 19612 6200 19616
rect 6136 19556 6140 19612
rect 6140 19556 6196 19612
rect 6196 19556 6200 19612
rect 6136 19552 6200 19556
rect 10841 19612 10905 19616
rect 10841 19556 10845 19612
rect 10845 19556 10901 19612
rect 10901 19556 10905 19612
rect 10841 19552 10905 19556
rect 10921 19612 10985 19616
rect 10921 19556 10925 19612
rect 10925 19556 10981 19612
rect 10981 19556 10985 19612
rect 10921 19552 10985 19556
rect 11001 19612 11065 19616
rect 11001 19556 11005 19612
rect 11005 19556 11061 19612
rect 11061 19556 11065 19612
rect 11001 19552 11065 19556
rect 11081 19612 11145 19616
rect 11081 19556 11085 19612
rect 11085 19556 11141 19612
rect 11141 19556 11145 19612
rect 11081 19552 11145 19556
rect 15786 19612 15850 19616
rect 15786 19556 15790 19612
rect 15790 19556 15846 19612
rect 15846 19556 15850 19612
rect 15786 19552 15850 19556
rect 15866 19612 15930 19616
rect 15866 19556 15870 19612
rect 15870 19556 15926 19612
rect 15926 19556 15930 19612
rect 15866 19552 15930 19556
rect 15946 19612 16010 19616
rect 15946 19556 15950 19612
rect 15950 19556 16006 19612
rect 16006 19556 16010 19612
rect 15946 19552 16010 19556
rect 16026 19612 16090 19616
rect 16026 19556 16030 19612
rect 16030 19556 16086 19612
rect 16086 19556 16090 19612
rect 16026 19552 16090 19556
rect 20731 19612 20795 19616
rect 20731 19556 20735 19612
rect 20735 19556 20791 19612
rect 20791 19556 20795 19612
rect 20731 19552 20795 19556
rect 20811 19612 20875 19616
rect 20811 19556 20815 19612
rect 20815 19556 20871 19612
rect 20871 19556 20875 19612
rect 20811 19552 20875 19556
rect 20891 19612 20955 19616
rect 20891 19556 20895 19612
rect 20895 19556 20951 19612
rect 20951 19556 20955 19612
rect 20891 19552 20955 19556
rect 20971 19612 21035 19616
rect 20971 19556 20975 19612
rect 20975 19556 21031 19612
rect 21031 19556 21035 19612
rect 20971 19552 21035 19556
rect 3424 19068 3488 19072
rect 3424 19012 3428 19068
rect 3428 19012 3484 19068
rect 3484 19012 3488 19068
rect 3424 19008 3488 19012
rect 3504 19068 3568 19072
rect 3504 19012 3508 19068
rect 3508 19012 3564 19068
rect 3564 19012 3568 19068
rect 3504 19008 3568 19012
rect 3584 19068 3648 19072
rect 3584 19012 3588 19068
rect 3588 19012 3644 19068
rect 3644 19012 3648 19068
rect 3584 19008 3648 19012
rect 3664 19068 3728 19072
rect 3664 19012 3668 19068
rect 3668 19012 3724 19068
rect 3724 19012 3728 19068
rect 3664 19008 3728 19012
rect 8369 19068 8433 19072
rect 8369 19012 8373 19068
rect 8373 19012 8429 19068
rect 8429 19012 8433 19068
rect 8369 19008 8433 19012
rect 8449 19068 8513 19072
rect 8449 19012 8453 19068
rect 8453 19012 8509 19068
rect 8509 19012 8513 19068
rect 8449 19008 8513 19012
rect 8529 19068 8593 19072
rect 8529 19012 8533 19068
rect 8533 19012 8589 19068
rect 8589 19012 8593 19068
rect 8529 19008 8593 19012
rect 8609 19068 8673 19072
rect 8609 19012 8613 19068
rect 8613 19012 8669 19068
rect 8669 19012 8673 19068
rect 8609 19008 8673 19012
rect 13314 19068 13378 19072
rect 13314 19012 13318 19068
rect 13318 19012 13374 19068
rect 13374 19012 13378 19068
rect 13314 19008 13378 19012
rect 13394 19068 13458 19072
rect 13394 19012 13398 19068
rect 13398 19012 13454 19068
rect 13454 19012 13458 19068
rect 13394 19008 13458 19012
rect 13474 19068 13538 19072
rect 13474 19012 13478 19068
rect 13478 19012 13534 19068
rect 13534 19012 13538 19068
rect 13474 19008 13538 19012
rect 13554 19068 13618 19072
rect 13554 19012 13558 19068
rect 13558 19012 13614 19068
rect 13614 19012 13618 19068
rect 13554 19008 13618 19012
rect 18259 19068 18323 19072
rect 18259 19012 18263 19068
rect 18263 19012 18319 19068
rect 18319 19012 18323 19068
rect 18259 19008 18323 19012
rect 18339 19068 18403 19072
rect 18339 19012 18343 19068
rect 18343 19012 18399 19068
rect 18399 19012 18403 19068
rect 18339 19008 18403 19012
rect 18419 19068 18483 19072
rect 18419 19012 18423 19068
rect 18423 19012 18479 19068
rect 18479 19012 18483 19068
rect 18419 19008 18483 19012
rect 18499 19068 18563 19072
rect 18499 19012 18503 19068
rect 18503 19012 18559 19068
rect 18559 19012 18563 19068
rect 18499 19008 18563 19012
rect 5896 18524 5960 18528
rect 5896 18468 5900 18524
rect 5900 18468 5956 18524
rect 5956 18468 5960 18524
rect 5896 18464 5960 18468
rect 5976 18524 6040 18528
rect 5976 18468 5980 18524
rect 5980 18468 6036 18524
rect 6036 18468 6040 18524
rect 5976 18464 6040 18468
rect 6056 18524 6120 18528
rect 6056 18468 6060 18524
rect 6060 18468 6116 18524
rect 6116 18468 6120 18524
rect 6056 18464 6120 18468
rect 6136 18524 6200 18528
rect 6136 18468 6140 18524
rect 6140 18468 6196 18524
rect 6196 18468 6200 18524
rect 6136 18464 6200 18468
rect 10841 18524 10905 18528
rect 10841 18468 10845 18524
rect 10845 18468 10901 18524
rect 10901 18468 10905 18524
rect 10841 18464 10905 18468
rect 10921 18524 10985 18528
rect 10921 18468 10925 18524
rect 10925 18468 10981 18524
rect 10981 18468 10985 18524
rect 10921 18464 10985 18468
rect 11001 18524 11065 18528
rect 11001 18468 11005 18524
rect 11005 18468 11061 18524
rect 11061 18468 11065 18524
rect 11001 18464 11065 18468
rect 11081 18524 11145 18528
rect 11081 18468 11085 18524
rect 11085 18468 11141 18524
rect 11141 18468 11145 18524
rect 11081 18464 11145 18468
rect 15786 18524 15850 18528
rect 15786 18468 15790 18524
rect 15790 18468 15846 18524
rect 15846 18468 15850 18524
rect 15786 18464 15850 18468
rect 15866 18524 15930 18528
rect 15866 18468 15870 18524
rect 15870 18468 15926 18524
rect 15926 18468 15930 18524
rect 15866 18464 15930 18468
rect 15946 18524 16010 18528
rect 15946 18468 15950 18524
rect 15950 18468 16006 18524
rect 16006 18468 16010 18524
rect 15946 18464 16010 18468
rect 16026 18524 16090 18528
rect 16026 18468 16030 18524
rect 16030 18468 16086 18524
rect 16086 18468 16090 18524
rect 16026 18464 16090 18468
rect 20731 18524 20795 18528
rect 20731 18468 20735 18524
rect 20735 18468 20791 18524
rect 20791 18468 20795 18524
rect 20731 18464 20795 18468
rect 20811 18524 20875 18528
rect 20811 18468 20815 18524
rect 20815 18468 20871 18524
rect 20871 18468 20875 18524
rect 20811 18464 20875 18468
rect 20891 18524 20955 18528
rect 20891 18468 20895 18524
rect 20895 18468 20951 18524
rect 20951 18468 20955 18524
rect 20891 18464 20955 18468
rect 20971 18524 21035 18528
rect 20971 18468 20975 18524
rect 20975 18468 21031 18524
rect 21031 18468 21035 18524
rect 20971 18464 21035 18468
rect 3424 17980 3488 17984
rect 3424 17924 3428 17980
rect 3428 17924 3484 17980
rect 3484 17924 3488 17980
rect 3424 17920 3488 17924
rect 3504 17980 3568 17984
rect 3504 17924 3508 17980
rect 3508 17924 3564 17980
rect 3564 17924 3568 17980
rect 3504 17920 3568 17924
rect 3584 17980 3648 17984
rect 3584 17924 3588 17980
rect 3588 17924 3644 17980
rect 3644 17924 3648 17980
rect 3584 17920 3648 17924
rect 3664 17980 3728 17984
rect 3664 17924 3668 17980
rect 3668 17924 3724 17980
rect 3724 17924 3728 17980
rect 3664 17920 3728 17924
rect 8369 17980 8433 17984
rect 8369 17924 8373 17980
rect 8373 17924 8429 17980
rect 8429 17924 8433 17980
rect 8369 17920 8433 17924
rect 8449 17980 8513 17984
rect 8449 17924 8453 17980
rect 8453 17924 8509 17980
rect 8509 17924 8513 17980
rect 8449 17920 8513 17924
rect 8529 17980 8593 17984
rect 8529 17924 8533 17980
rect 8533 17924 8589 17980
rect 8589 17924 8593 17980
rect 8529 17920 8593 17924
rect 8609 17980 8673 17984
rect 8609 17924 8613 17980
rect 8613 17924 8669 17980
rect 8669 17924 8673 17980
rect 8609 17920 8673 17924
rect 13314 17980 13378 17984
rect 13314 17924 13318 17980
rect 13318 17924 13374 17980
rect 13374 17924 13378 17980
rect 13314 17920 13378 17924
rect 13394 17980 13458 17984
rect 13394 17924 13398 17980
rect 13398 17924 13454 17980
rect 13454 17924 13458 17980
rect 13394 17920 13458 17924
rect 13474 17980 13538 17984
rect 13474 17924 13478 17980
rect 13478 17924 13534 17980
rect 13534 17924 13538 17980
rect 13474 17920 13538 17924
rect 13554 17980 13618 17984
rect 13554 17924 13558 17980
rect 13558 17924 13614 17980
rect 13614 17924 13618 17980
rect 13554 17920 13618 17924
rect 18259 17980 18323 17984
rect 18259 17924 18263 17980
rect 18263 17924 18319 17980
rect 18319 17924 18323 17980
rect 18259 17920 18323 17924
rect 18339 17980 18403 17984
rect 18339 17924 18343 17980
rect 18343 17924 18399 17980
rect 18399 17924 18403 17980
rect 18339 17920 18403 17924
rect 18419 17980 18483 17984
rect 18419 17924 18423 17980
rect 18423 17924 18479 17980
rect 18479 17924 18483 17980
rect 18419 17920 18483 17924
rect 18499 17980 18563 17984
rect 18499 17924 18503 17980
rect 18503 17924 18559 17980
rect 18559 17924 18563 17980
rect 18499 17920 18563 17924
rect 5896 17436 5960 17440
rect 5896 17380 5900 17436
rect 5900 17380 5956 17436
rect 5956 17380 5960 17436
rect 5896 17376 5960 17380
rect 5976 17436 6040 17440
rect 5976 17380 5980 17436
rect 5980 17380 6036 17436
rect 6036 17380 6040 17436
rect 5976 17376 6040 17380
rect 6056 17436 6120 17440
rect 6056 17380 6060 17436
rect 6060 17380 6116 17436
rect 6116 17380 6120 17436
rect 6056 17376 6120 17380
rect 6136 17436 6200 17440
rect 6136 17380 6140 17436
rect 6140 17380 6196 17436
rect 6196 17380 6200 17436
rect 6136 17376 6200 17380
rect 10841 17436 10905 17440
rect 10841 17380 10845 17436
rect 10845 17380 10901 17436
rect 10901 17380 10905 17436
rect 10841 17376 10905 17380
rect 10921 17436 10985 17440
rect 10921 17380 10925 17436
rect 10925 17380 10981 17436
rect 10981 17380 10985 17436
rect 10921 17376 10985 17380
rect 11001 17436 11065 17440
rect 11001 17380 11005 17436
rect 11005 17380 11061 17436
rect 11061 17380 11065 17436
rect 11001 17376 11065 17380
rect 11081 17436 11145 17440
rect 11081 17380 11085 17436
rect 11085 17380 11141 17436
rect 11141 17380 11145 17436
rect 11081 17376 11145 17380
rect 15786 17436 15850 17440
rect 15786 17380 15790 17436
rect 15790 17380 15846 17436
rect 15846 17380 15850 17436
rect 15786 17376 15850 17380
rect 15866 17436 15930 17440
rect 15866 17380 15870 17436
rect 15870 17380 15926 17436
rect 15926 17380 15930 17436
rect 15866 17376 15930 17380
rect 15946 17436 16010 17440
rect 15946 17380 15950 17436
rect 15950 17380 16006 17436
rect 16006 17380 16010 17436
rect 15946 17376 16010 17380
rect 16026 17436 16090 17440
rect 16026 17380 16030 17436
rect 16030 17380 16086 17436
rect 16086 17380 16090 17436
rect 16026 17376 16090 17380
rect 20731 17436 20795 17440
rect 20731 17380 20735 17436
rect 20735 17380 20791 17436
rect 20791 17380 20795 17436
rect 20731 17376 20795 17380
rect 20811 17436 20875 17440
rect 20811 17380 20815 17436
rect 20815 17380 20871 17436
rect 20871 17380 20875 17436
rect 20811 17376 20875 17380
rect 20891 17436 20955 17440
rect 20891 17380 20895 17436
rect 20895 17380 20951 17436
rect 20951 17380 20955 17436
rect 20891 17376 20955 17380
rect 20971 17436 21035 17440
rect 20971 17380 20975 17436
rect 20975 17380 21031 17436
rect 21031 17380 21035 17436
rect 20971 17376 21035 17380
rect 3424 16892 3488 16896
rect 3424 16836 3428 16892
rect 3428 16836 3484 16892
rect 3484 16836 3488 16892
rect 3424 16832 3488 16836
rect 3504 16892 3568 16896
rect 3504 16836 3508 16892
rect 3508 16836 3564 16892
rect 3564 16836 3568 16892
rect 3504 16832 3568 16836
rect 3584 16892 3648 16896
rect 3584 16836 3588 16892
rect 3588 16836 3644 16892
rect 3644 16836 3648 16892
rect 3584 16832 3648 16836
rect 3664 16892 3728 16896
rect 3664 16836 3668 16892
rect 3668 16836 3724 16892
rect 3724 16836 3728 16892
rect 3664 16832 3728 16836
rect 8369 16892 8433 16896
rect 8369 16836 8373 16892
rect 8373 16836 8429 16892
rect 8429 16836 8433 16892
rect 8369 16832 8433 16836
rect 8449 16892 8513 16896
rect 8449 16836 8453 16892
rect 8453 16836 8509 16892
rect 8509 16836 8513 16892
rect 8449 16832 8513 16836
rect 8529 16892 8593 16896
rect 8529 16836 8533 16892
rect 8533 16836 8589 16892
rect 8589 16836 8593 16892
rect 8529 16832 8593 16836
rect 8609 16892 8673 16896
rect 8609 16836 8613 16892
rect 8613 16836 8669 16892
rect 8669 16836 8673 16892
rect 8609 16832 8673 16836
rect 13314 16892 13378 16896
rect 13314 16836 13318 16892
rect 13318 16836 13374 16892
rect 13374 16836 13378 16892
rect 13314 16832 13378 16836
rect 13394 16892 13458 16896
rect 13394 16836 13398 16892
rect 13398 16836 13454 16892
rect 13454 16836 13458 16892
rect 13394 16832 13458 16836
rect 13474 16892 13538 16896
rect 13474 16836 13478 16892
rect 13478 16836 13534 16892
rect 13534 16836 13538 16892
rect 13474 16832 13538 16836
rect 13554 16892 13618 16896
rect 13554 16836 13558 16892
rect 13558 16836 13614 16892
rect 13614 16836 13618 16892
rect 13554 16832 13618 16836
rect 18259 16892 18323 16896
rect 18259 16836 18263 16892
rect 18263 16836 18319 16892
rect 18319 16836 18323 16892
rect 18259 16832 18323 16836
rect 18339 16892 18403 16896
rect 18339 16836 18343 16892
rect 18343 16836 18399 16892
rect 18399 16836 18403 16892
rect 18339 16832 18403 16836
rect 18419 16892 18483 16896
rect 18419 16836 18423 16892
rect 18423 16836 18479 16892
rect 18479 16836 18483 16892
rect 18419 16832 18483 16836
rect 18499 16892 18563 16896
rect 18499 16836 18503 16892
rect 18503 16836 18559 16892
rect 18559 16836 18563 16892
rect 18499 16832 18563 16836
rect 5896 16348 5960 16352
rect 5896 16292 5900 16348
rect 5900 16292 5956 16348
rect 5956 16292 5960 16348
rect 5896 16288 5960 16292
rect 5976 16348 6040 16352
rect 5976 16292 5980 16348
rect 5980 16292 6036 16348
rect 6036 16292 6040 16348
rect 5976 16288 6040 16292
rect 6056 16348 6120 16352
rect 6056 16292 6060 16348
rect 6060 16292 6116 16348
rect 6116 16292 6120 16348
rect 6056 16288 6120 16292
rect 6136 16348 6200 16352
rect 6136 16292 6140 16348
rect 6140 16292 6196 16348
rect 6196 16292 6200 16348
rect 6136 16288 6200 16292
rect 10841 16348 10905 16352
rect 10841 16292 10845 16348
rect 10845 16292 10901 16348
rect 10901 16292 10905 16348
rect 10841 16288 10905 16292
rect 10921 16348 10985 16352
rect 10921 16292 10925 16348
rect 10925 16292 10981 16348
rect 10981 16292 10985 16348
rect 10921 16288 10985 16292
rect 11001 16348 11065 16352
rect 11001 16292 11005 16348
rect 11005 16292 11061 16348
rect 11061 16292 11065 16348
rect 11001 16288 11065 16292
rect 11081 16348 11145 16352
rect 11081 16292 11085 16348
rect 11085 16292 11141 16348
rect 11141 16292 11145 16348
rect 11081 16288 11145 16292
rect 15786 16348 15850 16352
rect 15786 16292 15790 16348
rect 15790 16292 15846 16348
rect 15846 16292 15850 16348
rect 15786 16288 15850 16292
rect 15866 16348 15930 16352
rect 15866 16292 15870 16348
rect 15870 16292 15926 16348
rect 15926 16292 15930 16348
rect 15866 16288 15930 16292
rect 15946 16348 16010 16352
rect 15946 16292 15950 16348
rect 15950 16292 16006 16348
rect 16006 16292 16010 16348
rect 15946 16288 16010 16292
rect 16026 16348 16090 16352
rect 16026 16292 16030 16348
rect 16030 16292 16086 16348
rect 16086 16292 16090 16348
rect 16026 16288 16090 16292
rect 20731 16348 20795 16352
rect 20731 16292 20735 16348
rect 20735 16292 20791 16348
rect 20791 16292 20795 16348
rect 20731 16288 20795 16292
rect 20811 16348 20875 16352
rect 20811 16292 20815 16348
rect 20815 16292 20871 16348
rect 20871 16292 20875 16348
rect 20811 16288 20875 16292
rect 20891 16348 20955 16352
rect 20891 16292 20895 16348
rect 20895 16292 20951 16348
rect 20951 16292 20955 16348
rect 20891 16288 20955 16292
rect 20971 16348 21035 16352
rect 20971 16292 20975 16348
rect 20975 16292 21031 16348
rect 21031 16292 21035 16348
rect 20971 16288 21035 16292
rect 3424 15804 3488 15808
rect 3424 15748 3428 15804
rect 3428 15748 3484 15804
rect 3484 15748 3488 15804
rect 3424 15744 3488 15748
rect 3504 15804 3568 15808
rect 3504 15748 3508 15804
rect 3508 15748 3564 15804
rect 3564 15748 3568 15804
rect 3504 15744 3568 15748
rect 3584 15804 3648 15808
rect 3584 15748 3588 15804
rect 3588 15748 3644 15804
rect 3644 15748 3648 15804
rect 3584 15744 3648 15748
rect 3664 15804 3728 15808
rect 3664 15748 3668 15804
rect 3668 15748 3724 15804
rect 3724 15748 3728 15804
rect 3664 15744 3728 15748
rect 8369 15804 8433 15808
rect 8369 15748 8373 15804
rect 8373 15748 8429 15804
rect 8429 15748 8433 15804
rect 8369 15744 8433 15748
rect 8449 15804 8513 15808
rect 8449 15748 8453 15804
rect 8453 15748 8509 15804
rect 8509 15748 8513 15804
rect 8449 15744 8513 15748
rect 8529 15804 8593 15808
rect 8529 15748 8533 15804
rect 8533 15748 8589 15804
rect 8589 15748 8593 15804
rect 8529 15744 8593 15748
rect 8609 15804 8673 15808
rect 8609 15748 8613 15804
rect 8613 15748 8669 15804
rect 8669 15748 8673 15804
rect 8609 15744 8673 15748
rect 13314 15804 13378 15808
rect 13314 15748 13318 15804
rect 13318 15748 13374 15804
rect 13374 15748 13378 15804
rect 13314 15744 13378 15748
rect 13394 15804 13458 15808
rect 13394 15748 13398 15804
rect 13398 15748 13454 15804
rect 13454 15748 13458 15804
rect 13394 15744 13458 15748
rect 13474 15804 13538 15808
rect 13474 15748 13478 15804
rect 13478 15748 13534 15804
rect 13534 15748 13538 15804
rect 13474 15744 13538 15748
rect 13554 15804 13618 15808
rect 13554 15748 13558 15804
rect 13558 15748 13614 15804
rect 13614 15748 13618 15804
rect 13554 15744 13618 15748
rect 18259 15804 18323 15808
rect 18259 15748 18263 15804
rect 18263 15748 18319 15804
rect 18319 15748 18323 15804
rect 18259 15744 18323 15748
rect 18339 15804 18403 15808
rect 18339 15748 18343 15804
rect 18343 15748 18399 15804
rect 18399 15748 18403 15804
rect 18339 15744 18403 15748
rect 18419 15804 18483 15808
rect 18419 15748 18423 15804
rect 18423 15748 18479 15804
rect 18479 15748 18483 15804
rect 18419 15744 18483 15748
rect 18499 15804 18563 15808
rect 18499 15748 18503 15804
rect 18503 15748 18559 15804
rect 18559 15748 18563 15804
rect 18499 15744 18563 15748
rect 5896 15260 5960 15264
rect 5896 15204 5900 15260
rect 5900 15204 5956 15260
rect 5956 15204 5960 15260
rect 5896 15200 5960 15204
rect 5976 15260 6040 15264
rect 5976 15204 5980 15260
rect 5980 15204 6036 15260
rect 6036 15204 6040 15260
rect 5976 15200 6040 15204
rect 6056 15260 6120 15264
rect 6056 15204 6060 15260
rect 6060 15204 6116 15260
rect 6116 15204 6120 15260
rect 6056 15200 6120 15204
rect 6136 15260 6200 15264
rect 6136 15204 6140 15260
rect 6140 15204 6196 15260
rect 6196 15204 6200 15260
rect 6136 15200 6200 15204
rect 10841 15260 10905 15264
rect 10841 15204 10845 15260
rect 10845 15204 10901 15260
rect 10901 15204 10905 15260
rect 10841 15200 10905 15204
rect 10921 15260 10985 15264
rect 10921 15204 10925 15260
rect 10925 15204 10981 15260
rect 10981 15204 10985 15260
rect 10921 15200 10985 15204
rect 11001 15260 11065 15264
rect 11001 15204 11005 15260
rect 11005 15204 11061 15260
rect 11061 15204 11065 15260
rect 11001 15200 11065 15204
rect 11081 15260 11145 15264
rect 11081 15204 11085 15260
rect 11085 15204 11141 15260
rect 11141 15204 11145 15260
rect 11081 15200 11145 15204
rect 15786 15260 15850 15264
rect 15786 15204 15790 15260
rect 15790 15204 15846 15260
rect 15846 15204 15850 15260
rect 15786 15200 15850 15204
rect 15866 15260 15930 15264
rect 15866 15204 15870 15260
rect 15870 15204 15926 15260
rect 15926 15204 15930 15260
rect 15866 15200 15930 15204
rect 15946 15260 16010 15264
rect 15946 15204 15950 15260
rect 15950 15204 16006 15260
rect 16006 15204 16010 15260
rect 15946 15200 16010 15204
rect 16026 15260 16090 15264
rect 16026 15204 16030 15260
rect 16030 15204 16086 15260
rect 16086 15204 16090 15260
rect 16026 15200 16090 15204
rect 20731 15260 20795 15264
rect 20731 15204 20735 15260
rect 20735 15204 20791 15260
rect 20791 15204 20795 15260
rect 20731 15200 20795 15204
rect 20811 15260 20875 15264
rect 20811 15204 20815 15260
rect 20815 15204 20871 15260
rect 20871 15204 20875 15260
rect 20811 15200 20875 15204
rect 20891 15260 20955 15264
rect 20891 15204 20895 15260
rect 20895 15204 20951 15260
rect 20951 15204 20955 15260
rect 20891 15200 20955 15204
rect 20971 15260 21035 15264
rect 20971 15204 20975 15260
rect 20975 15204 21031 15260
rect 21031 15204 21035 15260
rect 20971 15200 21035 15204
rect 3424 14716 3488 14720
rect 3424 14660 3428 14716
rect 3428 14660 3484 14716
rect 3484 14660 3488 14716
rect 3424 14656 3488 14660
rect 3504 14716 3568 14720
rect 3504 14660 3508 14716
rect 3508 14660 3564 14716
rect 3564 14660 3568 14716
rect 3504 14656 3568 14660
rect 3584 14716 3648 14720
rect 3584 14660 3588 14716
rect 3588 14660 3644 14716
rect 3644 14660 3648 14716
rect 3584 14656 3648 14660
rect 3664 14716 3728 14720
rect 3664 14660 3668 14716
rect 3668 14660 3724 14716
rect 3724 14660 3728 14716
rect 3664 14656 3728 14660
rect 8369 14716 8433 14720
rect 8369 14660 8373 14716
rect 8373 14660 8429 14716
rect 8429 14660 8433 14716
rect 8369 14656 8433 14660
rect 8449 14716 8513 14720
rect 8449 14660 8453 14716
rect 8453 14660 8509 14716
rect 8509 14660 8513 14716
rect 8449 14656 8513 14660
rect 8529 14716 8593 14720
rect 8529 14660 8533 14716
rect 8533 14660 8589 14716
rect 8589 14660 8593 14716
rect 8529 14656 8593 14660
rect 8609 14716 8673 14720
rect 8609 14660 8613 14716
rect 8613 14660 8669 14716
rect 8669 14660 8673 14716
rect 8609 14656 8673 14660
rect 13314 14716 13378 14720
rect 13314 14660 13318 14716
rect 13318 14660 13374 14716
rect 13374 14660 13378 14716
rect 13314 14656 13378 14660
rect 13394 14716 13458 14720
rect 13394 14660 13398 14716
rect 13398 14660 13454 14716
rect 13454 14660 13458 14716
rect 13394 14656 13458 14660
rect 13474 14716 13538 14720
rect 13474 14660 13478 14716
rect 13478 14660 13534 14716
rect 13534 14660 13538 14716
rect 13474 14656 13538 14660
rect 13554 14716 13618 14720
rect 13554 14660 13558 14716
rect 13558 14660 13614 14716
rect 13614 14660 13618 14716
rect 13554 14656 13618 14660
rect 18259 14716 18323 14720
rect 18259 14660 18263 14716
rect 18263 14660 18319 14716
rect 18319 14660 18323 14716
rect 18259 14656 18323 14660
rect 18339 14716 18403 14720
rect 18339 14660 18343 14716
rect 18343 14660 18399 14716
rect 18399 14660 18403 14716
rect 18339 14656 18403 14660
rect 18419 14716 18483 14720
rect 18419 14660 18423 14716
rect 18423 14660 18479 14716
rect 18479 14660 18483 14716
rect 18419 14656 18483 14660
rect 18499 14716 18563 14720
rect 18499 14660 18503 14716
rect 18503 14660 18559 14716
rect 18559 14660 18563 14716
rect 18499 14656 18563 14660
rect 5896 14172 5960 14176
rect 5896 14116 5900 14172
rect 5900 14116 5956 14172
rect 5956 14116 5960 14172
rect 5896 14112 5960 14116
rect 5976 14172 6040 14176
rect 5976 14116 5980 14172
rect 5980 14116 6036 14172
rect 6036 14116 6040 14172
rect 5976 14112 6040 14116
rect 6056 14172 6120 14176
rect 6056 14116 6060 14172
rect 6060 14116 6116 14172
rect 6116 14116 6120 14172
rect 6056 14112 6120 14116
rect 6136 14172 6200 14176
rect 6136 14116 6140 14172
rect 6140 14116 6196 14172
rect 6196 14116 6200 14172
rect 6136 14112 6200 14116
rect 10841 14172 10905 14176
rect 10841 14116 10845 14172
rect 10845 14116 10901 14172
rect 10901 14116 10905 14172
rect 10841 14112 10905 14116
rect 10921 14172 10985 14176
rect 10921 14116 10925 14172
rect 10925 14116 10981 14172
rect 10981 14116 10985 14172
rect 10921 14112 10985 14116
rect 11001 14172 11065 14176
rect 11001 14116 11005 14172
rect 11005 14116 11061 14172
rect 11061 14116 11065 14172
rect 11001 14112 11065 14116
rect 11081 14172 11145 14176
rect 11081 14116 11085 14172
rect 11085 14116 11141 14172
rect 11141 14116 11145 14172
rect 11081 14112 11145 14116
rect 15786 14172 15850 14176
rect 15786 14116 15790 14172
rect 15790 14116 15846 14172
rect 15846 14116 15850 14172
rect 15786 14112 15850 14116
rect 15866 14172 15930 14176
rect 15866 14116 15870 14172
rect 15870 14116 15926 14172
rect 15926 14116 15930 14172
rect 15866 14112 15930 14116
rect 15946 14172 16010 14176
rect 15946 14116 15950 14172
rect 15950 14116 16006 14172
rect 16006 14116 16010 14172
rect 15946 14112 16010 14116
rect 16026 14172 16090 14176
rect 16026 14116 16030 14172
rect 16030 14116 16086 14172
rect 16086 14116 16090 14172
rect 16026 14112 16090 14116
rect 20731 14172 20795 14176
rect 20731 14116 20735 14172
rect 20735 14116 20791 14172
rect 20791 14116 20795 14172
rect 20731 14112 20795 14116
rect 20811 14172 20875 14176
rect 20811 14116 20815 14172
rect 20815 14116 20871 14172
rect 20871 14116 20875 14172
rect 20811 14112 20875 14116
rect 20891 14172 20955 14176
rect 20891 14116 20895 14172
rect 20895 14116 20951 14172
rect 20951 14116 20955 14172
rect 20891 14112 20955 14116
rect 20971 14172 21035 14176
rect 20971 14116 20975 14172
rect 20975 14116 21031 14172
rect 21031 14116 21035 14172
rect 20971 14112 21035 14116
rect 3424 13628 3488 13632
rect 3424 13572 3428 13628
rect 3428 13572 3484 13628
rect 3484 13572 3488 13628
rect 3424 13568 3488 13572
rect 3504 13628 3568 13632
rect 3504 13572 3508 13628
rect 3508 13572 3564 13628
rect 3564 13572 3568 13628
rect 3504 13568 3568 13572
rect 3584 13628 3648 13632
rect 3584 13572 3588 13628
rect 3588 13572 3644 13628
rect 3644 13572 3648 13628
rect 3584 13568 3648 13572
rect 3664 13628 3728 13632
rect 3664 13572 3668 13628
rect 3668 13572 3724 13628
rect 3724 13572 3728 13628
rect 3664 13568 3728 13572
rect 8369 13628 8433 13632
rect 8369 13572 8373 13628
rect 8373 13572 8429 13628
rect 8429 13572 8433 13628
rect 8369 13568 8433 13572
rect 8449 13628 8513 13632
rect 8449 13572 8453 13628
rect 8453 13572 8509 13628
rect 8509 13572 8513 13628
rect 8449 13568 8513 13572
rect 8529 13628 8593 13632
rect 8529 13572 8533 13628
rect 8533 13572 8589 13628
rect 8589 13572 8593 13628
rect 8529 13568 8593 13572
rect 8609 13628 8673 13632
rect 8609 13572 8613 13628
rect 8613 13572 8669 13628
rect 8669 13572 8673 13628
rect 8609 13568 8673 13572
rect 13314 13628 13378 13632
rect 13314 13572 13318 13628
rect 13318 13572 13374 13628
rect 13374 13572 13378 13628
rect 13314 13568 13378 13572
rect 13394 13628 13458 13632
rect 13394 13572 13398 13628
rect 13398 13572 13454 13628
rect 13454 13572 13458 13628
rect 13394 13568 13458 13572
rect 13474 13628 13538 13632
rect 13474 13572 13478 13628
rect 13478 13572 13534 13628
rect 13534 13572 13538 13628
rect 13474 13568 13538 13572
rect 13554 13628 13618 13632
rect 13554 13572 13558 13628
rect 13558 13572 13614 13628
rect 13614 13572 13618 13628
rect 13554 13568 13618 13572
rect 18259 13628 18323 13632
rect 18259 13572 18263 13628
rect 18263 13572 18319 13628
rect 18319 13572 18323 13628
rect 18259 13568 18323 13572
rect 18339 13628 18403 13632
rect 18339 13572 18343 13628
rect 18343 13572 18399 13628
rect 18399 13572 18403 13628
rect 18339 13568 18403 13572
rect 18419 13628 18483 13632
rect 18419 13572 18423 13628
rect 18423 13572 18479 13628
rect 18479 13572 18483 13628
rect 18419 13568 18483 13572
rect 18499 13628 18563 13632
rect 18499 13572 18503 13628
rect 18503 13572 18559 13628
rect 18559 13572 18563 13628
rect 18499 13568 18563 13572
rect 5896 13084 5960 13088
rect 5896 13028 5900 13084
rect 5900 13028 5956 13084
rect 5956 13028 5960 13084
rect 5896 13024 5960 13028
rect 5976 13084 6040 13088
rect 5976 13028 5980 13084
rect 5980 13028 6036 13084
rect 6036 13028 6040 13084
rect 5976 13024 6040 13028
rect 6056 13084 6120 13088
rect 6056 13028 6060 13084
rect 6060 13028 6116 13084
rect 6116 13028 6120 13084
rect 6056 13024 6120 13028
rect 6136 13084 6200 13088
rect 6136 13028 6140 13084
rect 6140 13028 6196 13084
rect 6196 13028 6200 13084
rect 6136 13024 6200 13028
rect 10841 13084 10905 13088
rect 10841 13028 10845 13084
rect 10845 13028 10901 13084
rect 10901 13028 10905 13084
rect 10841 13024 10905 13028
rect 10921 13084 10985 13088
rect 10921 13028 10925 13084
rect 10925 13028 10981 13084
rect 10981 13028 10985 13084
rect 10921 13024 10985 13028
rect 11001 13084 11065 13088
rect 11001 13028 11005 13084
rect 11005 13028 11061 13084
rect 11061 13028 11065 13084
rect 11001 13024 11065 13028
rect 11081 13084 11145 13088
rect 11081 13028 11085 13084
rect 11085 13028 11141 13084
rect 11141 13028 11145 13084
rect 11081 13024 11145 13028
rect 15786 13084 15850 13088
rect 15786 13028 15790 13084
rect 15790 13028 15846 13084
rect 15846 13028 15850 13084
rect 15786 13024 15850 13028
rect 15866 13084 15930 13088
rect 15866 13028 15870 13084
rect 15870 13028 15926 13084
rect 15926 13028 15930 13084
rect 15866 13024 15930 13028
rect 15946 13084 16010 13088
rect 15946 13028 15950 13084
rect 15950 13028 16006 13084
rect 16006 13028 16010 13084
rect 15946 13024 16010 13028
rect 16026 13084 16090 13088
rect 16026 13028 16030 13084
rect 16030 13028 16086 13084
rect 16086 13028 16090 13084
rect 16026 13024 16090 13028
rect 20731 13084 20795 13088
rect 20731 13028 20735 13084
rect 20735 13028 20791 13084
rect 20791 13028 20795 13084
rect 20731 13024 20795 13028
rect 20811 13084 20875 13088
rect 20811 13028 20815 13084
rect 20815 13028 20871 13084
rect 20871 13028 20875 13084
rect 20811 13024 20875 13028
rect 20891 13084 20955 13088
rect 20891 13028 20895 13084
rect 20895 13028 20951 13084
rect 20951 13028 20955 13084
rect 20891 13024 20955 13028
rect 20971 13084 21035 13088
rect 20971 13028 20975 13084
rect 20975 13028 21031 13084
rect 21031 13028 21035 13084
rect 20971 13024 21035 13028
rect 3424 12540 3488 12544
rect 3424 12484 3428 12540
rect 3428 12484 3484 12540
rect 3484 12484 3488 12540
rect 3424 12480 3488 12484
rect 3504 12540 3568 12544
rect 3504 12484 3508 12540
rect 3508 12484 3564 12540
rect 3564 12484 3568 12540
rect 3504 12480 3568 12484
rect 3584 12540 3648 12544
rect 3584 12484 3588 12540
rect 3588 12484 3644 12540
rect 3644 12484 3648 12540
rect 3584 12480 3648 12484
rect 3664 12540 3728 12544
rect 3664 12484 3668 12540
rect 3668 12484 3724 12540
rect 3724 12484 3728 12540
rect 3664 12480 3728 12484
rect 8369 12540 8433 12544
rect 8369 12484 8373 12540
rect 8373 12484 8429 12540
rect 8429 12484 8433 12540
rect 8369 12480 8433 12484
rect 8449 12540 8513 12544
rect 8449 12484 8453 12540
rect 8453 12484 8509 12540
rect 8509 12484 8513 12540
rect 8449 12480 8513 12484
rect 8529 12540 8593 12544
rect 8529 12484 8533 12540
rect 8533 12484 8589 12540
rect 8589 12484 8593 12540
rect 8529 12480 8593 12484
rect 8609 12540 8673 12544
rect 8609 12484 8613 12540
rect 8613 12484 8669 12540
rect 8669 12484 8673 12540
rect 8609 12480 8673 12484
rect 13314 12540 13378 12544
rect 13314 12484 13318 12540
rect 13318 12484 13374 12540
rect 13374 12484 13378 12540
rect 13314 12480 13378 12484
rect 13394 12540 13458 12544
rect 13394 12484 13398 12540
rect 13398 12484 13454 12540
rect 13454 12484 13458 12540
rect 13394 12480 13458 12484
rect 13474 12540 13538 12544
rect 13474 12484 13478 12540
rect 13478 12484 13534 12540
rect 13534 12484 13538 12540
rect 13474 12480 13538 12484
rect 13554 12540 13618 12544
rect 13554 12484 13558 12540
rect 13558 12484 13614 12540
rect 13614 12484 13618 12540
rect 13554 12480 13618 12484
rect 18259 12540 18323 12544
rect 18259 12484 18263 12540
rect 18263 12484 18319 12540
rect 18319 12484 18323 12540
rect 18259 12480 18323 12484
rect 18339 12540 18403 12544
rect 18339 12484 18343 12540
rect 18343 12484 18399 12540
rect 18399 12484 18403 12540
rect 18339 12480 18403 12484
rect 18419 12540 18483 12544
rect 18419 12484 18423 12540
rect 18423 12484 18479 12540
rect 18479 12484 18483 12540
rect 18419 12480 18483 12484
rect 18499 12540 18563 12544
rect 18499 12484 18503 12540
rect 18503 12484 18559 12540
rect 18559 12484 18563 12540
rect 18499 12480 18563 12484
rect 5896 11996 5960 12000
rect 5896 11940 5900 11996
rect 5900 11940 5956 11996
rect 5956 11940 5960 11996
rect 5896 11936 5960 11940
rect 5976 11996 6040 12000
rect 5976 11940 5980 11996
rect 5980 11940 6036 11996
rect 6036 11940 6040 11996
rect 5976 11936 6040 11940
rect 6056 11996 6120 12000
rect 6056 11940 6060 11996
rect 6060 11940 6116 11996
rect 6116 11940 6120 11996
rect 6056 11936 6120 11940
rect 6136 11996 6200 12000
rect 6136 11940 6140 11996
rect 6140 11940 6196 11996
rect 6196 11940 6200 11996
rect 6136 11936 6200 11940
rect 10841 11996 10905 12000
rect 10841 11940 10845 11996
rect 10845 11940 10901 11996
rect 10901 11940 10905 11996
rect 10841 11936 10905 11940
rect 10921 11996 10985 12000
rect 10921 11940 10925 11996
rect 10925 11940 10981 11996
rect 10981 11940 10985 11996
rect 10921 11936 10985 11940
rect 11001 11996 11065 12000
rect 11001 11940 11005 11996
rect 11005 11940 11061 11996
rect 11061 11940 11065 11996
rect 11001 11936 11065 11940
rect 11081 11996 11145 12000
rect 11081 11940 11085 11996
rect 11085 11940 11141 11996
rect 11141 11940 11145 11996
rect 11081 11936 11145 11940
rect 15786 11996 15850 12000
rect 15786 11940 15790 11996
rect 15790 11940 15846 11996
rect 15846 11940 15850 11996
rect 15786 11936 15850 11940
rect 15866 11996 15930 12000
rect 15866 11940 15870 11996
rect 15870 11940 15926 11996
rect 15926 11940 15930 11996
rect 15866 11936 15930 11940
rect 15946 11996 16010 12000
rect 15946 11940 15950 11996
rect 15950 11940 16006 11996
rect 16006 11940 16010 11996
rect 15946 11936 16010 11940
rect 16026 11996 16090 12000
rect 16026 11940 16030 11996
rect 16030 11940 16086 11996
rect 16086 11940 16090 11996
rect 16026 11936 16090 11940
rect 20731 11996 20795 12000
rect 20731 11940 20735 11996
rect 20735 11940 20791 11996
rect 20791 11940 20795 11996
rect 20731 11936 20795 11940
rect 20811 11996 20875 12000
rect 20811 11940 20815 11996
rect 20815 11940 20871 11996
rect 20871 11940 20875 11996
rect 20811 11936 20875 11940
rect 20891 11996 20955 12000
rect 20891 11940 20895 11996
rect 20895 11940 20951 11996
rect 20951 11940 20955 11996
rect 20891 11936 20955 11940
rect 20971 11996 21035 12000
rect 20971 11940 20975 11996
rect 20975 11940 21031 11996
rect 21031 11940 21035 11996
rect 20971 11936 21035 11940
rect 3424 11452 3488 11456
rect 3424 11396 3428 11452
rect 3428 11396 3484 11452
rect 3484 11396 3488 11452
rect 3424 11392 3488 11396
rect 3504 11452 3568 11456
rect 3504 11396 3508 11452
rect 3508 11396 3564 11452
rect 3564 11396 3568 11452
rect 3504 11392 3568 11396
rect 3584 11452 3648 11456
rect 3584 11396 3588 11452
rect 3588 11396 3644 11452
rect 3644 11396 3648 11452
rect 3584 11392 3648 11396
rect 3664 11452 3728 11456
rect 3664 11396 3668 11452
rect 3668 11396 3724 11452
rect 3724 11396 3728 11452
rect 3664 11392 3728 11396
rect 8369 11452 8433 11456
rect 8369 11396 8373 11452
rect 8373 11396 8429 11452
rect 8429 11396 8433 11452
rect 8369 11392 8433 11396
rect 8449 11452 8513 11456
rect 8449 11396 8453 11452
rect 8453 11396 8509 11452
rect 8509 11396 8513 11452
rect 8449 11392 8513 11396
rect 8529 11452 8593 11456
rect 8529 11396 8533 11452
rect 8533 11396 8589 11452
rect 8589 11396 8593 11452
rect 8529 11392 8593 11396
rect 8609 11452 8673 11456
rect 8609 11396 8613 11452
rect 8613 11396 8669 11452
rect 8669 11396 8673 11452
rect 8609 11392 8673 11396
rect 13314 11452 13378 11456
rect 13314 11396 13318 11452
rect 13318 11396 13374 11452
rect 13374 11396 13378 11452
rect 13314 11392 13378 11396
rect 13394 11452 13458 11456
rect 13394 11396 13398 11452
rect 13398 11396 13454 11452
rect 13454 11396 13458 11452
rect 13394 11392 13458 11396
rect 13474 11452 13538 11456
rect 13474 11396 13478 11452
rect 13478 11396 13534 11452
rect 13534 11396 13538 11452
rect 13474 11392 13538 11396
rect 13554 11452 13618 11456
rect 13554 11396 13558 11452
rect 13558 11396 13614 11452
rect 13614 11396 13618 11452
rect 13554 11392 13618 11396
rect 18259 11452 18323 11456
rect 18259 11396 18263 11452
rect 18263 11396 18319 11452
rect 18319 11396 18323 11452
rect 18259 11392 18323 11396
rect 18339 11452 18403 11456
rect 18339 11396 18343 11452
rect 18343 11396 18399 11452
rect 18399 11396 18403 11452
rect 18339 11392 18403 11396
rect 18419 11452 18483 11456
rect 18419 11396 18423 11452
rect 18423 11396 18479 11452
rect 18479 11396 18483 11452
rect 18419 11392 18483 11396
rect 18499 11452 18563 11456
rect 18499 11396 18503 11452
rect 18503 11396 18559 11452
rect 18559 11396 18563 11452
rect 18499 11392 18563 11396
rect 5896 10908 5960 10912
rect 5896 10852 5900 10908
rect 5900 10852 5956 10908
rect 5956 10852 5960 10908
rect 5896 10848 5960 10852
rect 5976 10908 6040 10912
rect 5976 10852 5980 10908
rect 5980 10852 6036 10908
rect 6036 10852 6040 10908
rect 5976 10848 6040 10852
rect 6056 10908 6120 10912
rect 6056 10852 6060 10908
rect 6060 10852 6116 10908
rect 6116 10852 6120 10908
rect 6056 10848 6120 10852
rect 6136 10908 6200 10912
rect 6136 10852 6140 10908
rect 6140 10852 6196 10908
rect 6196 10852 6200 10908
rect 6136 10848 6200 10852
rect 10841 10908 10905 10912
rect 10841 10852 10845 10908
rect 10845 10852 10901 10908
rect 10901 10852 10905 10908
rect 10841 10848 10905 10852
rect 10921 10908 10985 10912
rect 10921 10852 10925 10908
rect 10925 10852 10981 10908
rect 10981 10852 10985 10908
rect 10921 10848 10985 10852
rect 11001 10908 11065 10912
rect 11001 10852 11005 10908
rect 11005 10852 11061 10908
rect 11061 10852 11065 10908
rect 11001 10848 11065 10852
rect 11081 10908 11145 10912
rect 11081 10852 11085 10908
rect 11085 10852 11141 10908
rect 11141 10852 11145 10908
rect 11081 10848 11145 10852
rect 15786 10908 15850 10912
rect 15786 10852 15790 10908
rect 15790 10852 15846 10908
rect 15846 10852 15850 10908
rect 15786 10848 15850 10852
rect 15866 10908 15930 10912
rect 15866 10852 15870 10908
rect 15870 10852 15926 10908
rect 15926 10852 15930 10908
rect 15866 10848 15930 10852
rect 15946 10908 16010 10912
rect 15946 10852 15950 10908
rect 15950 10852 16006 10908
rect 16006 10852 16010 10908
rect 15946 10848 16010 10852
rect 16026 10908 16090 10912
rect 16026 10852 16030 10908
rect 16030 10852 16086 10908
rect 16086 10852 16090 10908
rect 16026 10848 16090 10852
rect 20731 10908 20795 10912
rect 20731 10852 20735 10908
rect 20735 10852 20791 10908
rect 20791 10852 20795 10908
rect 20731 10848 20795 10852
rect 20811 10908 20875 10912
rect 20811 10852 20815 10908
rect 20815 10852 20871 10908
rect 20871 10852 20875 10908
rect 20811 10848 20875 10852
rect 20891 10908 20955 10912
rect 20891 10852 20895 10908
rect 20895 10852 20951 10908
rect 20951 10852 20955 10908
rect 20891 10848 20955 10852
rect 20971 10908 21035 10912
rect 20971 10852 20975 10908
rect 20975 10852 21031 10908
rect 21031 10852 21035 10908
rect 20971 10848 21035 10852
rect 3424 10364 3488 10368
rect 3424 10308 3428 10364
rect 3428 10308 3484 10364
rect 3484 10308 3488 10364
rect 3424 10304 3488 10308
rect 3504 10364 3568 10368
rect 3504 10308 3508 10364
rect 3508 10308 3564 10364
rect 3564 10308 3568 10364
rect 3504 10304 3568 10308
rect 3584 10364 3648 10368
rect 3584 10308 3588 10364
rect 3588 10308 3644 10364
rect 3644 10308 3648 10364
rect 3584 10304 3648 10308
rect 3664 10364 3728 10368
rect 3664 10308 3668 10364
rect 3668 10308 3724 10364
rect 3724 10308 3728 10364
rect 3664 10304 3728 10308
rect 8369 10364 8433 10368
rect 8369 10308 8373 10364
rect 8373 10308 8429 10364
rect 8429 10308 8433 10364
rect 8369 10304 8433 10308
rect 8449 10364 8513 10368
rect 8449 10308 8453 10364
rect 8453 10308 8509 10364
rect 8509 10308 8513 10364
rect 8449 10304 8513 10308
rect 8529 10364 8593 10368
rect 8529 10308 8533 10364
rect 8533 10308 8589 10364
rect 8589 10308 8593 10364
rect 8529 10304 8593 10308
rect 8609 10364 8673 10368
rect 8609 10308 8613 10364
rect 8613 10308 8669 10364
rect 8669 10308 8673 10364
rect 8609 10304 8673 10308
rect 13314 10364 13378 10368
rect 13314 10308 13318 10364
rect 13318 10308 13374 10364
rect 13374 10308 13378 10364
rect 13314 10304 13378 10308
rect 13394 10364 13458 10368
rect 13394 10308 13398 10364
rect 13398 10308 13454 10364
rect 13454 10308 13458 10364
rect 13394 10304 13458 10308
rect 13474 10364 13538 10368
rect 13474 10308 13478 10364
rect 13478 10308 13534 10364
rect 13534 10308 13538 10364
rect 13474 10304 13538 10308
rect 13554 10364 13618 10368
rect 13554 10308 13558 10364
rect 13558 10308 13614 10364
rect 13614 10308 13618 10364
rect 13554 10304 13618 10308
rect 18259 10364 18323 10368
rect 18259 10308 18263 10364
rect 18263 10308 18319 10364
rect 18319 10308 18323 10364
rect 18259 10304 18323 10308
rect 18339 10364 18403 10368
rect 18339 10308 18343 10364
rect 18343 10308 18399 10364
rect 18399 10308 18403 10364
rect 18339 10304 18403 10308
rect 18419 10364 18483 10368
rect 18419 10308 18423 10364
rect 18423 10308 18479 10364
rect 18479 10308 18483 10364
rect 18419 10304 18483 10308
rect 18499 10364 18563 10368
rect 18499 10308 18503 10364
rect 18503 10308 18559 10364
rect 18559 10308 18563 10364
rect 18499 10304 18563 10308
rect 5896 9820 5960 9824
rect 5896 9764 5900 9820
rect 5900 9764 5956 9820
rect 5956 9764 5960 9820
rect 5896 9760 5960 9764
rect 5976 9820 6040 9824
rect 5976 9764 5980 9820
rect 5980 9764 6036 9820
rect 6036 9764 6040 9820
rect 5976 9760 6040 9764
rect 6056 9820 6120 9824
rect 6056 9764 6060 9820
rect 6060 9764 6116 9820
rect 6116 9764 6120 9820
rect 6056 9760 6120 9764
rect 6136 9820 6200 9824
rect 6136 9764 6140 9820
rect 6140 9764 6196 9820
rect 6196 9764 6200 9820
rect 6136 9760 6200 9764
rect 10841 9820 10905 9824
rect 10841 9764 10845 9820
rect 10845 9764 10901 9820
rect 10901 9764 10905 9820
rect 10841 9760 10905 9764
rect 10921 9820 10985 9824
rect 10921 9764 10925 9820
rect 10925 9764 10981 9820
rect 10981 9764 10985 9820
rect 10921 9760 10985 9764
rect 11001 9820 11065 9824
rect 11001 9764 11005 9820
rect 11005 9764 11061 9820
rect 11061 9764 11065 9820
rect 11001 9760 11065 9764
rect 11081 9820 11145 9824
rect 11081 9764 11085 9820
rect 11085 9764 11141 9820
rect 11141 9764 11145 9820
rect 11081 9760 11145 9764
rect 15786 9820 15850 9824
rect 15786 9764 15790 9820
rect 15790 9764 15846 9820
rect 15846 9764 15850 9820
rect 15786 9760 15850 9764
rect 15866 9820 15930 9824
rect 15866 9764 15870 9820
rect 15870 9764 15926 9820
rect 15926 9764 15930 9820
rect 15866 9760 15930 9764
rect 15946 9820 16010 9824
rect 15946 9764 15950 9820
rect 15950 9764 16006 9820
rect 16006 9764 16010 9820
rect 15946 9760 16010 9764
rect 16026 9820 16090 9824
rect 16026 9764 16030 9820
rect 16030 9764 16086 9820
rect 16086 9764 16090 9820
rect 16026 9760 16090 9764
rect 20731 9820 20795 9824
rect 20731 9764 20735 9820
rect 20735 9764 20791 9820
rect 20791 9764 20795 9820
rect 20731 9760 20795 9764
rect 20811 9820 20875 9824
rect 20811 9764 20815 9820
rect 20815 9764 20871 9820
rect 20871 9764 20875 9820
rect 20811 9760 20875 9764
rect 20891 9820 20955 9824
rect 20891 9764 20895 9820
rect 20895 9764 20951 9820
rect 20951 9764 20955 9820
rect 20891 9760 20955 9764
rect 20971 9820 21035 9824
rect 20971 9764 20975 9820
rect 20975 9764 21031 9820
rect 21031 9764 21035 9820
rect 20971 9760 21035 9764
rect 3424 9276 3488 9280
rect 3424 9220 3428 9276
rect 3428 9220 3484 9276
rect 3484 9220 3488 9276
rect 3424 9216 3488 9220
rect 3504 9276 3568 9280
rect 3504 9220 3508 9276
rect 3508 9220 3564 9276
rect 3564 9220 3568 9276
rect 3504 9216 3568 9220
rect 3584 9276 3648 9280
rect 3584 9220 3588 9276
rect 3588 9220 3644 9276
rect 3644 9220 3648 9276
rect 3584 9216 3648 9220
rect 3664 9276 3728 9280
rect 3664 9220 3668 9276
rect 3668 9220 3724 9276
rect 3724 9220 3728 9276
rect 3664 9216 3728 9220
rect 8369 9276 8433 9280
rect 8369 9220 8373 9276
rect 8373 9220 8429 9276
rect 8429 9220 8433 9276
rect 8369 9216 8433 9220
rect 8449 9276 8513 9280
rect 8449 9220 8453 9276
rect 8453 9220 8509 9276
rect 8509 9220 8513 9276
rect 8449 9216 8513 9220
rect 8529 9276 8593 9280
rect 8529 9220 8533 9276
rect 8533 9220 8589 9276
rect 8589 9220 8593 9276
rect 8529 9216 8593 9220
rect 8609 9276 8673 9280
rect 8609 9220 8613 9276
rect 8613 9220 8669 9276
rect 8669 9220 8673 9276
rect 8609 9216 8673 9220
rect 13314 9276 13378 9280
rect 13314 9220 13318 9276
rect 13318 9220 13374 9276
rect 13374 9220 13378 9276
rect 13314 9216 13378 9220
rect 13394 9276 13458 9280
rect 13394 9220 13398 9276
rect 13398 9220 13454 9276
rect 13454 9220 13458 9276
rect 13394 9216 13458 9220
rect 13474 9276 13538 9280
rect 13474 9220 13478 9276
rect 13478 9220 13534 9276
rect 13534 9220 13538 9276
rect 13474 9216 13538 9220
rect 13554 9276 13618 9280
rect 13554 9220 13558 9276
rect 13558 9220 13614 9276
rect 13614 9220 13618 9276
rect 13554 9216 13618 9220
rect 18259 9276 18323 9280
rect 18259 9220 18263 9276
rect 18263 9220 18319 9276
rect 18319 9220 18323 9276
rect 18259 9216 18323 9220
rect 18339 9276 18403 9280
rect 18339 9220 18343 9276
rect 18343 9220 18399 9276
rect 18399 9220 18403 9276
rect 18339 9216 18403 9220
rect 18419 9276 18483 9280
rect 18419 9220 18423 9276
rect 18423 9220 18479 9276
rect 18479 9220 18483 9276
rect 18419 9216 18483 9220
rect 18499 9276 18563 9280
rect 18499 9220 18503 9276
rect 18503 9220 18559 9276
rect 18559 9220 18563 9276
rect 18499 9216 18563 9220
rect 5896 8732 5960 8736
rect 5896 8676 5900 8732
rect 5900 8676 5956 8732
rect 5956 8676 5960 8732
rect 5896 8672 5960 8676
rect 5976 8732 6040 8736
rect 5976 8676 5980 8732
rect 5980 8676 6036 8732
rect 6036 8676 6040 8732
rect 5976 8672 6040 8676
rect 6056 8732 6120 8736
rect 6056 8676 6060 8732
rect 6060 8676 6116 8732
rect 6116 8676 6120 8732
rect 6056 8672 6120 8676
rect 6136 8732 6200 8736
rect 6136 8676 6140 8732
rect 6140 8676 6196 8732
rect 6196 8676 6200 8732
rect 6136 8672 6200 8676
rect 10841 8732 10905 8736
rect 10841 8676 10845 8732
rect 10845 8676 10901 8732
rect 10901 8676 10905 8732
rect 10841 8672 10905 8676
rect 10921 8732 10985 8736
rect 10921 8676 10925 8732
rect 10925 8676 10981 8732
rect 10981 8676 10985 8732
rect 10921 8672 10985 8676
rect 11001 8732 11065 8736
rect 11001 8676 11005 8732
rect 11005 8676 11061 8732
rect 11061 8676 11065 8732
rect 11001 8672 11065 8676
rect 11081 8732 11145 8736
rect 11081 8676 11085 8732
rect 11085 8676 11141 8732
rect 11141 8676 11145 8732
rect 11081 8672 11145 8676
rect 15786 8732 15850 8736
rect 15786 8676 15790 8732
rect 15790 8676 15846 8732
rect 15846 8676 15850 8732
rect 15786 8672 15850 8676
rect 15866 8732 15930 8736
rect 15866 8676 15870 8732
rect 15870 8676 15926 8732
rect 15926 8676 15930 8732
rect 15866 8672 15930 8676
rect 15946 8732 16010 8736
rect 15946 8676 15950 8732
rect 15950 8676 16006 8732
rect 16006 8676 16010 8732
rect 15946 8672 16010 8676
rect 16026 8732 16090 8736
rect 16026 8676 16030 8732
rect 16030 8676 16086 8732
rect 16086 8676 16090 8732
rect 16026 8672 16090 8676
rect 20731 8732 20795 8736
rect 20731 8676 20735 8732
rect 20735 8676 20791 8732
rect 20791 8676 20795 8732
rect 20731 8672 20795 8676
rect 20811 8732 20875 8736
rect 20811 8676 20815 8732
rect 20815 8676 20871 8732
rect 20871 8676 20875 8732
rect 20811 8672 20875 8676
rect 20891 8732 20955 8736
rect 20891 8676 20895 8732
rect 20895 8676 20951 8732
rect 20951 8676 20955 8732
rect 20891 8672 20955 8676
rect 20971 8732 21035 8736
rect 20971 8676 20975 8732
rect 20975 8676 21031 8732
rect 21031 8676 21035 8732
rect 20971 8672 21035 8676
rect 3424 8188 3488 8192
rect 3424 8132 3428 8188
rect 3428 8132 3484 8188
rect 3484 8132 3488 8188
rect 3424 8128 3488 8132
rect 3504 8188 3568 8192
rect 3504 8132 3508 8188
rect 3508 8132 3564 8188
rect 3564 8132 3568 8188
rect 3504 8128 3568 8132
rect 3584 8188 3648 8192
rect 3584 8132 3588 8188
rect 3588 8132 3644 8188
rect 3644 8132 3648 8188
rect 3584 8128 3648 8132
rect 3664 8188 3728 8192
rect 3664 8132 3668 8188
rect 3668 8132 3724 8188
rect 3724 8132 3728 8188
rect 3664 8128 3728 8132
rect 8369 8188 8433 8192
rect 8369 8132 8373 8188
rect 8373 8132 8429 8188
rect 8429 8132 8433 8188
rect 8369 8128 8433 8132
rect 8449 8188 8513 8192
rect 8449 8132 8453 8188
rect 8453 8132 8509 8188
rect 8509 8132 8513 8188
rect 8449 8128 8513 8132
rect 8529 8188 8593 8192
rect 8529 8132 8533 8188
rect 8533 8132 8589 8188
rect 8589 8132 8593 8188
rect 8529 8128 8593 8132
rect 8609 8188 8673 8192
rect 8609 8132 8613 8188
rect 8613 8132 8669 8188
rect 8669 8132 8673 8188
rect 8609 8128 8673 8132
rect 13314 8188 13378 8192
rect 13314 8132 13318 8188
rect 13318 8132 13374 8188
rect 13374 8132 13378 8188
rect 13314 8128 13378 8132
rect 13394 8188 13458 8192
rect 13394 8132 13398 8188
rect 13398 8132 13454 8188
rect 13454 8132 13458 8188
rect 13394 8128 13458 8132
rect 13474 8188 13538 8192
rect 13474 8132 13478 8188
rect 13478 8132 13534 8188
rect 13534 8132 13538 8188
rect 13474 8128 13538 8132
rect 13554 8188 13618 8192
rect 13554 8132 13558 8188
rect 13558 8132 13614 8188
rect 13614 8132 13618 8188
rect 13554 8128 13618 8132
rect 18259 8188 18323 8192
rect 18259 8132 18263 8188
rect 18263 8132 18319 8188
rect 18319 8132 18323 8188
rect 18259 8128 18323 8132
rect 18339 8188 18403 8192
rect 18339 8132 18343 8188
rect 18343 8132 18399 8188
rect 18399 8132 18403 8188
rect 18339 8128 18403 8132
rect 18419 8188 18483 8192
rect 18419 8132 18423 8188
rect 18423 8132 18479 8188
rect 18479 8132 18483 8188
rect 18419 8128 18483 8132
rect 18499 8188 18563 8192
rect 18499 8132 18503 8188
rect 18503 8132 18559 8188
rect 18559 8132 18563 8188
rect 18499 8128 18563 8132
rect 5896 7644 5960 7648
rect 5896 7588 5900 7644
rect 5900 7588 5956 7644
rect 5956 7588 5960 7644
rect 5896 7584 5960 7588
rect 5976 7644 6040 7648
rect 5976 7588 5980 7644
rect 5980 7588 6036 7644
rect 6036 7588 6040 7644
rect 5976 7584 6040 7588
rect 6056 7644 6120 7648
rect 6056 7588 6060 7644
rect 6060 7588 6116 7644
rect 6116 7588 6120 7644
rect 6056 7584 6120 7588
rect 6136 7644 6200 7648
rect 6136 7588 6140 7644
rect 6140 7588 6196 7644
rect 6196 7588 6200 7644
rect 6136 7584 6200 7588
rect 10841 7644 10905 7648
rect 10841 7588 10845 7644
rect 10845 7588 10901 7644
rect 10901 7588 10905 7644
rect 10841 7584 10905 7588
rect 10921 7644 10985 7648
rect 10921 7588 10925 7644
rect 10925 7588 10981 7644
rect 10981 7588 10985 7644
rect 10921 7584 10985 7588
rect 11001 7644 11065 7648
rect 11001 7588 11005 7644
rect 11005 7588 11061 7644
rect 11061 7588 11065 7644
rect 11001 7584 11065 7588
rect 11081 7644 11145 7648
rect 11081 7588 11085 7644
rect 11085 7588 11141 7644
rect 11141 7588 11145 7644
rect 11081 7584 11145 7588
rect 15786 7644 15850 7648
rect 15786 7588 15790 7644
rect 15790 7588 15846 7644
rect 15846 7588 15850 7644
rect 15786 7584 15850 7588
rect 15866 7644 15930 7648
rect 15866 7588 15870 7644
rect 15870 7588 15926 7644
rect 15926 7588 15930 7644
rect 15866 7584 15930 7588
rect 15946 7644 16010 7648
rect 15946 7588 15950 7644
rect 15950 7588 16006 7644
rect 16006 7588 16010 7644
rect 15946 7584 16010 7588
rect 16026 7644 16090 7648
rect 16026 7588 16030 7644
rect 16030 7588 16086 7644
rect 16086 7588 16090 7644
rect 16026 7584 16090 7588
rect 20731 7644 20795 7648
rect 20731 7588 20735 7644
rect 20735 7588 20791 7644
rect 20791 7588 20795 7644
rect 20731 7584 20795 7588
rect 20811 7644 20875 7648
rect 20811 7588 20815 7644
rect 20815 7588 20871 7644
rect 20871 7588 20875 7644
rect 20811 7584 20875 7588
rect 20891 7644 20955 7648
rect 20891 7588 20895 7644
rect 20895 7588 20951 7644
rect 20951 7588 20955 7644
rect 20891 7584 20955 7588
rect 20971 7644 21035 7648
rect 20971 7588 20975 7644
rect 20975 7588 21031 7644
rect 21031 7588 21035 7644
rect 20971 7584 21035 7588
rect 3424 7100 3488 7104
rect 3424 7044 3428 7100
rect 3428 7044 3484 7100
rect 3484 7044 3488 7100
rect 3424 7040 3488 7044
rect 3504 7100 3568 7104
rect 3504 7044 3508 7100
rect 3508 7044 3564 7100
rect 3564 7044 3568 7100
rect 3504 7040 3568 7044
rect 3584 7100 3648 7104
rect 3584 7044 3588 7100
rect 3588 7044 3644 7100
rect 3644 7044 3648 7100
rect 3584 7040 3648 7044
rect 3664 7100 3728 7104
rect 3664 7044 3668 7100
rect 3668 7044 3724 7100
rect 3724 7044 3728 7100
rect 3664 7040 3728 7044
rect 8369 7100 8433 7104
rect 8369 7044 8373 7100
rect 8373 7044 8429 7100
rect 8429 7044 8433 7100
rect 8369 7040 8433 7044
rect 8449 7100 8513 7104
rect 8449 7044 8453 7100
rect 8453 7044 8509 7100
rect 8509 7044 8513 7100
rect 8449 7040 8513 7044
rect 8529 7100 8593 7104
rect 8529 7044 8533 7100
rect 8533 7044 8589 7100
rect 8589 7044 8593 7100
rect 8529 7040 8593 7044
rect 8609 7100 8673 7104
rect 8609 7044 8613 7100
rect 8613 7044 8669 7100
rect 8669 7044 8673 7100
rect 8609 7040 8673 7044
rect 13314 7100 13378 7104
rect 13314 7044 13318 7100
rect 13318 7044 13374 7100
rect 13374 7044 13378 7100
rect 13314 7040 13378 7044
rect 13394 7100 13458 7104
rect 13394 7044 13398 7100
rect 13398 7044 13454 7100
rect 13454 7044 13458 7100
rect 13394 7040 13458 7044
rect 13474 7100 13538 7104
rect 13474 7044 13478 7100
rect 13478 7044 13534 7100
rect 13534 7044 13538 7100
rect 13474 7040 13538 7044
rect 13554 7100 13618 7104
rect 13554 7044 13558 7100
rect 13558 7044 13614 7100
rect 13614 7044 13618 7100
rect 13554 7040 13618 7044
rect 18259 7100 18323 7104
rect 18259 7044 18263 7100
rect 18263 7044 18319 7100
rect 18319 7044 18323 7100
rect 18259 7040 18323 7044
rect 18339 7100 18403 7104
rect 18339 7044 18343 7100
rect 18343 7044 18399 7100
rect 18399 7044 18403 7100
rect 18339 7040 18403 7044
rect 18419 7100 18483 7104
rect 18419 7044 18423 7100
rect 18423 7044 18479 7100
rect 18479 7044 18483 7100
rect 18419 7040 18483 7044
rect 18499 7100 18563 7104
rect 18499 7044 18503 7100
rect 18503 7044 18559 7100
rect 18559 7044 18563 7100
rect 18499 7040 18563 7044
rect 5896 6556 5960 6560
rect 5896 6500 5900 6556
rect 5900 6500 5956 6556
rect 5956 6500 5960 6556
rect 5896 6496 5960 6500
rect 5976 6556 6040 6560
rect 5976 6500 5980 6556
rect 5980 6500 6036 6556
rect 6036 6500 6040 6556
rect 5976 6496 6040 6500
rect 6056 6556 6120 6560
rect 6056 6500 6060 6556
rect 6060 6500 6116 6556
rect 6116 6500 6120 6556
rect 6056 6496 6120 6500
rect 6136 6556 6200 6560
rect 6136 6500 6140 6556
rect 6140 6500 6196 6556
rect 6196 6500 6200 6556
rect 6136 6496 6200 6500
rect 10841 6556 10905 6560
rect 10841 6500 10845 6556
rect 10845 6500 10901 6556
rect 10901 6500 10905 6556
rect 10841 6496 10905 6500
rect 10921 6556 10985 6560
rect 10921 6500 10925 6556
rect 10925 6500 10981 6556
rect 10981 6500 10985 6556
rect 10921 6496 10985 6500
rect 11001 6556 11065 6560
rect 11001 6500 11005 6556
rect 11005 6500 11061 6556
rect 11061 6500 11065 6556
rect 11001 6496 11065 6500
rect 11081 6556 11145 6560
rect 11081 6500 11085 6556
rect 11085 6500 11141 6556
rect 11141 6500 11145 6556
rect 11081 6496 11145 6500
rect 15786 6556 15850 6560
rect 15786 6500 15790 6556
rect 15790 6500 15846 6556
rect 15846 6500 15850 6556
rect 15786 6496 15850 6500
rect 15866 6556 15930 6560
rect 15866 6500 15870 6556
rect 15870 6500 15926 6556
rect 15926 6500 15930 6556
rect 15866 6496 15930 6500
rect 15946 6556 16010 6560
rect 15946 6500 15950 6556
rect 15950 6500 16006 6556
rect 16006 6500 16010 6556
rect 15946 6496 16010 6500
rect 16026 6556 16090 6560
rect 16026 6500 16030 6556
rect 16030 6500 16086 6556
rect 16086 6500 16090 6556
rect 16026 6496 16090 6500
rect 20731 6556 20795 6560
rect 20731 6500 20735 6556
rect 20735 6500 20791 6556
rect 20791 6500 20795 6556
rect 20731 6496 20795 6500
rect 20811 6556 20875 6560
rect 20811 6500 20815 6556
rect 20815 6500 20871 6556
rect 20871 6500 20875 6556
rect 20811 6496 20875 6500
rect 20891 6556 20955 6560
rect 20891 6500 20895 6556
rect 20895 6500 20951 6556
rect 20951 6500 20955 6556
rect 20891 6496 20955 6500
rect 20971 6556 21035 6560
rect 20971 6500 20975 6556
rect 20975 6500 21031 6556
rect 21031 6500 21035 6556
rect 20971 6496 21035 6500
rect 3424 6012 3488 6016
rect 3424 5956 3428 6012
rect 3428 5956 3484 6012
rect 3484 5956 3488 6012
rect 3424 5952 3488 5956
rect 3504 6012 3568 6016
rect 3504 5956 3508 6012
rect 3508 5956 3564 6012
rect 3564 5956 3568 6012
rect 3504 5952 3568 5956
rect 3584 6012 3648 6016
rect 3584 5956 3588 6012
rect 3588 5956 3644 6012
rect 3644 5956 3648 6012
rect 3584 5952 3648 5956
rect 3664 6012 3728 6016
rect 3664 5956 3668 6012
rect 3668 5956 3724 6012
rect 3724 5956 3728 6012
rect 3664 5952 3728 5956
rect 8369 6012 8433 6016
rect 8369 5956 8373 6012
rect 8373 5956 8429 6012
rect 8429 5956 8433 6012
rect 8369 5952 8433 5956
rect 8449 6012 8513 6016
rect 8449 5956 8453 6012
rect 8453 5956 8509 6012
rect 8509 5956 8513 6012
rect 8449 5952 8513 5956
rect 8529 6012 8593 6016
rect 8529 5956 8533 6012
rect 8533 5956 8589 6012
rect 8589 5956 8593 6012
rect 8529 5952 8593 5956
rect 8609 6012 8673 6016
rect 8609 5956 8613 6012
rect 8613 5956 8669 6012
rect 8669 5956 8673 6012
rect 8609 5952 8673 5956
rect 13314 6012 13378 6016
rect 13314 5956 13318 6012
rect 13318 5956 13374 6012
rect 13374 5956 13378 6012
rect 13314 5952 13378 5956
rect 13394 6012 13458 6016
rect 13394 5956 13398 6012
rect 13398 5956 13454 6012
rect 13454 5956 13458 6012
rect 13394 5952 13458 5956
rect 13474 6012 13538 6016
rect 13474 5956 13478 6012
rect 13478 5956 13534 6012
rect 13534 5956 13538 6012
rect 13474 5952 13538 5956
rect 13554 6012 13618 6016
rect 13554 5956 13558 6012
rect 13558 5956 13614 6012
rect 13614 5956 13618 6012
rect 13554 5952 13618 5956
rect 18259 6012 18323 6016
rect 18259 5956 18263 6012
rect 18263 5956 18319 6012
rect 18319 5956 18323 6012
rect 18259 5952 18323 5956
rect 18339 6012 18403 6016
rect 18339 5956 18343 6012
rect 18343 5956 18399 6012
rect 18399 5956 18403 6012
rect 18339 5952 18403 5956
rect 18419 6012 18483 6016
rect 18419 5956 18423 6012
rect 18423 5956 18479 6012
rect 18479 5956 18483 6012
rect 18419 5952 18483 5956
rect 18499 6012 18563 6016
rect 18499 5956 18503 6012
rect 18503 5956 18559 6012
rect 18559 5956 18563 6012
rect 18499 5952 18563 5956
rect 5896 5468 5960 5472
rect 5896 5412 5900 5468
rect 5900 5412 5956 5468
rect 5956 5412 5960 5468
rect 5896 5408 5960 5412
rect 5976 5468 6040 5472
rect 5976 5412 5980 5468
rect 5980 5412 6036 5468
rect 6036 5412 6040 5468
rect 5976 5408 6040 5412
rect 6056 5468 6120 5472
rect 6056 5412 6060 5468
rect 6060 5412 6116 5468
rect 6116 5412 6120 5468
rect 6056 5408 6120 5412
rect 6136 5468 6200 5472
rect 6136 5412 6140 5468
rect 6140 5412 6196 5468
rect 6196 5412 6200 5468
rect 6136 5408 6200 5412
rect 10841 5468 10905 5472
rect 10841 5412 10845 5468
rect 10845 5412 10901 5468
rect 10901 5412 10905 5468
rect 10841 5408 10905 5412
rect 10921 5468 10985 5472
rect 10921 5412 10925 5468
rect 10925 5412 10981 5468
rect 10981 5412 10985 5468
rect 10921 5408 10985 5412
rect 11001 5468 11065 5472
rect 11001 5412 11005 5468
rect 11005 5412 11061 5468
rect 11061 5412 11065 5468
rect 11001 5408 11065 5412
rect 11081 5468 11145 5472
rect 11081 5412 11085 5468
rect 11085 5412 11141 5468
rect 11141 5412 11145 5468
rect 11081 5408 11145 5412
rect 15786 5468 15850 5472
rect 15786 5412 15790 5468
rect 15790 5412 15846 5468
rect 15846 5412 15850 5468
rect 15786 5408 15850 5412
rect 15866 5468 15930 5472
rect 15866 5412 15870 5468
rect 15870 5412 15926 5468
rect 15926 5412 15930 5468
rect 15866 5408 15930 5412
rect 15946 5468 16010 5472
rect 15946 5412 15950 5468
rect 15950 5412 16006 5468
rect 16006 5412 16010 5468
rect 15946 5408 16010 5412
rect 16026 5468 16090 5472
rect 16026 5412 16030 5468
rect 16030 5412 16086 5468
rect 16086 5412 16090 5468
rect 16026 5408 16090 5412
rect 20731 5468 20795 5472
rect 20731 5412 20735 5468
rect 20735 5412 20791 5468
rect 20791 5412 20795 5468
rect 20731 5408 20795 5412
rect 20811 5468 20875 5472
rect 20811 5412 20815 5468
rect 20815 5412 20871 5468
rect 20871 5412 20875 5468
rect 20811 5408 20875 5412
rect 20891 5468 20955 5472
rect 20891 5412 20895 5468
rect 20895 5412 20951 5468
rect 20951 5412 20955 5468
rect 20891 5408 20955 5412
rect 20971 5468 21035 5472
rect 20971 5412 20975 5468
rect 20975 5412 21031 5468
rect 21031 5412 21035 5468
rect 20971 5408 21035 5412
rect 3424 4924 3488 4928
rect 3424 4868 3428 4924
rect 3428 4868 3484 4924
rect 3484 4868 3488 4924
rect 3424 4864 3488 4868
rect 3504 4924 3568 4928
rect 3504 4868 3508 4924
rect 3508 4868 3564 4924
rect 3564 4868 3568 4924
rect 3504 4864 3568 4868
rect 3584 4924 3648 4928
rect 3584 4868 3588 4924
rect 3588 4868 3644 4924
rect 3644 4868 3648 4924
rect 3584 4864 3648 4868
rect 3664 4924 3728 4928
rect 3664 4868 3668 4924
rect 3668 4868 3724 4924
rect 3724 4868 3728 4924
rect 3664 4864 3728 4868
rect 8369 4924 8433 4928
rect 8369 4868 8373 4924
rect 8373 4868 8429 4924
rect 8429 4868 8433 4924
rect 8369 4864 8433 4868
rect 8449 4924 8513 4928
rect 8449 4868 8453 4924
rect 8453 4868 8509 4924
rect 8509 4868 8513 4924
rect 8449 4864 8513 4868
rect 8529 4924 8593 4928
rect 8529 4868 8533 4924
rect 8533 4868 8589 4924
rect 8589 4868 8593 4924
rect 8529 4864 8593 4868
rect 8609 4924 8673 4928
rect 8609 4868 8613 4924
rect 8613 4868 8669 4924
rect 8669 4868 8673 4924
rect 8609 4864 8673 4868
rect 13314 4924 13378 4928
rect 13314 4868 13318 4924
rect 13318 4868 13374 4924
rect 13374 4868 13378 4924
rect 13314 4864 13378 4868
rect 13394 4924 13458 4928
rect 13394 4868 13398 4924
rect 13398 4868 13454 4924
rect 13454 4868 13458 4924
rect 13394 4864 13458 4868
rect 13474 4924 13538 4928
rect 13474 4868 13478 4924
rect 13478 4868 13534 4924
rect 13534 4868 13538 4924
rect 13474 4864 13538 4868
rect 13554 4924 13618 4928
rect 13554 4868 13558 4924
rect 13558 4868 13614 4924
rect 13614 4868 13618 4924
rect 13554 4864 13618 4868
rect 18259 4924 18323 4928
rect 18259 4868 18263 4924
rect 18263 4868 18319 4924
rect 18319 4868 18323 4924
rect 18259 4864 18323 4868
rect 18339 4924 18403 4928
rect 18339 4868 18343 4924
rect 18343 4868 18399 4924
rect 18399 4868 18403 4924
rect 18339 4864 18403 4868
rect 18419 4924 18483 4928
rect 18419 4868 18423 4924
rect 18423 4868 18479 4924
rect 18479 4868 18483 4924
rect 18419 4864 18483 4868
rect 18499 4924 18563 4928
rect 18499 4868 18503 4924
rect 18503 4868 18559 4924
rect 18559 4868 18563 4924
rect 18499 4864 18563 4868
rect 5896 4380 5960 4384
rect 5896 4324 5900 4380
rect 5900 4324 5956 4380
rect 5956 4324 5960 4380
rect 5896 4320 5960 4324
rect 5976 4380 6040 4384
rect 5976 4324 5980 4380
rect 5980 4324 6036 4380
rect 6036 4324 6040 4380
rect 5976 4320 6040 4324
rect 6056 4380 6120 4384
rect 6056 4324 6060 4380
rect 6060 4324 6116 4380
rect 6116 4324 6120 4380
rect 6056 4320 6120 4324
rect 6136 4380 6200 4384
rect 6136 4324 6140 4380
rect 6140 4324 6196 4380
rect 6196 4324 6200 4380
rect 6136 4320 6200 4324
rect 10841 4380 10905 4384
rect 10841 4324 10845 4380
rect 10845 4324 10901 4380
rect 10901 4324 10905 4380
rect 10841 4320 10905 4324
rect 10921 4380 10985 4384
rect 10921 4324 10925 4380
rect 10925 4324 10981 4380
rect 10981 4324 10985 4380
rect 10921 4320 10985 4324
rect 11001 4380 11065 4384
rect 11001 4324 11005 4380
rect 11005 4324 11061 4380
rect 11061 4324 11065 4380
rect 11001 4320 11065 4324
rect 11081 4380 11145 4384
rect 11081 4324 11085 4380
rect 11085 4324 11141 4380
rect 11141 4324 11145 4380
rect 11081 4320 11145 4324
rect 15786 4380 15850 4384
rect 15786 4324 15790 4380
rect 15790 4324 15846 4380
rect 15846 4324 15850 4380
rect 15786 4320 15850 4324
rect 15866 4380 15930 4384
rect 15866 4324 15870 4380
rect 15870 4324 15926 4380
rect 15926 4324 15930 4380
rect 15866 4320 15930 4324
rect 15946 4380 16010 4384
rect 15946 4324 15950 4380
rect 15950 4324 16006 4380
rect 16006 4324 16010 4380
rect 15946 4320 16010 4324
rect 16026 4380 16090 4384
rect 16026 4324 16030 4380
rect 16030 4324 16086 4380
rect 16086 4324 16090 4380
rect 16026 4320 16090 4324
rect 20731 4380 20795 4384
rect 20731 4324 20735 4380
rect 20735 4324 20791 4380
rect 20791 4324 20795 4380
rect 20731 4320 20795 4324
rect 20811 4380 20875 4384
rect 20811 4324 20815 4380
rect 20815 4324 20871 4380
rect 20871 4324 20875 4380
rect 20811 4320 20875 4324
rect 20891 4380 20955 4384
rect 20891 4324 20895 4380
rect 20895 4324 20951 4380
rect 20951 4324 20955 4380
rect 20891 4320 20955 4324
rect 20971 4380 21035 4384
rect 20971 4324 20975 4380
rect 20975 4324 21031 4380
rect 21031 4324 21035 4380
rect 20971 4320 21035 4324
rect 3424 3836 3488 3840
rect 3424 3780 3428 3836
rect 3428 3780 3484 3836
rect 3484 3780 3488 3836
rect 3424 3776 3488 3780
rect 3504 3836 3568 3840
rect 3504 3780 3508 3836
rect 3508 3780 3564 3836
rect 3564 3780 3568 3836
rect 3504 3776 3568 3780
rect 3584 3836 3648 3840
rect 3584 3780 3588 3836
rect 3588 3780 3644 3836
rect 3644 3780 3648 3836
rect 3584 3776 3648 3780
rect 3664 3836 3728 3840
rect 3664 3780 3668 3836
rect 3668 3780 3724 3836
rect 3724 3780 3728 3836
rect 3664 3776 3728 3780
rect 8369 3836 8433 3840
rect 8369 3780 8373 3836
rect 8373 3780 8429 3836
rect 8429 3780 8433 3836
rect 8369 3776 8433 3780
rect 8449 3836 8513 3840
rect 8449 3780 8453 3836
rect 8453 3780 8509 3836
rect 8509 3780 8513 3836
rect 8449 3776 8513 3780
rect 8529 3836 8593 3840
rect 8529 3780 8533 3836
rect 8533 3780 8589 3836
rect 8589 3780 8593 3836
rect 8529 3776 8593 3780
rect 8609 3836 8673 3840
rect 8609 3780 8613 3836
rect 8613 3780 8669 3836
rect 8669 3780 8673 3836
rect 8609 3776 8673 3780
rect 13314 3836 13378 3840
rect 13314 3780 13318 3836
rect 13318 3780 13374 3836
rect 13374 3780 13378 3836
rect 13314 3776 13378 3780
rect 13394 3836 13458 3840
rect 13394 3780 13398 3836
rect 13398 3780 13454 3836
rect 13454 3780 13458 3836
rect 13394 3776 13458 3780
rect 13474 3836 13538 3840
rect 13474 3780 13478 3836
rect 13478 3780 13534 3836
rect 13534 3780 13538 3836
rect 13474 3776 13538 3780
rect 13554 3836 13618 3840
rect 13554 3780 13558 3836
rect 13558 3780 13614 3836
rect 13614 3780 13618 3836
rect 13554 3776 13618 3780
rect 18259 3836 18323 3840
rect 18259 3780 18263 3836
rect 18263 3780 18319 3836
rect 18319 3780 18323 3836
rect 18259 3776 18323 3780
rect 18339 3836 18403 3840
rect 18339 3780 18343 3836
rect 18343 3780 18399 3836
rect 18399 3780 18403 3836
rect 18339 3776 18403 3780
rect 18419 3836 18483 3840
rect 18419 3780 18423 3836
rect 18423 3780 18479 3836
rect 18479 3780 18483 3836
rect 18419 3776 18483 3780
rect 18499 3836 18563 3840
rect 18499 3780 18503 3836
rect 18503 3780 18559 3836
rect 18559 3780 18563 3836
rect 18499 3776 18563 3780
rect 5896 3292 5960 3296
rect 5896 3236 5900 3292
rect 5900 3236 5956 3292
rect 5956 3236 5960 3292
rect 5896 3232 5960 3236
rect 5976 3292 6040 3296
rect 5976 3236 5980 3292
rect 5980 3236 6036 3292
rect 6036 3236 6040 3292
rect 5976 3232 6040 3236
rect 6056 3292 6120 3296
rect 6056 3236 6060 3292
rect 6060 3236 6116 3292
rect 6116 3236 6120 3292
rect 6056 3232 6120 3236
rect 6136 3292 6200 3296
rect 6136 3236 6140 3292
rect 6140 3236 6196 3292
rect 6196 3236 6200 3292
rect 6136 3232 6200 3236
rect 10841 3292 10905 3296
rect 10841 3236 10845 3292
rect 10845 3236 10901 3292
rect 10901 3236 10905 3292
rect 10841 3232 10905 3236
rect 10921 3292 10985 3296
rect 10921 3236 10925 3292
rect 10925 3236 10981 3292
rect 10981 3236 10985 3292
rect 10921 3232 10985 3236
rect 11001 3292 11065 3296
rect 11001 3236 11005 3292
rect 11005 3236 11061 3292
rect 11061 3236 11065 3292
rect 11001 3232 11065 3236
rect 11081 3292 11145 3296
rect 11081 3236 11085 3292
rect 11085 3236 11141 3292
rect 11141 3236 11145 3292
rect 11081 3232 11145 3236
rect 15786 3292 15850 3296
rect 15786 3236 15790 3292
rect 15790 3236 15846 3292
rect 15846 3236 15850 3292
rect 15786 3232 15850 3236
rect 15866 3292 15930 3296
rect 15866 3236 15870 3292
rect 15870 3236 15926 3292
rect 15926 3236 15930 3292
rect 15866 3232 15930 3236
rect 15946 3292 16010 3296
rect 15946 3236 15950 3292
rect 15950 3236 16006 3292
rect 16006 3236 16010 3292
rect 15946 3232 16010 3236
rect 16026 3292 16090 3296
rect 16026 3236 16030 3292
rect 16030 3236 16086 3292
rect 16086 3236 16090 3292
rect 16026 3232 16090 3236
rect 20731 3292 20795 3296
rect 20731 3236 20735 3292
rect 20735 3236 20791 3292
rect 20791 3236 20795 3292
rect 20731 3232 20795 3236
rect 20811 3292 20875 3296
rect 20811 3236 20815 3292
rect 20815 3236 20871 3292
rect 20871 3236 20875 3292
rect 20811 3232 20875 3236
rect 20891 3292 20955 3296
rect 20891 3236 20895 3292
rect 20895 3236 20951 3292
rect 20951 3236 20955 3292
rect 20891 3232 20955 3236
rect 20971 3292 21035 3296
rect 20971 3236 20975 3292
rect 20975 3236 21031 3292
rect 21031 3236 21035 3292
rect 20971 3232 21035 3236
rect 3424 2748 3488 2752
rect 3424 2692 3428 2748
rect 3428 2692 3484 2748
rect 3484 2692 3488 2748
rect 3424 2688 3488 2692
rect 3504 2748 3568 2752
rect 3504 2692 3508 2748
rect 3508 2692 3564 2748
rect 3564 2692 3568 2748
rect 3504 2688 3568 2692
rect 3584 2748 3648 2752
rect 3584 2692 3588 2748
rect 3588 2692 3644 2748
rect 3644 2692 3648 2748
rect 3584 2688 3648 2692
rect 3664 2748 3728 2752
rect 3664 2692 3668 2748
rect 3668 2692 3724 2748
rect 3724 2692 3728 2748
rect 3664 2688 3728 2692
rect 8369 2748 8433 2752
rect 8369 2692 8373 2748
rect 8373 2692 8429 2748
rect 8429 2692 8433 2748
rect 8369 2688 8433 2692
rect 8449 2748 8513 2752
rect 8449 2692 8453 2748
rect 8453 2692 8509 2748
rect 8509 2692 8513 2748
rect 8449 2688 8513 2692
rect 8529 2748 8593 2752
rect 8529 2692 8533 2748
rect 8533 2692 8589 2748
rect 8589 2692 8593 2748
rect 8529 2688 8593 2692
rect 8609 2748 8673 2752
rect 8609 2692 8613 2748
rect 8613 2692 8669 2748
rect 8669 2692 8673 2748
rect 8609 2688 8673 2692
rect 13314 2748 13378 2752
rect 13314 2692 13318 2748
rect 13318 2692 13374 2748
rect 13374 2692 13378 2748
rect 13314 2688 13378 2692
rect 13394 2748 13458 2752
rect 13394 2692 13398 2748
rect 13398 2692 13454 2748
rect 13454 2692 13458 2748
rect 13394 2688 13458 2692
rect 13474 2748 13538 2752
rect 13474 2692 13478 2748
rect 13478 2692 13534 2748
rect 13534 2692 13538 2748
rect 13474 2688 13538 2692
rect 13554 2748 13618 2752
rect 13554 2692 13558 2748
rect 13558 2692 13614 2748
rect 13614 2692 13618 2748
rect 13554 2688 13618 2692
rect 18259 2748 18323 2752
rect 18259 2692 18263 2748
rect 18263 2692 18319 2748
rect 18319 2692 18323 2748
rect 18259 2688 18323 2692
rect 18339 2748 18403 2752
rect 18339 2692 18343 2748
rect 18343 2692 18399 2748
rect 18399 2692 18403 2748
rect 18339 2688 18403 2692
rect 18419 2748 18483 2752
rect 18419 2692 18423 2748
rect 18423 2692 18479 2748
rect 18479 2692 18483 2748
rect 18419 2688 18483 2692
rect 18499 2748 18563 2752
rect 18499 2692 18503 2748
rect 18503 2692 18559 2748
rect 18559 2692 18563 2748
rect 18499 2688 18563 2692
rect 5896 2204 5960 2208
rect 5896 2148 5900 2204
rect 5900 2148 5956 2204
rect 5956 2148 5960 2204
rect 5896 2144 5960 2148
rect 5976 2204 6040 2208
rect 5976 2148 5980 2204
rect 5980 2148 6036 2204
rect 6036 2148 6040 2204
rect 5976 2144 6040 2148
rect 6056 2204 6120 2208
rect 6056 2148 6060 2204
rect 6060 2148 6116 2204
rect 6116 2148 6120 2204
rect 6056 2144 6120 2148
rect 6136 2204 6200 2208
rect 6136 2148 6140 2204
rect 6140 2148 6196 2204
rect 6196 2148 6200 2204
rect 6136 2144 6200 2148
rect 10841 2204 10905 2208
rect 10841 2148 10845 2204
rect 10845 2148 10901 2204
rect 10901 2148 10905 2204
rect 10841 2144 10905 2148
rect 10921 2204 10985 2208
rect 10921 2148 10925 2204
rect 10925 2148 10981 2204
rect 10981 2148 10985 2204
rect 10921 2144 10985 2148
rect 11001 2204 11065 2208
rect 11001 2148 11005 2204
rect 11005 2148 11061 2204
rect 11061 2148 11065 2204
rect 11001 2144 11065 2148
rect 11081 2204 11145 2208
rect 11081 2148 11085 2204
rect 11085 2148 11141 2204
rect 11141 2148 11145 2204
rect 11081 2144 11145 2148
rect 15786 2204 15850 2208
rect 15786 2148 15790 2204
rect 15790 2148 15846 2204
rect 15846 2148 15850 2204
rect 15786 2144 15850 2148
rect 15866 2204 15930 2208
rect 15866 2148 15870 2204
rect 15870 2148 15926 2204
rect 15926 2148 15930 2204
rect 15866 2144 15930 2148
rect 15946 2204 16010 2208
rect 15946 2148 15950 2204
rect 15950 2148 16006 2204
rect 16006 2148 16010 2204
rect 15946 2144 16010 2148
rect 16026 2204 16090 2208
rect 16026 2148 16030 2204
rect 16030 2148 16086 2204
rect 16086 2148 16090 2204
rect 16026 2144 16090 2148
rect 20731 2204 20795 2208
rect 20731 2148 20735 2204
rect 20735 2148 20791 2204
rect 20791 2148 20795 2204
rect 20731 2144 20795 2148
rect 20811 2204 20875 2208
rect 20811 2148 20815 2204
rect 20815 2148 20871 2204
rect 20871 2148 20875 2204
rect 20811 2144 20875 2148
rect 20891 2204 20955 2208
rect 20891 2148 20895 2204
rect 20895 2148 20951 2204
rect 20951 2148 20955 2204
rect 20891 2144 20955 2148
rect 20971 2204 21035 2208
rect 20971 2148 20975 2204
rect 20975 2148 21031 2204
rect 21031 2148 21035 2204
rect 20971 2144 21035 2148
<< metal4 >>
rect 3416 19072 3736 19632
rect 3416 19008 3424 19072
rect 3488 19008 3504 19072
rect 3568 19008 3584 19072
rect 3648 19008 3664 19072
rect 3728 19008 3736 19072
rect 3416 17984 3736 19008
rect 3416 17920 3424 17984
rect 3488 17920 3504 17984
rect 3568 17920 3584 17984
rect 3648 17920 3664 17984
rect 3728 17920 3736 17984
rect 3416 16896 3736 17920
rect 3416 16832 3424 16896
rect 3488 16832 3504 16896
rect 3568 16832 3584 16896
rect 3648 16832 3664 16896
rect 3728 16832 3736 16896
rect 3416 15808 3736 16832
rect 3416 15744 3424 15808
rect 3488 15744 3504 15808
rect 3568 15744 3584 15808
rect 3648 15744 3664 15808
rect 3728 15744 3736 15808
rect 3416 14720 3736 15744
rect 3416 14656 3424 14720
rect 3488 14656 3504 14720
rect 3568 14656 3584 14720
rect 3648 14656 3664 14720
rect 3728 14656 3736 14720
rect 3416 13632 3736 14656
rect 3416 13568 3424 13632
rect 3488 13568 3504 13632
rect 3568 13568 3584 13632
rect 3648 13568 3664 13632
rect 3728 13568 3736 13632
rect 3416 12544 3736 13568
rect 3416 12480 3424 12544
rect 3488 12480 3504 12544
rect 3568 12480 3584 12544
rect 3648 12480 3664 12544
rect 3728 12480 3736 12544
rect 3416 11456 3736 12480
rect 3416 11392 3424 11456
rect 3488 11392 3504 11456
rect 3568 11392 3584 11456
rect 3648 11392 3664 11456
rect 3728 11392 3736 11456
rect 3416 10368 3736 11392
rect 3416 10304 3424 10368
rect 3488 10304 3504 10368
rect 3568 10304 3584 10368
rect 3648 10304 3664 10368
rect 3728 10304 3736 10368
rect 3416 9280 3736 10304
rect 3416 9216 3424 9280
rect 3488 9216 3504 9280
rect 3568 9216 3584 9280
rect 3648 9216 3664 9280
rect 3728 9216 3736 9280
rect 3416 8192 3736 9216
rect 3416 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3584 8192
rect 3648 8128 3664 8192
rect 3728 8128 3736 8192
rect 3416 7104 3736 8128
rect 3416 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3584 7104
rect 3648 7040 3664 7104
rect 3728 7040 3736 7104
rect 3416 6016 3736 7040
rect 3416 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3584 6016
rect 3648 5952 3664 6016
rect 3728 5952 3736 6016
rect 3416 4928 3736 5952
rect 3416 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3584 4928
rect 3648 4864 3664 4928
rect 3728 4864 3736 4928
rect 3416 3840 3736 4864
rect 3416 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3584 3840
rect 3648 3776 3664 3840
rect 3728 3776 3736 3840
rect 3416 2752 3736 3776
rect 3416 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3584 2752
rect 3648 2688 3664 2752
rect 3728 2688 3736 2752
rect 3416 2128 3736 2688
rect 5888 19616 6208 19632
rect 5888 19552 5896 19616
rect 5960 19552 5976 19616
rect 6040 19552 6056 19616
rect 6120 19552 6136 19616
rect 6200 19552 6208 19616
rect 5888 18528 6208 19552
rect 5888 18464 5896 18528
rect 5960 18464 5976 18528
rect 6040 18464 6056 18528
rect 6120 18464 6136 18528
rect 6200 18464 6208 18528
rect 5888 17440 6208 18464
rect 5888 17376 5896 17440
rect 5960 17376 5976 17440
rect 6040 17376 6056 17440
rect 6120 17376 6136 17440
rect 6200 17376 6208 17440
rect 5888 16352 6208 17376
rect 5888 16288 5896 16352
rect 5960 16288 5976 16352
rect 6040 16288 6056 16352
rect 6120 16288 6136 16352
rect 6200 16288 6208 16352
rect 5888 15264 6208 16288
rect 5888 15200 5896 15264
rect 5960 15200 5976 15264
rect 6040 15200 6056 15264
rect 6120 15200 6136 15264
rect 6200 15200 6208 15264
rect 5888 14176 6208 15200
rect 5888 14112 5896 14176
rect 5960 14112 5976 14176
rect 6040 14112 6056 14176
rect 6120 14112 6136 14176
rect 6200 14112 6208 14176
rect 5888 13088 6208 14112
rect 5888 13024 5896 13088
rect 5960 13024 5976 13088
rect 6040 13024 6056 13088
rect 6120 13024 6136 13088
rect 6200 13024 6208 13088
rect 5888 12000 6208 13024
rect 5888 11936 5896 12000
rect 5960 11936 5976 12000
rect 6040 11936 6056 12000
rect 6120 11936 6136 12000
rect 6200 11936 6208 12000
rect 5888 10912 6208 11936
rect 5888 10848 5896 10912
rect 5960 10848 5976 10912
rect 6040 10848 6056 10912
rect 6120 10848 6136 10912
rect 6200 10848 6208 10912
rect 5888 9824 6208 10848
rect 5888 9760 5896 9824
rect 5960 9760 5976 9824
rect 6040 9760 6056 9824
rect 6120 9760 6136 9824
rect 6200 9760 6208 9824
rect 5888 8736 6208 9760
rect 5888 8672 5896 8736
rect 5960 8672 5976 8736
rect 6040 8672 6056 8736
rect 6120 8672 6136 8736
rect 6200 8672 6208 8736
rect 5888 7648 6208 8672
rect 5888 7584 5896 7648
rect 5960 7584 5976 7648
rect 6040 7584 6056 7648
rect 6120 7584 6136 7648
rect 6200 7584 6208 7648
rect 5888 6560 6208 7584
rect 5888 6496 5896 6560
rect 5960 6496 5976 6560
rect 6040 6496 6056 6560
rect 6120 6496 6136 6560
rect 6200 6496 6208 6560
rect 5888 5472 6208 6496
rect 5888 5408 5896 5472
rect 5960 5408 5976 5472
rect 6040 5408 6056 5472
rect 6120 5408 6136 5472
rect 6200 5408 6208 5472
rect 5888 4384 6208 5408
rect 5888 4320 5896 4384
rect 5960 4320 5976 4384
rect 6040 4320 6056 4384
rect 6120 4320 6136 4384
rect 6200 4320 6208 4384
rect 5888 3296 6208 4320
rect 5888 3232 5896 3296
rect 5960 3232 5976 3296
rect 6040 3232 6056 3296
rect 6120 3232 6136 3296
rect 6200 3232 6208 3296
rect 5888 2208 6208 3232
rect 5888 2144 5896 2208
rect 5960 2144 5976 2208
rect 6040 2144 6056 2208
rect 6120 2144 6136 2208
rect 6200 2144 6208 2208
rect 5888 2128 6208 2144
rect 8361 19072 8681 19632
rect 8361 19008 8369 19072
rect 8433 19008 8449 19072
rect 8513 19008 8529 19072
rect 8593 19008 8609 19072
rect 8673 19008 8681 19072
rect 8361 17984 8681 19008
rect 8361 17920 8369 17984
rect 8433 17920 8449 17984
rect 8513 17920 8529 17984
rect 8593 17920 8609 17984
rect 8673 17920 8681 17984
rect 8361 16896 8681 17920
rect 8361 16832 8369 16896
rect 8433 16832 8449 16896
rect 8513 16832 8529 16896
rect 8593 16832 8609 16896
rect 8673 16832 8681 16896
rect 8361 15808 8681 16832
rect 8361 15744 8369 15808
rect 8433 15744 8449 15808
rect 8513 15744 8529 15808
rect 8593 15744 8609 15808
rect 8673 15744 8681 15808
rect 8361 14720 8681 15744
rect 8361 14656 8369 14720
rect 8433 14656 8449 14720
rect 8513 14656 8529 14720
rect 8593 14656 8609 14720
rect 8673 14656 8681 14720
rect 8361 13632 8681 14656
rect 8361 13568 8369 13632
rect 8433 13568 8449 13632
rect 8513 13568 8529 13632
rect 8593 13568 8609 13632
rect 8673 13568 8681 13632
rect 8361 12544 8681 13568
rect 8361 12480 8369 12544
rect 8433 12480 8449 12544
rect 8513 12480 8529 12544
rect 8593 12480 8609 12544
rect 8673 12480 8681 12544
rect 8361 11456 8681 12480
rect 8361 11392 8369 11456
rect 8433 11392 8449 11456
rect 8513 11392 8529 11456
rect 8593 11392 8609 11456
rect 8673 11392 8681 11456
rect 8361 10368 8681 11392
rect 8361 10304 8369 10368
rect 8433 10304 8449 10368
rect 8513 10304 8529 10368
rect 8593 10304 8609 10368
rect 8673 10304 8681 10368
rect 8361 9280 8681 10304
rect 8361 9216 8369 9280
rect 8433 9216 8449 9280
rect 8513 9216 8529 9280
rect 8593 9216 8609 9280
rect 8673 9216 8681 9280
rect 8361 8192 8681 9216
rect 8361 8128 8369 8192
rect 8433 8128 8449 8192
rect 8513 8128 8529 8192
rect 8593 8128 8609 8192
rect 8673 8128 8681 8192
rect 8361 7104 8681 8128
rect 8361 7040 8369 7104
rect 8433 7040 8449 7104
rect 8513 7040 8529 7104
rect 8593 7040 8609 7104
rect 8673 7040 8681 7104
rect 8361 6016 8681 7040
rect 8361 5952 8369 6016
rect 8433 5952 8449 6016
rect 8513 5952 8529 6016
rect 8593 5952 8609 6016
rect 8673 5952 8681 6016
rect 8361 4928 8681 5952
rect 8361 4864 8369 4928
rect 8433 4864 8449 4928
rect 8513 4864 8529 4928
rect 8593 4864 8609 4928
rect 8673 4864 8681 4928
rect 8361 3840 8681 4864
rect 8361 3776 8369 3840
rect 8433 3776 8449 3840
rect 8513 3776 8529 3840
rect 8593 3776 8609 3840
rect 8673 3776 8681 3840
rect 8361 2752 8681 3776
rect 8361 2688 8369 2752
rect 8433 2688 8449 2752
rect 8513 2688 8529 2752
rect 8593 2688 8609 2752
rect 8673 2688 8681 2752
rect 8361 2128 8681 2688
rect 10833 19616 11153 19632
rect 10833 19552 10841 19616
rect 10905 19552 10921 19616
rect 10985 19552 11001 19616
rect 11065 19552 11081 19616
rect 11145 19552 11153 19616
rect 10833 18528 11153 19552
rect 10833 18464 10841 18528
rect 10905 18464 10921 18528
rect 10985 18464 11001 18528
rect 11065 18464 11081 18528
rect 11145 18464 11153 18528
rect 10833 17440 11153 18464
rect 10833 17376 10841 17440
rect 10905 17376 10921 17440
rect 10985 17376 11001 17440
rect 11065 17376 11081 17440
rect 11145 17376 11153 17440
rect 10833 16352 11153 17376
rect 10833 16288 10841 16352
rect 10905 16288 10921 16352
rect 10985 16288 11001 16352
rect 11065 16288 11081 16352
rect 11145 16288 11153 16352
rect 10833 15264 11153 16288
rect 10833 15200 10841 15264
rect 10905 15200 10921 15264
rect 10985 15200 11001 15264
rect 11065 15200 11081 15264
rect 11145 15200 11153 15264
rect 10833 14176 11153 15200
rect 10833 14112 10841 14176
rect 10905 14112 10921 14176
rect 10985 14112 11001 14176
rect 11065 14112 11081 14176
rect 11145 14112 11153 14176
rect 10833 13088 11153 14112
rect 10833 13024 10841 13088
rect 10905 13024 10921 13088
rect 10985 13024 11001 13088
rect 11065 13024 11081 13088
rect 11145 13024 11153 13088
rect 10833 12000 11153 13024
rect 10833 11936 10841 12000
rect 10905 11936 10921 12000
rect 10985 11936 11001 12000
rect 11065 11936 11081 12000
rect 11145 11936 11153 12000
rect 10833 10912 11153 11936
rect 10833 10848 10841 10912
rect 10905 10848 10921 10912
rect 10985 10848 11001 10912
rect 11065 10848 11081 10912
rect 11145 10848 11153 10912
rect 10833 9824 11153 10848
rect 10833 9760 10841 9824
rect 10905 9760 10921 9824
rect 10985 9760 11001 9824
rect 11065 9760 11081 9824
rect 11145 9760 11153 9824
rect 10833 8736 11153 9760
rect 10833 8672 10841 8736
rect 10905 8672 10921 8736
rect 10985 8672 11001 8736
rect 11065 8672 11081 8736
rect 11145 8672 11153 8736
rect 10833 7648 11153 8672
rect 10833 7584 10841 7648
rect 10905 7584 10921 7648
rect 10985 7584 11001 7648
rect 11065 7584 11081 7648
rect 11145 7584 11153 7648
rect 10833 6560 11153 7584
rect 10833 6496 10841 6560
rect 10905 6496 10921 6560
rect 10985 6496 11001 6560
rect 11065 6496 11081 6560
rect 11145 6496 11153 6560
rect 10833 5472 11153 6496
rect 10833 5408 10841 5472
rect 10905 5408 10921 5472
rect 10985 5408 11001 5472
rect 11065 5408 11081 5472
rect 11145 5408 11153 5472
rect 10833 4384 11153 5408
rect 10833 4320 10841 4384
rect 10905 4320 10921 4384
rect 10985 4320 11001 4384
rect 11065 4320 11081 4384
rect 11145 4320 11153 4384
rect 10833 3296 11153 4320
rect 10833 3232 10841 3296
rect 10905 3232 10921 3296
rect 10985 3232 11001 3296
rect 11065 3232 11081 3296
rect 11145 3232 11153 3296
rect 10833 2208 11153 3232
rect 10833 2144 10841 2208
rect 10905 2144 10921 2208
rect 10985 2144 11001 2208
rect 11065 2144 11081 2208
rect 11145 2144 11153 2208
rect 10833 2128 11153 2144
rect 13306 19072 13626 19632
rect 13306 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13554 19072
rect 13618 19008 13626 19072
rect 13306 17984 13626 19008
rect 13306 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13554 17984
rect 13618 17920 13626 17984
rect 13306 16896 13626 17920
rect 13306 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13554 16896
rect 13618 16832 13626 16896
rect 13306 15808 13626 16832
rect 13306 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13554 15808
rect 13618 15744 13626 15808
rect 13306 14720 13626 15744
rect 13306 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13554 14720
rect 13618 14656 13626 14720
rect 13306 13632 13626 14656
rect 13306 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13554 13632
rect 13618 13568 13626 13632
rect 13306 12544 13626 13568
rect 13306 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13554 12544
rect 13618 12480 13626 12544
rect 13306 11456 13626 12480
rect 13306 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13554 11456
rect 13618 11392 13626 11456
rect 13306 10368 13626 11392
rect 13306 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13554 10368
rect 13618 10304 13626 10368
rect 13306 9280 13626 10304
rect 13306 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13554 9280
rect 13618 9216 13626 9280
rect 13306 8192 13626 9216
rect 13306 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13554 8192
rect 13618 8128 13626 8192
rect 13306 7104 13626 8128
rect 13306 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13554 7104
rect 13618 7040 13626 7104
rect 13306 6016 13626 7040
rect 13306 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13554 6016
rect 13618 5952 13626 6016
rect 13306 4928 13626 5952
rect 13306 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13554 4928
rect 13618 4864 13626 4928
rect 13306 3840 13626 4864
rect 13306 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13554 3840
rect 13618 3776 13626 3840
rect 13306 2752 13626 3776
rect 13306 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13554 2752
rect 13618 2688 13626 2752
rect 13306 2128 13626 2688
rect 15778 19616 16098 19632
rect 15778 19552 15786 19616
rect 15850 19552 15866 19616
rect 15930 19552 15946 19616
rect 16010 19552 16026 19616
rect 16090 19552 16098 19616
rect 15778 18528 16098 19552
rect 15778 18464 15786 18528
rect 15850 18464 15866 18528
rect 15930 18464 15946 18528
rect 16010 18464 16026 18528
rect 16090 18464 16098 18528
rect 15778 17440 16098 18464
rect 15778 17376 15786 17440
rect 15850 17376 15866 17440
rect 15930 17376 15946 17440
rect 16010 17376 16026 17440
rect 16090 17376 16098 17440
rect 15778 16352 16098 17376
rect 15778 16288 15786 16352
rect 15850 16288 15866 16352
rect 15930 16288 15946 16352
rect 16010 16288 16026 16352
rect 16090 16288 16098 16352
rect 15778 15264 16098 16288
rect 15778 15200 15786 15264
rect 15850 15200 15866 15264
rect 15930 15200 15946 15264
rect 16010 15200 16026 15264
rect 16090 15200 16098 15264
rect 15778 14176 16098 15200
rect 15778 14112 15786 14176
rect 15850 14112 15866 14176
rect 15930 14112 15946 14176
rect 16010 14112 16026 14176
rect 16090 14112 16098 14176
rect 15778 13088 16098 14112
rect 15778 13024 15786 13088
rect 15850 13024 15866 13088
rect 15930 13024 15946 13088
rect 16010 13024 16026 13088
rect 16090 13024 16098 13088
rect 15778 12000 16098 13024
rect 15778 11936 15786 12000
rect 15850 11936 15866 12000
rect 15930 11936 15946 12000
rect 16010 11936 16026 12000
rect 16090 11936 16098 12000
rect 15778 10912 16098 11936
rect 15778 10848 15786 10912
rect 15850 10848 15866 10912
rect 15930 10848 15946 10912
rect 16010 10848 16026 10912
rect 16090 10848 16098 10912
rect 15778 9824 16098 10848
rect 15778 9760 15786 9824
rect 15850 9760 15866 9824
rect 15930 9760 15946 9824
rect 16010 9760 16026 9824
rect 16090 9760 16098 9824
rect 15778 8736 16098 9760
rect 15778 8672 15786 8736
rect 15850 8672 15866 8736
rect 15930 8672 15946 8736
rect 16010 8672 16026 8736
rect 16090 8672 16098 8736
rect 15778 7648 16098 8672
rect 15778 7584 15786 7648
rect 15850 7584 15866 7648
rect 15930 7584 15946 7648
rect 16010 7584 16026 7648
rect 16090 7584 16098 7648
rect 15778 6560 16098 7584
rect 15778 6496 15786 6560
rect 15850 6496 15866 6560
rect 15930 6496 15946 6560
rect 16010 6496 16026 6560
rect 16090 6496 16098 6560
rect 15778 5472 16098 6496
rect 15778 5408 15786 5472
rect 15850 5408 15866 5472
rect 15930 5408 15946 5472
rect 16010 5408 16026 5472
rect 16090 5408 16098 5472
rect 15778 4384 16098 5408
rect 15778 4320 15786 4384
rect 15850 4320 15866 4384
rect 15930 4320 15946 4384
rect 16010 4320 16026 4384
rect 16090 4320 16098 4384
rect 15778 3296 16098 4320
rect 15778 3232 15786 3296
rect 15850 3232 15866 3296
rect 15930 3232 15946 3296
rect 16010 3232 16026 3296
rect 16090 3232 16098 3296
rect 15778 2208 16098 3232
rect 15778 2144 15786 2208
rect 15850 2144 15866 2208
rect 15930 2144 15946 2208
rect 16010 2144 16026 2208
rect 16090 2144 16098 2208
rect 15778 2128 16098 2144
rect 18251 19072 18571 19632
rect 18251 19008 18259 19072
rect 18323 19008 18339 19072
rect 18403 19008 18419 19072
rect 18483 19008 18499 19072
rect 18563 19008 18571 19072
rect 18251 17984 18571 19008
rect 18251 17920 18259 17984
rect 18323 17920 18339 17984
rect 18403 17920 18419 17984
rect 18483 17920 18499 17984
rect 18563 17920 18571 17984
rect 18251 16896 18571 17920
rect 18251 16832 18259 16896
rect 18323 16832 18339 16896
rect 18403 16832 18419 16896
rect 18483 16832 18499 16896
rect 18563 16832 18571 16896
rect 18251 15808 18571 16832
rect 18251 15744 18259 15808
rect 18323 15744 18339 15808
rect 18403 15744 18419 15808
rect 18483 15744 18499 15808
rect 18563 15744 18571 15808
rect 18251 14720 18571 15744
rect 18251 14656 18259 14720
rect 18323 14656 18339 14720
rect 18403 14656 18419 14720
rect 18483 14656 18499 14720
rect 18563 14656 18571 14720
rect 18251 13632 18571 14656
rect 18251 13568 18259 13632
rect 18323 13568 18339 13632
rect 18403 13568 18419 13632
rect 18483 13568 18499 13632
rect 18563 13568 18571 13632
rect 18251 12544 18571 13568
rect 18251 12480 18259 12544
rect 18323 12480 18339 12544
rect 18403 12480 18419 12544
rect 18483 12480 18499 12544
rect 18563 12480 18571 12544
rect 18251 11456 18571 12480
rect 18251 11392 18259 11456
rect 18323 11392 18339 11456
rect 18403 11392 18419 11456
rect 18483 11392 18499 11456
rect 18563 11392 18571 11456
rect 18251 10368 18571 11392
rect 18251 10304 18259 10368
rect 18323 10304 18339 10368
rect 18403 10304 18419 10368
rect 18483 10304 18499 10368
rect 18563 10304 18571 10368
rect 18251 9280 18571 10304
rect 18251 9216 18259 9280
rect 18323 9216 18339 9280
rect 18403 9216 18419 9280
rect 18483 9216 18499 9280
rect 18563 9216 18571 9280
rect 18251 8192 18571 9216
rect 18251 8128 18259 8192
rect 18323 8128 18339 8192
rect 18403 8128 18419 8192
rect 18483 8128 18499 8192
rect 18563 8128 18571 8192
rect 18251 7104 18571 8128
rect 18251 7040 18259 7104
rect 18323 7040 18339 7104
rect 18403 7040 18419 7104
rect 18483 7040 18499 7104
rect 18563 7040 18571 7104
rect 18251 6016 18571 7040
rect 18251 5952 18259 6016
rect 18323 5952 18339 6016
rect 18403 5952 18419 6016
rect 18483 5952 18499 6016
rect 18563 5952 18571 6016
rect 18251 4928 18571 5952
rect 18251 4864 18259 4928
rect 18323 4864 18339 4928
rect 18403 4864 18419 4928
rect 18483 4864 18499 4928
rect 18563 4864 18571 4928
rect 18251 3840 18571 4864
rect 18251 3776 18259 3840
rect 18323 3776 18339 3840
rect 18403 3776 18419 3840
rect 18483 3776 18499 3840
rect 18563 3776 18571 3840
rect 18251 2752 18571 3776
rect 18251 2688 18259 2752
rect 18323 2688 18339 2752
rect 18403 2688 18419 2752
rect 18483 2688 18499 2752
rect 18563 2688 18571 2752
rect 18251 2128 18571 2688
rect 20723 19616 21043 19632
rect 20723 19552 20731 19616
rect 20795 19552 20811 19616
rect 20875 19552 20891 19616
rect 20955 19552 20971 19616
rect 21035 19552 21043 19616
rect 20723 18528 21043 19552
rect 20723 18464 20731 18528
rect 20795 18464 20811 18528
rect 20875 18464 20891 18528
rect 20955 18464 20971 18528
rect 21035 18464 21043 18528
rect 20723 17440 21043 18464
rect 20723 17376 20731 17440
rect 20795 17376 20811 17440
rect 20875 17376 20891 17440
rect 20955 17376 20971 17440
rect 21035 17376 21043 17440
rect 20723 16352 21043 17376
rect 20723 16288 20731 16352
rect 20795 16288 20811 16352
rect 20875 16288 20891 16352
rect 20955 16288 20971 16352
rect 21035 16288 21043 16352
rect 20723 15264 21043 16288
rect 20723 15200 20731 15264
rect 20795 15200 20811 15264
rect 20875 15200 20891 15264
rect 20955 15200 20971 15264
rect 21035 15200 21043 15264
rect 20723 14176 21043 15200
rect 20723 14112 20731 14176
rect 20795 14112 20811 14176
rect 20875 14112 20891 14176
rect 20955 14112 20971 14176
rect 21035 14112 21043 14176
rect 20723 13088 21043 14112
rect 20723 13024 20731 13088
rect 20795 13024 20811 13088
rect 20875 13024 20891 13088
rect 20955 13024 20971 13088
rect 21035 13024 21043 13088
rect 20723 12000 21043 13024
rect 20723 11936 20731 12000
rect 20795 11936 20811 12000
rect 20875 11936 20891 12000
rect 20955 11936 20971 12000
rect 21035 11936 21043 12000
rect 20723 10912 21043 11936
rect 20723 10848 20731 10912
rect 20795 10848 20811 10912
rect 20875 10848 20891 10912
rect 20955 10848 20971 10912
rect 21035 10848 21043 10912
rect 20723 9824 21043 10848
rect 20723 9760 20731 9824
rect 20795 9760 20811 9824
rect 20875 9760 20891 9824
rect 20955 9760 20971 9824
rect 21035 9760 21043 9824
rect 20723 8736 21043 9760
rect 20723 8672 20731 8736
rect 20795 8672 20811 8736
rect 20875 8672 20891 8736
rect 20955 8672 20971 8736
rect 21035 8672 21043 8736
rect 20723 7648 21043 8672
rect 20723 7584 20731 7648
rect 20795 7584 20811 7648
rect 20875 7584 20891 7648
rect 20955 7584 20971 7648
rect 21035 7584 21043 7648
rect 20723 6560 21043 7584
rect 20723 6496 20731 6560
rect 20795 6496 20811 6560
rect 20875 6496 20891 6560
rect 20955 6496 20971 6560
rect 21035 6496 21043 6560
rect 20723 5472 21043 6496
rect 20723 5408 20731 5472
rect 20795 5408 20811 5472
rect 20875 5408 20891 5472
rect 20955 5408 20971 5472
rect 21035 5408 21043 5472
rect 20723 4384 21043 5408
rect 20723 4320 20731 4384
rect 20795 4320 20811 4384
rect 20875 4320 20891 4384
rect 20955 4320 20971 4384
rect 21035 4320 21043 4384
rect 20723 3296 21043 4320
rect 20723 3232 20731 3296
rect 20795 3232 20811 3296
rect 20875 3232 20891 3296
rect 20955 3232 20971 3296
rect 21035 3232 21043 3296
rect 20723 2208 21043 3232
rect 20723 2144 20731 2208
rect 20795 2144 20811 2208
rect 20875 2144 20891 2208
rect 20955 2144 20971 2208
rect 21035 2144 21043 2208
rect 20723 2128 21043 2144
use sky130_fd_sc_hd__decap_3  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36
timestamp 1676037725
transform 1 0 4416 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1676037725
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127
timestamp 1676037725
transform 1 0 12788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1676037725
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 1676037725
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1676037725
transform 1 0 15456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1676037725
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_36
timestamp 1676037725
transform 1 0 4416 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_44
timestamp 1676037725
transform 1 0 5152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_65
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_103
timestamp 1676037725
transform 1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_133
timestamp 1676037725
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1676037725
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_150
timestamp 1676037725
transform 1 0 14904 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1676037725
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_179
timestamp 1676037725
transform 1 0 17572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_191
timestamp 1676037725
transform 1 0 18676 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_203
timestamp 1676037725
transform 1 0 19780 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_211
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1676037725
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_35
timestamp 1676037725
transform 1 0 4324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_47
timestamp 1676037725
transform 1 0 5428 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_59
timestamp 1676037725
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1676037725
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1676037725
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1676037725
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_128
timestamp 1676037725
transform 1 0 12880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1676037725
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_151
timestamp 1676037725
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_158
timestamp 1676037725
transform 1 0 15640 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_166
timestamp 1676037725
transform 1 0 16376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_176
timestamp 1676037725
transform 1 0 17296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1676037725
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_10
timestamp 1676037725
transform 1 0 2024 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_34
timestamp 1676037725
transform 1 0 4232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1676037725
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_148
timestamp 1676037725
transform 1 0 14720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1676037725
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_211
timestamp 1676037725
transform 1 0 20516 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_116
timestamp 1676037725
transform 1 0 11776 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_128
timestamp 1676037725
transform 1 0 12880 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_146
timestamp 1676037725
transform 1 0 14536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_150
timestamp 1676037725
transform 1 0 14904 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_154
timestamp 1676037725
transform 1 0 15272 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_166
timestamp 1676037725
transform 1 0 16376 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_175
timestamp 1676037725
transform 1 0 17204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_182
timestamp 1676037725
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_22
timestamp 1676037725
transform 1 0 3128 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_34
timestamp 1676037725
transform 1 0 4232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1676037725
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_138
timestamp 1676037725
transform 1 0 13800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_150
timestamp 1676037725
transform 1 0 14904 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_162
timestamp 1676037725
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1676037725
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_182
timestamp 1676037725
transform 1 0 17848 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_194
timestamp 1676037725
transform 1 0 18952 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_206
timestamp 1676037725
transform 1 0 20056 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_33
timestamp 1676037725
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1676037725
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1676037725
transform 1 0 9660 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_110
timestamp 1676037725
transform 1 0 11224 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_122
timestamp 1676037725
transform 1 0 12328 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_175
timestamp 1676037725
transform 1 0 17204 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_182
timestamp 1676037725
transform 1 0 17848 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_33
timestamp 1676037725
transform 1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1676037725
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_73
timestamp 1676037725
transform 1 0 7820 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_90
timestamp 1676037725
transform 1 0 9384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_140
timestamp 1676037725
transform 1 0 13984 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_156
timestamp 1676037725
transform 1 0 15456 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_177
timestamp 1676037725
transform 1 0 17388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1676037725
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_198
timestamp 1676037725
transform 1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_207
timestamp 1676037725
transform 1 0 20148 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_211
timestamp 1676037725
transform 1 0 20516 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1676037725
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_116
timestamp 1676037725
transform 1 0 11776 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_128
timestamp 1676037725
transform 1 0 12880 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_152
timestamp 1676037725
transform 1 0 15088 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_161
timestamp 1676037725
transform 1 0 15916 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_173
timestamp 1676037725
transform 1 0 17020 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_181
timestamp 1676037725
transform 1 0 17756 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1676037725
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_207
timestamp 1676037725
transform 1 0 20148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_211
timestamp 1676037725
transform 1 0 20516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_36
timestamp 1676037725
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1676037725
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_144
timestamp 1676037725
transform 1 0 14352 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_156
timestamp 1676037725
transform 1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1676037725
transform 1 0 17480 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_189
timestamp 1676037725
transform 1 0 18492 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_196
timestamp 1676037725
transform 1 0 19136 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_208
timestamp 1676037725
transform 1 0 20240 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1676037725
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_54
timestamp 1676037725
transform 1 0 6072 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1676037725
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_117
timestamp 1676037725
transform 1 0 11868 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_157
timestamp 1676037725
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_167
timestamp 1676037725
transform 1 0 16468 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_179
timestamp 1676037725
transform 1 0 17572 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_183
timestamp 1676037725
transform 1 0 17940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_77
timestamp 1676037725
transform 1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_96
timestamp 1676037725
transform 1 0 9936 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1676037725
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_133
timestamp 1676037725
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_144
timestamp 1676037725
transform 1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_151
timestamp 1676037725
transform 1 0 14996 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_176
timestamp 1676037725
transform 1 0 17296 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_184
timestamp 1676037725
transform 1 0 18032 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_200
timestamp 1676037725
transform 1 0 19504 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_35
timestamp 1676037725
transform 1 0 4324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_74
timestamp 1676037725
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1676037725
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_119
timestamp 1676037725
transform 1 0 12052 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_131
timestamp 1676037725
transform 1 0 13156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_148
timestamp 1676037725
transform 1 0 14720 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_176
timestamp 1676037725
transform 1 0 17296 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_184
timestamp 1676037725
transform 1 0 18032 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1676037725
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_33
timestamp 1676037725
transform 1 0 4140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_78
timestamp 1676037725
transform 1 0 8280 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_90
timestamp 1676037725
transform 1 0 9384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1676037725
transform 1 0 15456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1676037725
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_210
timestamp 1676037725
transform 1 0 20424 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1676037725
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_119
timestamp 1676037725
transform 1 0 12052 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_131
timestamp 1676037725
transform 1 0 13156 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_149
timestamp 1676037725
transform 1 0 14812 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_157
timestamp 1676037725
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_163
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_171
timestamp 1676037725
transform 1 0 16836 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_11
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_133
timestamp 1676037725
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_144
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_156
timestamp 1676037725
transform 1 0 15456 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1676037725
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_177
timestamp 1676037725
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_185
timestamp 1676037725
transform 1 0 18124 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_11
timestamp 1676037725
transform 1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1676037725
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_48
timestamp 1676037725
transform 1 0 5520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_56
timestamp 1676037725
transform 1 0 6256 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_68
timestamp 1676037725
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1676037725
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_94
timestamp 1676037725
transform 1 0 9752 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_106
timestamp 1676037725
transform 1 0 10856 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_119
timestamp 1676037725
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1676037725
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_146
timestamp 1676037725
transform 1 0 14536 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_158
timestamp 1676037725
transform 1 0 15640 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_178
timestamp 1676037725
transform 1 0 17480 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_184
timestamp 1676037725
transform 1 0 18032 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_14
timestamp 1676037725
transform 1 0 2392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_18
timestamp 1676037725
transform 1 0 2760 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_40
timestamp 1676037725
transform 1 0 4784 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 1676037725
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_71
timestamp 1676037725
transform 1 0 7636 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_79
timestamp 1676037725
transform 1 0 8372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_90
timestamp 1676037725
transform 1 0 9384 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_98
timestamp 1676037725
transform 1 0 10120 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1676037725
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_123
timestamp 1676037725
transform 1 0 12420 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_154
timestamp 1676037725
transform 1 0 15272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_175
timestamp 1676037725
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_179
timestamp 1676037725
transform 1 0 17572 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_185
timestamp 1676037725
transform 1 0 18124 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_194
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_204
timestamp 1676037725
transform 1 0 19872 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_11
timestamp 1676037725
transform 1 0 2116 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1676037725
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_44
timestamp 1676037725
transform 1 0 5152 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_56
timestamp 1676037725
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_116
timestamp 1676037725
transform 1 0 11776 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_120
timestamp 1676037725
transform 1 0 12144 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_132
timestamp 1676037725
transform 1 0 13248 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_150
timestamp 1676037725
transform 1 0 14904 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_157
timestamp 1676037725
transform 1 0 15548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_169
timestamp 1676037725
transform 1 0 16652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1676037725
transform 1 0 17296 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_188
timestamp 1676037725
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1676037725
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1676037725
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_25
timestamp 1676037725
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_37
timestamp 1676037725
transform 1 0 4508 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1676037725
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_76
timestamp 1676037725
transform 1 0 8096 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_88
timestamp 1676037725
transform 1 0 9200 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_100
timestamp 1676037725
transform 1 0 10304 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1676037725
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_129
timestamp 1676037725
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_176
timestamp 1676037725
transform 1 0 17296 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_189
timestamp 1676037725
transform 1 0 18492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_198
timestamp 1676037725
transform 1 0 19320 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1676037725
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1676037725
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_17
timestamp 1676037725
transform 1 0 2668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1676037725
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_34
timestamp 1676037725
transform 1 0 4232 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_40
timestamp 1676037725
transform 1 0 4784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_50
timestamp 1676037725
transform 1 0 5704 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_66
timestamp 1676037725
transform 1 0 7176 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_78
timestamp 1676037725
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_94
timestamp 1676037725
transform 1 0 9752 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_105
timestamp 1676037725
transform 1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_118
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_126
timestamp 1676037725
transform 1 0 12696 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1676037725
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_158
timestamp 1676037725
transform 1 0 15640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_169
timestamp 1676037725
transform 1 0 16652 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_206
timestamp 1676037725
transform 1 0 20056 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_14
timestamp 1676037725
transform 1 0 2392 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_22
timestamp 1676037725
transform 1 0 3128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_32
timestamp 1676037725
transform 1 0 4048 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_40
timestamp 1676037725
transform 1 0 4784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1676037725
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_77
timestamp 1676037725
transform 1 0 8188 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_82
timestamp 1676037725
transform 1 0 8648 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_94
timestamp 1676037725
transform 1 0 9752 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_102
timestamp 1676037725
transform 1 0 10488 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_123
timestamp 1676037725
transform 1 0 12420 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_134
timestamp 1676037725
transform 1 0 13432 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_177
timestamp 1676037725
transform 1 0 17388 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_186
timestamp 1676037725
transform 1 0 18216 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_210
timestamp 1676037725
transform 1 0 20424 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_61
timestamp 1676037725
transform 1 0 6716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1676037725
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_95
timestamp 1676037725
transform 1 0 9844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1676037725
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_112
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_120
timestamp 1676037725
transform 1 0 12144 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1676037725
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1676037725
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_152
timestamp 1676037725
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_159
timestamp 1676037725
transform 1 0 15732 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_171
timestamp 1676037725
transform 1 0 16836 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_180
timestamp 1676037725
transform 1 0 17664 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_207
timestamp 1676037725
transform 1 0 20148 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_211
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_35
timestamp 1676037725
transform 1 0 4324 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_43
timestamp 1676037725
transform 1 0 5060 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1676037725
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_67
timestamp 1676037725
transform 1 0 7268 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_79
timestamp 1676037725
transform 1 0 8372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_91
timestamp 1676037725
transform 1 0 9476 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_99
timestamp 1676037725
transform 1 0 10212 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_124
timestamp 1676037725
transform 1 0 12512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_128
timestamp 1676037725
transform 1 0 12880 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_133
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_145
timestamp 1676037725
transform 1 0 14444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_150
timestamp 1676037725
transform 1 0 14904 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1676037725
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_180
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_188
timestamp 1676037725
transform 1 0 18400 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_198
timestamp 1676037725
transform 1 0 19320 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_210
timestamp 1676037725
transform 1 0 20424 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1676037725
transform 1 0 2116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_16
timestamp 1676037725
transform 1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1676037725
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_44
timestamp 1676037725
transform 1 0 5152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_54
timestamp 1676037725
transform 1 0 6072 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_64
timestamp 1676037725
transform 1 0 6992 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_71
timestamp 1676037725
transform 1 0 7636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1676037725
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_102
timestamp 1676037725
transform 1 0 10488 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1676037725
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_123
timestamp 1676037725
transform 1 0 12420 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1676037725
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1676037725
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1676037725
transform 1 0 14812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1676037725
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_175
timestamp 1676037725
transform 1 0 17204 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_187
timestamp 1676037725
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_71
timestamp 1676037725
transform 1 0 7636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_95
timestamp 1676037725
transform 1 0 9844 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_103
timestamp 1676037725
transform 1 0 10580 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_121
timestamp 1676037725
transform 1 0 12236 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_134
timestamp 1676037725
transform 1 0 13432 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_154
timestamp 1676037725
transform 1 0 15272 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_211
timestamp 1676037725
transform 1 0 20516 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_35
timestamp 1676037725
transform 1 0 4324 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_54
timestamp 1676037725
transform 1 0 6072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_58
timestamp 1676037725
transform 1 0 6440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1676037725
transform 1 0 7452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_78
timestamp 1676037725
transform 1 0 8280 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_116
timestamp 1676037725
transform 1 0 11776 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_128
timestamp 1676037725
transform 1 0 12880 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_23
timestamp 1676037725
transform 1 0 3220 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_29
timestamp 1676037725
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1676037725
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1676037725
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_72
timestamp 1676037725
transform 1 0 7728 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_84
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_96
timestamp 1676037725
transform 1 0 9936 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1676037725
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_205
timestamp 1676037725
transform 1 0 19964 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_211
timestamp 1676037725
transform 1 0 20516 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_205
timestamp 1676037725
transform 1 0 19964 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_211
timestamp 1676037725
transform 1 0 20516 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_11
timestamp 1676037725
transform 1 0 2116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1676037725
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_29
timestamp 1676037725
transform 1 0 3772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1676037725
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_85
timestamp 1676037725
transform 1 0 8924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_97
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1676037725
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_141
timestamp 1676037725
transform 1 0 14076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_153
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1676037725
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_197
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_209
timestamp 1676037725
transform 1 0 20332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 20884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 20884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 20884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 20884 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 20884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 20884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 20884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 20884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 20884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 3680 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 8832 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 13984 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17572 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1676037725
transform -1 0 20056 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1676037725
transform -1 0 12144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1676037725
transform 1 0 15180 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1676037725
transform -1 0 15272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1676037725
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2300 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5152 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and4_4  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5244 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12972 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14904 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _211_
timestamp 1676037725
transform 1 0 14628 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_2  _213_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13800 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_2  _214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15272 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19688 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15456 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16376 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1676037725
transform 1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17296 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17204 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1676037725
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18952 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_4  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17296 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_4  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20424 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_4  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20332 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1676037725
transform -1 0 17296 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _229_
timestamp 1676037725
transform 1 0 15272 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20240 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18860 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18308 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_4  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18952 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__and2_2  _234_
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _235_
timestamp 1676037725
transform -1 0 15272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _236_
timestamp 1676037725
transform -1 0 18952 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12420 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _239_
timestamp 1676037725
transform 1 0 10580 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1676037725
transform -1 0 11776 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _241_
timestamp 1676037725
transform -1 0 16376 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _242_
timestamp 1676037725
transform 1 0 12880 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20332 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _244_
timestamp 1676037725
transform -1 0 18124 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _245_
timestamp 1676037725
transform 1 0 11408 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10304 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12052 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _249_
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _250_
timestamp 1676037725
transform 1 0 15640 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _252_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _253_
timestamp 1676037725
transform 1 0 8740 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _254_
timestamp 1676037725
transform -1 0 9844 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1676037725
transform -1 0 14536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _260_
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18952 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _262_
timestamp 1676037725
transform -1 0 18492 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 1676037725
transform -1 0 13432 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13064 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _266_
timestamp 1676037725
transform -1 0 13340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _268_
timestamp 1676037725
transform -1 0 13800 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14812 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _270_
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12788 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _274_
timestamp 1676037725
transform -1 0 18124 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _275_
timestamp 1676037725
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _276_
timestamp 1676037725
transform 1 0 14536 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12512 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11040 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10212 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _280_
timestamp 1676037725
transform -1 0 15732 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1676037725
transform 1 0 15824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _283_
timestamp 1676037725
transform -1 0 19320 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _284_
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16376 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _287_
timestamp 1676037725
transform 1 0 16468 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _288_
timestamp 1676037725
transform -1 0 17296 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _289_
timestamp 1676037725
transform 1 0 15732 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _290_
timestamp 1676037725
transform -1 0 14904 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _291_
timestamp 1676037725
transform 1 0 14536 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _292_
timestamp 1676037725
transform 1 0 15272 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _293_
timestamp 1676037725
transform 1 0 17112 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _294_
timestamp 1676037725
transform -1 0 18400 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _295_
timestamp 1676037725
transform -1 0 18676 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _296_
timestamp 1676037725
transform 1 0 17664 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _297_
timestamp 1676037725
transform 1 0 17664 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16652 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _300_
timestamp 1676037725
transform -1 0 17664 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15088 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15640 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _304_
timestamp 1676037725
transform 1 0 12788 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _305_
timestamp 1676037725
transform 1 0 8004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _306_
timestamp 1676037725
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _307_
timestamp 1676037725
transform -1 0 13340 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _308_
timestamp 1676037725
transform 1 0 9844 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _309_
timestamp 1676037725
transform 1 0 8740 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _310_
timestamp 1676037725
transform 1 0 8464 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _311_
timestamp 1676037725
transform 1 0 8372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _312_
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _313_
timestamp 1676037725
transform 1 0 9108 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _314_
timestamp 1676037725
transform -1 0 2944 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18860 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _316_
timestamp 1676037725
transform -1 0 14996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13800 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _318_
timestamp 1676037725
transform 1 0 13156 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _319_
timestamp 1676037725
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _320_
timestamp 1676037725
transform -1 0 14720 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13616 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _322_
timestamp 1676037725
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _323_
timestamp 1676037725
transform 1 0 16836 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _324_
timestamp 1676037725
transform 1 0 16836 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _325_
timestamp 1676037725
transform 1 0 15640 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _326_
timestamp 1676037725
transform 1 0 15088 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _327_
timestamp 1676037725
transform 1 0 14352 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _328_
timestamp 1676037725
transform 1 0 12972 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _329_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18584 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _331_
timestamp 1676037725
transform 1 0 1748 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _332_
timestamp 1676037725
transform 1 0 6348 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_4  _333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_1  _334_
timestamp 1676037725
transform -1 0 2392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _335_
timestamp 1676037725
transform 1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _336_
timestamp 1676037725
transform 1 0 7360 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _337_
timestamp 1676037725
transform -1 0 3772 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _338_
timestamp 1676037725
transform -1 0 8188 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8280 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _340_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3496 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1676037725
transform 1 0 1656 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _343_
timestamp 1676037725
transform -1 0 5520 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _344_
timestamp 1676037725
transform 1 0 4416 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _345_
timestamp 1676037725
transform 1 0 5428 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _346_
timestamp 1676037725
transform -1 0 7360 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _347_
timestamp 1676037725
transform 1 0 6440 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1676037725
transform 1 0 1840 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _349_
timestamp 1676037725
transform -1 0 7728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _350_
timestamp 1676037725
transform 1 0 6624 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7636 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1676037725
transform 1 0 6808 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1676037725
transform 1 0 6532 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _354_
timestamp 1676037725
transform 1 0 3128 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _355_
timestamp 1676037725
transform 1 0 2300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _356_
timestamp 1676037725
transform 1 0 3680 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1676037725
transform 1 0 4324 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1676037725
transform 1 0 3956 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _359_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7268 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _360_
timestamp 1676037725
transform -1 0 5152 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _361_
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1676037725
transform 1 0 4600 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _364_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7452 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _365_
timestamp 1676037725
transform 1 0 5428 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _366_
timestamp 1676037725
transform -1 0 5336 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _367_
timestamp 1676037725
transform 1 0 4968 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _368_
timestamp 1676037725
transform 1 0 5152 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2944 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _370_
timestamp 1676037725
transform -1 0 4232 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _371_
timestamp 1676037725
transform 1 0 3036 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _372_
timestamp 1676037725
transform 1 0 3312 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _373_
timestamp 1676037725
transform -1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1676037725
transform 1 0 12512 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _375_
timestamp 1676037725
transform 1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _376_
timestamp 1676037725
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _377_
timestamp 1676037725
transform 1 0 2392 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _378_
timestamp 1676037725
transform -1 0 4416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _379_
timestamp 1676037725
transform -1 0 4324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _380_
timestamp 1676037725
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _381_
timestamp 1676037725
transform -1 0 7084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _382_
timestamp 1676037725
transform -1 0 8648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _383_
timestamp 1676037725
transform 1 0 10028 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _384_
timestamp 1676037725
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _385_
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _386_
timestamp 1676037725
transform 1 0 15364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _387_
timestamp 1676037725
transform 1 0 13524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _388_
timestamp 1676037725
transform 1 0 15548 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _389_
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _390_
timestamp 1676037725
transform -1 0 14904 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17848 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1676037725
transform 1 0 18216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _393_
timestamp 1676037725
transform 1 0 16652 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _394_
timestamp 1676037725
transform -1 0 17848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1676037725
transform 1 0 16376 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _396_
timestamp 1676037725
transform 1 0 17112 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16928 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _398_
timestamp 1676037725
transform -1 0 18308 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _399_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10304 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1676037725
transform 1 0 9752 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4508 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _402_
timestamp 1676037725
transform -1 0 7912 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _403_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8280 0 -1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _404_
timestamp 1676037725
transform 1 0 2668 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1676037725
transform 1 0 7084 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1676037725
transform 1 0 9752 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1676037725
transform 1 0 7912 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1676037725
transform 1 0 9752 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1676037725
transform 1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _410_
timestamp 1676037725
transform 1 0 10304 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _411_
timestamp 1676037725
transform 1 0 10304 0 1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _412_
timestamp 1676037725
transform 1 0 8464 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _413_
timestamp 1676037725
transform 1 0 6808 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1676037725
transform 1 0 7176 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1676037725
transform 1 0 4508 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _416_
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _418_
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1676037725
transform 1 0 4508 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1676037725
transform 1 0 2668 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _421_
timestamp 1676037725
transform 1 0 4508 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _422_
timestamp 1676037725
transform 1 0 4416 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _423_
timestamp 1676037725
transform 1 0 2024 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _424_
timestamp 1676037725
transform 1 0 9752 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _425_
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _426_
timestamp 1676037725
transform 1 0 1748 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _427_
timestamp 1676037725
transform 1 0 2760 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _428_
timestamp 1676037725
transform 1 0 4600 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _429_
timestamp 1676037725
transform 1 0 7084 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _430_
timestamp 1676037725
transform 1 0 6808 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _431_
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _432_
timestamp 1676037725
transform 1 0 9108 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _433_
timestamp 1676037725
transform 1 0 4600 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _434_
timestamp 1676037725
transform 1 0 10304 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _435_
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _436_
timestamp 1676037725
transform 1 0 9752 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _437_
timestamp 1676037725
transform 1 0 11040 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _438_
timestamp 1676037725
transform 1 0 4232 0 1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout4
timestamp 1676037725
transform -1 0 12236 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6072 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout7
timestamp 1676037725
transform 1 0 12972 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  fanout8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output2
timestamp 1676037725
transform -1 0 2116 0 1 18496
box -38 -48 590 592
<< labels >>
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 OP
port 0 nsew signal tristate
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 clk
port 1 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 rst
port 2 nsew signal input
flabel metal4 s 3416 2128 3736 19632 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 8361 2128 8681 19632 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 13306 2128 13626 19632 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 18251 2128 18571 19632 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 5888 2128 6208 19632 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 10833 2128 11153 19632 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 15778 2128 16098 19632 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 20723 2128 21043 19632 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 22000 22000
<< end >>
