magic
tech sky130B
magscale 1 2
timestamp 1686562148
<< viali >>
rect 26249 37417 26283 37451
rect 32597 37417 32631 37451
rect 33241 37417 33275 37451
rect 7021 37281 7055 37315
rect 9689 37281 9723 37315
rect 12357 37281 12391 37315
rect 13553 37281 13587 37315
rect 19717 37281 19751 37315
rect 32413 37281 32447 37315
rect 33701 37281 33735 37315
rect 1961 37213 1995 37247
rect 3249 37213 3283 37247
rect 3433 37213 3467 37247
rect 4537 37213 4571 37247
rect 4721 37213 4755 37247
rect 5273 37213 5307 37247
rect 7205 37213 7239 37247
rect 7941 37213 7975 37247
rect 10517 37213 10551 37247
rect 14381 37213 14415 37247
rect 14565 37213 14599 37247
rect 15117 37213 15151 37247
rect 17049 37213 17083 37247
rect 17969 37213 18003 37247
rect 19441 37213 19475 37247
rect 22109 37213 22143 37247
rect 23581 37213 23615 37247
rect 25145 37213 25179 37247
rect 26249 37213 26283 37247
rect 26433 37213 26467 37247
rect 27169 37213 27203 37247
rect 28181 37213 28215 37247
rect 29009 37213 29043 37247
rect 29193 37213 29227 37247
rect 30297 37213 30331 37247
rect 30564 37213 30598 37247
rect 32328 37213 32362 37247
rect 32597 37213 32631 37247
rect 33425 37213 33459 37247
rect 33609 37213 33643 37247
rect 34161 37213 34195 37247
rect 34253 37213 34287 37247
rect 35449 37213 35483 37247
rect 37657 37213 37691 37247
rect 2513 37145 2547 37179
rect 3341 37145 3375 37179
rect 5825 37145 5859 37179
rect 8493 37145 8527 37179
rect 11069 37145 11103 37179
rect 12173 37145 12207 37179
rect 15945 37145 15979 37179
rect 17325 37145 17359 37179
rect 18797 37145 18831 37179
rect 22661 37145 22695 37179
rect 23857 37145 23891 37179
rect 25513 37145 25547 37179
rect 27445 37145 27479 37179
rect 35716 37145 35750 37179
rect 38025 37145 38059 37179
rect 4169 37077 4203 37111
rect 4721 37077 4755 37111
rect 7389 37077 7423 37111
rect 9137 37077 9171 37111
rect 9505 37077 9539 37111
rect 9597 37077 9631 37111
rect 11805 37077 11839 37111
rect 12265 37077 12299 37111
rect 13001 37077 13035 37111
rect 13369 37077 13403 37111
rect 13461 37077 13495 37111
rect 14565 37077 14599 37111
rect 21189 37077 21223 37111
rect 26617 37077 26651 37111
rect 28273 37077 28307 37111
rect 29101 37077 29135 37111
rect 31677 37077 31711 37111
rect 32781 37077 32815 37111
rect 36829 37077 36863 37111
rect 3065 36873 3099 36907
rect 3709 36873 3743 36907
rect 4445 36873 4479 36907
rect 5089 36873 5123 36907
rect 6009 36873 6043 36907
rect 9321 36873 9355 36907
rect 14381 36873 14415 36907
rect 4997 36805 5031 36839
rect 7297 36805 7331 36839
rect 12357 36805 12391 36839
rect 22569 36805 22603 36839
rect 24317 36805 24351 36839
rect 27721 36805 27755 36839
rect 28733 36805 28767 36839
rect 35716 36805 35750 36839
rect 37841 36805 37875 36839
rect 1685 36737 1719 36771
rect 2329 36737 2363 36771
rect 2973 36737 3007 36771
rect 3617 36737 3651 36771
rect 4261 36737 4295 36771
rect 4445 36737 4479 36771
rect 5733 36737 5767 36771
rect 5825 36737 5859 36771
rect 7113 36737 7147 36771
rect 8208 36737 8242 36771
rect 9781 36737 9815 36771
rect 10048 36737 10082 36771
rect 12173 36737 12207 36771
rect 13001 36737 13035 36771
rect 13257 36737 13291 36771
rect 14841 36737 14875 36771
rect 15097 36737 15131 36771
rect 17141 36737 17175 36771
rect 17408 36737 17442 36771
rect 18981 36737 19015 36771
rect 19165 36737 19199 36771
rect 19257 36737 19291 36771
rect 24777 36737 24811 36771
rect 27353 36737 27387 36771
rect 28457 36737 28491 36771
rect 31125 36737 31159 36771
rect 32321 36737 32355 36771
rect 32588 36737 32622 36771
rect 33977 36737 34011 36771
rect 34529 36737 34563 36771
rect 37473 36737 37507 36771
rect 37657 36737 37691 36771
rect 37933 36737 37967 36771
rect 7481 36669 7515 36703
rect 7941 36669 7975 36703
rect 12449 36669 12483 36703
rect 19717 36669 19751 36703
rect 19993 36669 20027 36703
rect 22293 36669 22327 36703
rect 25053 36669 25087 36703
rect 26525 36669 26559 36703
rect 30205 36669 30239 36703
rect 31585 36669 31619 36703
rect 34621 36669 34655 36703
rect 35449 36669 35483 36703
rect 1777 36533 1811 36567
rect 2421 36533 2455 36567
rect 11161 36533 11195 36567
rect 11897 36533 11931 36567
rect 16221 36533 16255 36567
rect 18521 36533 18555 36567
rect 18981 36533 19015 36567
rect 21465 36533 21499 36567
rect 33701 36533 33735 36567
rect 34805 36533 34839 36567
rect 36829 36533 36863 36567
rect 2605 36329 2639 36363
rect 3341 36329 3375 36363
rect 5273 36329 5307 36363
rect 6745 36329 6779 36363
rect 7757 36329 7791 36363
rect 10517 36329 10551 36363
rect 23351 36329 23385 36363
rect 30849 36329 30883 36363
rect 38025 36329 38059 36363
rect 8585 36261 8619 36295
rect 9321 36261 9355 36295
rect 13093 36261 13127 36295
rect 14749 36261 14783 36295
rect 19441 36261 19475 36295
rect 34069 36261 34103 36295
rect 38117 36261 38151 36295
rect 9781 36193 9815 36227
rect 9873 36193 9907 36227
rect 11069 36193 11103 36227
rect 11713 36193 11747 36227
rect 15209 36193 15243 36227
rect 15301 36193 15335 36227
rect 19901 36193 19935 36227
rect 19993 36193 20027 36227
rect 21557 36193 21591 36227
rect 21925 36193 21959 36227
rect 25421 36193 25455 36227
rect 25789 36193 25823 36227
rect 30021 36193 30055 36227
rect 31861 36193 31895 36227
rect 38301 36193 38335 36227
rect 2605 36125 2639 36159
rect 2789 36125 2823 36159
rect 3249 36125 3283 36159
rect 4353 36125 4387 36159
rect 5181 36125 5215 36159
rect 5917 36125 5951 36159
rect 6561 36125 6595 36159
rect 6654 36125 6688 36159
rect 7481 36125 7515 36159
rect 7573 36125 7607 36159
rect 11969 36125 12003 36159
rect 13553 36125 13587 36159
rect 13737 36125 13771 36159
rect 15945 36125 15979 36159
rect 18153 36125 18187 36159
rect 18245 36125 18279 36159
rect 18429 36125 18463 36159
rect 20637 36125 20671 36159
rect 20913 36125 20947 36159
rect 23857 36125 23891 36159
rect 24041 36125 24075 36159
rect 24593 36125 24627 36159
rect 24777 36125 24811 36159
rect 26893 36125 26927 36159
rect 28641 36125 28675 36159
rect 28733 36125 28767 36159
rect 28825 36125 28859 36159
rect 29009 36125 29043 36159
rect 29745 36125 29779 36159
rect 33885 36125 33919 36159
rect 34897 36125 34931 36159
rect 36093 36125 36127 36159
rect 36349 36125 36383 36159
rect 38025 36125 38059 36159
rect 4445 36057 4479 36091
rect 6101 36057 6135 36091
rect 8217 36057 8251 36091
rect 8401 36057 8435 36091
rect 10885 36057 10919 36091
rect 16212 36057 16246 36091
rect 18889 36057 18923 36091
rect 25906 36057 25940 36091
rect 27629 36057 27663 36091
rect 30757 36057 30791 36091
rect 32106 36057 32140 36091
rect 35173 36057 35207 36091
rect 9689 35989 9723 36023
rect 10977 35989 11011 36023
rect 13645 35989 13679 36023
rect 15117 35989 15151 36023
rect 17325 35989 17359 36023
rect 19809 35989 19843 36023
rect 23949 35989 23983 36023
rect 24869 35989 24903 36023
rect 25697 35989 25731 36023
rect 26065 35989 26099 36023
rect 28365 35989 28399 36023
rect 33241 35989 33275 36023
rect 37473 35989 37507 36023
rect 4445 35785 4479 35819
rect 6009 35785 6043 35819
rect 6653 35785 6687 35819
rect 9413 35785 9447 35819
rect 10333 35785 10367 35819
rect 14473 35785 14507 35819
rect 17417 35785 17451 35819
rect 32873 35785 32907 35819
rect 37565 35785 37599 35819
rect 10241 35717 10275 35751
rect 13645 35717 13679 35751
rect 21281 35717 21315 35751
rect 22293 35717 22327 35751
rect 23029 35717 23063 35751
rect 26479 35717 26513 35751
rect 33517 35717 33551 35751
rect 38025 35717 38059 35751
rect 3709 35649 3743 35683
rect 3893 35649 3927 35683
rect 4353 35649 4387 35683
rect 4537 35649 4571 35683
rect 4813 35649 4847 35683
rect 4997 35649 5031 35683
rect 5089 35649 5123 35683
rect 5733 35649 5767 35683
rect 6561 35649 6595 35683
rect 7297 35649 7331 35683
rect 7389 35649 7423 35683
rect 8300 35649 8334 35683
rect 11989 35649 12023 35683
rect 12081 35649 12115 35683
rect 12265 35649 12299 35683
rect 13277 35649 13311 35683
rect 13461 35649 13495 35683
rect 15669 35649 15703 35683
rect 15853 35649 15887 35683
rect 17509 35649 17543 35683
rect 21005 35649 21039 35683
rect 22017 35649 22051 35683
rect 23857 35649 23891 35683
rect 24409 35649 24443 35683
rect 24869 35649 24903 35683
rect 25513 35649 25547 35683
rect 26157 35649 26191 35683
rect 26249 35649 26283 35683
rect 26341 35649 26375 35683
rect 27905 35649 27939 35683
rect 29837 35649 29871 35683
rect 29929 35649 29963 35683
rect 31217 35649 31251 35683
rect 32321 35649 32355 35683
rect 33149 35649 33183 35683
rect 33333 35649 33367 35683
rect 34417 35649 34451 35683
rect 36645 35649 36679 35683
rect 37933 35649 37967 35683
rect 5457 35581 5491 35615
rect 6009 35581 6043 35615
rect 8033 35581 8067 35615
rect 10425 35581 10459 35615
rect 12725 35581 12759 35615
rect 14565 35581 14599 35615
rect 14749 35581 14783 35615
rect 15577 35581 15611 35615
rect 16313 35581 16347 35615
rect 17417 35581 17451 35615
rect 18521 35581 18555 35615
rect 18797 35581 18831 35615
rect 24133 35581 24167 35615
rect 26617 35581 26651 35615
rect 27813 35581 27847 35615
rect 28365 35581 28399 35615
rect 30389 35581 30423 35615
rect 31401 35581 31435 35615
rect 32597 35581 32631 35615
rect 34161 35581 34195 35615
rect 36921 35581 36955 35615
rect 38117 35581 38151 35615
rect 4813 35513 4847 35547
rect 5825 35513 5859 35547
rect 7573 35513 7607 35547
rect 33701 35513 33735 35547
rect 3709 35445 3743 35479
rect 9873 35445 9907 35479
rect 14105 35445 14139 35479
rect 16957 35445 16991 35479
rect 19901 35445 19935 35479
rect 23121 35445 23155 35479
rect 25973 35445 26007 35479
rect 28273 35445 28307 35479
rect 28641 35445 28675 35479
rect 30297 35445 30331 35479
rect 30481 35445 30515 35479
rect 32689 35445 32723 35479
rect 35541 35445 35575 35479
rect 36461 35445 36495 35479
rect 36829 35445 36863 35479
rect 5089 35241 5123 35275
rect 8401 35241 8435 35275
rect 9137 35241 9171 35275
rect 11529 35241 11563 35275
rect 14473 35241 14507 35275
rect 16589 35241 16623 35275
rect 18521 35241 18555 35275
rect 26801 35241 26835 35275
rect 27261 35241 27295 35275
rect 28457 35241 28491 35275
rect 30251 35241 30285 35275
rect 33057 35241 33091 35275
rect 33241 35241 33275 35275
rect 4813 35173 4847 35207
rect 18889 35173 18923 35207
rect 25145 35173 25179 35207
rect 26065 35173 26099 35207
rect 28089 35173 28123 35207
rect 28549 35173 28583 35207
rect 30389 35173 30423 35207
rect 5733 35105 5767 35139
rect 9597 35105 9631 35139
rect 9689 35105 9723 35139
rect 10885 35105 10919 35139
rect 17141 35105 17175 35139
rect 17877 35105 17911 35139
rect 18061 35105 18095 35139
rect 23673 35105 23707 35139
rect 24685 35105 24719 35139
rect 25237 35105 25271 35139
rect 28641 35105 28675 35139
rect 30481 35105 30515 35139
rect 31861 35105 31895 35139
rect 33885 35105 33919 35139
rect 34345 35105 34379 35139
rect 4261 35037 4295 35071
rect 4445 35037 4479 35071
rect 5917 35037 5951 35071
rect 6653 35037 6687 35071
rect 6837 35037 6871 35071
rect 7481 35037 7515 35071
rect 7665 35037 7699 35071
rect 8217 35037 8251 35071
rect 8401 35037 8435 35071
rect 10333 35037 10367 35071
rect 10425 35037 10459 35071
rect 11529 35037 11563 35071
rect 12357 35037 12391 35071
rect 13277 35037 13311 35071
rect 13553 35037 13587 35071
rect 15485 35037 15519 35071
rect 15669 35037 15703 35071
rect 15761 35037 15795 35071
rect 17049 35037 17083 35071
rect 17785 35037 17819 35071
rect 18521 35037 18555 35071
rect 18613 35037 18647 35071
rect 19625 35037 19659 35071
rect 19993 35037 20027 35071
rect 20637 35037 20671 35071
rect 20729 35037 20763 35071
rect 20821 35037 20855 35071
rect 21373 35037 21407 35071
rect 21649 35037 21683 35071
rect 22569 35037 22603 35071
rect 23489 35037 23523 35071
rect 24777 35037 24811 35071
rect 26341 35037 26375 35071
rect 26985 35037 27019 35071
rect 27077 35037 27111 35071
rect 31493 35037 31527 35071
rect 33977 35037 34011 35071
rect 34897 35037 34931 35071
rect 35081 35037 35115 35071
rect 35541 35037 35575 35071
rect 37473 35037 37507 35071
rect 37749 35037 37783 35071
rect 37841 35037 37875 35071
rect 4905 34969 4939 35003
rect 6929 34969 6963 35003
rect 7757 34969 7791 35003
rect 14381 34969 14415 35003
rect 16957 34969 16991 35003
rect 19441 34969 19475 35003
rect 21925 34969 21959 35003
rect 22845 34969 22879 35003
rect 25605 34969 25639 35003
rect 26065 34969 26099 35003
rect 30113 34969 30147 35003
rect 31309 34969 31343 35003
rect 32873 34969 32907 35003
rect 35786 34969 35820 35003
rect 37657 34969 37691 35003
rect 4353 34901 4387 34935
rect 5105 34901 5139 34935
rect 5273 34901 5307 34935
rect 6101 34901 6135 34935
rect 8585 34901 8619 34935
rect 9505 34901 9539 34935
rect 15301 34901 15335 34935
rect 18061 34901 18095 34935
rect 20453 34901 20487 34935
rect 26249 34901 26283 34935
rect 28917 34901 28951 34935
rect 30757 34901 30791 34935
rect 33057 34901 33091 34935
rect 35081 34901 35115 34935
rect 36921 34901 36955 34935
rect 38025 34901 38059 34935
rect 3617 34697 3651 34731
rect 4353 34697 4387 34731
rect 14657 34697 14691 34731
rect 15485 34697 15519 34731
rect 19993 34697 20027 34731
rect 21097 34697 21131 34731
rect 22661 34697 22695 34731
rect 34161 34697 34195 34731
rect 35357 34697 35391 34731
rect 36921 34697 36955 34731
rect 37473 34697 37507 34731
rect 11713 34629 11747 34663
rect 20453 34629 20487 34663
rect 23213 34629 23247 34663
rect 27905 34629 27939 34663
rect 33793 34629 33827 34663
rect 34989 34629 35023 34663
rect 3249 34561 3283 34595
rect 3525 34561 3559 34595
rect 4169 34561 4203 34595
rect 4353 34561 4387 34595
rect 4905 34561 4939 34595
rect 5089 34561 5123 34595
rect 5733 34561 5767 34595
rect 5825 34561 5859 34595
rect 6653 34561 6687 34595
rect 6837 34561 6871 34595
rect 7389 34561 7423 34595
rect 7573 34561 7607 34595
rect 8217 34561 8251 34595
rect 8401 34561 8435 34595
rect 9321 34561 9355 34595
rect 9505 34561 9539 34595
rect 10057 34561 10091 34595
rect 10149 34561 10183 34595
rect 11897 34561 11931 34595
rect 12173 34561 12207 34595
rect 13461 34561 13495 34595
rect 14197 34561 14231 34595
rect 14381 34561 14415 34595
rect 14473 34561 14507 34595
rect 15209 34561 15243 34595
rect 15393 34561 15427 34595
rect 17233 34561 17267 34595
rect 17325 34561 17359 34595
rect 17509 34561 17543 34595
rect 17601 34561 17635 34595
rect 18245 34561 18279 34595
rect 19625 34561 19659 34595
rect 19717 34561 19751 34595
rect 19809 34561 19843 34595
rect 20913 34561 20947 34595
rect 22017 34561 22051 34595
rect 22477 34561 22511 34595
rect 23121 34561 23155 34595
rect 23305 34561 23339 34595
rect 23857 34561 23891 34595
rect 24225 34561 24259 34595
rect 25697 34561 25731 34595
rect 25789 34561 25823 34595
rect 25973 34561 26007 34595
rect 26065 34561 26099 34595
rect 27445 34561 27479 34595
rect 27537 34561 27571 34595
rect 28549 34561 28583 34595
rect 30757 34561 30791 34595
rect 32505 34561 32539 34595
rect 33517 34561 33551 34595
rect 33610 34561 33644 34595
rect 33885 34561 33919 34595
rect 33982 34561 34016 34595
rect 34713 34561 34747 34595
rect 34806 34561 34840 34595
rect 35081 34561 35115 34595
rect 35178 34561 35212 34595
rect 36277 34561 36311 34595
rect 36370 34561 36404 34595
rect 36553 34561 36587 34595
rect 36645 34561 36679 34595
rect 36742 34561 36776 34595
rect 37841 34561 37875 34595
rect 5181 34493 5215 34527
rect 5917 34493 5951 34527
rect 9137 34493 9171 34527
rect 13737 34493 13771 34527
rect 20821 34493 20855 34527
rect 22293 34493 22327 34527
rect 27813 34493 27847 34527
rect 29561 34493 29595 34527
rect 31033 34493 31067 34527
rect 32689 34493 32723 34527
rect 32781 34493 32815 34527
rect 37933 34493 37967 34527
rect 38117 34493 38151 34527
rect 6653 34425 6687 34459
rect 8585 34425 8619 34459
rect 11989 34425 12023 34459
rect 12081 34425 12115 34459
rect 17049 34425 17083 34459
rect 18429 34425 18463 34459
rect 7481 34357 7515 34391
rect 10333 34357 10367 34391
rect 13277 34357 13311 34391
rect 13645 34357 13679 34391
rect 14197 34357 14231 34391
rect 20821 34357 20855 34391
rect 22109 34357 22143 34391
rect 25513 34357 25547 34391
rect 27261 34357 27295 34391
rect 30849 34357 30883 34391
rect 32321 34357 32355 34391
rect 5181 34153 5215 34187
rect 5917 34153 5951 34187
rect 7573 34153 7607 34187
rect 9597 34153 9631 34187
rect 14565 34153 14599 34187
rect 14749 34153 14783 34187
rect 21281 34153 21315 34187
rect 21925 34153 21959 34187
rect 23857 34153 23891 34187
rect 24041 34153 24075 34187
rect 24869 34153 24903 34187
rect 33701 34153 33735 34187
rect 5089 34085 5123 34119
rect 9873 34085 9907 34119
rect 17417 34085 17451 34119
rect 19809 34085 19843 34119
rect 25237 34085 25271 34119
rect 27905 34085 27939 34119
rect 30573 34085 30607 34119
rect 5273 34017 5307 34051
rect 8585 34017 8619 34051
rect 14381 34017 14415 34051
rect 15761 34017 15795 34051
rect 15853 34017 15887 34051
rect 16221 34017 16255 34051
rect 19441 34017 19475 34051
rect 21097 34017 21131 34051
rect 22109 34017 22143 34051
rect 22937 34017 22971 34051
rect 23121 34017 23155 34051
rect 23765 34017 23799 34051
rect 31953 34017 31987 34051
rect 34253 34017 34287 34051
rect 36829 34017 36863 34051
rect 4077 33949 4111 33983
rect 4353 33949 4387 33983
rect 4537 33949 4571 33983
rect 4997 33949 5031 33983
rect 5733 33949 5767 33983
rect 5917 33949 5951 33983
rect 7389 33949 7423 33983
rect 7481 33949 7515 33983
rect 8401 33949 8435 33983
rect 9505 33949 9539 33983
rect 9597 33949 9631 33983
rect 10333 33949 10367 33983
rect 10701 33949 10735 33983
rect 11069 33949 11103 33983
rect 11989 33949 12023 33983
rect 12357 33949 12391 33983
rect 12541 33949 12575 33983
rect 13369 33949 13403 33983
rect 13461 33949 13495 33983
rect 13645 33949 13679 33983
rect 13737 33949 13771 33983
rect 14565 33949 14599 33983
rect 15485 33949 15519 33983
rect 15669 33949 15703 33983
rect 16037 33949 16071 33983
rect 16681 33949 16715 33983
rect 17785 33949 17819 33983
rect 18521 33949 18555 33983
rect 18705 33949 18739 33983
rect 19625 33949 19659 33983
rect 19717 33949 19751 33983
rect 19901 33949 19935 33983
rect 21281 33949 21315 33983
rect 21925 33949 21959 33983
rect 22201 33949 22235 33983
rect 22845 33949 22879 33983
rect 23857 33949 23891 33983
rect 24961 33949 24995 33983
rect 25053 33949 25087 33983
rect 26065 33949 26099 33983
rect 26157 33949 26191 33983
rect 26249 33949 26283 33983
rect 26341 33949 26375 33983
rect 27077 33949 27111 33983
rect 27261 33949 27295 33983
rect 27353 33949 27387 33983
rect 28089 33949 28123 33983
rect 28181 33949 28215 33983
rect 28549 33949 28583 33983
rect 29009 33949 29043 33983
rect 29193 33949 29227 33983
rect 29837 33949 29871 33983
rect 30297 33949 30331 33983
rect 31401 33949 31435 33983
rect 33057 33949 33091 33983
rect 33195 33949 33229 33983
rect 33333 33949 33367 33983
rect 33425 33949 33459 33983
rect 33522 33949 33556 33983
rect 34161 33949 34195 33983
rect 34345 33949 34379 33983
rect 34897 33949 34931 33983
rect 35045 33949 35079 33983
rect 35362 33949 35396 33983
rect 36001 33949 36035 33983
rect 36185 33949 36219 33983
rect 37096 33949 37130 33983
rect 6561 33881 6595 33915
rect 6745 33881 6779 33915
rect 6929 33881 6963 33915
rect 8217 33881 8251 33915
rect 13185 33881 13219 33915
rect 14289 33881 14323 33915
rect 17601 33881 17635 33915
rect 21005 33881 21039 33915
rect 23581 33881 23615 33915
rect 24593 33881 24627 33915
rect 28457 33881 28491 33915
rect 30021 33881 30055 33915
rect 35173 33881 35207 33915
rect 35265 33881 35299 33915
rect 4445 33813 4479 33847
rect 6101 33813 6135 33847
rect 7757 33813 7791 33847
rect 16865 33813 16899 33847
rect 17693 33813 17727 33847
rect 17969 33813 18003 33847
rect 18889 33813 18923 33847
rect 21465 33813 21499 33847
rect 22385 33813 22419 33847
rect 23121 33813 23155 33847
rect 25881 33813 25915 33847
rect 26893 33813 26927 33847
rect 29101 33813 29135 33847
rect 35541 33813 35575 33847
rect 36093 33813 36127 33847
rect 38209 33813 38243 33847
rect 4537 33609 4571 33643
rect 9597 33609 9631 33643
rect 9965 33609 9999 33643
rect 13553 33609 13587 33643
rect 15117 33609 15151 33643
rect 16957 33609 16991 33643
rect 17417 33609 17451 33643
rect 21465 33609 21499 33643
rect 28549 33609 28583 33643
rect 30205 33609 30239 33643
rect 30573 33609 30607 33643
rect 35633 33609 35667 33643
rect 7932 33541 7966 33575
rect 10793 33541 10827 33575
rect 11161 33541 11195 33575
rect 12449 33541 12483 33575
rect 15485 33541 15519 33575
rect 15577 33541 15611 33575
rect 17325 33541 17359 33575
rect 23673 33541 23707 33575
rect 25697 33541 25731 33575
rect 27169 33541 27203 33575
rect 29377 33541 29411 33575
rect 33149 33541 33183 33575
rect 35357 33541 35391 33575
rect 3893 33473 3927 33507
rect 4077 33473 4111 33507
rect 4353 33473 4387 33507
rect 4537 33473 4571 33507
rect 5181 33473 5215 33507
rect 5365 33473 5399 33507
rect 5825 33473 5859 33507
rect 6009 33473 6043 33507
rect 6837 33473 6871 33507
rect 7021 33473 7055 33507
rect 7573 33473 7607 33507
rect 10977 33473 11011 33507
rect 11713 33473 11747 33507
rect 11989 33473 12023 33507
rect 12633 33473 12667 33507
rect 13737 33473 13771 33507
rect 13921 33473 13955 33507
rect 14013 33473 14047 33507
rect 15393 33473 15427 33507
rect 15761 33473 15795 33507
rect 15853 33473 15887 33507
rect 17233 33473 17267 33507
rect 18521 33473 18555 33507
rect 19809 33473 19843 33507
rect 21005 33473 21039 33507
rect 21281 33473 21315 33507
rect 22017 33495 22051 33529
rect 22201 33473 22235 33507
rect 22293 33473 22327 33507
rect 22385 33473 22419 33507
rect 22569 33473 22603 33507
rect 23949 33473 23983 33507
rect 24593 33473 24627 33507
rect 24961 33473 24995 33507
rect 25053 33473 25087 33507
rect 26157 33473 26191 33507
rect 27445 33473 27479 33507
rect 28181 33473 28215 33507
rect 29561 33473 29595 33507
rect 30849 33473 30883 33507
rect 30941 33473 30975 33507
rect 31033 33473 31067 33507
rect 31217 33473 31251 33507
rect 32873 33473 32907 33507
rect 33021 33473 33055 33507
rect 33249 33473 33283 33507
rect 33338 33473 33372 33507
rect 33977 33473 34011 33507
rect 34125 33473 34159 33507
rect 34253 33473 34287 33507
rect 34345 33473 34379 33507
rect 34442 33473 34476 33507
rect 35081 33473 35115 33507
rect 35265 33473 35299 33507
rect 35449 33473 35483 33507
rect 36093 33473 36127 33507
rect 36241 33473 36275 33507
rect 36369 33473 36403 33507
rect 36461 33473 36495 33507
rect 36599 33473 36633 33507
rect 37473 33473 37507 33507
rect 37657 33473 37691 33507
rect 37749 33473 37783 33507
rect 37841 33473 37875 33507
rect 7665 33405 7699 33439
rect 10057 33405 10091 33439
rect 10149 33405 10183 33439
rect 13829 33405 13863 33439
rect 17693 33405 17727 33439
rect 18613 33405 18647 33439
rect 19993 33405 20027 33439
rect 21097 33405 21131 33439
rect 23765 33405 23799 33439
rect 25973 33405 26007 33439
rect 27261 33405 27295 33439
rect 28273 33405 28307 33439
rect 7205 33337 7239 33371
rect 9045 33337 9079 33371
rect 11805 33337 11839 33371
rect 27629 33337 27663 33371
rect 33517 33337 33551 33371
rect 3893 33269 3927 33303
rect 4813 33269 4847 33303
rect 5273 33269 5307 33303
rect 5825 33269 5859 33303
rect 11713 33269 11747 33303
rect 12725 33269 12759 33303
rect 17601 33269 17635 33303
rect 18705 33269 18739 33303
rect 18889 33269 18923 33303
rect 21189 33269 21223 33303
rect 22753 33269 22787 33303
rect 23949 33269 23983 33303
rect 24133 33269 24167 33303
rect 25053 33269 25087 33303
rect 25237 33269 25271 33303
rect 25789 33269 25823 33303
rect 26341 33269 26375 33303
rect 27169 33269 27203 33303
rect 28181 33269 28215 33303
rect 29653 33269 29687 33303
rect 34621 33269 34655 33303
rect 36737 33269 36771 33303
rect 38025 33269 38059 33303
rect 8125 33065 8159 33099
rect 12633 33065 12667 33099
rect 13277 33065 13311 33099
rect 14381 33065 14415 33099
rect 15301 33065 15335 33099
rect 15577 33065 15611 33099
rect 16037 33065 16071 33099
rect 16497 33065 16531 33099
rect 17417 33065 17451 33099
rect 17601 33065 17635 33099
rect 20361 33065 20395 33099
rect 22385 33065 22419 33099
rect 23581 33065 23615 33099
rect 24041 33065 24075 33099
rect 26433 33065 26467 33099
rect 27629 33065 27663 33099
rect 31401 33065 31435 33099
rect 33609 33065 33643 33099
rect 5825 32997 5859 33031
rect 7665 32997 7699 33031
rect 11713 32997 11747 33031
rect 12817 32997 12851 33031
rect 21603 32997 21637 33031
rect 24593 32997 24627 33031
rect 26341 32997 26375 33031
rect 27813 32997 27847 33031
rect 34253 32997 34287 33031
rect 5273 32929 5307 32963
rect 8585 32929 8619 32963
rect 9413 32929 9447 32963
rect 11345 32929 11379 32963
rect 12449 32929 12483 32963
rect 14381 32929 14415 32963
rect 15209 32929 15243 32963
rect 16129 32929 16163 32963
rect 22753 32929 22787 32963
rect 23765 32929 23799 32963
rect 30021 32929 30055 32963
rect 30389 32929 30423 32963
rect 34345 32929 34379 32963
rect 4537 32861 4571 32895
rect 4721 32861 4755 32895
rect 5181 32861 5215 32895
rect 5365 32861 5399 32895
rect 5825 32861 5859 32895
rect 6009 32861 6043 32895
rect 6561 32861 6595 32895
rect 7297 32861 7331 32895
rect 8309 32861 8343 32895
rect 8493 32861 8527 32895
rect 9321 32861 9355 32895
rect 9505 32861 9539 32895
rect 9597 32861 9631 32895
rect 10425 32861 10459 32895
rect 10701 32861 10735 32895
rect 11529 32861 11563 32895
rect 11621 32861 11655 32895
rect 11805 32861 11839 32895
rect 12633 32861 12667 32895
rect 13461 32861 13495 32895
rect 13737 32861 13771 32895
rect 14289 32861 14323 32895
rect 15393 32861 15427 32895
rect 16037 32861 16071 32895
rect 16313 32861 16347 32895
rect 17049 32861 17083 32895
rect 18061 32861 18095 32895
rect 19809 32861 19843 32895
rect 20177 32861 20211 32895
rect 20821 32861 20855 32895
rect 21005 32861 21039 32895
rect 21454 32861 21488 32895
rect 21741 32861 21775 32895
rect 21937 32855 21971 32889
rect 22569 32861 22603 32895
rect 22845 32861 22879 32895
rect 23581 32861 23615 32895
rect 23857 32861 23891 32895
rect 24869 32861 24903 32895
rect 24961 32861 24995 32895
rect 25053 32861 25087 32895
rect 25237 32861 25271 32895
rect 25973 32861 26007 32895
rect 27445 32861 27479 32895
rect 27537 32861 27571 32895
rect 28365 32861 28399 32895
rect 28825 32861 28859 32895
rect 29929 32861 29963 32895
rect 30205 32861 30239 32895
rect 31953 32861 31987 32895
rect 32045 32861 32079 32895
rect 32321 32861 32355 32895
rect 32505 32861 32539 32895
rect 32965 32861 32999 32895
rect 33058 32861 33092 32895
rect 33241 32861 33275 32895
rect 33333 32861 33367 32895
rect 33430 32861 33464 32895
rect 34069 32861 34103 32895
rect 34161 32861 34195 32895
rect 34897 32861 34931 32895
rect 35081 32861 35115 32895
rect 35541 32861 35575 32895
rect 35634 32861 35668 32895
rect 36047 32861 36081 32895
rect 36829 32861 36863 32895
rect 7481 32793 7515 32827
rect 12357 32793 12391 32827
rect 15117 32793 15151 32827
rect 18337 32793 18371 32827
rect 19993 32793 20027 32827
rect 20085 32793 20119 32827
rect 35817 32793 35851 32827
rect 35909 32793 35943 32827
rect 37096 32793 37130 32827
rect 4629 32725 4663 32759
rect 6745 32725 6779 32759
rect 9137 32725 9171 32759
rect 13645 32725 13679 32759
rect 14657 32725 14691 32759
rect 17417 32725 17451 32759
rect 20913 32725 20947 32759
rect 21833 32725 21867 32759
rect 28457 32725 28491 32759
rect 34989 32725 35023 32759
rect 36185 32725 36219 32759
rect 38209 32725 38243 32759
rect 4169 32521 4203 32555
rect 19625 32521 19659 32555
rect 20269 32521 20303 32555
rect 22293 32521 22327 32555
rect 25513 32521 25547 32555
rect 37473 32521 37507 32555
rect 37841 32521 37875 32555
rect 7840 32453 7874 32487
rect 10057 32453 10091 32487
rect 11805 32453 11839 32487
rect 11989 32453 12023 32487
rect 15209 32453 15243 32487
rect 17969 32453 18003 32487
rect 18061 32453 18095 32487
rect 20821 32453 20855 32487
rect 27905 32453 27939 32487
rect 34161 32453 34195 32487
rect 37933 32453 37967 32487
rect 4077 32385 4111 32419
rect 4721 32385 4755 32419
rect 4905 32385 4939 32419
rect 5825 32385 5859 32419
rect 5917 32385 5951 32419
rect 6009 32385 6043 32419
rect 6745 32385 6779 32419
rect 6929 32385 6963 32419
rect 9781 32385 9815 32419
rect 9965 32385 9999 32419
rect 10149 32385 10183 32419
rect 10977 32395 11011 32429
rect 11161 32385 11195 32419
rect 12265 32385 12299 32419
rect 12909 32385 12943 32419
rect 13921 32385 13955 32419
rect 15485 32385 15519 32419
rect 16957 32385 16991 32419
rect 17141 32385 17175 32419
rect 17785 32385 17819 32419
rect 18153 32385 18187 32419
rect 19441 32385 19475 32419
rect 19717 32385 19751 32419
rect 20177 32385 20211 32419
rect 20361 32385 20395 32419
rect 21005 32385 21039 32419
rect 21097 32385 21131 32419
rect 22477 32385 22511 32419
rect 22661 32385 22695 32419
rect 22937 32385 22971 32419
rect 23857 32385 23891 32419
rect 24961 32385 24995 32419
rect 25329 32385 25363 32419
rect 26157 32385 26191 32419
rect 27629 32385 27663 32419
rect 28549 32385 28583 32419
rect 28696 32385 28730 32419
rect 29745 32385 29779 32419
rect 29929 32385 29963 32419
rect 30665 32385 30699 32419
rect 31033 32385 31067 32419
rect 31585 32385 31619 32419
rect 31769 32385 31803 32419
rect 32321 32385 32355 32419
rect 32505 32385 32539 32419
rect 33057 32385 33091 32419
rect 33885 32385 33919 32419
rect 34069 32385 34103 32419
rect 34253 32385 34287 32419
rect 35081 32385 35115 32419
rect 35909 32385 35943 32419
rect 36093 32385 36127 32419
rect 36185 32385 36219 32419
rect 36277 32385 36311 32419
rect 7573 32317 7607 32351
rect 13093 32317 13127 32351
rect 14197 32317 14231 32351
rect 15301 32317 15335 32351
rect 22753 32317 22787 32351
rect 24133 32317 24167 32351
rect 24869 32317 24903 32351
rect 26433 32317 26467 32351
rect 28917 32317 28951 32351
rect 29009 32317 29043 32351
rect 32781 32317 32815 32351
rect 34989 32317 35023 32351
rect 38025 32317 38059 32351
rect 7113 32249 7147 32283
rect 10701 32249 10735 32283
rect 21281 32249 21315 32283
rect 22569 32249 22603 32283
rect 28825 32249 28859 32283
rect 34437 32249 34471 32283
rect 4721 32181 4755 32215
rect 8953 32181 8987 32215
rect 10333 32181 10367 32215
rect 11069 32181 11103 32215
rect 11955 32181 11989 32215
rect 15209 32181 15243 32215
rect 15669 32181 15703 32215
rect 16957 32181 16991 32215
rect 17325 32181 17359 32215
rect 18337 32181 18371 32215
rect 19257 32181 19291 32215
rect 21005 32181 21039 32215
rect 25329 32181 25363 32215
rect 30113 32181 30147 32215
rect 32413 32181 32447 32215
rect 33149 32181 33183 32215
rect 35449 32181 35483 32215
rect 36461 32181 36495 32215
rect 7665 31977 7699 32011
rect 8401 31977 8435 32011
rect 11805 31977 11839 32011
rect 14933 31977 14967 32011
rect 16221 31977 16255 32011
rect 17141 31977 17175 32011
rect 19993 31977 20027 32011
rect 20361 31977 20395 32011
rect 21189 31977 21223 32011
rect 24777 31977 24811 32011
rect 28457 31977 28491 32011
rect 33609 31977 33643 32011
rect 6837 31909 6871 31943
rect 13461 31909 13495 31943
rect 15393 31909 15427 31943
rect 16497 31909 16531 31943
rect 18521 31909 18555 31943
rect 21373 31909 21407 31943
rect 26157 31909 26191 31943
rect 26249 31909 26283 31943
rect 29009 31909 29043 31943
rect 34069 31909 34103 31943
rect 36277 31909 36311 31943
rect 36645 31909 36679 31943
rect 4445 31841 4479 31875
rect 8217 31841 8251 31875
rect 9413 31841 9447 31875
rect 9505 31841 9539 31875
rect 15025 31841 15059 31875
rect 20085 31841 20119 31875
rect 23305 31841 23339 31875
rect 24961 31841 24995 31875
rect 25053 31841 25087 31875
rect 25145 31841 25179 31875
rect 25237 31841 25271 31875
rect 25789 31841 25823 31875
rect 26341 31841 26375 31875
rect 29837 31841 29871 31875
rect 30389 31841 30423 31875
rect 31125 31841 31159 31875
rect 34897 31841 34931 31875
rect 36829 31841 36863 31875
rect 4353 31773 4387 31807
rect 4537 31773 4571 31807
rect 4905 31773 4939 31807
rect 5181 31773 5215 31807
rect 5365 31773 5399 31807
rect 5825 31773 5859 31807
rect 6009 31773 6043 31807
rect 6561 31773 6595 31807
rect 6653 31773 6687 31807
rect 7297 31773 7331 31807
rect 8401 31773 8435 31807
rect 9597 31773 9631 31807
rect 9689 31773 9723 31807
rect 10425 31773 10459 31807
rect 10609 31773 10643 31807
rect 10701 31773 10735 31807
rect 10793 31773 10827 31807
rect 11529 31773 11563 31807
rect 11713 31773 11747 31807
rect 12449 31773 12483 31807
rect 13277 31773 13311 31807
rect 14289 31773 14323 31807
rect 14473 31773 14507 31807
rect 15209 31773 15243 31807
rect 16129 31773 16163 31807
rect 16313 31773 16347 31807
rect 17969 31773 18003 31807
rect 18337 31773 18371 31807
rect 19809 31773 19843 31807
rect 21005 31773 21039 31807
rect 21097 31773 21131 31807
rect 21925 31773 21959 31807
rect 22109 31773 22143 31807
rect 22753 31773 22787 31807
rect 22937 31773 22971 31807
rect 23949 31773 23983 31807
rect 27445 31773 27479 31807
rect 28641 31773 28675 31807
rect 28825 31773 28859 31807
rect 29745 31773 29779 31807
rect 30021 31773 30055 31807
rect 31493 31773 31527 31807
rect 32137 31773 32171 31807
rect 32965 31773 32999 31807
rect 33058 31773 33092 31807
rect 33430 31773 33464 31807
rect 34345 31773 34379 31807
rect 35164 31773 35198 31807
rect 37096 31773 37130 31807
rect 5273 31705 5307 31739
rect 7481 31705 7515 31739
rect 8125 31705 8159 31739
rect 14933 31705 14967 31739
rect 16957 31705 16991 31739
rect 18153 31705 18187 31739
rect 18245 31705 18279 31739
rect 27721 31705 27755 31739
rect 28365 31705 28399 31739
rect 33241 31705 33275 31739
rect 33333 31705 33367 31739
rect 34069 31705 34103 31739
rect 34253 31705 34287 31739
rect 5917 31637 5951 31671
rect 8585 31637 8619 31671
rect 9229 31637 9263 31671
rect 10977 31637 11011 31671
rect 14381 31637 14415 31671
rect 17157 31637 17191 31671
rect 17325 31637 17359 31671
rect 22293 31637 22327 31671
rect 23949 31637 23983 31671
rect 26617 31637 26651 31671
rect 31886 31637 31920 31671
rect 38209 31637 38243 31671
rect 37473 31433 37507 31467
rect 7389 31365 7423 31399
rect 16129 31365 16163 31399
rect 18398 31365 18432 31399
rect 30113 31365 30147 31399
rect 30297 31365 30331 31399
rect 33149 31365 33183 31399
rect 33241 31365 33275 31399
rect 34253 31365 34287 31399
rect 35357 31365 35391 31399
rect 37841 31365 37875 31399
rect 5181 31297 5215 31331
rect 5365 31297 5399 31331
rect 5825 31297 5859 31331
rect 6009 31297 6043 31331
rect 7113 31297 7147 31331
rect 7297 31297 7331 31331
rect 7941 31297 7975 31331
rect 8033 31297 8067 31331
rect 8217 31297 8251 31331
rect 8861 31297 8895 31331
rect 9045 31297 9079 31331
rect 9689 31297 9723 31331
rect 10149 31297 10183 31331
rect 10885 31297 10919 31331
rect 11069 31297 11103 31331
rect 12357 31297 12391 31331
rect 12541 31297 12575 31331
rect 12909 31297 12943 31331
rect 13369 31297 13403 31331
rect 13645 31297 13679 31331
rect 13921 31297 13955 31331
rect 14013 31297 14047 31331
rect 14841 31297 14875 31331
rect 15301 31297 15335 31331
rect 16865 31297 16899 31331
rect 20260 31297 20294 31331
rect 22477 31297 22511 31331
rect 22661 31297 22695 31331
rect 23305 31297 23339 31331
rect 25513 31297 25547 31331
rect 25605 31297 25639 31331
rect 25973 31297 26007 31331
rect 27261 31297 27295 31331
rect 28089 31297 28123 31331
rect 31033 31297 31067 31331
rect 31493 31297 31527 31331
rect 32873 31297 32907 31331
rect 32966 31297 33000 31331
rect 33338 31297 33372 31331
rect 33977 31297 34011 31331
rect 34125 31297 34159 31331
rect 34345 31297 34379 31331
rect 34442 31297 34476 31331
rect 35081 31297 35115 31331
rect 35265 31297 35299 31331
rect 35449 31297 35483 31331
rect 36185 31297 36219 31331
rect 36333 31297 36367 31331
rect 36461 31297 36495 31331
rect 36553 31297 36587 31331
rect 36650 31297 36684 31331
rect 37933 31297 37967 31331
rect 5917 31229 5951 31263
rect 8677 31229 8711 31263
rect 9873 31229 9907 31263
rect 9965 31229 9999 31263
rect 11161 31229 11195 31263
rect 14197 31229 14231 31263
rect 15393 31229 15427 31263
rect 17049 31229 17083 31263
rect 18153 31229 18187 31263
rect 19993 31229 20027 31263
rect 23765 31229 23799 31263
rect 27537 31229 27571 31263
rect 28549 31229 28583 31263
rect 31585 31229 31619 31263
rect 38117 31229 38151 31263
rect 9781 31161 9815 31195
rect 33517 31161 33551 31195
rect 5181 31093 5215 31127
rect 9505 31093 9539 31127
rect 16221 31093 16255 31127
rect 19533 31093 19567 31127
rect 21373 31093 21407 31127
rect 22753 31093 22787 31127
rect 25973 31093 26007 31127
rect 26157 31093 26191 31127
rect 30297 31093 30331 31127
rect 30481 31093 30515 31127
rect 34621 31093 34655 31127
rect 35633 31093 35667 31127
rect 36829 31093 36863 31127
rect 5917 30889 5951 30923
rect 6469 30889 6503 30923
rect 8585 30889 8619 30923
rect 11529 30889 11563 30923
rect 14657 30889 14691 30923
rect 19625 30889 19659 30923
rect 20177 30889 20211 30923
rect 31217 30889 31251 30923
rect 36553 30889 36587 30923
rect 38117 30889 38151 30923
rect 11713 30821 11747 30855
rect 13001 30821 13035 30855
rect 23029 30821 23063 30855
rect 26249 30821 26283 30855
rect 28549 30821 28583 30855
rect 4905 30753 4939 30787
rect 9597 30753 9631 30787
rect 10425 30753 10459 30787
rect 13645 30753 13679 30787
rect 15669 30753 15703 30787
rect 20637 30753 20671 30787
rect 20729 30753 20763 30787
rect 23581 30753 23615 30787
rect 24593 30753 24627 30787
rect 24777 30753 24811 30787
rect 25053 30753 25087 30787
rect 27261 30753 27295 30787
rect 29745 30753 29779 30787
rect 30205 30753 30239 30787
rect 30297 30753 30331 30787
rect 32229 30753 32263 30787
rect 34253 30753 34287 30787
rect 37105 30753 37139 30787
rect 37565 30753 37599 30787
rect 38301 30753 38335 30787
rect 5181 30685 5215 30719
rect 5365 30685 5399 30719
rect 5825 30685 5859 30719
rect 6469 30685 6503 30719
rect 6745 30685 6779 30719
rect 7205 30685 7239 30719
rect 7472 30685 7506 30719
rect 9229 30685 9263 30719
rect 9413 30685 9447 30719
rect 10057 30685 10091 30719
rect 10241 30685 10275 30719
rect 10333 30685 10367 30719
rect 10609 30685 10643 30719
rect 12357 30685 12391 30719
rect 12541 30685 12575 30719
rect 13185 30685 13219 30719
rect 13369 30685 13403 30719
rect 13487 30685 13521 30719
rect 15301 30685 15335 30719
rect 15485 30685 15519 30719
rect 16129 30685 16163 30719
rect 18705 30685 18739 30719
rect 20545 30685 20579 30719
rect 21833 30685 21867 30719
rect 21925 30685 21959 30719
rect 22017 30685 22051 30719
rect 22109 30685 22143 30719
rect 22661 30685 22695 30719
rect 23213 30685 23247 30719
rect 23673 30685 23707 30719
rect 25145 30685 25179 30719
rect 26065 30685 26099 30719
rect 26341 30685 26375 30719
rect 27169 30685 27203 30719
rect 27353 30685 27387 30719
rect 27445 30685 27479 30719
rect 27537 30685 27571 30719
rect 28457 30685 28491 30719
rect 28733 30685 28767 30719
rect 31769 30685 31803 30719
rect 31861 30685 31895 30719
rect 32137 30685 32171 30719
rect 32781 30685 32815 30719
rect 32874 30685 32908 30719
rect 33246 30685 33280 30719
rect 34069 30685 34103 30719
rect 34345 30685 34379 30719
rect 34897 30685 34931 30719
rect 35173 30685 35207 30719
rect 35265 30685 35299 30719
rect 35909 30685 35943 30719
rect 36057 30685 36091 30719
rect 36415 30685 36449 30719
rect 37197 30685 37231 30719
rect 38025 30685 38059 30719
rect 5733 30617 5767 30651
rect 11345 30617 11379 30651
rect 11545 30617 11579 30651
rect 12173 30617 12207 30651
rect 13277 30617 13311 30651
rect 14473 30617 14507 30651
rect 16396 30617 16430 30651
rect 17969 30617 18003 30651
rect 19533 30617 19567 30651
rect 33057 30617 33091 30651
rect 33149 30617 33183 30651
rect 35081 30617 35115 30651
rect 36185 30617 36219 30651
rect 36277 30617 36311 30651
rect 5273 30549 5307 30583
rect 6653 30549 6687 30583
rect 10793 30549 10827 30583
rect 14673 30549 14707 30583
rect 14841 30549 14875 30583
rect 17509 30549 17543 30583
rect 21649 30549 21683 30583
rect 25881 30549 25915 30583
rect 26893 30549 26927 30583
rect 28917 30549 28951 30583
rect 29929 30549 29963 30583
rect 33425 30549 33459 30583
rect 33885 30549 33919 30583
rect 35449 30549 35483 30583
rect 38301 30549 38335 30583
rect 22109 30345 22143 30379
rect 34161 30345 34195 30379
rect 37841 30345 37875 30379
rect 10977 30277 11011 30311
rect 11805 30277 11839 30311
rect 13369 30277 13403 30311
rect 14381 30277 14415 30311
rect 17141 30277 17175 30311
rect 24593 30277 24627 30311
rect 25145 30277 25179 30311
rect 31217 30277 31251 30311
rect 32321 30277 32355 30311
rect 33793 30277 33827 30311
rect 37933 30277 37967 30311
rect 6745 30209 6779 30243
rect 6929 30209 6963 30243
rect 7656 30209 7690 30243
rect 9689 30209 9723 30243
rect 9781 30209 9815 30243
rect 9965 30209 9999 30243
rect 10149 30209 10183 30243
rect 11713 30209 11747 30243
rect 11897 30209 11931 30243
rect 13645 30209 13679 30243
rect 14289 30209 14323 30243
rect 14933 30209 14967 30243
rect 15200 30209 15234 30243
rect 16865 30209 16899 30243
rect 17049 30209 17083 30243
rect 17233 30209 17267 30243
rect 18153 30209 18187 30243
rect 20269 30209 20303 30243
rect 20913 30209 20947 30243
rect 21005 30209 21039 30243
rect 21281 30209 21315 30243
rect 21373 30209 21407 30243
rect 22293 30209 22327 30243
rect 22477 30209 22511 30243
rect 23029 30209 23063 30243
rect 23213 30209 23247 30243
rect 23949 30209 23983 30243
rect 24777 30209 24811 30243
rect 27445 30209 27479 30243
rect 27537 30209 27571 30243
rect 29745 30209 29779 30243
rect 31493 30209 31527 30243
rect 33517 30209 33551 30243
rect 33665 30209 33699 30243
rect 33885 30209 33919 30243
rect 34023 30209 34057 30243
rect 35081 30209 35115 30243
rect 35348 30209 35382 30243
rect 7389 30141 7423 30175
rect 10609 30141 10643 30175
rect 12541 30141 12575 30175
rect 12633 30141 12667 30175
rect 12725 30141 12759 30175
rect 12817 30141 12851 30175
rect 13553 30141 13587 30175
rect 18429 30141 18463 30175
rect 25605 30141 25639 30175
rect 26065 30141 26099 30175
rect 27353 30141 27387 30175
rect 27629 30141 27663 30175
rect 28181 30141 28215 30175
rect 28733 30141 28767 30175
rect 29101 30141 29135 30175
rect 29653 30141 29687 30175
rect 30205 30141 30239 30175
rect 31401 30141 31435 30175
rect 32689 30141 32723 30175
rect 38117 30141 38151 30175
rect 17417 30073 17451 30107
rect 25881 30073 25915 30107
rect 28549 30073 28583 30107
rect 28641 30073 28675 30107
rect 30113 30073 30147 30107
rect 32597 30073 32631 30107
rect 6745 30005 6779 30039
rect 8769 30005 8803 30039
rect 9413 30005 9447 30039
rect 9873 30005 9907 30039
rect 10977 30005 11011 30039
rect 11161 30005 11195 30039
rect 12357 30005 12391 30039
rect 13369 30005 13403 30039
rect 13829 30005 13863 30039
rect 16313 30005 16347 30039
rect 19717 30005 19751 30039
rect 24041 30005 24075 30039
rect 27169 30005 27203 30039
rect 30481 30005 30515 30039
rect 31217 30005 31251 30039
rect 31677 30005 31711 30039
rect 32459 30005 32493 30039
rect 32781 30005 32815 30039
rect 36461 30005 36495 30039
rect 37473 30005 37507 30039
rect 8125 29801 8159 29835
rect 10333 29801 10367 29835
rect 11437 29801 11471 29835
rect 13553 29801 13587 29835
rect 16221 29801 16255 29835
rect 27353 29801 27387 29835
rect 30297 29801 30331 29835
rect 34989 29801 35023 29835
rect 38209 29801 38243 29835
rect 6837 29733 6871 29767
rect 10885 29733 10919 29767
rect 13737 29733 13771 29767
rect 23581 29733 23615 29767
rect 30757 29733 30791 29767
rect 8585 29665 8619 29699
rect 9137 29665 9171 29699
rect 9597 29665 9631 29699
rect 10517 29665 10551 29699
rect 11621 29665 11655 29699
rect 11713 29665 11747 29699
rect 12817 29665 12851 29699
rect 21925 29665 21959 29699
rect 30389 29665 30423 29699
rect 34253 29665 34287 29699
rect 34989 29665 35023 29699
rect 6837 29597 6871 29631
rect 7021 29597 7055 29631
rect 7481 29597 7515 29631
rect 7665 29597 7699 29631
rect 8309 29597 8343 29631
rect 8493 29597 8527 29631
rect 9505 29597 9539 29631
rect 10241 29597 10275 29631
rect 10701 29597 10735 29631
rect 11805 29597 11839 29631
rect 11897 29597 11931 29631
rect 15669 29597 15703 29631
rect 15945 29597 15979 29631
rect 16037 29597 16071 29631
rect 17233 29597 17267 29631
rect 19441 29597 19475 29631
rect 21189 29597 21223 29631
rect 21741 29597 21775 29631
rect 22201 29597 22235 29631
rect 22753 29597 22787 29631
rect 23489 29597 23523 29631
rect 23673 29597 23707 29631
rect 23765 29597 23799 29631
rect 23949 29597 23983 29631
rect 24593 29597 24627 29631
rect 25053 29597 25087 29631
rect 26065 29597 26099 29631
rect 27537 29597 27571 29631
rect 27629 29597 27663 29631
rect 28733 29597 28767 29631
rect 29009 29597 29043 29631
rect 30573 29597 30607 29631
rect 31309 29597 31343 29631
rect 31953 29597 31987 29631
rect 33057 29597 33091 29631
rect 33150 29597 33184 29631
rect 33333 29597 33367 29631
rect 33522 29597 33556 29631
rect 34161 29597 34195 29631
rect 34897 29597 34931 29631
rect 35725 29597 35759 29631
rect 35818 29597 35852 29631
rect 36093 29597 36127 29631
rect 36231 29597 36265 29631
rect 36829 29597 36863 29631
rect 37096 29597 37130 29631
rect 7573 29529 7607 29563
rect 12449 29529 12483 29563
rect 12633 29529 12667 29563
rect 13369 29529 13403 29563
rect 14289 29529 14323 29563
rect 15025 29529 15059 29563
rect 15853 29529 15887 29563
rect 17478 29529 17512 29563
rect 20269 29529 20303 29563
rect 26249 29529 26283 29563
rect 26617 29529 26651 29563
rect 26801 29529 26835 29563
rect 27353 29529 27387 29563
rect 30113 29529 30147 29563
rect 33425 29529 33459 29563
rect 36001 29529 36035 29563
rect 9781 29461 9815 29495
rect 13569 29461 13603 29495
rect 18613 29461 18647 29495
rect 23305 29461 23339 29495
rect 24685 29461 24719 29495
rect 26709 29461 26743 29495
rect 27813 29461 27847 29495
rect 28549 29461 28583 29495
rect 29745 29461 29779 29495
rect 32321 29461 32355 29495
rect 33701 29461 33735 29495
rect 35265 29461 35299 29495
rect 36369 29461 36403 29495
rect 7481 29257 7515 29291
rect 8125 29257 8159 29291
rect 20545 29257 20579 29291
rect 21005 29257 21039 29291
rect 21373 29257 21407 29291
rect 22477 29257 22511 29291
rect 23765 29257 23799 29291
rect 24133 29257 24167 29291
rect 24685 29257 24719 29291
rect 26525 29257 26559 29291
rect 34345 29257 34379 29291
rect 37933 29257 37967 29291
rect 12909 29189 12943 29223
rect 15761 29189 15795 29223
rect 25697 29189 25731 29223
rect 26065 29189 26099 29223
rect 28549 29189 28583 29223
rect 29101 29189 29135 29223
rect 31585 29189 31619 29223
rect 33057 29189 33091 29223
rect 33977 29189 34011 29223
rect 34069 29189 34103 29223
rect 37841 29189 37875 29223
rect 7297 29121 7331 29155
rect 7481 29121 7515 29155
rect 7941 29121 7975 29155
rect 8125 29121 8159 29155
rect 8585 29121 8619 29155
rect 8769 29121 8803 29155
rect 9505 29121 9539 29155
rect 9689 29121 9723 29155
rect 10425 29121 10459 29155
rect 10701 29121 10735 29155
rect 11989 29121 12023 29155
rect 13093 29121 13127 29155
rect 13185 29121 13219 29155
rect 13645 29121 13679 29155
rect 13901 29121 13935 29155
rect 15485 29121 15519 29155
rect 15669 29121 15703 29155
rect 15853 29121 15887 29155
rect 16865 29121 16899 29155
rect 18153 29121 18187 29155
rect 18337 29121 18371 29155
rect 18429 29121 18463 29155
rect 19165 29121 19199 29155
rect 19421 29121 19455 29155
rect 21189 29121 21223 29155
rect 21465 29121 21499 29155
rect 22385 29121 22419 29155
rect 23949 29121 23983 29155
rect 24225 29121 24259 29155
rect 24869 29121 24903 29155
rect 24961 29121 24995 29155
rect 25053 29121 25087 29155
rect 25145 29121 25179 29155
rect 25329 29121 25363 29155
rect 26341 29121 26375 29155
rect 27169 29121 27203 29155
rect 27353 29121 27387 29155
rect 28181 29121 28215 29155
rect 28365 29121 28399 29155
rect 29377 29121 29411 29155
rect 29469 29121 29503 29155
rect 29561 29121 29595 29155
rect 29745 29121 29779 29155
rect 30481 29121 30515 29155
rect 30573 29121 30607 29155
rect 30665 29121 30699 29155
rect 30849 29121 30883 29155
rect 31309 29121 31343 29155
rect 32597 29121 32631 29155
rect 33701 29121 33735 29155
rect 33794 29121 33828 29155
rect 34166 29121 34200 29155
rect 34989 29121 35023 29155
rect 35081 29121 35115 29155
rect 35265 29121 35299 29155
rect 35357 29121 35391 29155
rect 35817 29121 35851 29155
rect 36001 29121 36035 29155
rect 9229 29053 9263 29087
rect 9413 29053 9447 29087
rect 9597 29053 9631 29087
rect 12173 29053 12207 29087
rect 17049 29053 17083 29087
rect 22661 29053 22695 29087
rect 26249 29053 26283 29087
rect 34805 29053 34839 29087
rect 38117 29053 38151 29087
rect 8677 28985 8711 29019
rect 10609 28985 10643 29019
rect 12909 28985 12943 29019
rect 18613 28985 18647 29019
rect 27445 28985 27479 29019
rect 10241 28917 10275 28951
rect 15025 28917 15059 28951
rect 16037 28917 16071 28951
rect 18153 28917 18187 28951
rect 22017 28917 22051 28951
rect 26065 28917 26099 28951
rect 28457 28917 28491 28951
rect 30205 28917 30239 28951
rect 36093 28917 36127 28951
rect 37473 28917 37507 28951
rect 10425 28713 10459 28747
rect 12449 28713 12483 28747
rect 20085 28713 20119 28747
rect 26157 28713 26191 28747
rect 26985 28713 27019 28747
rect 27077 28713 27111 28747
rect 30849 28713 30883 28747
rect 33517 28713 33551 28747
rect 36277 28713 36311 28747
rect 38209 28713 38243 28747
rect 10701 28645 10735 28679
rect 17049 28645 17083 28679
rect 11437 28577 11471 28611
rect 12633 28577 12667 28611
rect 15658 28577 15692 28611
rect 18153 28577 18187 28611
rect 19901 28577 19935 28611
rect 21925 28577 21959 28611
rect 23949 28577 23983 28611
rect 26065 28577 26099 28611
rect 26985 28577 27019 28611
rect 29193 28577 29227 28611
rect 32045 28577 32079 28611
rect 34897 28577 34931 28611
rect 7205 28509 7239 28543
rect 9321 28509 9355 28543
rect 9413 28509 9447 28543
rect 9597 28509 9631 28543
rect 9689 28509 9723 28543
rect 10609 28509 10643 28543
rect 10793 28509 10827 28543
rect 10885 28509 10919 28543
rect 11621 28509 11655 28543
rect 11713 28509 11747 28543
rect 12449 28509 12483 28543
rect 12725 28509 12759 28543
rect 13461 28509 13495 28543
rect 13553 28509 13587 28543
rect 14289 28509 14323 28543
rect 15936 28509 15970 28543
rect 17969 28509 18003 28543
rect 18705 28509 18739 28543
rect 19809 28509 19843 28543
rect 20913 28509 20947 28543
rect 21189 28509 21223 28543
rect 22201 28509 22235 28543
rect 22477 28509 22511 28543
rect 22661 28509 22695 28543
rect 22937 28509 22971 28543
rect 23857 28509 23891 28543
rect 24593 28509 24627 28543
rect 25145 28509 25179 28543
rect 26157 28509 26191 28543
rect 27169 28509 27203 28543
rect 28641 28509 28675 28543
rect 28825 28509 28859 28543
rect 30297 28509 30331 28543
rect 30665 28509 30699 28543
rect 31585 28509 31619 28543
rect 33425 28509 33459 28543
rect 33977 28509 34011 28543
rect 36829 28509 36863 28543
rect 37096 28509 37130 28543
rect 7472 28441 7506 28475
rect 11805 28441 11839 28475
rect 11989 28441 12023 28475
rect 13737 28441 13771 28475
rect 15117 28441 15151 28475
rect 20637 28441 20671 28475
rect 21005 28441 21039 28475
rect 23397 28441 23431 28475
rect 25881 28441 25915 28475
rect 26801 28441 26835 28475
rect 27721 28441 27755 28475
rect 29101 28441 29135 28475
rect 35164 28441 35198 28475
rect 8585 28373 8619 28407
rect 9137 28373 9171 28407
rect 12909 28373 12943 28407
rect 13461 28373 13495 28407
rect 17509 28373 17543 28407
rect 17877 28373 17911 28407
rect 18797 28373 18831 28407
rect 20821 28373 20855 28407
rect 24685 28373 24719 28407
rect 26341 28373 26375 28407
rect 27997 28373 28031 28407
rect 8033 28169 8067 28203
rect 8493 28169 8527 28203
rect 9965 28169 9999 28203
rect 10701 28169 10735 28203
rect 11805 28169 11839 28203
rect 17877 28169 17911 28203
rect 18705 28169 18739 28203
rect 22477 28169 22511 28203
rect 36921 28169 36955 28203
rect 15577 28101 15611 28135
rect 15669 28101 15703 28135
rect 20637 28101 20671 28135
rect 33057 28101 33091 28135
rect 35808 28101 35842 28135
rect 8401 28033 8435 28067
rect 9781 28033 9815 28067
rect 10057 28033 10091 28067
rect 10885 28033 10919 28067
rect 11069 28033 11103 28067
rect 11161 28033 11195 28067
rect 12061 28033 12095 28067
rect 12173 28033 12207 28067
rect 12265 28033 12299 28067
rect 12449 28033 12483 28067
rect 13176 28033 13210 28067
rect 14749 28033 14783 28067
rect 14933 28033 14967 28067
rect 15393 28033 15427 28067
rect 15761 28033 15795 28067
rect 16865 28033 16899 28067
rect 17969 28033 18003 28067
rect 19073 28033 19107 28067
rect 20269 28033 20303 28067
rect 20453 28033 20487 28067
rect 21097 28033 21131 28067
rect 21281 28033 21315 28067
rect 22385 28033 22419 28067
rect 23397 28033 23431 28067
rect 23581 28033 23615 28067
rect 23673 28033 23707 28067
rect 24685 28033 24719 28067
rect 24961 28033 24995 28067
rect 25421 28033 25455 28067
rect 25605 28033 25639 28067
rect 25697 28033 25731 28067
rect 25973 28033 26007 28067
rect 27261 28033 27295 28067
rect 28365 28033 28399 28067
rect 29009 28033 29043 28067
rect 29377 28033 29411 28067
rect 29653 28033 29687 28067
rect 30665 28033 30699 28067
rect 31585 28033 31619 28067
rect 32321 28033 32355 28067
rect 33701 28033 33735 28067
rect 33794 28033 33828 28067
rect 33977 28033 34011 28067
rect 34069 28033 34103 28067
rect 34207 28033 34241 28067
rect 34897 28033 34931 28067
rect 35081 28033 35115 28067
rect 35541 28033 35575 28067
rect 37565 28033 37599 28067
rect 8585 27965 8619 27999
rect 12909 27965 12943 27999
rect 18153 27965 18187 27999
rect 19165 27965 19199 27999
rect 19257 27965 19291 27999
rect 22661 27965 22695 27999
rect 25789 27965 25823 27999
rect 27997 27965 28031 27999
rect 31769 27965 31803 27999
rect 38025 27965 38059 27999
rect 14289 27897 14323 27931
rect 16957 27897 16991 27931
rect 21373 27897 21407 27931
rect 23489 27897 23523 27931
rect 24869 27897 24903 27931
rect 29469 27897 29503 27931
rect 9597 27829 9631 27863
rect 14749 27829 14783 27863
rect 15945 27829 15979 27863
rect 17509 27829 17543 27863
rect 22017 27829 22051 27863
rect 23213 27829 23247 27863
rect 24501 27829 24535 27863
rect 26157 27829 26191 27863
rect 34345 27829 34379 27863
rect 34897 27829 34931 27863
rect 9137 27625 9171 27659
rect 10057 27625 10091 27659
rect 13277 27625 13311 27659
rect 17877 27625 17911 27659
rect 23121 27625 23155 27659
rect 24685 27625 24719 27659
rect 35541 27625 35575 27659
rect 17049 27557 17083 27591
rect 23397 27557 23431 27591
rect 36001 27557 36035 27591
rect 7113 27489 7147 27523
rect 11897 27489 11931 27523
rect 11989 27489 12023 27523
rect 12173 27489 12207 27523
rect 18337 27489 18371 27523
rect 18429 27489 18463 27523
rect 19809 27489 19843 27523
rect 22293 27489 22327 27523
rect 22477 27489 22511 27523
rect 24869 27489 24903 27523
rect 26157 27489 26191 27523
rect 26249 27489 26283 27523
rect 27997 27489 28031 27523
rect 32229 27489 32263 27523
rect 9137 27421 9171 27455
rect 9321 27421 9355 27455
rect 9965 27421 9999 27455
rect 10793 27421 10827 27455
rect 10977 27421 11011 27455
rect 11069 27421 11103 27455
rect 12081 27421 12115 27455
rect 12725 27421 12759 27455
rect 12909 27421 12943 27455
rect 13093 27421 13127 27455
rect 14289 27421 14323 27455
rect 14473 27421 14507 27455
rect 14565 27421 14599 27455
rect 14657 27421 14691 27455
rect 15669 27421 15703 27455
rect 15936 27421 15970 27455
rect 19901 27421 19935 27455
rect 20821 27421 20855 27455
rect 20913 27421 20947 27455
rect 23029 27421 23063 27455
rect 23121 27421 23155 27455
rect 23857 27421 23891 27455
rect 24041 27421 24075 27455
rect 25053 27421 25087 27455
rect 25881 27421 25915 27455
rect 27537 27421 27571 27455
rect 27721 27421 27755 27455
rect 28825 27421 28859 27455
rect 28917 27421 28951 27455
rect 29009 27421 29043 27455
rect 29101 27421 29135 27455
rect 29929 27421 29963 27455
rect 30389 27421 30423 27455
rect 30573 27421 30607 27455
rect 32781 27421 32815 27455
rect 34161 27421 34195 27455
rect 34345 27421 34379 27455
rect 34897 27421 34931 27455
rect 34990 27421 35024 27455
rect 35362 27421 35396 27455
rect 36277 27421 36311 27455
rect 36737 27421 36771 27455
rect 7380 27353 7414 27387
rect 13001 27353 13035 27387
rect 20177 27353 20211 27387
rect 20269 27353 20303 27387
rect 21097 27353 21131 27387
rect 22201 27353 22235 27387
rect 24593 27353 24627 27387
rect 26366 27353 26400 27387
rect 31401 27353 31435 27387
rect 33517 27353 33551 27387
rect 35173 27353 35207 27387
rect 35265 27353 35299 27387
rect 36001 27353 36035 27387
rect 37004 27353 37038 27387
rect 8493 27285 8527 27319
rect 10609 27285 10643 27319
rect 11713 27285 11747 27319
rect 14841 27285 14875 27319
rect 18245 27285 18279 27319
rect 19625 27285 19659 27319
rect 21833 27285 21867 27319
rect 23949 27285 23983 27319
rect 25237 27285 25271 27319
rect 26525 27285 26559 27319
rect 28641 27285 28675 27319
rect 29837 27285 29871 27319
rect 34253 27285 34287 27319
rect 36185 27285 36219 27319
rect 38117 27285 38151 27319
rect 8033 27081 8067 27115
rect 8493 27081 8527 27115
rect 15961 27081 15995 27115
rect 18889 27081 18923 27115
rect 26617 27081 26651 27115
rect 37473 27081 37507 27115
rect 37933 27081 37967 27115
rect 8401 27013 8435 27047
rect 14188 27013 14222 27047
rect 15761 27013 15795 27047
rect 20545 27013 20579 27047
rect 20637 27013 20671 27047
rect 20755 27013 20789 27047
rect 23397 27013 23431 27047
rect 24685 27013 24719 27047
rect 27629 27013 27663 27047
rect 27721 27013 27755 27047
rect 31401 27013 31435 27047
rect 35173 27013 35207 27047
rect 35265 27013 35299 27047
rect 9597 26945 9631 26979
rect 9781 26945 9815 26979
rect 9873 26945 9907 26979
rect 9965 26945 9999 26979
rect 10793 26945 10827 26979
rect 12449 26945 12483 26979
rect 12633 26945 12667 26979
rect 12725 26945 12759 26979
rect 13277 26945 13311 26979
rect 13461 26945 13495 26979
rect 16957 26945 16991 26979
rect 17224 26945 17258 26979
rect 19073 26945 19107 26979
rect 19165 26945 19199 26979
rect 19441 26945 19475 26979
rect 20453 26945 20487 26979
rect 22385 26945 22419 26979
rect 22569 26945 22603 26979
rect 22937 26945 22971 26979
rect 23581 26945 23615 26979
rect 24409 26945 24443 26979
rect 24777 26945 24811 26979
rect 25605 26945 25639 26979
rect 26341 26945 26375 26979
rect 26525 26945 26559 26979
rect 27261 26945 27295 26979
rect 28549 26945 28583 26979
rect 29193 26945 29227 26979
rect 31033 26945 31067 26979
rect 32597 26945 32631 26979
rect 32689 26945 32723 26979
rect 32873 26945 32907 26979
rect 33333 26945 33367 26979
rect 33793 26945 33827 26979
rect 33885 26945 33919 26979
rect 34069 26945 34103 26979
rect 34989 26945 35023 26979
rect 35357 26945 35391 26979
rect 36001 26945 36035 26979
rect 36185 26945 36219 26979
rect 36277 26945 36311 26979
rect 36461 26945 36495 26979
rect 36553 26945 36587 26979
rect 37841 26945 37875 26979
rect 8677 26877 8711 26911
rect 10609 26877 10643 26911
rect 13921 26877 13955 26911
rect 19349 26877 19383 26911
rect 20913 26877 20947 26911
rect 24225 26877 24259 26911
rect 29285 26877 29319 26911
rect 30941 26877 30975 26911
rect 31309 26877 31343 26911
rect 34529 26877 34563 26911
rect 38025 26877 38059 26911
rect 10977 26809 11011 26843
rect 10149 26741 10183 26775
rect 12265 26741 12299 26775
rect 13277 26741 13311 26775
rect 15301 26741 15335 26775
rect 15945 26741 15979 26775
rect 16129 26741 16163 26775
rect 18337 26741 18371 26775
rect 20269 26741 20303 26775
rect 23765 26741 23799 26775
rect 30757 26741 30791 26775
rect 35541 26741 35575 26775
rect 11345 26537 11379 26571
rect 18521 26537 18555 26571
rect 36461 26537 36495 26571
rect 13185 26469 13219 26503
rect 15301 26469 15335 26503
rect 18889 26469 18923 26503
rect 23857 26469 23891 26503
rect 32045 26469 32079 26503
rect 35449 26469 35483 26503
rect 9965 26401 9999 26435
rect 15761 26401 15795 26435
rect 18061 26401 18095 26435
rect 18613 26401 18647 26435
rect 22477 26401 22511 26435
rect 27813 26401 27847 26435
rect 28181 26401 28215 26435
rect 28273 26401 28307 26435
rect 28365 26401 28399 26435
rect 34069 26401 34103 26435
rect 11805 26333 11839 26367
rect 14749 26333 14783 26367
rect 15025 26333 15059 26367
rect 15117 26333 15151 26367
rect 16017 26333 16051 26367
rect 17785 26333 17819 26367
rect 17877 26333 17911 26367
rect 18521 26333 18555 26367
rect 19993 26333 20027 26367
rect 20177 26333 20211 26367
rect 20499 26333 20533 26367
rect 20637 26333 20671 26367
rect 21649 26333 21683 26367
rect 21833 26333 21867 26367
rect 22744 26333 22778 26367
rect 24685 26333 24719 26367
rect 24869 26333 24903 26367
rect 26433 26333 26467 26367
rect 29009 26333 29043 26367
rect 29193 26333 29227 26367
rect 30113 26333 30147 26367
rect 30573 26333 30607 26367
rect 30721 26333 30755 26367
rect 30941 26333 30975 26367
rect 31079 26333 31113 26367
rect 31861 26333 31895 26367
rect 33885 26333 33919 26367
rect 34897 26333 34931 26367
rect 35265 26333 35299 26367
rect 35909 26333 35943 26367
rect 36093 26333 36127 26367
rect 36185 26333 36219 26367
rect 36277 26333 36311 26367
rect 36921 26333 36955 26367
rect 10232 26265 10266 26299
rect 12072 26265 12106 26299
rect 14933 26265 14967 26299
rect 20269 26265 20303 26299
rect 20361 26265 20395 26299
rect 22017 26265 22051 26299
rect 25237 26265 25271 26299
rect 26157 26265 26191 26299
rect 26341 26265 26375 26299
rect 26525 26265 26559 26299
rect 26893 26265 26927 26299
rect 29101 26265 29135 26299
rect 29745 26265 29779 26299
rect 29929 26265 29963 26299
rect 30849 26265 30883 26299
rect 31677 26265 31711 26299
rect 32505 26265 32539 26299
rect 33241 26265 33275 26299
rect 35081 26265 35115 26299
rect 35173 26265 35207 26299
rect 37188 26265 37222 26299
rect 17141 26197 17175 26231
rect 31217 26197 31251 26231
rect 38301 26197 38335 26231
rect 10977 25993 11011 26027
rect 13093 25993 13127 26027
rect 18797 25993 18831 26027
rect 22201 25993 22235 26027
rect 22937 25993 22971 26027
rect 37473 25993 37507 26027
rect 8668 25925 8702 25959
rect 13645 25925 13679 25959
rect 19257 25925 19291 25959
rect 20453 25925 20487 25959
rect 20913 25925 20947 25959
rect 22017 25925 22051 25959
rect 23765 25925 23799 25959
rect 24685 25925 24719 25959
rect 29101 25925 29135 25959
rect 32413 25925 32447 25959
rect 37841 25925 37875 25959
rect 8401 25857 8435 25891
rect 10425 25857 10459 25891
rect 10609 25857 10643 25891
rect 10701 25857 10735 25891
rect 10793 25857 10827 25891
rect 11713 25857 11747 25891
rect 11980 25857 12014 25891
rect 13553 25857 13587 25891
rect 14197 25857 14231 25891
rect 14381 25857 14415 25891
rect 15108 25857 15142 25891
rect 17601 25857 17635 25891
rect 17785 25857 17819 25891
rect 17877 25857 17911 25891
rect 18613 25857 18647 25891
rect 19441 25857 19475 25891
rect 19625 25857 19659 25891
rect 20177 25857 20211 25891
rect 20361 25857 20395 25891
rect 21189 25857 21223 25891
rect 22293 25857 22327 25891
rect 23949 25857 23983 25891
rect 26065 25857 26099 25891
rect 27169 25857 27203 25891
rect 27629 25857 27663 25891
rect 27997 25857 28031 25891
rect 28825 25857 28859 25891
rect 29009 25857 29043 25891
rect 29193 25857 29227 25891
rect 30021 25857 30055 25891
rect 30849 25857 30883 25891
rect 33793 25857 33827 25891
rect 34069 25857 34103 25891
rect 35449 25857 35483 25891
rect 35716 25857 35750 25891
rect 37933 25857 37967 25891
rect 14841 25789 14875 25823
rect 18429 25789 18463 25823
rect 21005 25789 21039 25823
rect 22753 25789 22787 25823
rect 23121 25789 23155 25823
rect 24225 25789 24259 25823
rect 24869 25789 24903 25823
rect 25053 25789 25087 25823
rect 26249 25789 26283 25823
rect 28181 25789 28215 25823
rect 30757 25789 30791 25823
rect 31309 25789 31343 25823
rect 33241 25789 33275 25823
rect 34437 25789 34471 25823
rect 38025 25789 38059 25823
rect 9781 25721 9815 25755
rect 14289 25721 14323 25755
rect 21373 25721 21407 25755
rect 22017 25721 22051 25755
rect 24133 25721 24167 25755
rect 24685 25721 24719 25755
rect 33885 25721 33919 25755
rect 16221 25653 16255 25687
rect 17417 25653 17451 25687
rect 20913 25653 20947 25687
rect 23121 25653 23155 25687
rect 24961 25653 24995 25687
rect 29377 25653 29411 25687
rect 36829 25653 36863 25687
rect 13277 25449 13311 25483
rect 15577 25449 15611 25483
rect 16589 25449 16623 25483
rect 17049 25449 17083 25483
rect 18797 25449 18831 25483
rect 23765 25449 23799 25483
rect 25881 25449 25915 25483
rect 30297 25449 30331 25483
rect 33793 25449 33827 25483
rect 23949 25381 23983 25415
rect 25145 25381 25179 25415
rect 26709 25381 26743 25415
rect 28733 25381 28767 25415
rect 33682 25381 33716 25415
rect 9597 25313 9631 25347
rect 9781 25313 9815 25347
rect 16681 25313 16715 25347
rect 18153 25313 18187 25347
rect 19441 25313 19475 25347
rect 21465 25313 21499 25347
rect 21649 25313 21683 25347
rect 22661 25313 22695 25347
rect 23581 25313 23615 25347
rect 24685 25313 24719 25347
rect 30849 25313 30883 25347
rect 33885 25313 33919 25347
rect 36921 25313 36955 25347
rect 10425 25245 10459 25279
rect 10609 25245 10643 25279
rect 11529 25245 11563 25279
rect 11713 25245 11747 25279
rect 13277 25245 13311 25279
rect 13461 25245 13495 25279
rect 14381 25245 14415 25279
rect 14565 25245 14599 25279
rect 15025 25245 15059 25279
rect 15301 25245 15335 25279
rect 15393 25245 15427 25279
rect 16589 25245 16623 25279
rect 16865 25245 16899 25279
rect 17969 25245 18003 25279
rect 18705 25245 18739 25279
rect 18889 25245 18923 25279
rect 19625 25245 19659 25279
rect 19790 25245 19824 25279
rect 19886 25245 19920 25279
rect 19993 25245 20027 25279
rect 22385 25245 22419 25279
rect 22477 25245 22511 25279
rect 22753 25245 22787 25279
rect 23765 25245 23799 25279
rect 24777 25245 24811 25279
rect 25789 25245 25823 25279
rect 26525 25245 26559 25279
rect 26617 25245 26651 25279
rect 27445 25245 27479 25279
rect 27629 25245 27663 25279
rect 27721 25245 27755 25279
rect 28181 25245 28215 25279
rect 28457 25245 28491 25279
rect 28549 25245 28583 25279
rect 29745 25245 29779 25279
rect 30021 25245 30055 25279
rect 30113 25245 30147 25279
rect 31033 25245 31067 25279
rect 32229 25245 32263 25279
rect 32413 25245 32447 25279
rect 32781 25245 32815 25279
rect 34897 25245 34931 25279
rect 35265 25245 35299 25279
rect 36093 25245 36127 25279
rect 36185 25245 36219 25279
rect 36369 25245 36403 25279
rect 36461 25245 36495 25279
rect 14473 25177 14507 25211
rect 15209 25177 15243 25211
rect 17877 25177 17911 25211
rect 22201 25177 22235 25211
rect 23489 25177 23523 25211
rect 25605 25177 25639 25211
rect 28365 25177 28399 25211
rect 29929 25177 29963 25211
rect 31217 25177 31251 25211
rect 31309 25177 31343 25211
rect 33517 25177 33551 25211
rect 34253 25177 34287 25211
rect 35081 25177 35115 25211
rect 35173 25177 35207 25211
rect 35909 25177 35943 25211
rect 37188 25177 37222 25211
rect 9137 25109 9171 25143
rect 9505 25109 9539 25143
rect 10517 25109 10551 25143
rect 11621 25109 11655 25143
rect 17509 25109 17543 25143
rect 21005 25109 21039 25143
rect 21373 25109 21407 25143
rect 27261 25109 27295 25143
rect 33057 25109 33091 25143
rect 35449 25109 35483 25143
rect 38301 25109 38335 25143
rect 9597 24905 9631 24939
rect 14289 24905 14323 24939
rect 15117 24905 15151 24939
rect 16957 24905 16991 24939
rect 17785 24905 17819 24939
rect 21005 24905 21039 24939
rect 30573 24905 30607 24939
rect 37841 24905 37875 24939
rect 8484 24837 8518 24871
rect 18705 24837 18739 24871
rect 19809 24837 19843 24871
rect 24216 24837 24250 24871
rect 32873 24837 32907 24871
rect 34069 24837 34103 24871
rect 36093 24837 36127 24871
rect 10241 24769 10275 24803
rect 10333 24769 10367 24803
rect 10609 24769 10643 24803
rect 11713 24769 11747 24803
rect 11897 24769 11931 24803
rect 11989 24769 12023 24803
rect 12081 24769 12115 24803
rect 13176 24769 13210 24803
rect 16129 24769 16163 24803
rect 16313 24769 16347 24803
rect 17693 24769 17727 24803
rect 18981 24769 19015 24803
rect 19073 24769 19107 24803
rect 19441 24769 19475 24803
rect 20913 24769 20947 24803
rect 22273 24769 22307 24803
rect 23949 24769 23983 24803
rect 25973 24769 26007 24803
rect 26157 24769 26191 24803
rect 26249 24769 26283 24803
rect 26346 24769 26380 24803
rect 27445 24769 27479 24803
rect 27629 24769 27663 24803
rect 27721 24769 27755 24803
rect 27813 24769 27847 24803
rect 28273 24769 28307 24803
rect 29377 24769 29411 24803
rect 29561 24769 29595 24803
rect 29653 24769 29687 24803
rect 29745 24769 29779 24803
rect 30389 24769 30423 24803
rect 30665 24769 30699 24803
rect 31401 24769 31435 24803
rect 31493 24769 31527 24803
rect 31677 24769 31711 24803
rect 31769 24769 31803 24803
rect 32597 24769 32631 24803
rect 33701 24769 33735 24803
rect 34621 24769 34655 24803
rect 34769 24769 34803 24803
rect 34897 24769 34931 24803
rect 34997 24769 35031 24803
rect 35127 24769 35161 24803
rect 35725 24769 35759 24803
rect 35818 24769 35852 24803
rect 36001 24769 36035 24803
rect 36231 24769 36265 24803
rect 8217 24701 8251 24735
rect 10701 24701 10735 24735
rect 12909 24701 12943 24735
rect 15209 24701 15243 24735
rect 15301 24701 15335 24735
rect 17969 24701 18003 24735
rect 21097 24701 21131 24735
rect 22017 24701 22051 24735
rect 28549 24701 28583 24735
rect 32505 24701 32539 24735
rect 32965 24701 32999 24735
rect 33609 24701 33643 24735
rect 33977 24701 34011 24735
rect 37933 24701 37967 24735
rect 38025 24701 38059 24735
rect 14749 24633 14783 24667
rect 19993 24633 20027 24667
rect 32321 24633 32355 24667
rect 37473 24633 37507 24667
rect 10057 24565 10091 24599
rect 12265 24565 12299 24599
rect 16129 24565 16163 24599
rect 17325 24565 17359 24599
rect 20545 24565 20579 24599
rect 23397 24565 23431 24599
rect 25329 24565 25363 24599
rect 26525 24565 26559 24599
rect 27997 24565 28031 24599
rect 29101 24565 29135 24599
rect 29929 24565 29963 24599
rect 30389 24565 30423 24599
rect 31217 24565 31251 24599
rect 33425 24565 33459 24599
rect 35265 24565 35299 24599
rect 36369 24565 36403 24599
rect 14473 24361 14507 24395
rect 18613 24361 18647 24395
rect 18705 24361 18739 24395
rect 21005 24361 21039 24395
rect 21925 24361 21959 24395
rect 31769 24361 31803 24395
rect 32689 24361 32723 24395
rect 12173 24293 12207 24327
rect 16405 24293 16439 24327
rect 28917 24293 28951 24327
rect 30757 24293 30791 24327
rect 34897 24293 34931 24327
rect 36093 24293 36127 24327
rect 15025 24225 15059 24259
rect 17325 24225 17359 24259
rect 17417 24225 17451 24259
rect 18521 24225 18555 24259
rect 22569 24225 22603 24259
rect 23765 24225 23799 24259
rect 24593 24225 24627 24259
rect 36921 24225 36955 24259
rect 10793 24157 10827 24191
rect 13218 24157 13252 24191
rect 13645 24157 13679 24191
rect 13737 24157 13771 24191
rect 14381 24157 14415 24191
rect 18429 24157 18463 24191
rect 18889 24157 18923 24191
rect 19625 24157 19659 24191
rect 23489 24157 23523 24191
rect 24777 24157 24811 24191
rect 25053 24157 25087 24191
rect 25237 24157 25271 24191
rect 26341 24157 26375 24191
rect 26433 24157 26467 24191
rect 26525 24157 26559 24191
rect 26617 24157 26651 24191
rect 26801 24157 26835 24191
rect 27905 24157 27939 24191
rect 27997 24157 28031 24191
rect 28273 24157 28307 24191
rect 28457 24157 28491 24191
rect 29193 24157 29227 24191
rect 29745 24157 29779 24191
rect 30113 24157 30147 24191
rect 30757 24157 30791 24191
rect 31033 24157 31067 24191
rect 31677 24157 31711 24191
rect 33333 24157 33367 24191
rect 33609 24157 33643 24191
rect 33793 24157 33827 24191
rect 33977 24157 34011 24191
rect 34897 24157 34931 24191
rect 35173 24157 35207 24191
rect 35817 24157 35851 24191
rect 35909 24157 35943 24191
rect 36185 24157 36219 24191
rect 11060 24089 11094 24123
rect 15292 24089 15326 24123
rect 19892 24089 19926 24123
rect 22293 24089 22327 24123
rect 27261 24089 27295 24123
rect 28917 24089 28951 24123
rect 29929 24089 29963 24123
rect 30021 24089 30055 24123
rect 31493 24089 31527 24123
rect 32505 24089 32539 24123
rect 32705 24089 32739 24123
rect 34161 24089 34195 24123
rect 35633 24089 35667 24123
rect 37188 24089 37222 24123
rect 13093 24021 13127 24055
rect 13277 24021 13311 24055
rect 16865 24021 16899 24055
rect 17233 24021 17267 24055
rect 18153 24021 18187 24055
rect 22385 24021 22419 24055
rect 23121 24021 23155 24055
rect 23581 24021 23615 24055
rect 26157 24021 26191 24055
rect 29101 24021 29135 24055
rect 30297 24021 30331 24055
rect 30941 24021 30975 24055
rect 32873 24021 32907 24055
rect 35081 24021 35115 24055
rect 38301 24021 38335 24055
rect 10885 23817 10919 23851
rect 12449 23817 12483 23851
rect 15945 23817 15979 23851
rect 18153 23817 18187 23851
rect 19901 23817 19935 23851
rect 20453 23817 20487 23851
rect 27169 23817 27203 23851
rect 27537 23817 27571 23851
rect 35633 23817 35667 23851
rect 37473 23817 37507 23851
rect 37841 23817 37875 23851
rect 9772 23749 9806 23783
rect 13706 23749 13740 23783
rect 15577 23749 15611 23783
rect 22385 23749 22419 23783
rect 30113 23749 30147 23783
rect 31033 23749 31067 23783
rect 34161 23749 34195 23783
rect 9505 23681 9539 23715
rect 12357 23681 12391 23715
rect 13461 23681 13495 23715
rect 15393 23681 15427 23715
rect 15669 23681 15703 23715
rect 15761 23681 15795 23715
rect 17141 23681 17175 23715
rect 17325 23681 17359 23715
rect 18245 23681 18279 23715
rect 19717 23681 19751 23715
rect 19993 23681 20027 23715
rect 20637 23681 20671 23715
rect 20913 23681 20947 23715
rect 22017 23681 22051 23715
rect 22293 23681 22327 23715
rect 22845 23681 22879 23715
rect 25513 23681 25547 23715
rect 25605 23681 25639 23715
rect 25881 23681 25915 23715
rect 26157 23681 26191 23715
rect 26341 23681 26375 23715
rect 27353 23681 27387 23715
rect 27629 23681 27663 23715
rect 28549 23681 28583 23715
rect 28888 23681 28922 23715
rect 29745 23681 29779 23715
rect 29893 23681 29927 23715
rect 30021 23681 30055 23715
rect 30210 23681 30244 23715
rect 30849 23681 30883 23715
rect 31125 23681 31159 23715
rect 31217 23681 31251 23715
rect 32689 23681 32723 23715
rect 33241 23681 33275 23715
rect 33885 23681 33919 23715
rect 34033 23681 34067 23715
rect 34253 23681 34287 23715
rect 34391 23681 34425 23715
rect 34989 23681 35023 23715
rect 35137 23681 35171 23715
rect 35265 23681 35299 23715
rect 35357 23681 35391 23715
rect 35454 23681 35488 23715
rect 36277 23681 36311 23715
rect 36369 23681 36403 23715
rect 36645 23681 36679 23715
rect 12633 23613 12667 23647
rect 18429 23613 18463 23647
rect 20821 23613 20855 23647
rect 29285 23613 29319 23647
rect 32413 23613 32447 23647
rect 33425 23613 33459 23647
rect 36093 23613 36127 23647
rect 37933 23613 37967 23647
rect 38025 23613 38059 23647
rect 24317 23545 24351 23579
rect 36553 23545 36587 23579
rect 11989 23477 12023 23511
rect 14841 23477 14875 23511
rect 17233 23477 17267 23511
rect 17785 23477 17819 23511
rect 19533 23477 19567 23511
rect 25145 23477 25179 23511
rect 28687 23477 28721 23511
rect 28825 23477 28859 23511
rect 30389 23477 30423 23511
rect 31401 23477 31435 23511
rect 34529 23477 34563 23511
rect 12817 23273 12851 23307
rect 15025 23273 15059 23307
rect 23305 23273 23339 23307
rect 30849 23273 30883 23307
rect 35541 23273 35575 23307
rect 37565 23273 37599 23307
rect 18889 23205 18923 23239
rect 22109 23205 22143 23239
rect 28457 23205 28491 23239
rect 28917 23205 28951 23239
rect 11437 23137 11471 23171
rect 19441 23137 19475 23171
rect 23949 23137 23983 23171
rect 26709 23137 26743 23171
rect 11704 23069 11738 23103
rect 14841 23069 14875 23103
rect 15117 23069 15151 23103
rect 15577 23069 15611 23103
rect 17509 23069 17543 23103
rect 19625 23069 19659 23103
rect 20729 23069 20763 23103
rect 24593 23069 24627 23103
rect 25421 23069 25455 23103
rect 25605 23069 25639 23103
rect 26157 23069 26191 23103
rect 26341 23069 26375 23103
rect 27169 23069 27203 23103
rect 28917 23069 28951 23103
rect 29193 23069 29227 23103
rect 29745 23069 29779 23103
rect 29893 23069 29927 23103
rect 30021 23069 30055 23103
rect 30210 23069 30244 23103
rect 30849 23069 30883 23103
rect 31125 23069 31159 23103
rect 31861 23069 31895 23103
rect 32137 23069 32171 23103
rect 32321 23069 32355 23103
rect 32781 23069 32815 23103
rect 32919 23069 32953 23103
rect 33287 23069 33321 23103
rect 34069 23069 34103 23103
rect 34253 23069 34287 23103
rect 34345 23069 34379 23103
rect 34897 23069 34931 23103
rect 34990 23069 35024 23103
rect 35173 23069 35207 23103
rect 35362 23069 35396 23103
rect 36185 23069 36219 23103
rect 38117 23069 38151 23103
rect 38301 23069 38335 23103
rect 15844 23001 15878 23035
rect 17765 23001 17799 23035
rect 20974 23001 21008 23035
rect 23673 23001 23707 23035
rect 27445 23001 27479 23035
rect 28089 23001 28123 23035
rect 28273 23001 28307 23035
rect 30113 23001 30147 23035
rect 33057 23001 33091 23035
rect 33149 23001 33183 23035
rect 35265 23001 35299 23035
rect 36452 23001 36486 23035
rect 14657 22933 14691 22967
rect 16957 22933 16991 22967
rect 19809 22933 19843 22967
rect 23029 22933 23063 22967
rect 23765 22933 23799 22967
rect 24685 22933 24719 22967
rect 26341 22933 26375 22967
rect 29101 22933 29135 22967
rect 30389 22933 30423 22967
rect 31033 22933 31067 22967
rect 33425 22933 33459 22967
rect 33885 22933 33919 22967
rect 38209 22933 38243 22967
rect 14197 22729 14231 22763
rect 18613 22729 18647 22763
rect 20453 22729 20487 22763
rect 21373 22729 21407 22763
rect 27353 22729 27387 22763
rect 28641 22729 28675 22763
rect 32781 22729 32815 22763
rect 33701 22729 33735 22763
rect 13084 22661 13118 22695
rect 14749 22661 14783 22695
rect 17417 22661 17451 22695
rect 34345 22661 34379 22695
rect 37749 22661 37783 22695
rect 12817 22593 12851 22627
rect 16129 22593 16163 22627
rect 16313 22593 16347 22627
rect 17141 22593 17175 22627
rect 17234 22593 17268 22627
rect 17509 22593 17543 22627
rect 17606 22593 17640 22627
rect 18429 22593 18463 22627
rect 19073 22593 19107 22627
rect 21281 22593 21315 22627
rect 21465 22593 21499 22627
rect 22201 22593 22235 22627
rect 22569 22593 22603 22627
rect 23673 22593 23707 22627
rect 25145 22593 25179 22627
rect 25513 22593 25547 22627
rect 25973 22593 26007 22627
rect 26157 22593 26191 22627
rect 26249 22593 26283 22627
rect 26393 22593 26427 22627
rect 27537 22593 27571 22627
rect 27813 22593 27847 22627
rect 28273 22593 28307 22627
rect 28457 22593 28491 22627
rect 29101 22593 29135 22627
rect 29377 22593 29411 22627
rect 30297 22593 30331 22627
rect 30849 22593 30883 22627
rect 31217 22593 31251 22627
rect 31677 22593 31711 22627
rect 32779 22593 32813 22627
rect 33886 22593 33920 22627
rect 33978 22593 34012 22627
rect 34253 22593 34287 22627
rect 35357 22593 35391 22627
rect 35449 22593 35483 22627
rect 35725 22593 35759 22627
rect 36369 22593 36403 22627
rect 37473 22593 37507 22627
rect 15577 22525 15611 22559
rect 18245 22525 18279 22559
rect 19349 22525 19383 22559
rect 22845 22525 22879 22559
rect 24961 22525 24995 22559
rect 31309 22525 31343 22559
rect 33241 22525 33275 22559
rect 36277 22525 36311 22559
rect 36737 22525 36771 22559
rect 22293 22457 22327 22491
rect 25421 22457 25455 22491
rect 29377 22457 29411 22491
rect 33149 22457 33183 22491
rect 35173 22457 35207 22491
rect 16129 22389 16163 22423
rect 17785 22389 17819 22423
rect 23765 22389 23799 22423
rect 26525 22389 26559 22423
rect 27721 22389 27755 22423
rect 32597 22389 32631 22423
rect 35633 22389 35667 22423
rect 17325 22185 17359 22219
rect 18797 22185 18831 22219
rect 19441 22185 19475 22219
rect 33241 22185 33275 22219
rect 35541 22185 35575 22219
rect 19809 22117 19843 22151
rect 21373 22117 21407 22151
rect 24869 22117 24903 22151
rect 26525 22117 26559 22151
rect 13553 22049 13587 22083
rect 14749 22049 14783 22083
rect 15301 22049 15335 22083
rect 16037 22049 16071 22083
rect 18429 22049 18463 22083
rect 22109 22049 22143 22083
rect 23305 22049 23339 22083
rect 25053 22049 25087 22083
rect 26065 22049 26099 22083
rect 27629 22049 27663 22083
rect 27813 22049 27847 22083
rect 28529 22049 28563 22083
rect 30021 22049 30055 22083
rect 33793 22049 33827 22083
rect 33885 22049 33919 22083
rect 36277 22049 36311 22083
rect 36921 22049 36955 22083
rect 10977 21981 11011 22015
rect 12817 21981 12851 22015
rect 14841 21981 14875 22015
rect 15761 21981 15795 22015
rect 18521 21981 18555 22015
rect 19625 21981 19659 22015
rect 19901 21981 19935 22015
rect 20361 21981 20395 22015
rect 21281 21981 21315 22015
rect 21649 21981 21683 22015
rect 23029 21981 23063 22015
rect 23857 21981 23891 22015
rect 24041 21981 24075 22015
rect 26157 21981 26191 22015
rect 27537 21981 27571 22015
rect 28641 21981 28675 22015
rect 29009 21981 29043 22015
rect 29837 21981 29871 22015
rect 29929 21981 29963 22015
rect 31033 21981 31067 22015
rect 31126 21981 31160 22015
rect 31309 21981 31343 22015
rect 31498 21981 31532 22015
rect 32137 21981 32171 22015
rect 32285 21981 32319 22015
rect 32413 21981 32447 22015
rect 32643 21981 32677 22015
rect 33425 21981 33459 22015
rect 33517 21981 33551 22015
rect 34897 21981 34931 22015
rect 35045 21981 35079 22015
rect 35173 21981 35207 22015
rect 35403 21981 35437 22015
rect 36001 21981 36035 22015
rect 11244 21913 11278 21947
rect 24593 21913 24627 21947
rect 28917 21913 28951 21947
rect 31401 21913 31435 21947
rect 32505 21913 32539 21947
rect 35265 21913 35299 21947
rect 37188 21913 37222 21947
rect 12357 21845 12391 21879
rect 20453 21845 20487 21879
rect 22661 21845 22695 21879
rect 23121 21845 23155 21879
rect 23949 21845 23983 21879
rect 27169 21845 27203 21879
rect 28365 21845 28399 21879
rect 31677 21845 31711 21879
rect 32781 21845 32815 21879
rect 38301 21845 38335 21879
rect 11805 21641 11839 21675
rect 12265 21641 12299 21675
rect 14749 21641 14783 21675
rect 18245 21641 18279 21675
rect 20269 21641 20303 21675
rect 21373 21641 21407 21675
rect 23857 21641 23891 21675
rect 23949 21641 23983 21675
rect 25053 21641 25087 21675
rect 28089 21641 28123 21675
rect 31401 21641 31435 21675
rect 37473 21641 37507 21675
rect 37841 21641 37875 21675
rect 18705 21573 18739 21607
rect 19441 21573 19475 21607
rect 24133 21573 24167 21607
rect 26157 21573 26191 21607
rect 26249 21573 26283 21607
rect 30113 21573 30147 21607
rect 30297 21573 30331 21607
rect 32505 21573 32539 21607
rect 32597 21573 32631 21607
rect 35633 21573 35667 21607
rect 12173 21505 12207 21539
rect 13369 21505 13403 21539
rect 14381 21505 14415 21539
rect 15485 21505 15519 21539
rect 15577 21505 15611 21539
rect 16865 21505 16899 21539
rect 17049 21505 17083 21539
rect 20210 21505 20244 21539
rect 21189 21505 21223 21539
rect 21465 21505 21499 21539
rect 22293 21505 22327 21539
rect 22385 21505 22419 21539
rect 22477 21505 22511 21539
rect 22661 21505 22695 21539
rect 23765 21505 23799 21539
rect 24593 21505 24627 21539
rect 24869 21505 24903 21539
rect 25973 21505 26007 21539
rect 26393 21505 26427 21539
rect 27261 21505 27295 21539
rect 28365 21505 28399 21539
rect 28457 21505 28491 21539
rect 28549 21505 28583 21539
rect 29101 21505 29135 21539
rect 30389 21505 30423 21539
rect 30849 21505 30883 21539
rect 31033 21505 31067 21539
rect 31125 21505 31159 21539
rect 31217 21505 31251 21539
rect 32321 21505 32355 21539
rect 32689 21505 32723 21539
rect 33333 21505 33367 21539
rect 33517 21505 33551 21539
rect 34529 21505 34563 21539
rect 34622 21505 34656 21539
rect 34805 21505 34839 21539
rect 34897 21505 34931 21539
rect 35035 21505 35069 21539
rect 35817 21505 35851 21539
rect 36461 21505 36495 21539
rect 12357 21437 12391 21471
rect 13461 21437 13495 21471
rect 14289 21437 14323 21471
rect 15761 21437 15795 21471
rect 17785 21437 17819 21471
rect 20729 21437 20763 21471
rect 24685 21437 24719 21471
rect 27353 21437 27387 21471
rect 28273 21437 28307 21471
rect 29377 21437 29411 21471
rect 36737 21437 36771 21471
rect 37933 21437 37967 21471
rect 38117 21437 38151 21471
rect 13737 21369 13771 21403
rect 18153 21369 18187 21403
rect 21189 21369 21223 21403
rect 23581 21369 23615 21403
rect 27629 21369 27663 21403
rect 29653 21369 29687 21403
rect 36001 21369 36035 21403
rect 17233 21301 17267 21335
rect 20085 21301 20119 21335
rect 20637 21301 20671 21335
rect 22017 21301 22051 21335
rect 24593 21301 24627 21335
rect 26525 21301 26559 21335
rect 27445 21301 27479 21335
rect 29193 21301 29227 21335
rect 30113 21301 30147 21335
rect 32873 21301 32907 21335
rect 33517 21301 33551 21335
rect 33701 21301 33735 21335
rect 35173 21301 35207 21335
rect 13645 21097 13679 21131
rect 22569 21097 22603 21131
rect 24593 21097 24627 21131
rect 25973 21097 26007 21131
rect 26801 21097 26835 21131
rect 12633 21029 12667 21063
rect 17601 21029 17635 21063
rect 23029 21029 23063 21063
rect 26157 21029 26191 21063
rect 31125 21029 31159 21063
rect 33425 21029 33459 21063
rect 34069 21029 34103 21063
rect 13185 20961 13219 20995
rect 15485 20961 15519 20995
rect 18889 20961 18923 20995
rect 20913 20961 20947 20995
rect 21925 20961 21959 20995
rect 22293 20961 22327 20995
rect 22385 20961 22419 20995
rect 23213 20961 23247 20995
rect 25237 20961 25271 20995
rect 29009 20961 29043 20995
rect 35541 20961 35575 20995
rect 35817 20961 35851 20995
rect 11253 20893 11287 20927
rect 13277 20893 13311 20927
rect 14657 20893 14691 20927
rect 15025 20893 15059 20927
rect 15761 20893 15795 20927
rect 17601 20893 17635 20927
rect 17877 20893 17911 20927
rect 18337 20893 18371 20927
rect 18521 20893 18555 20927
rect 19533 20893 19567 20927
rect 19809 20893 19843 20927
rect 20269 20893 20303 20927
rect 20545 20893 20579 20927
rect 23305 20893 23339 20927
rect 23397 20893 23431 20927
rect 23489 20893 23523 20927
rect 27445 20893 27479 20927
rect 27629 20893 27663 20927
rect 28699 20893 28733 20927
rect 29101 20893 29135 20927
rect 30113 20893 30147 20927
rect 30297 20893 30331 20927
rect 30481 20893 30515 20927
rect 31401 20893 31435 20927
rect 32137 20893 32171 20927
rect 32229 20893 32263 20927
rect 32321 20893 32355 20927
rect 32413 20893 32447 20927
rect 33241 20893 33275 20927
rect 33333 20893 33367 20927
rect 33517 20893 33551 20927
rect 34069 20893 34103 20927
rect 34345 20893 34379 20927
rect 35449 20893 35483 20927
rect 36277 20893 36311 20927
rect 11520 20825 11554 20859
rect 14841 20825 14875 20859
rect 17141 20825 17175 20859
rect 25789 20825 25823 20859
rect 26617 20825 26651 20859
rect 30389 20825 30423 20859
rect 31125 20825 31159 20859
rect 36522 20825 36556 20859
rect 17785 20757 17819 20791
rect 18521 20757 18555 20791
rect 24961 20757 24995 20791
rect 25053 20757 25087 20791
rect 25989 20757 26023 20791
rect 26817 20757 26851 20791
rect 26985 20757 27019 20791
rect 27721 20757 27755 20791
rect 28549 20757 28583 20791
rect 30665 20757 30699 20791
rect 31309 20757 31343 20791
rect 31953 20757 31987 20791
rect 33057 20757 33091 20791
rect 34253 20757 34287 20791
rect 37657 20757 37691 20791
rect 16221 20553 16255 20587
rect 20637 20553 20671 20587
rect 21373 20553 21407 20587
rect 24685 20553 24719 20587
rect 25605 20553 25639 20587
rect 28549 20553 28583 20587
rect 30849 20553 30883 20587
rect 36829 20553 36863 20587
rect 19165 20485 19199 20519
rect 24041 20485 24075 20519
rect 26433 20485 26467 20519
rect 28365 20485 28399 20519
rect 30481 20485 30515 20519
rect 36645 20485 36679 20519
rect 37933 20485 37967 20519
rect 12357 20417 12391 20451
rect 12541 20417 12575 20451
rect 15117 20417 15151 20451
rect 16037 20417 16071 20451
rect 16313 20417 16347 20451
rect 16865 20417 16899 20451
rect 17049 20417 17083 20451
rect 17693 20417 17727 20451
rect 17785 20417 17819 20451
rect 18429 20417 18463 20451
rect 18705 20417 18739 20451
rect 18797 20417 18831 20451
rect 21281 20417 21315 20451
rect 21465 20417 21499 20451
rect 22477 20417 22511 20451
rect 22753 20417 22787 20451
rect 22845 20417 22879 20451
rect 23121 20417 23155 20451
rect 23305 20417 23339 20451
rect 24501 20417 24535 20451
rect 26065 20417 26099 20451
rect 26158 20417 26192 20451
rect 27905 20417 27939 20451
rect 28641 20417 28675 20451
rect 29285 20417 29319 20451
rect 30297 20417 30331 20451
rect 30573 20417 30607 20451
rect 30665 20417 30699 20451
rect 32689 20417 32723 20451
rect 32781 20417 32815 20451
rect 33885 20417 33919 20451
rect 33977 20417 34011 20451
rect 34161 20417 34195 20451
rect 34253 20417 34287 20451
rect 34713 20417 34747 20451
rect 34989 20417 35023 20451
rect 35817 20417 35851 20451
rect 35909 20417 35943 20451
rect 36185 20417 36219 20451
rect 36921 20417 36955 20451
rect 37841 20417 37875 20451
rect 13001 20349 13035 20383
rect 13277 20349 13311 20383
rect 14381 20349 14415 20383
rect 15393 20349 15427 20383
rect 15485 20349 15519 20383
rect 17969 20349 18003 20383
rect 20545 20349 20579 20383
rect 20729 20349 20763 20383
rect 24409 20349 24443 20383
rect 25145 20349 25179 20383
rect 27629 20349 27663 20383
rect 29377 20349 29411 20383
rect 31309 20349 31343 20383
rect 32505 20349 32539 20383
rect 33057 20349 33091 20383
rect 36093 20349 36127 20383
rect 38117 20349 38151 20383
rect 17877 20281 17911 20315
rect 19441 20281 19475 20315
rect 20177 20281 20211 20315
rect 22109 20281 22143 20315
rect 25513 20281 25547 20315
rect 27813 20281 27847 20315
rect 28365 20281 28399 20315
rect 31585 20281 31619 20315
rect 12449 20213 12483 20247
rect 15209 20213 15243 20247
rect 15301 20213 15335 20247
rect 16037 20213 16071 20247
rect 17233 20213 17267 20247
rect 27445 20213 27479 20247
rect 29653 20213 29687 20247
rect 31769 20213 31803 20247
rect 32965 20213 32999 20247
rect 33701 20213 33735 20247
rect 35633 20213 35667 20247
rect 36645 20213 36679 20247
rect 37473 20213 37507 20247
rect 12633 20009 12667 20043
rect 13277 20009 13311 20043
rect 16589 20009 16623 20043
rect 20453 20009 20487 20043
rect 21925 20009 21959 20043
rect 23949 20009 23983 20043
rect 31125 20009 31159 20043
rect 32137 20009 32171 20043
rect 33977 20009 34011 20043
rect 19993 19941 20027 19975
rect 25053 19941 25087 19975
rect 35633 19941 35667 19975
rect 17233 19873 17267 19907
rect 22937 19873 22971 19907
rect 24041 19873 24075 19907
rect 26249 19873 26283 19907
rect 28641 19873 28675 19907
rect 11253 19805 11287 19839
rect 13461 19805 13495 19839
rect 13737 19805 13771 19839
rect 14749 19805 14783 19839
rect 14841 19805 14875 19839
rect 15025 19805 15059 19839
rect 15117 19805 15151 19839
rect 15577 19805 15611 19839
rect 16957 19805 16991 19839
rect 17969 19805 18003 19839
rect 19625 19805 19659 19839
rect 20729 19805 20763 19839
rect 20821 19805 20855 19839
rect 20913 19805 20947 19839
rect 21097 19805 21131 19839
rect 22109 19805 22143 19839
rect 22201 19805 22235 19839
rect 22385 19805 22419 19839
rect 22477 19805 22511 19839
rect 23121 19805 23155 19839
rect 23765 19805 23799 19839
rect 23857 19805 23891 19839
rect 25329 19805 25363 19839
rect 26157 19805 26191 19839
rect 26709 19805 26743 19839
rect 26985 19805 27019 19839
rect 27353 19805 27387 19839
rect 28089 19805 28123 19839
rect 28273 19805 28307 19839
rect 29745 19805 29779 19839
rect 32321 19805 32355 19839
rect 32413 19805 32447 19839
rect 33425 19805 33459 19839
rect 33793 19805 33827 19839
rect 34989 19805 35023 19839
rect 35082 19805 35116 19839
rect 35265 19805 35299 19839
rect 35495 19805 35529 19839
rect 36093 19805 36127 19839
rect 36277 19805 36311 19839
rect 36921 19805 36955 19839
rect 37188 19805 37222 19839
rect 11520 19737 11554 19771
rect 15853 19737 15887 19771
rect 18705 19737 18739 19771
rect 19809 19737 19843 19771
rect 25513 19737 25547 19771
rect 25605 19737 25639 19771
rect 29990 19737 30024 19771
rect 32689 19737 32723 19771
rect 32781 19737 32815 19771
rect 33609 19737 33643 19771
rect 33701 19737 33735 19771
rect 35357 19737 35391 19771
rect 13645 19669 13679 19703
rect 14565 19669 14599 19703
rect 17049 19669 17083 19703
rect 23305 19669 23339 19703
rect 28273 19669 28307 19703
rect 36369 19669 36403 19703
rect 38301 19669 38335 19703
rect 13829 19465 13863 19499
rect 15025 19465 15059 19499
rect 20729 19465 20763 19499
rect 21189 19465 21223 19499
rect 25421 19465 25455 19499
rect 31493 19465 31527 19499
rect 32873 19465 32907 19499
rect 35357 19465 35391 19499
rect 14933 19397 14967 19431
rect 19349 19397 19383 19431
rect 22017 19397 22051 19431
rect 28825 19397 28859 19431
rect 29009 19397 29043 19431
rect 33517 19397 33551 19431
rect 33977 19397 34011 19431
rect 35081 19397 35115 19431
rect 38117 19397 38151 19431
rect 12449 19329 12483 19363
rect 14841 19329 14875 19363
rect 15853 19329 15887 19363
rect 17141 19329 17175 19363
rect 17325 19329 17359 19363
rect 18153 19329 18187 19363
rect 21097 19329 21131 19363
rect 23305 19329 23339 19363
rect 24317 19329 24351 19363
rect 24501 19329 24535 19363
rect 24593 19329 24627 19363
rect 24685 19329 24719 19363
rect 25329 19329 25363 19363
rect 25973 19329 26007 19363
rect 26157 19329 26191 19363
rect 26249 19329 26283 19363
rect 26393 19329 26427 19363
rect 27169 19329 27203 19363
rect 27353 19329 27387 19363
rect 27445 19329 27479 19363
rect 27565 19329 27599 19363
rect 29929 19329 29963 19363
rect 30205 19329 30239 19363
rect 30941 19329 30975 19363
rect 31125 19329 31159 19363
rect 31213 19329 31247 19363
rect 31355 19329 31389 19363
rect 33149 19329 33183 19363
rect 34161 19329 34195 19363
rect 34253 19329 34287 19363
rect 34713 19329 34747 19363
rect 34861 19329 34895 19363
rect 34989 19329 35023 19363
rect 35219 19329 35253 19363
rect 35817 19329 35851 19363
rect 36093 19329 36127 19363
rect 36737 19329 36771 19363
rect 36921 19329 36955 19363
rect 37841 19329 37875 19363
rect 12725 19261 12759 19295
rect 14565 19261 14599 19295
rect 15209 19261 15243 19295
rect 15301 19261 15335 19295
rect 15945 19261 15979 19295
rect 18245 19261 18279 19295
rect 18429 19261 18463 19295
rect 19441 19261 19475 19295
rect 19625 19261 19659 19295
rect 21373 19261 21407 19295
rect 23121 19261 23155 19295
rect 23581 19261 23615 19295
rect 29101 19261 29135 19295
rect 30113 19261 30147 19295
rect 33057 19261 33091 19295
rect 33425 19261 33459 19295
rect 36829 19261 36863 19295
rect 17141 19193 17175 19227
rect 17785 19193 17819 19227
rect 22385 19193 22419 19227
rect 27721 19193 27755 19227
rect 29745 19193 29779 19227
rect 33977 19193 34011 19227
rect 16037 19125 16071 19159
rect 16221 19125 16255 19159
rect 18981 19125 19015 19159
rect 22477 19125 22511 19159
rect 23489 19125 23523 19159
rect 24869 19125 24903 19159
rect 26525 19125 26559 19159
rect 28549 19125 28583 19159
rect 12909 18921 12943 18955
rect 13645 18921 13679 18955
rect 21189 18921 21223 18955
rect 21741 18921 21775 18955
rect 21833 18921 21867 18955
rect 23949 18921 23983 18955
rect 25881 18921 25915 18955
rect 27997 18921 28031 18955
rect 37933 18921 37967 18955
rect 15577 18853 15611 18887
rect 24685 18853 24719 18887
rect 27261 18853 27295 18887
rect 30481 18853 30515 18887
rect 35541 18853 35575 18887
rect 14565 18785 14599 18819
rect 16221 18785 16255 18819
rect 16681 18785 16715 18819
rect 18613 18785 18647 18819
rect 18797 18785 18831 18819
rect 21005 18785 21039 18819
rect 21925 18785 21959 18819
rect 25145 18785 25179 18819
rect 30932 18785 30966 18819
rect 31033 18785 31067 18819
rect 33241 18785 33275 18819
rect 33793 18785 33827 18819
rect 34345 18785 34379 18819
rect 12909 18717 12943 18751
rect 13093 18717 13127 18751
rect 13553 18717 13587 18751
rect 14749 18717 14783 18751
rect 15025 18717 15059 18751
rect 15761 18717 15795 18751
rect 16589 18717 16623 18751
rect 17325 18717 17359 18751
rect 17509 18717 17543 18751
rect 19625 18717 19659 18751
rect 20545 18717 20579 18751
rect 20913 18717 20947 18751
rect 21649 18717 21683 18751
rect 22937 18717 22971 18751
rect 23213 18717 23247 18751
rect 23857 18717 23891 18751
rect 25881 18717 25915 18751
rect 26065 18717 26099 18751
rect 26709 18717 26743 18751
rect 26893 18717 26927 18751
rect 27082 18717 27116 18751
rect 28181 18717 28215 18751
rect 28365 18717 28399 18751
rect 28457 18717 28491 18751
rect 29101 18717 29135 18751
rect 29193 18717 29227 18751
rect 29929 18717 29963 18751
rect 30113 18717 30147 18751
rect 30343 18717 30377 18751
rect 31217 18717 31251 18751
rect 31493 18717 31527 18751
rect 31677 18717 31711 18751
rect 32781 18717 32815 18751
rect 32873 18717 32907 18751
rect 33977 18717 34011 18751
rect 34897 18717 34931 18751
rect 34990 18717 35024 18751
rect 35173 18717 35207 18751
rect 35362 18717 35396 18751
rect 36553 18717 36587 18751
rect 14933 18649 14967 18683
rect 15485 18649 15519 18683
rect 15669 18649 15703 18683
rect 17693 18649 17727 18683
rect 18521 18649 18555 18683
rect 19441 18649 19475 18683
rect 19993 18649 20027 18683
rect 23673 18649 23707 18683
rect 25145 18649 25179 18683
rect 25237 18649 25271 18683
rect 26985 18649 27019 18683
rect 28917 18649 28951 18683
rect 30205 18649 30239 18683
rect 33149 18649 33183 18683
rect 35265 18649 35299 18683
rect 36798 18649 36832 18683
rect 16865 18581 16899 18615
rect 18153 18581 18187 18615
rect 22753 18581 22787 18615
rect 23121 18581 23155 18615
rect 26249 18581 26283 18615
rect 29015 18581 29049 18615
rect 32597 18581 32631 18615
rect 33977 18581 34011 18615
rect 14381 18377 14415 18411
rect 15577 18377 15611 18411
rect 19625 18377 19659 18411
rect 23121 18377 23155 18411
rect 24685 18377 24719 18411
rect 16037 18309 16071 18343
rect 20729 18309 20763 18343
rect 27353 18309 27387 18343
rect 35173 18309 35207 18343
rect 14105 18241 14139 18275
rect 14197 18241 14231 18275
rect 15393 18241 15427 18275
rect 16221 18241 16255 18275
rect 16313 18241 16347 18275
rect 17325 18241 17359 18275
rect 18337 18241 18371 18275
rect 18429 18241 18463 18275
rect 18613 18241 18647 18275
rect 18705 18241 18739 18275
rect 19533 18241 19567 18275
rect 22293 18241 22327 18275
rect 22385 18241 22419 18275
rect 22661 18241 22695 18275
rect 23305 18241 23339 18275
rect 23397 18241 23431 18275
rect 23673 18241 23707 18275
rect 24133 18241 24167 18275
rect 25697 18241 25731 18275
rect 25881 18241 25915 18275
rect 26433 18241 26467 18275
rect 26617 18241 26651 18275
rect 27169 18241 27203 18275
rect 27446 18241 27480 18275
rect 27565 18241 27599 18275
rect 29101 18241 29135 18275
rect 29285 18241 29319 18275
rect 29377 18241 29411 18275
rect 30021 18241 30055 18275
rect 30389 18241 30423 18275
rect 30849 18241 30883 18275
rect 32597 18263 32631 18297
rect 32965 18241 32999 18275
rect 33425 18241 33459 18275
rect 33518 18241 33552 18275
rect 33701 18241 33735 18275
rect 33793 18241 33827 18275
rect 33890 18241 33924 18275
rect 34805 18241 34839 18275
rect 34898 18241 34932 18275
rect 35081 18241 35115 18275
rect 35270 18241 35304 18275
rect 36093 18241 36127 18275
rect 36185 18241 36219 18275
rect 36461 18241 36495 18275
rect 37841 18241 37875 18275
rect 15209 18173 15243 18207
rect 17601 18173 17635 18207
rect 19809 18173 19843 18207
rect 20821 18173 20855 18207
rect 21005 18173 21039 18207
rect 24409 18173 24443 18207
rect 25973 18173 26007 18207
rect 30205 18173 30239 18207
rect 31585 18173 31619 18207
rect 32505 18173 32539 18207
rect 32873 18173 32907 18207
rect 35909 18173 35943 18207
rect 37933 18173 37967 18207
rect 38117 18173 38151 18207
rect 16129 18105 16163 18139
rect 17509 18105 17543 18139
rect 22569 18105 22603 18139
rect 28917 18105 28951 18139
rect 30021 18105 30055 18139
rect 35449 18105 35483 18139
rect 17141 18037 17175 18071
rect 18153 18037 18187 18071
rect 19165 18037 19199 18071
rect 20361 18037 20395 18071
rect 22109 18037 22143 18071
rect 23581 18037 23615 18071
rect 24225 18037 24259 18071
rect 25513 18037 25547 18071
rect 26525 18037 26559 18071
rect 27721 18037 27755 18071
rect 32321 18037 32355 18071
rect 34069 18037 34103 18071
rect 36369 18037 36403 18071
rect 37473 18037 37507 18071
rect 15025 17833 15059 17867
rect 17877 17833 17911 17867
rect 18705 17833 18739 17867
rect 22661 17833 22695 17867
rect 23581 17833 23615 17867
rect 23949 17833 23983 17867
rect 30113 17833 30147 17867
rect 32321 17833 32355 17867
rect 35357 17833 35391 17867
rect 36461 17833 36495 17867
rect 38301 17833 38335 17867
rect 20361 17765 20395 17799
rect 24777 17765 24811 17799
rect 27721 17765 27755 17799
rect 28365 17765 28399 17799
rect 33977 17765 34011 17799
rect 24869 17697 24903 17731
rect 32321 17697 32355 17731
rect 34897 17697 34931 17731
rect 36001 17697 36035 17731
rect 15209 17629 15243 17663
rect 15393 17629 15427 17663
rect 15485 17629 15519 17663
rect 15945 17629 15979 17663
rect 16773 17629 16807 17663
rect 17233 17629 17267 17663
rect 17785 17629 17819 17663
rect 18245 17629 18279 17663
rect 18705 17629 18739 17663
rect 18889 17629 18923 17663
rect 19533 17629 19567 17663
rect 19625 17629 19659 17663
rect 20637 17629 20671 17663
rect 20913 17629 20947 17663
rect 22845 17629 22879 17663
rect 23121 17629 23155 17663
rect 23765 17629 23799 17663
rect 24041 17629 24075 17663
rect 24593 17629 24627 17663
rect 24685 17629 24719 17663
rect 25789 17629 25823 17663
rect 27169 17629 27203 17663
rect 27589 17629 27623 17663
rect 29745 17629 29779 17663
rect 30573 17629 30607 17663
rect 31401 17629 31435 17663
rect 31953 17629 31987 17663
rect 33333 17629 33367 17663
rect 33426 17629 33460 17663
rect 33798 17629 33832 17663
rect 35081 17629 35115 17663
rect 35173 17629 35207 17663
rect 35449 17629 35483 17663
rect 36093 17629 36127 17663
rect 36921 17629 36955 17663
rect 37188 17629 37222 17663
rect 16405 17561 16439 17595
rect 20821 17561 20855 17595
rect 21465 17561 21499 17595
rect 21649 17561 21683 17595
rect 23029 17561 23063 17595
rect 26617 17561 26651 17595
rect 27353 17561 27387 17595
rect 27445 17561 27479 17595
rect 28641 17561 28675 17595
rect 28917 17561 28951 17595
rect 29929 17561 29963 17595
rect 33609 17561 33643 17595
rect 33701 17561 33735 17595
rect 19533 17493 19567 17527
rect 21833 17493 21867 17527
rect 28825 17493 28859 17527
rect 32137 17493 32171 17527
rect 15209 17289 15243 17323
rect 22115 17289 22149 17323
rect 23029 17289 23063 17323
rect 24869 17289 24903 17323
rect 30021 17289 30055 17323
rect 33885 17289 33919 17323
rect 37841 17289 37875 17323
rect 19625 17221 19659 17255
rect 22017 17221 22051 17255
rect 22201 17221 22235 17255
rect 33517 17221 33551 17255
rect 33609 17221 33643 17255
rect 34345 17221 34379 17255
rect 37933 17221 37967 17255
rect 14933 17153 14967 17187
rect 15025 17153 15059 17187
rect 15669 17153 15703 17187
rect 15853 17153 15887 17187
rect 15945 17153 15979 17187
rect 16129 17153 16163 17187
rect 16221 17153 16255 17187
rect 17233 17153 17267 17187
rect 17969 17153 18003 17187
rect 18705 17153 18739 17187
rect 19809 17153 19843 17187
rect 19901 17153 19935 17187
rect 20177 17153 20211 17187
rect 20637 17153 20671 17187
rect 20821 17153 20855 17187
rect 22293 17153 22327 17187
rect 22753 17153 22787 17187
rect 23489 17153 23523 17187
rect 23745 17153 23779 17187
rect 25697 17153 25731 17187
rect 27353 17153 27387 17187
rect 27445 17153 27479 17187
rect 28641 17153 28675 17187
rect 28908 17153 28942 17187
rect 30665 17153 30699 17187
rect 30758 17153 30792 17187
rect 30941 17153 30975 17187
rect 31033 17153 31067 17187
rect 31171 17153 31205 17187
rect 32505 17153 32539 17187
rect 33333 17153 33367 17187
rect 33701 17153 33735 17187
rect 34529 17153 34563 17187
rect 34621 17153 34655 17187
rect 34897 17153 34931 17187
rect 35541 17153 35575 17187
rect 36461 17153 36495 17187
rect 17509 17085 17543 17119
rect 18797 17085 18831 17119
rect 23029 17085 23063 17119
rect 25585 17085 25619 17119
rect 25973 17085 26007 17119
rect 26065 17085 26099 17119
rect 27169 17085 27203 17119
rect 27537 17085 27571 17119
rect 27629 17085 27663 17119
rect 32413 17085 32447 17119
rect 35817 17085 35851 17119
rect 36737 17085 36771 17119
rect 38117 17085 38151 17119
rect 18245 17017 18279 17051
rect 20085 17017 20119 17051
rect 25421 17017 25455 17051
rect 34805 17017 34839 17051
rect 17049 16949 17083 16983
rect 17417 16949 17451 16983
rect 20913 16949 20947 16983
rect 22845 16949 22879 16983
rect 31309 16949 31343 16983
rect 32781 16949 32815 16983
rect 37473 16949 37507 16983
rect 15025 16745 15059 16779
rect 23857 16745 23891 16779
rect 24961 16745 24995 16779
rect 30205 16745 30239 16779
rect 34345 16745 34379 16779
rect 36093 16745 36127 16779
rect 38209 16745 38243 16779
rect 16405 16677 16439 16711
rect 17693 16677 17727 16711
rect 26065 16677 26099 16711
rect 28457 16677 28491 16711
rect 32229 16677 32263 16711
rect 16497 16609 16531 16643
rect 18429 16609 18463 16643
rect 20269 16609 20303 16643
rect 22017 16609 22051 16643
rect 27353 16609 27387 16643
rect 27997 16609 28031 16643
rect 29837 16609 29871 16643
rect 30849 16609 30883 16643
rect 32965 16609 32999 16643
rect 34805 16609 34839 16643
rect 35265 16609 35299 16643
rect 36829 16609 36863 16643
rect 15853 16541 15887 16575
rect 16221 16541 16255 16575
rect 16773 16541 16807 16575
rect 17601 16541 17635 16575
rect 18153 16541 18187 16575
rect 20361 16541 20395 16575
rect 20545 16541 20579 16575
rect 21741 16541 21775 16575
rect 23857 16541 23891 16575
rect 24041 16541 24075 16575
rect 24593 16541 24627 16575
rect 25789 16541 25823 16575
rect 25881 16541 25915 16575
rect 26525 16541 26559 16575
rect 28089 16541 28123 16575
rect 28917 16541 28951 16575
rect 29101 16541 29135 16575
rect 29929 16541 29963 16575
rect 31116 16541 31150 16575
rect 34897 16541 34931 16575
rect 35633 16541 35667 16575
rect 35909 16541 35943 16575
rect 36001 16541 36035 16575
rect 37096 16541 37130 16575
rect 14841 16473 14875 16507
rect 21005 16473 21039 16507
rect 24777 16473 24811 16507
rect 29009 16473 29043 16507
rect 33232 16473 33266 16507
rect 15041 16405 15075 16439
rect 15209 16405 15243 16439
rect 23121 16405 23155 16439
rect 25421 16405 25455 16439
rect 36277 16405 36311 16439
rect 15393 16201 15427 16235
rect 21373 16201 21407 16235
rect 25881 16201 25915 16235
rect 27721 16201 27755 16235
rect 30849 16201 30883 16235
rect 33609 16201 33643 16235
rect 33977 16201 34011 16235
rect 36369 16201 36403 16235
rect 15945 16133 15979 16167
rect 23673 16133 23707 16167
rect 24501 16133 24535 16167
rect 35256 16133 35290 16167
rect 37933 16133 37967 16167
rect 15301 16065 15335 16099
rect 15485 16065 15519 16099
rect 16129 16065 16163 16099
rect 16865 16065 16899 16099
rect 16957 16065 16991 16099
rect 18521 16065 18555 16099
rect 18613 16065 18647 16099
rect 20361 16065 20395 16099
rect 20821 16065 20855 16099
rect 21281 16065 21315 16099
rect 22017 16065 22051 16099
rect 24317 16065 24351 16099
rect 24593 16065 24627 16099
rect 25789 16065 25823 16099
rect 27629 16065 27663 16099
rect 28549 16065 28583 16099
rect 28816 16065 28850 16099
rect 30757 16065 30791 16099
rect 31585 16065 31619 16099
rect 31769 16065 31803 16099
rect 32321 16065 32355 16099
rect 32689 16065 32723 16099
rect 32965 16065 32999 16099
rect 34069 16065 34103 16099
rect 37841 16065 37875 16099
rect 16313 15997 16347 16031
rect 19257 15997 19291 16031
rect 22293 15997 22327 16031
rect 25973 15997 26007 16031
rect 27813 15997 27847 16031
rect 31033 15997 31067 16031
rect 32597 15997 32631 16031
rect 34253 15997 34287 16031
rect 34989 15997 35023 16031
rect 38025 15997 38059 16031
rect 24133 15929 24167 15963
rect 20177 15861 20211 15895
rect 25421 15861 25455 15895
rect 27261 15861 27295 15895
rect 29929 15861 29963 15895
rect 30389 15861 30423 15895
rect 31677 15861 31711 15895
rect 37473 15861 37507 15895
rect 17693 15657 17727 15691
rect 18429 15657 18463 15691
rect 28457 15657 28491 15691
rect 29009 15657 29043 15691
rect 37381 15657 37415 15691
rect 20177 15589 20211 15623
rect 21557 15589 21591 15623
rect 31953 15589 31987 15623
rect 16313 15521 16347 15555
rect 18797 15521 18831 15555
rect 21741 15521 21775 15555
rect 23581 15521 23615 15555
rect 27077 15521 27111 15555
rect 31585 15521 31619 15555
rect 38117 15521 38151 15555
rect 16589 15453 16623 15487
rect 18613 15453 18647 15487
rect 18889 15453 18923 15487
rect 19533 15453 19567 15487
rect 19993 15453 20027 15487
rect 20269 15453 20303 15487
rect 20637 15453 20671 15487
rect 21557 15453 21591 15487
rect 21925 15453 21959 15487
rect 23397 15453 23431 15487
rect 27344 15453 27378 15487
rect 28917 15453 28951 15487
rect 29101 15453 29135 15487
rect 29745 15453 29779 15487
rect 32505 15453 32539 15487
rect 36001 15453 36035 15487
rect 36268 15453 36302 15487
rect 37841 15453 37875 15487
rect 23305 15385 23339 15419
rect 24593 15385 24627 15419
rect 30012 15385 30046 15419
rect 32750 15385 32784 15419
rect 35173 15385 35207 15419
rect 35357 15385 35391 15419
rect 22937 15317 22971 15351
rect 25881 15317 25915 15351
rect 31125 15317 31159 15351
rect 32045 15317 32079 15351
rect 33885 15317 33919 15351
rect 35541 15317 35575 15351
rect 21189 15113 21223 15147
rect 27629 15113 27663 15147
rect 29653 15113 29687 15147
rect 30021 15113 30055 15147
rect 30113 15113 30147 15147
rect 31033 15113 31067 15147
rect 32597 15113 32631 15147
rect 34713 15113 34747 15147
rect 36461 15113 36495 15147
rect 17877 15045 17911 15079
rect 31401 15045 31435 15079
rect 36093 15045 36127 15079
rect 36277 15045 36311 15079
rect 38117 15045 38151 15079
rect 17693 14977 17727 15011
rect 18153 14977 18187 15011
rect 19165 14977 19199 15011
rect 19809 14977 19843 15011
rect 21097 14977 21131 15011
rect 22385 14977 22419 15011
rect 22652 14977 22686 15011
rect 25044 14977 25078 15011
rect 27353 14977 27387 15011
rect 28181 14977 28215 15011
rect 28641 14977 28675 15011
rect 32321 14977 32355 15011
rect 33149 14977 33183 15011
rect 33517 14977 33551 15011
rect 33609 14977 33643 15011
rect 34621 14977 34655 15011
rect 34805 14977 34839 15011
rect 35357 14977 35391 15011
rect 35449 14977 35483 15011
rect 37841 14977 37875 15011
rect 19257 14909 19291 14943
rect 19533 14909 19567 14943
rect 21373 14909 21407 14943
rect 24777 14909 24811 14943
rect 28365 14909 28399 14943
rect 28549 14909 28583 14943
rect 30205 14909 30239 14943
rect 31493 14909 31527 14943
rect 31677 14909 31711 14943
rect 33333 14909 33367 14943
rect 19349 14841 19383 14875
rect 20729 14773 20763 14807
rect 23765 14773 23799 14807
rect 26157 14773 26191 14807
rect 35633 14773 35667 14807
rect 18889 14569 18923 14603
rect 23213 14569 23247 14603
rect 23857 14569 23891 14603
rect 25053 14569 25087 14603
rect 37105 14569 37139 14603
rect 18797 14501 18831 14535
rect 27537 14501 27571 14535
rect 28457 14433 28491 14467
rect 28549 14433 28583 14467
rect 38117 14433 38151 14467
rect 19533 14365 19567 14399
rect 20085 14365 20119 14399
rect 21833 14365 21867 14399
rect 25329 14365 25363 14399
rect 25421 14365 25455 14399
rect 25513 14365 25547 14399
rect 25697 14365 25731 14399
rect 26157 14365 26191 14399
rect 28365 14365 28399 14399
rect 30757 14365 30791 14399
rect 30849 14365 30883 14399
rect 31953 14365 31987 14399
rect 34897 14365 34931 14399
rect 36921 14365 36955 14399
rect 37841 14365 37875 14399
rect 23903 14331 23937 14365
rect 18429 14297 18463 14331
rect 22100 14297 22134 14331
rect 23673 14297 23707 14331
rect 26424 14297 26458 14331
rect 32198 14297 32232 14331
rect 33977 14297 34011 14331
rect 34161 14297 34195 14331
rect 34345 14297 34379 14331
rect 35142 14297 35176 14331
rect 36737 14297 36771 14331
rect 37565 14297 37599 14331
rect 24041 14229 24075 14263
rect 27997 14229 28031 14263
rect 30389 14229 30423 14263
rect 33333 14229 33367 14263
rect 36277 14229 36311 14263
rect 18981 14025 19015 14059
rect 21281 14025 21315 14059
rect 22477 14025 22511 14059
rect 27813 14025 27847 14059
rect 31677 14025 31711 14059
rect 32689 14025 32723 14059
rect 36093 14025 36127 14059
rect 36461 14025 36495 14059
rect 36829 14025 36863 14059
rect 38133 14025 38167 14059
rect 38301 14025 38335 14059
rect 23949 13957 23983 13991
rect 24041 13957 24075 13991
rect 29653 13957 29687 13991
rect 29837 13957 29871 13991
rect 30021 13957 30055 13991
rect 34958 13957 34992 13991
rect 37933 13957 37967 13991
rect 18797 13889 18831 13923
rect 18981 13889 19015 13923
rect 19993 13889 20027 13923
rect 22385 13889 22419 13923
rect 24777 13889 24811 13923
rect 25044 13889 25078 13923
rect 28365 13889 28399 13923
rect 28457 13889 28491 13923
rect 30757 13889 30791 13923
rect 30849 13889 30883 13923
rect 30941 13889 30975 13923
rect 31125 13889 31159 13923
rect 31585 13889 31619 13923
rect 32413 13889 32447 13923
rect 33241 13889 33275 13923
rect 33609 13889 33643 13923
rect 33885 13889 33919 13923
rect 34713 13889 34747 13923
rect 36277 13889 36311 13923
rect 37657 13889 37691 13923
rect 19717 13821 19751 13855
rect 22661 13821 22695 13855
rect 23949 13821 23983 13855
rect 33425 13821 33459 13855
rect 23489 13753 23523 13787
rect 30481 13753 30515 13787
rect 22017 13685 22051 13719
rect 26157 13685 26191 13719
rect 38117 13685 38151 13719
rect 19441 13481 19475 13515
rect 20269 13481 20303 13515
rect 22201 13481 22235 13515
rect 24593 13481 24627 13515
rect 25329 13481 25363 13515
rect 31953 13481 31987 13515
rect 33609 13481 33643 13515
rect 34897 13481 34931 13515
rect 36829 13481 36863 13515
rect 38301 13481 38335 13515
rect 24041 13413 24075 13447
rect 36093 13413 36127 13447
rect 20361 13345 20395 13379
rect 22661 13345 22695 13379
rect 25973 13345 26007 13379
rect 27813 13345 27847 13379
rect 29837 13345 29871 13379
rect 32413 13345 32447 13379
rect 32505 13345 32539 13379
rect 34161 13345 34195 13379
rect 35449 13345 35483 13379
rect 37473 13345 37507 13379
rect 19441 13277 19475 13311
rect 19625 13277 19659 13311
rect 20085 13277 20119 13311
rect 20177 13277 20211 13311
rect 20821 13277 20855 13311
rect 24593 13277 24627 13311
rect 24777 13277 24811 13311
rect 24869 13277 24903 13311
rect 25697 13277 25731 13311
rect 26617 13277 26651 13311
rect 26893 13277 26927 13311
rect 34069 13277 34103 13311
rect 35357 13277 35391 13311
rect 36093 13277 36127 13311
rect 36277 13277 36311 13311
rect 36737 13277 36771 13311
rect 36921 13277 36955 13311
rect 37381 13277 37415 13311
rect 37565 13277 37599 13311
rect 21088 13209 21122 13243
rect 22928 13209 22962 13243
rect 26801 13209 26835 13243
rect 27353 13209 27387 13243
rect 28080 13209 28114 13243
rect 30104 13209 30138 13243
rect 25789 13141 25823 13175
rect 29193 13141 29227 13175
rect 31217 13141 31251 13175
rect 32321 13141 32355 13175
rect 33977 13141 34011 13175
rect 35265 13141 35299 13175
rect 23581 12937 23615 12971
rect 23949 12937 23983 12971
rect 28641 12937 28675 12971
rect 29101 12937 29135 12971
rect 30297 12937 30331 12971
rect 30665 12937 30699 12971
rect 30757 12937 30791 12971
rect 31677 12937 31711 12971
rect 35909 12937 35943 12971
rect 36553 12937 36587 12971
rect 20453 12869 20487 12903
rect 21281 12869 21315 12903
rect 24041 12869 24075 12903
rect 25329 12869 25363 12903
rect 20269 12801 20303 12835
rect 20545 12801 20579 12835
rect 21005 12801 21039 12835
rect 22661 12801 22695 12835
rect 24777 12801 24811 12835
rect 24869 12801 24903 12835
rect 26157 12801 26191 12835
rect 26617 12801 26651 12835
rect 27537 12801 27571 12835
rect 27629 12801 27663 12835
rect 27721 12801 27755 12835
rect 29009 12801 29043 12835
rect 31585 12801 31619 12835
rect 31769 12801 31803 12835
rect 32321 12801 32355 12835
rect 32873 12801 32907 12835
rect 33149 12801 33183 12835
rect 33517 12801 33551 12835
rect 33701 12801 33735 12835
rect 34989 12801 35023 12835
rect 35817 12801 35851 12835
rect 36001 12801 36035 12835
rect 36461 12801 36495 12835
rect 36645 12801 36679 12835
rect 22569 12733 22603 12767
rect 24225 12733 24259 12767
rect 26065 12733 26099 12767
rect 29193 12733 29227 12767
rect 30849 12733 30883 12767
rect 33241 12733 33275 12767
rect 35081 12733 35115 12767
rect 35173 12733 35207 12767
rect 20269 12597 20303 12631
rect 22845 12597 22879 12631
rect 27905 12597 27939 12631
rect 34621 12597 34655 12631
rect 38301 12597 38335 12631
rect 23857 12393 23891 12427
rect 28549 12393 28583 12427
rect 36277 12393 36311 12427
rect 20821 12325 20855 12359
rect 22569 12325 22603 12359
rect 24041 12325 24075 12359
rect 30573 12325 30607 12359
rect 32689 12325 32723 12359
rect 19441 12257 19475 12291
rect 21833 12257 21867 12291
rect 23121 12257 23155 12291
rect 25605 12257 25639 12291
rect 27353 12257 27387 12291
rect 30113 12257 30147 12291
rect 33425 12257 33459 12291
rect 33609 12257 33643 12291
rect 22845 12189 22879 12223
rect 26617 12189 26651 12223
rect 26709 12189 26743 12223
rect 26893 12189 26927 12223
rect 28825 12189 28859 12223
rect 28917 12189 28951 12223
rect 29009 12189 29043 12223
rect 29193 12189 29227 12223
rect 29929 12189 29963 12223
rect 30849 12189 30883 12223
rect 30941 12189 30975 12223
rect 31033 12189 31067 12223
rect 31217 12189 31251 12223
rect 31677 12189 31711 12223
rect 31861 12189 31895 12223
rect 32413 12189 32447 12223
rect 33333 12189 33367 12223
rect 33885 12189 33919 12223
rect 34897 12189 34931 12223
rect 35153 12189 35187 12223
rect 19708 12121 19742 12155
rect 21649 12121 21683 12155
rect 23673 12121 23707 12155
rect 23889 12121 23923 12155
rect 25421 12121 25455 12155
rect 29745 12121 29779 12155
rect 21281 12053 21315 12087
rect 21741 12053 21775 12087
rect 23029 12053 23063 12087
rect 24961 12053 24995 12087
rect 25329 12053 25363 12087
rect 31769 12053 31803 12087
rect 21005 11849 21039 11883
rect 21097 11849 21131 11883
rect 25697 11849 25731 11883
rect 26525 11849 26559 11883
rect 27169 11849 27203 11883
rect 28365 11849 28399 11883
rect 33701 11849 33735 11883
rect 35633 11849 35667 11883
rect 22477 11781 22511 11815
rect 24584 11781 24618 11815
rect 26157 11781 26191 11815
rect 27537 11781 27571 11815
rect 22385 11713 22419 11747
rect 23213 11713 23247 11747
rect 26341 11713 26375 11747
rect 28733 11713 28767 11747
rect 29929 11713 29963 11747
rect 31125 11713 31159 11747
rect 32781 11713 32815 11747
rect 33609 11713 33643 11747
rect 33793 11713 33827 11747
rect 34520 11713 34554 11747
rect 21281 11645 21315 11679
rect 22661 11645 22695 11679
rect 23397 11645 23431 11679
rect 24317 11645 24351 11679
rect 27629 11645 27663 11679
rect 27813 11645 27847 11679
rect 28825 11645 28859 11679
rect 28917 11645 28951 11679
rect 30021 11645 30055 11679
rect 30205 11645 30239 11679
rect 31217 11645 31251 11679
rect 31309 11645 31343 11679
rect 32873 11645 32907 11679
rect 32965 11645 32999 11679
rect 34253 11645 34287 11679
rect 20637 11509 20671 11543
rect 22017 11509 22051 11543
rect 29561 11509 29595 11543
rect 30757 11509 30791 11543
rect 32413 11509 32447 11543
rect 22385 11305 22419 11339
rect 25973 11305 26007 11339
rect 29193 11305 29227 11339
rect 31769 11305 31803 11339
rect 33609 11305 33643 11339
rect 34897 11305 34931 11339
rect 21005 11169 21039 11203
rect 23765 11169 23799 11203
rect 23949 11169 23983 11203
rect 24593 11169 24627 11203
rect 26893 11169 26927 11203
rect 27077 11169 27111 11203
rect 27813 11169 27847 11203
rect 30389 11169 30423 11203
rect 35449 11169 35483 11203
rect 21272 11101 21306 11135
rect 24860 11101 24894 11135
rect 26801 11101 26835 11135
rect 28080 11101 28114 11135
rect 32229 11101 32263 11135
rect 32496 11101 32530 11135
rect 35265 11101 35299 11135
rect 37841 11101 37875 11135
rect 30645 11033 30679 11067
rect 38117 11033 38151 11067
rect 23305 10965 23339 10999
rect 23673 10965 23707 10999
rect 26433 10965 26467 10999
rect 35357 10965 35391 10999
rect 21097 10761 21131 10795
rect 22293 10761 22327 10795
rect 26617 10761 26651 10795
rect 31309 10761 31343 10795
rect 33701 10761 33735 10795
rect 19984 10693 20018 10727
rect 19717 10625 19751 10659
rect 22017 10625 22051 10659
rect 22753 10625 22787 10659
rect 23020 10625 23054 10659
rect 25237 10625 25271 10659
rect 25504 10625 25538 10659
rect 28089 10625 28123 10659
rect 28356 10625 28390 10659
rect 29929 10625 29963 10659
rect 30196 10625 30230 10659
rect 32321 10625 32355 10659
rect 32577 10625 32611 10659
rect 22109 10557 22143 10591
rect 22293 10557 22327 10591
rect 24133 10421 24167 10455
rect 29469 10421 29503 10455
rect 22109 10217 22143 10251
rect 23121 10217 23155 10251
rect 27537 10217 27571 10251
rect 27997 10217 28031 10251
rect 30205 10217 30239 10251
rect 32413 10217 32447 10251
rect 28457 10081 28491 10115
rect 28641 10081 28675 10115
rect 30757 10081 30791 10115
rect 32873 10081 32907 10115
rect 32965 10081 32999 10115
rect 22017 10013 22051 10047
rect 22201 10013 22235 10047
rect 23305 10013 23339 10047
rect 23581 10013 23615 10047
rect 26157 10013 26191 10047
rect 28365 10013 28399 10047
rect 30573 10013 30607 10047
rect 31585 10013 31619 10047
rect 32781 10013 32815 10047
rect 37841 10013 37875 10047
rect 26424 9945 26458 9979
rect 31401 9945 31435 9979
rect 38117 9945 38151 9979
rect 23489 9877 23523 9911
rect 30665 9877 30699 9911
rect 31769 9877 31803 9911
rect 27169 9673 27203 9707
rect 27537 9673 27571 9707
rect 27629 9673 27663 9707
rect 28549 9673 28583 9707
rect 29009 9673 29043 9707
rect 28917 9605 28951 9639
rect 29929 9605 29963 9639
rect 30757 9605 30791 9639
rect 29745 9537 29779 9571
rect 31033 9537 31067 9571
rect 31125 9537 31159 9571
rect 31217 9537 31251 9571
rect 31401 9537 31435 9571
rect 27721 9469 27755 9503
rect 29101 9469 29135 9503
rect 30113 9469 30147 9503
rect 37841 8449 37875 8483
rect 38117 8381 38151 8415
rect 37841 7361 37875 7395
rect 38117 7293 38151 7327
rect 37841 5661 37875 5695
rect 38117 5593 38151 5627
rect 37841 4573 37875 4607
rect 38117 4505 38151 4539
rect 37841 3009 37875 3043
rect 38117 2941 38151 2975
rect 37841 2397 37875 2431
rect 38117 2329 38151 2363
<< metal1 >>
rect 4982 39244 4988 39296
rect 5040 39284 5046 39296
rect 5040 39256 31616 39284
rect 5040 39244 5046 39256
rect 5902 39176 5908 39228
rect 5960 39216 5966 39228
rect 5960 39188 28304 39216
rect 5960 39176 5966 39188
rect 28276 39160 28304 39188
rect 31588 39160 31616 39256
rect 10502 39108 10508 39160
rect 10560 39148 10566 39160
rect 11698 39148 11704 39160
rect 10560 39120 11704 39148
rect 10560 39108 10566 39120
rect 11698 39108 11704 39120
rect 11756 39108 11762 39160
rect 21634 39108 21640 39160
rect 21692 39148 21698 39160
rect 22094 39148 22100 39160
rect 21692 39120 22100 39148
rect 21692 39108 21698 39120
rect 22094 39108 22100 39120
rect 22152 39108 22158 39160
rect 28258 39108 28264 39160
rect 28316 39108 28322 39160
rect 31570 39108 31576 39160
rect 31628 39108 31634 39160
rect 3970 38972 3976 39024
rect 4028 39012 4034 39024
rect 23290 39012 23296 39024
rect 4028 38984 23296 39012
rect 4028 38972 4034 38984
rect 23290 38972 23296 38984
rect 23348 38972 23354 39024
rect 5258 38904 5264 38956
rect 5316 38944 5322 38956
rect 18598 38944 18604 38956
rect 5316 38916 18604 38944
rect 5316 38904 5322 38916
rect 18598 38904 18604 38916
rect 18656 38904 18662 38956
rect 3326 38836 3332 38888
rect 3384 38876 3390 38888
rect 23382 38876 23388 38888
rect 3384 38848 23388 38876
rect 3384 38836 3390 38848
rect 23382 38836 23388 38848
rect 23440 38836 23446 38888
rect 5534 38768 5540 38820
rect 5592 38808 5598 38820
rect 16942 38808 16948 38820
rect 5592 38780 16948 38808
rect 5592 38768 5598 38780
rect 16942 38768 16948 38780
rect 17000 38768 17006 38820
rect 18138 38768 18144 38820
rect 18196 38808 18202 38820
rect 20162 38808 20168 38820
rect 18196 38780 20168 38808
rect 18196 38768 18202 38780
rect 20162 38768 20168 38780
rect 20220 38808 20226 38820
rect 26878 38808 26884 38820
rect 20220 38780 26884 38808
rect 20220 38768 20226 38780
rect 26878 38768 26884 38780
rect 26936 38768 26942 38820
rect 6638 38700 6644 38752
rect 6696 38740 6702 38752
rect 22278 38740 22284 38752
rect 6696 38712 22284 38740
rect 6696 38700 6702 38712
rect 22278 38700 22284 38712
rect 22336 38700 22342 38752
rect 23198 38700 23204 38752
rect 23256 38740 23262 38752
rect 34238 38740 34244 38752
rect 23256 38712 34244 38740
rect 23256 38700 23262 38712
rect 34238 38700 34244 38712
rect 34296 38700 34302 38752
rect 13722 38632 13728 38684
rect 13780 38672 13786 38684
rect 26786 38672 26792 38684
rect 13780 38644 26792 38672
rect 13780 38632 13786 38644
rect 26786 38632 26792 38644
rect 26844 38632 26850 38684
rect 6178 38564 6184 38616
rect 6236 38604 6242 38616
rect 31938 38604 31944 38616
rect 6236 38576 31944 38604
rect 6236 38564 6242 38576
rect 31938 38564 31944 38576
rect 31996 38564 32002 38616
rect 3050 38496 3056 38548
rect 3108 38536 3114 38548
rect 23658 38536 23664 38548
rect 3108 38508 23664 38536
rect 3108 38496 3114 38508
rect 23658 38496 23664 38508
rect 23716 38496 23722 38548
rect 6270 38428 6276 38480
rect 6328 38468 6334 38480
rect 17954 38468 17960 38480
rect 6328 38440 17960 38468
rect 6328 38428 6334 38440
rect 17954 38428 17960 38440
rect 18012 38428 18018 38480
rect 18230 38428 18236 38480
rect 18288 38468 18294 38480
rect 32490 38468 32496 38480
rect 18288 38440 32496 38468
rect 18288 38428 18294 38440
rect 32490 38428 32496 38440
rect 32548 38428 32554 38480
rect 7742 38360 7748 38412
rect 7800 38400 7806 38412
rect 25958 38400 25964 38412
rect 7800 38372 25964 38400
rect 7800 38360 7806 38372
rect 25958 38360 25964 38372
rect 26016 38360 26022 38412
rect 7006 38292 7012 38344
rect 7064 38332 7070 38344
rect 18138 38332 18144 38344
rect 7064 38304 18144 38332
rect 7064 38292 7070 38304
rect 18138 38292 18144 38304
rect 18196 38292 18202 38344
rect 26142 38292 26148 38344
rect 26200 38332 26206 38344
rect 31754 38332 31760 38344
rect 26200 38304 31760 38332
rect 26200 38292 26206 38304
rect 31754 38292 31760 38304
rect 31812 38292 31818 38344
rect 5994 38224 6000 38276
rect 6052 38264 6058 38276
rect 35710 38264 35716 38276
rect 6052 38236 35716 38264
rect 6052 38224 6058 38236
rect 35710 38224 35716 38236
rect 35768 38224 35774 38276
rect 5810 38156 5816 38208
rect 5868 38196 5874 38208
rect 33686 38196 33692 38208
rect 5868 38168 33692 38196
rect 5868 38156 5874 38168
rect 33686 38156 33692 38168
rect 33744 38156 33750 38208
rect 6362 38088 6368 38140
rect 6420 38128 6426 38140
rect 16482 38128 16488 38140
rect 6420 38100 16488 38128
rect 6420 38088 6426 38100
rect 16482 38088 16488 38100
rect 16540 38088 16546 38140
rect 20898 38088 20904 38140
rect 20956 38128 20962 38140
rect 35342 38128 35348 38140
rect 20956 38100 35348 38128
rect 20956 38088 20962 38100
rect 35342 38088 35348 38100
rect 35400 38088 35406 38140
rect 4062 38020 4068 38072
rect 4120 38060 4126 38072
rect 23014 38060 23020 38072
rect 4120 38032 23020 38060
rect 4120 38020 4126 38032
rect 23014 38020 23020 38032
rect 23072 38020 23078 38072
rect 25498 38020 25504 38072
rect 25556 38060 25562 38072
rect 30558 38060 30564 38072
rect 25556 38032 30564 38060
rect 25556 38020 25562 38032
rect 30558 38020 30564 38032
rect 30616 38020 30622 38072
rect 30650 38020 30656 38072
rect 30708 38060 30714 38072
rect 32766 38060 32772 38072
rect 30708 38032 32772 38060
rect 30708 38020 30714 38032
rect 32766 38020 32772 38032
rect 32824 38020 32830 38072
rect 2590 37952 2596 38004
rect 2648 37992 2654 38004
rect 13722 37992 13728 38004
rect 2648 37964 13728 37992
rect 2648 37952 2654 37964
rect 13722 37952 13728 37964
rect 13780 37952 13786 38004
rect 21266 37952 21272 38004
rect 21324 37992 21330 38004
rect 35434 37992 35440 38004
rect 21324 37964 35440 37992
rect 21324 37952 21330 37964
rect 35434 37952 35440 37964
rect 35492 37952 35498 38004
rect 7282 37884 7288 37936
rect 7340 37924 7346 37936
rect 27522 37924 27528 37936
rect 7340 37896 27528 37924
rect 7340 37884 7346 37896
rect 27522 37884 27528 37896
rect 27580 37884 27586 37936
rect 4798 37816 4804 37868
rect 4856 37856 4862 37868
rect 26326 37856 26332 37868
rect 4856 37828 26332 37856
rect 4856 37816 4862 37828
rect 26326 37816 26332 37828
rect 26384 37816 26390 37868
rect 26970 37816 26976 37868
rect 27028 37856 27034 37868
rect 33318 37856 33324 37868
rect 27028 37828 33324 37856
rect 27028 37816 27034 37828
rect 33318 37816 33324 37828
rect 33376 37816 33382 37868
rect 6730 37748 6736 37800
rect 6788 37788 6794 37800
rect 31386 37788 31392 37800
rect 6788 37760 31392 37788
rect 6788 37748 6794 37760
rect 31386 37748 31392 37760
rect 31444 37748 31450 37800
rect 6914 37680 6920 37732
rect 6972 37720 6978 37732
rect 30650 37720 30656 37732
rect 6972 37692 30656 37720
rect 6972 37680 6978 37692
rect 30650 37680 30656 37692
rect 30708 37680 30714 37732
rect 3694 37612 3700 37664
rect 3752 37652 3758 37664
rect 20714 37652 20720 37664
rect 3752 37624 20720 37652
rect 3752 37612 3758 37624
rect 20714 37612 20720 37624
rect 20772 37612 20778 37664
rect 21910 37612 21916 37664
rect 21968 37652 21974 37664
rect 25498 37652 25504 37664
rect 21968 37624 25504 37652
rect 21968 37612 21974 37624
rect 25498 37612 25504 37624
rect 25556 37612 25562 37664
rect 26234 37612 26240 37664
rect 26292 37652 26298 37664
rect 34146 37652 34152 37664
rect 26292 37624 34152 37652
rect 26292 37612 26298 37624
rect 34146 37612 34152 37624
rect 34204 37612 34210 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 11054 37448 11060 37460
rect 7852 37420 11060 37448
rect 3160 37284 3556 37312
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 1949 37247 2007 37253
rect 1949 37244 1961 37247
rect 1820 37216 1961 37244
rect 1820 37204 1826 37216
rect 1949 37213 1961 37216
rect 1995 37213 2007 37247
rect 1949 37207 2007 37213
rect 2501 37179 2559 37185
rect 2501 37145 2513 37179
rect 2547 37176 2559 37179
rect 3160 37176 3188 37284
rect 3237 37247 3295 37253
rect 3237 37213 3249 37247
rect 3283 37213 3295 37247
rect 3237 37207 3295 37213
rect 2547 37148 3188 37176
rect 2547 37145 2559 37148
rect 2501 37139 2559 37145
rect 3252 37108 3280 37207
rect 3418 37204 3424 37256
rect 3476 37204 3482 37256
rect 3528 37244 3556 37284
rect 4448 37284 5396 37312
rect 4448 37244 4476 37284
rect 3528 37216 4476 37244
rect 4522 37204 4528 37256
rect 4580 37204 4586 37256
rect 4614 37204 4620 37256
rect 4672 37244 4678 37256
rect 4709 37247 4767 37253
rect 4709 37244 4721 37247
rect 4672 37216 4721 37244
rect 4672 37204 4678 37216
rect 4709 37213 4721 37216
rect 4755 37213 4767 37247
rect 4709 37207 4767 37213
rect 5074 37204 5080 37256
rect 5132 37244 5138 37256
rect 5261 37247 5319 37253
rect 5261 37244 5273 37247
rect 5132 37216 5273 37244
rect 5132 37204 5138 37216
rect 5261 37213 5273 37216
rect 5307 37213 5319 37247
rect 5368 37244 5396 37284
rect 7006 37272 7012 37324
rect 7064 37272 7070 37324
rect 5368 37216 7144 37244
rect 5261 37207 5319 37213
rect 3329 37179 3387 37185
rect 3329 37145 3341 37179
rect 3375 37176 3387 37179
rect 5718 37176 5724 37188
rect 3375 37148 5724 37176
rect 3375 37145 3387 37148
rect 3329 37139 3387 37145
rect 5718 37136 5724 37148
rect 5776 37136 5782 37188
rect 5813 37179 5871 37185
rect 5813 37145 5825 37179
rect 5859 37176 5871 37179
rect 6546 37176 6552 37188
rect 5859 37148 6552 37176
rect 5859 37145 5871 37148
rect 5813 37139 5871 37145
rect 6546 37136 6552 37148
rect 6604 37136 6610 37188
rect 7116 37176 7144 37216
rect 7190 37204 7196 37256
rect 7248 37244 7254 37256
rect 7852 37244 7880 37420
rect 11054 37408 11060 37420
rect 11112 37408 11118 37460
rect 15194 37408 15200 37460
rect 15252 37448 15258 37460
rect 15252 37420 20760 37448
rect 15252 37408 15258 37420
rect 8570 37340 8576 37392
rect 8628 37380 8634 37392
rect 16482 37380 16488 37392
rect 8628 37352 16488 37380
rect 8628 37340 8634 37352
rect 16482 37340 16488 37352
rect 16540 37340 16546 37392
rect 9490 37272 9496 37324
rect 9548 37312 9554 37324
rect 9677 37315 9735 37321
rect 9677 37312 9689 37315
rect 9548 37284 9689 37312
rect 9548 37272 9554 37284
rect 9677 37281 9689 37284
rect 9723 37312 9735 37315
rect 10962 37312 10968 37324
rect 9723 37284 10968 37312
rect 9723 37281 9735 37284
rect 9677 37275 9735 37281
rect 10962 37272 10968 37284
rect 11020 37312 11026 37324
rect 12345 37315 12403 37321
rect 12345 37312 12357 37315
rect 11020 37284 12357 37312
rect 11020 37272 11026 37284
rect 12345 37281 12357 37284
rect 12391 37312 12403 37315
rect 13541 37315 13599 37321
rect 13541 37312 13553 37315
rect 12391 37284 13553 37312
rect 12391 37281 12403 37284
rect 12345 37275 12403 37281
rect 13541 37281 13553 37284
rect 13587 37312 13599 37315
rect 14826 37312 14832 37324
rect 13587 37284 14832 37312
rect 13587 37281 13599 37284
rect 13541 37275 13599 37281
rect 14826 37272 14832 37284
rect 14884 37272 14890 37324
rect 19705 37315 19763 37321
rect 19705 37281 19717 37315
rect 19751 37312 19763 37315
rect 20070 37312 20076 37324
rect 19751 37284 20076 37312
rect 19751 37281 19763 37284
rect 19705 37275 19763 37281
rect 20070 37272 20076 37284
rect 20128 37272 20134 37324
rect 20732 37312 20760 37420
rect 20990 37408 20996 37460
rect 21048 37448 21054 37460
rect 22554 37448 22560 37460
rect 21048 37420 22560 37448
rect 21048 37408 21054 37420
rect 22554 37408 22560 37420
rect 22612 37408 22618 37460
rect 25774 37408 25780 37460
rect 25832 37448 25838 37460
rect 26237 37451 26295 37457
rect 26237 37448 26249 37451
rect 25832 37420 26249 37448
rect 25832 37408 25838 37420
rect 26237 37417 26249 37420
rect 26283 37417 26295 37451
rect 26237 37411 26295 37417
rect 27614 37408 27620 37460
rect 27672 37448 27678 37460
rect 32585 37451 32643 37457
rect 27672 37420 31754 37448
rect 27672 37408 27678 37420
rect 24302 37340 24308 37392
rect 24360 37380 24366 37392
rect 28442 37380 28448 37392
rect 24360 37352 28448 37380
rect 24360 37340 24366 37352
rect 28442 37340 28448 37352
rect 28500 37340 28506 37392
rect 31726 37380 31754 37420
rect 32585 37417 32597 37451
rect 32631 37448 32643 37451
rect 32950 37448 32956 37460
rect 32631 37420 32956 37448
rect 32631 37417 32643 37420
rect 32585 37411 32643 37417
rect 32950 37408 32956 37420
rect 33008 37408 33014 37460
rect 33229 37451 33287 37457
rect 33229 37417 33241 37451
rect 33275 37448 33287 37451
rect 38470 37448 38476 37460
rect 33275 37420 38476 37448
rect 33275 37417 33287 37420
rect 33229 37411 33287 37417
rect 38470 37408 38476 37420
rect 38528 37408 38534 37460
rect 34514 37380 34520 37392
rect 31726 37352 34520 37380
rect 34514 37340 34520 37352
rect 34572 37340 34578 37392
rect 26970 37312 26976 37324
rect 20732 37284 22232 37312
rect 7248 37216 7880 37244
rect 7929 37247 7987 37253
rect 7248 37204 7254 37216
rect 7929 37213 7941 37247
rect 7975 37244 7987 37247
rect 8202 37244 8208 37256
rect 7975 37216 8208 37244
rect 7975 37213 7987 37216
rect 7929 37207 7987 37213
rect 8202 37204 8208 37216
rect 8260 37204 8266 37256
rect 10502 37204 10508 37256
rect 10560 37204 10566 37256
rect 10612 37216 14228 37244
rect 7116 37148 8432 37176
rect 3510 37108 3516 37120
rect 3252 37080 3516 37108
rect 3510 37068 3516 37080
rect 3568 37068 3574 37120
rect 3786 37068 3792 37120
rect 3844 37108 3850 37120
rect 4157 37111 4215 37117
rect 4157 37108 4169 37111
rect 3844 37080 4169 37108
rect 3844 37068 3850 37080
rect 4157 37077 4169 37080
rect 4203 37108 4215 37111
rect 4614 37108 4620 37120
rect 4203 37080 4620 37108
rect 4203 37077 4215 37080
rect 4157 37071 4215 37077
rect 4614 37068 4620 37080
rect 4672 37068 4678 37120
rect 4706 37068 4712 37120
rect 4764 37068 4770 37120
rect 7282 37068 7288 37120
rect 7340 37108 7346 37120
rect 7377 37111 7435 37117
rect 7377 37108 7389 37111
rect 7340 37080 7389 37108
rect 7340 37068 7346 37080
rect 7377 37077 7389 37080
rect 7423 37077 7435 37111
rect 8404 37108 8432 37148
rect 8478 37136 8484 37188
rect 8536 37136 8542 37188
rect 9674 37176 9680 37188
rect 8588 37148 9680 37176
rect 8588 37108 8616 37148
rect 8404 37080 8616 37108
rect 7377 37071 7435 37077
rect 9122 37068 9128 37120
rect 9180 37068 9186 37120
rect 9508 37117 9536 37148
rect 9674 37136 9680 37148
rect 9732 37136 9738 37188
rect 9766 37136 9772 37188
rect 9824 37176 9830 37188
rect 10612 37176 10640 37216
rect 9824 37148 10640 37176
rect 11057 37179 11115 37185
rect 9824 37136 9830 37148
rect 11057 37145 11069 37179
rect 11103 37176 11115 37179
rect 12161 37179 12219 37185
rect 12161 37176 12173 37179
rect 11103 37148 12173 37176
rect 11103 37145 11115 37148
rect 11057 37139 11115 37145
rect 12161 37145 12173 37148
rect 12207 37176 12219 37179
rect 12434 37176 12440 37188
rect 12207 37148 12440 37176
rect 12207 37145 12219 37148
rect 12161 37139 12219 37145
rect 12434 37136 12440 37148
rect 12492 37136 12498 37188
rect 14200 37176 14228 37216
rect 14366 37204 14372 37256
rect 14424 37204 14430 37256
rect 14553 37247 14611 37253
rect 14553 37213 14565 37247
rect 14599 37244 14611 37247
rect 14642 37244 14648 37256
rect 14599 37216 14648 37244
rect 14599 37213 14611 37216
rect 14553 37207 14611 37213
rect 14642 37204 14648 37216
rect 14700 37204 14706 37256
rect 15010 37204 15016 37256
rect 15068 37244 15074 37256
rect 15105 37247 15163 37253
rect 15105 37244 15117 37247
rect 15068 37216 15117 37244
rect 15068 37204 15074 37216
rect 15105 37213 15117 37216
rect 15151 37213 15163 37247
rect 15105 37207 15163 37213
rect 17034 37204 17040 37256
rect 17092 37204 17098 37256
rect 17957 37247 18015 37253
rect 17957 37213 17969 37247
rect 18003 37244 18015 37247
rect 18322 37244 18328 37256
rect 18003 37216 18328 37244
rect 18003 37213 18015 37216
rect 17957 37207 18015 37213
rect 18322 37204 18328 37216
rect 18380 37204 18386 37256
rect 19242 37204 19248 37256
rect 19300 37244 19306 37256
rect 19429 37247 19487 37253
rect 19429 37244 19441 37247
rect 19300 37216 19441 37244
rect 19300 37204 19306 37216
rect 19429 37213 19441 37216
rect 19475 37213 19487 37247
rect 19429 37207 19487 37213
rect 22094 37204 22100 37256
rect 22152 37204 22158 37256
rect 22204 37244 22232 37284
rect 23492 37284 26976 37312
rect 23492 37244 23520 37284
rect 26970 37272 26976 37284
rect 27028 37272 27034 37324
rect 28074 37272 28080 37324
rect 28132 37312 28138 37324
rect 28132 37284 28212 37312
rect 28132 37272 28138 37284
rect 22204 37216 23520 37244
rect 23566 37204 23572 37256
rect 23624 37204 23630 37256
rect 24946 37204 24952 37256
rect 25004 37244 25010 37256
rect 25133 37247 25191 37253
rect 25133 37244 25145 37247
rect 25004 37216 25145 37244
rect 25004 37204 25010 37216
rect 25133 37213 25145 37216
rect 25179 37213 25191 37247
rect 26237 37247 26295 37253
rect 26237 37244 26249 37247
rect 25133 37207 25191 37213
rect 25240 37216 26249 37244
rect 15746 37176 15752 37188
rect 14200 37148 15752 37176
rect 15746 37136 15752 37148
rect 15804 37136 15810 37188
rect 15930 37136 15936 37188
rect 15988 37136 15994 37188
rect 17310 37136 17316 37188
rect 17368 37136 17374 37188
rect 18782 37136 18788 37188
rect 18840 37136 18846 37188
rect 20714 37136 20720 37188
rect 20772 37136 20778 37188
rect 22462 37176 22468 37188
rect 21100 37148 22468 37176
rect 9493 37111 9551 37117
rect 9493 37077 9505 37111
rect 9539 37077 9551 37111
rect 9493 37071 9551 37077
rect 9582 37068 9588 37120
rect 9640 37068 9646 37120
rect 11790 37068 11796 37120
rect 11848 37068 11854 37120
rect 12253 37111 12311 37117
rect 12253 37077 12265 37111
rect 12299 37108 12311 37111
rect 12710 37108 12716 37120
rect 12299 37080 12716 37108
rect 12299 37077 12311 37080
rect 12253 37071 12311 37077
rect 12710 37068 12716 37080
rect 12768 37068 12774 37120
rect 12989 37111 13047 37117
rect 12989 37077 13001 37111
rect 13035 37108 13047 37111
rect 13078 37108 13084 37120
rect 13035 37080 13084 37108
rect 13035 37077 13047 37080
rect 12989 37071 13047 37077
rect 13078 37068 13084 37080
rect 13136 37068 13142 37120
rect 13354 37068 13360 37120
rect 13412 37068 13418 37120
rect 13449 37111 13507 37117
rect 13449 37077 13461 37111
rect 13495 37108 13507 37111
rect 14274 37108 14280 37120
rect 13495 37080 14280 37108
rect 13495 37077 13507 37080
rect 13449 37071 13507 37077
rect 14274 37068 14280 37080
rect 14332 37068 14338 37120
rect 14550 37068 14556 37120
rect 14608 37068 14614 37120
rect 15010 37068 15016 37120
rect 15068 37108 15074 37120
rect 21100 37108 21128 37148
rect 22462 37136 22468 37148
rect 22520 37136 22526 37188
rect 22646 37136 22652 37188
rect 22704 37176 22710 37188
rect 22704 37148 23796 37176
rect 22704 37136 22710 37148
rect 15068 37080 21128 37108
rect 21177 37111 21235 37117
rect 15068 37068 15074 37080
rect 21177 37077 21189 37111
rect 21223 37108 21235 37111
rect 23474 37108 23480 37120
rect 21223 37080 23480 37108
rect 21223 37077 21235 37080
rect 21177 37071 21235 37077
rect 23474 37068 23480 37080
rect 23532 37068 23538 37120
rect 23768 37108 23796 37148
rect 23842 37136 23848 37188
rect 23900 37136 23906 37188
rect 24118 37136 24124 37188
rect 24176 37176 24182 37188
rect 25240 37176 25268 37216
rect 26237 37213 26249 37216
rect 26283 37213 26295 37247
rect 26237 37207 26295 37213
rect 26421 37247 26479 37253
rect 26421 37213 26433 37247
rect 26467 37244 26479 37247
rect 26602 37244 26608 37256
rect 26467 37216 26608 37244
rect 26467 37213 26479 37216
rect 26421 37207 26479 37213
rect 26602 37204 26608 37216
rect 26660 37204 26666 37256
rect 27157 37247 27215 37253
rect 27157 37213 27169 37247
rect 27203 37244 27215 37247
rect 27246 37244 27252 37256
rect 27203 37216 27252 37244
rect 27203 37213 27215 37216
rect 27157 37207 27215 37213
rect 27246 37204 27252 37216
rect 27304 37204 27310 37256
rect 28184 37253 28212 37284
rect 32398 37272 32404 37324
rect 32456 37272 32462 37324
rect 33686 37272 33692 37324
rect 33744 37272 33750 37324
rect 28169 37247 28227 37253
rect 28169 37213 28181 37247
rect 28215 37213 28227 37247
rect 28169 37207 28227 37213
rect 28258 37204 28264 37256
rect 28316 37244 28322 37256
rect 28997 37247 29055 37253
rect 28997 37244 29009 37247
rect 28316 37216 29009 37244
rect 28316 37204 28322 37216
rect 28997 37213 29009 37216
rect 29043 37213 29055 37247
rect 28997 37207 29055 37213
rect 29178 37204 29184 37256
rect 29236 37204 29242 37256
rect 30282 37204 30288 37256
rect 30340 37204 30346 37256
rect 30552 37247 30610 37253
rect 30552 37213 30564 37247
rect 30598 37244 30610 37247
rect 32030 37244 32036 37256
rect 30598 37216 32036 37244
rect 30598 37213 30610 37216
rect 30552 37207 30610 37213
rect 32030 37204 32036 37216
rect 32088 37204 32094 37256
rect 32306 37204 32312 37256
rect 32364 37253 32370 37256
rect 32364 37244 32374 37253
rect 32364 37216 32409 37244
rect 32364 37207 32374 37216
rect 32364 37204 32370 37207
rect 32582 37204 32588 37256
rect 32640 37204 32646 37256
rect 33134 37204 33140 37256
rect 33192 37244 33198 37256
rect 33413 37247 33471 37253
rect 33413 37244 33425 37247
rect 33192 37216 33425 37244
rect 33192 37204 33198 37216
rect 33413 37213 33425 37216
rect 33459 37213 33471 37247
rect 33413 37207 33471 37213
rect 33597 37247 33655 37253
rect 33597 37213 33609 37247
rect 33643 37213 33655 37247
rect 33597 37207 33655 37213
rect 24176 37148 25268 37176
rect 24176 37136 24182 37148
rect 25314 37136 25320 37188
rect 25372 37176 25378 37188
rect 25501 37179 25559 37185
rect 25501 37176 25513 37179
rect 25372 37148 25513 37176
rect 25372 37136 25378 37148
rect 25501 37145 25513 37148
rect 25547 37145 25559 37179
rect 25501 37139 25559 37145
rect 27433 37179 27491 37185
rect 27433 37145 27445 37179
rect 27479 37176 27491 37179
rect 29454 37176 29460 37188
rect 27479 37148 29460 37176
rect 27479 37145 27491 37148
rect 27433 37139 27491 37145
rect 29454 37136 29460 37148
rect 29512 37136 29518 37188
rect 31110 37136 31116 37188
rect 31168 37176 31174 37188
rect 33612 37176 33640 37207
rect 33778 37204 33784 37256
rect 33836 37244 33842 37256
rect 34149 37247 34207 37253
rect 34149 37244 34161 37247
rect 33836 37216 34161 37244
rect 33836 37204 33842 37216
rect 34149 37213 34161 37216
rect 34195 37213 34207 37247
rect 34149 37207 34207 37213
rect 34238 37204 34244 37256
rect 34296 37204 34302 37256
rect 35158 37204 35164 37256
rect 35216 37244 35222 37256
rect 35437 37247 35495 37253
rect 35437 37244 35449 37247
rect 35216 37216 35449 37244
rect 35216 37204 35222 37216
rect 35437 37213 35449 37216
rect 35483 37244 35495 37247
rect 35526 37244 35532 37256
rect 35483 37216 35532 37244
rect 35483 37213 35495 37216
rect 35437 37207 35495 37213
rect 35526 37204 35532 37216
rect 35584 37204 35590 37256
rect 37645 37247 37703 37253
rect 37645 37213 37657 37247
rect 37691 37244 37703 37247
rect 38102 37244 38108 37256
rect 37691 37216 38108 37244
rect 37691 37213 37703 37216
rect 37645 37207 37703 37213
rect 38102 37204 38108 37216
rect 38160 37204 38166 37256
rect 35704 37179 35762 37185
rect 31168 37148 34376 37176
rect 31168 37136 31174 37148
rect 26234 37108 26240 37120
rect 23768 37080 26240 37108
rect 26234 37068 26240 37080
rect 26292 37068 26298 37120
rect 26510 37068 26516 37120
rect 26568 37108 26574 37120
rect 26605 37111 26663 37117
rect 26605 37108 26617 37111
rect 26568 37080 26617 37108
rect 26568 37068 26574 37080
rect 26605 37077 26617 37080
rect 26651 37077 26663 37111
rect 26605 37071 26663 37077
rect 26878 37068 26884 37120
rect 26936 37108 26942 37120
rect 28261 37111 28319 37117
rect 28261 37108 28273 37111
rect 26936 37080 28273 37108
rect 26936 37068 26942 37080
rect 28261 37077 28273 37080
rect 28307 37108 28319 37111
rect 28350 37108 28356 37120
rect 28307 37080 28356 37108
rect 28307 37077 28319 37080
rect 28261 37071 28319 37077
rect 28350 37068 28356 37080
rect 28408 37068 28414 37120
rect 29086 37068 29092 37120
rect 29144 37068 29150 37120
rect 31680 37117 31708 37148
rect 31665 37111 31723 37117
rect 31665 37077 31677 37111
rect 31711 37108 31723 37111
rect 31711 37080 31745 37108
rect 31711 37077 31723 37080
rect 31665 37071 31723 37077
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32769 37111 32827 37117
rect 32769 37108 32781 37111
rect 32272 37080 32781 37108
rect 32272 37068 32278 37080
rect 32769 37077 32781 37080
rect 32815 37077 32827 37111
rect 34348 37108 34376 37148
rect 35704 37145 35716 37179
rect 35750 37176 35762 37179
rect 37550 37176 37556 37188
rect 35750 37148 37556 37176
rect 35750 37145 35762 37148
rect 35704 37139 35762 37145
rect 37550 37136 37556 37148
rect 37608 37136 37614 37188
rect 38010 37136 38016 37188
rect 38068 37136 38074 37188
rect 35802 37108 35808 37120
rect 34348 37080 35808 37108
rect 32769 37071 32827 37077
rect 35802 37068 35808 37080
rect 35860 37068 35866 37120
rect 36817 37111 36875 37117
rect 36817 37077 36829 37111
rect 36863 37108 36875 37111
rect 37366 37108 37372 37120
rect 36863 37080 37372 37108
rect 36863 37077 36875 37080
rect 36817 37071 36875 37077
rect 37366 37068 37372 37080
rect 37424 37068 37430 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 3050 36864 3056 36916
rect 3108 36864 3114 36916
rect 3694 36864 3700 36916
rect 3752 36864 3758 36916
rect 4433 36907 4491 36913
rect 4433 36873 4445 36907
rect 4479 36904 4491 36907
rect 4798 36904 4804 36916
rect 4479 36876 4804 36904
rect 4479 36873 4491 36876
rect 4433 36867 4491 36873
rect 4798 36864 4804 36876
rect 4856 36864 4862 36916
rect 5077 36907 5135 36913
rect 5077 36873 5089 36907
rect 5123 36904 5135 36907
rect 5442 36904 5448 36916
rect 5123 36876 5448 36904
rect 5123 36873 5135 36876
rect 5077 36867 5135 36873
rect 5442 36864 5448 36876
rect 5500 36864 5506 36916
rect 5994 36864 6000 36916
rect 6052 36864 6058 36916
rect 9309 36907 9367 36913
rect 9309 36873 9321 36907
rect 9355 36904 9367 36907
rect 9582 36904 9588 36916
rect 9355 36876 9588 36904
rect 9355 36873 9367 36876
rect 9309 36867 9367 36873
rect 9582 36864 9588 36876
rect 9640 36864 9646 36916
rect 12434 36904 12440 36916
rect 12176 36876 12440 36904
rect 4264 36808 4936 36836
rect 1670 36728 1676 36780
rect 1728 36728 1734 36780
rect 4264 36777 4292 36808
rect 2317 36771 2375 36777
rect 2317 36737 2329 36771
rect 2363 36768 2375 36771
rect 2961 36771 3019 36777
rect 2961 36768 2973 36771
rect 2363 36740 2973 36768
rect 2363 36737 2375 36740
rect 2317 36731 2375 36737
rect 2961 36737 2973 36740
rect 3007 36768 3019 36771
rect 3605 36771 3663 36777
rect 3605 36768 3617 36771
rect 3007 36740 3617 36768
rect 3007 36737 3019 36740
rect 2961 36731 3019 36737
rect 3605 36737 3617 36740
rect 3651 36737 3663 36771
rect 3605 36731 3663 36737
rect 4249 36771 4307 36777
rect 4249 36737 4261 36771
rect 4295 36737 4307 36771
rect 4249 36731 4307 36737
rect 4433 36771 4491 36777
rect 4433 36737 4445 36771
rect 4479 36737 4491 36771
rect 4908 36768 4936 36808
rect 4982 36796 4988 36848
rect 5040 36796 5046 36848
rect 5350 36796 5356 36848
rect 5408 36836 5414 36848
rect 7285 36839 7343 36845
rect 7285 36836 7297 36839
rect 5408 36808 7297 36836
rect 5408 36796 5414 36808
rect 7285 36805 7297 36808
rect 7331 36805 7343 36839
rect 11698 36836 11704 36848
rect 7285 36799 7343 36805
rect 7944 36808 11704 36836
rect 5626 36768 5632 36780
rect 4908 36740 5632 36768
rect 4433 36731 4491 36737
rect 1762 36524 1768 36576
rect 1820 36524 1826 36576
rect 2406 36524 2412 36576
rect 2464 36524 2470 36576
rect 3234 36524 3240 36576
rect 3292 36564 3298 36576
rect 3620 36564 3648 36731
rect 4448 36700 4476 36731
rect 5626 36728 5632 36740
rect 5684 36728 5690 36780
rect 5718 36728 5724 36780
rect 5776 36728 5782 36780
rect 5813 36771 5871 36777
rect 5813 36737 5825 36771
rect 5859 36737 5871 36771
rect 5813 36731 5871 36737
rect 5828 36700 5856 36731
rect 7006 36728 7012 36780
rect 7064 36768 7070 36780
rect 7101 36771 7159 36777
rect 7101 36768 7113 36771
rect 7064 36740 7113 36768
rect 7064 36728 7070 36740
rect 7101 36737 7113 36740
rect 7147 36737 7159 36771
rect 7101 36731 7159 36737
rect 7469 36703 7527 36709
rect 7469 36700 7481 36703
rect 4448 36672 5764 36700
rect 5828 36672 7481 36700
rect 4522 36592 4528 36644
rect 4580 36632 4586 36644
rect 4982 36632 4988 36644
rect 4580 36604 4988 36632
rect 4580 36592 4586 36604
rect 4982 36592 4988 36604
rect 5040 36592 5046 36644
rect 5736 36632 5764 36672
rect 7469 36669 7481 36672
rect 7515 36669 7527 36703
rect 7469 36663 7527 36669
rect 7650 36660 7656 36712
rect 7708 36700 7714 36712
rect 7944 36709 7972 36808
rect 8196 36771 8254 36777
rect 8196 36737 8208 36771
rect 8242 36768 8254 36771
rect 9122 36768 9128 36780
rect 8242 36740 9128 36768
rect 8242 36737 8254 36740
rect 8196 36731 8254 36737
rect 9122 36728 9128 36740
rect 9180 36728 9186 36780
rect 9784 36777 9812 36808
rect 11698 36796 11704 36808
rect 11756 36796 11762 36848
rect 9769 36771 9827 36777
rect 9769 36737 9781 36771
rect 9815 36737 9827 36771
rect 9769 36731 9827 36737
rect 10036 36771 10094 36777
rect 10036 36737 10048 36771
rect 10082 36768 10094 36771
rect 10502 36768 10508 36780
rect 10082 36740 10508 36768
rect 10082 36737 10094 36740
rect 10036 36731 10094 36737
rect 10502 36728 10508 36740
rect 10560 36728 10566 36780
rect 12176 36777 12204 36876
rect 12434 36864 12440 36876
rect 12492 36904 12498 36916
rect 13538 36904 13544 36916
rect 12492 36876 13544 36904
rect 12492 36864 12498 36876
rect 13538 36864 13544 36876
rect 13596 36864 13602 36916
rect 14274 36864 14280 36916
rect 14332 36904 14338 36916
rect 14369 36907 14427 36913
rect 14369 36904 14381 36907
rect 14332 36876 14381 36904
rect 14332 36864 14338 36876
rect 14369 36873 14381 36876
rect 14415 36873 14427 36907
rect 14369 36867 14427 36873
rect 15746 36864 15752 36916
rect 15804 36904 15810 36916
rect 23842 36904 23848 36916
rect 15804 36876 23848 36904
rect 15804 36864 15810 36876
rect 23842 36864 23848 36876
rect 23900 36864 23906 36916
rect 31846 36904 31852 36916
rect 24780 36876 31852 36904
rect 12345 36839 12403 36845
rect 12345 36805 12357 36839
rect 12391 36836 12403 36839
rect 12710 36836 12716 36848
rect 12391 36808 12716 36836
rect 12391 36805 12403 36808
rect 12345 36799 12403 36805
rect 12710 36796 12716 36808
rect 12768 36796 12774 36848
rect 18506 36836 18512 36848
rect 13004 36808 14872 36836
rect 13004 36777 13032 36808
rect 12161 36771 12219 36777
rect 12161 36737 12173 36771
rect 12207 36737 12219 36771
rect 12989 36771 13047 36777
rect 12989 36768 13001 36771
rect 12161 36731 12219 36737
rect 12268 36740 13001 36768
rect 7929 36703 7987 36709
rect 7929 36700 7941 36703
rect 7708 36672 7941 36700
rect 7708 36660 7714 36672
rect 7929 36669 7941 36672
rect 7975 36669 7987 36703
rect 7929 36663 7987 36669
rect 11698 36660 11704 36712
rect 11756 36700 11762 36712
rect 12268 36700 12296 36740
rect 12989 36737 13001 36740
rect 13035 36737 13047 36771
rect 12989 36731 13047 36737
rect 13078 36728 13084 36780
rect 13136 36768 13142 36780
rect 14844 36777 14872 36808
rect 17144 36808 18512 36836
rect 17144 36780 17172 36808
rect 18506 36796 18512 36808
rect 18564 36796 18570 36848
rect 18598 36796 18604 36848
rect 18656 36836 18662 36848
rect 18656 36808 20470 36836
rect 18656 36796 18662 36808
rect 22554 36796 22560 36848
rect 22612 36796 22618 36848
rect 24302 36796 24308 36848
rect 24360 36796 24366 36848
rect 13245 36771 13303 36777
rect 13245 36768 13257 36771
rect 13136 36740 13257 36768
rect 13136 36728 13142 36740
rect 13245 36737 13257 36740
rect 13291 36737 13303 36771
rect 13245 36731 13303 36737
rect 14829 36771 14887 36777
rect 14829 36737 14841 36771
rect 14875 36737 14887 36771
rect 14829 36731 14887 36737
rect 14918 36728 14924 36780
rect 14976 36768 14982 36780
rect 15085 36771 15143 36777
rect 15085 36768 15097 36771
rect 14976 36740 15097 36768
rect 14976 36728 14982 36740
rect 15085 36737 15097 36740
rect 15131 36737 15143 36771
rect 15085 36731 15143 36737
rect 17126 36728 17132 36780
rect 17184 36728 17190 36780
rect 17396 36771 17454 36777
rect 17396 36737 17408 36771
rect 17442 36768 17454 36771
rect 18414 36768 18420 36780
rect 17442 36740 18420 36768
rect 17442 36737 17454 36740
rect 17396 36731 17454 36737
rect 18414 36728 18420 36740
rect 18472 36728 18478 36780
rect 18874 36728 18880 36780
rect 18932 36768 18938 36780
rect 18969 36771 19027 36777
rect 18969 36768 18981 36771
rect 18932 36740 18981 36768
rect 18932 36728 18938 36740
rect 18969 36737 18981 36740
rect 19015 36737 19027 36771
rect 18969 36731 19027 36737
rect 19150 36728 19156 36780
rect 19208 36728 19214 36780
rect 19245 36771 19303 36777
rect 19245 36737 19257 36771
rect 19291 36737 19303 36771
rect 19245 36731 19303 36737
rect 11756 36672 12296 36700
rect 11756 36660 11762 36672
rect 12434 36660 12440 36712
rect 12492 36660 12498 36712
rect 7834 36632 7840 36644
rect 5736 36604 7840 36632
rect 7834 36592 7840 36604
rect 7892 36592 7898 36644
rect 9214 36592 9220 36644
rect 9272 36632 9278 36644
rect 9766 36632 9772 36644
rect 9272 36604 9772 36632
rect 9272 36592 9278 36604
rect 9766 36592 9772 36604
rect 9824 36592 9830 36644
rect 10704 36604 12434 36632
rect 5442 36564 5448 36576
rect 3292 36536 5448 36564
rect 3292 36524 3298 36536
rect 5442 36524 5448 36536
rect 5500 36524 5506 36576
rect 7466 36524 7472 36576
rect 7524 36564 7530 36576
rect 10704 36564 10732 36604
rect 7524 36536 10732 36564
rect 7524 36524 7530 36536
rect 11146 36524 11152 36576
rect 11204 36524 11210 36576
rect 11885 36567 11943 36573
rect 11885 36533 11897 36567
rect 11931 36564 11943 36567
rect 11974 36564 11980 36576
rect 11931 36536 11980 36564
rect 11931 36533 11943 36536
rect 11885 36527 11943 36533
rect 11974 36524 11980 36536
rect 12032 36524 12038 36576
rect 12406 36564 12434 36604
rect 15838 36592 15844 36644
rect 15896 36632 15902 36644
rect 19260 36632 19288 36731
rect 23658 36728 23664 36780
rect 23716 36728 23722 36780
rect 19705 36703 19763 36709
rect 19705 36669 19717 36703
rect 19751 36669 19763 36703
rect 19705 36663 19763 36669
rect 15896 36604 16344 36632
rect 15896 36592 15902 36604
rect 15010 36564 15016 36576
rect 12406 36536 15016 36564
rect 15010 36524 15016 36536
rect 15068 36524 15074 36576
rect 15194 36524 15200 36576
rect 15252 36564 15258 36576
rect 16209 36567 16267 36573
rect 16209 36564 16221 36567
rect 15252 36536 16221 36564
rect 15252 36524 15258 36536
rect 16209 36533 16221 36536
rect 16255 36533 16267 36567
rect 16316 36564 16344 36604
rect 18064 36604 19288 36632
rect 17402 36564 17408 36576
rect 16316 36536 17408 36564
rect 16209 36527 16267 36533
rect 17402 36524 17408 36536
rect 17460 36524 17466 36576
rect 17770 36524 17776 36576
rect 17828 36564 17834 36576
rect 18064 36564 18092 36604
rect 17828 36536 18092 36564
rect 18509 36567 18567 36573
rect 17828 36524 17834 36536
rect 18509 36533 18521 36567
rect 18555 36564 18567 36567
rect 18598 36564 18604 36576
rect 18555 36536 18604 36564
rect 18555 36533 18567 36536
rect 18509 36527 18567 36533
rect 18598 36524 18604 36536
rect 18656 36524 18662 36576
rect 18966 36524 18972 36576
rect 19024 36524 19030 36576
rect 19242 36524 19248 36576
rect 19300 36564 19306 36576
rect 19720 36564 19748 36663
rect 19978 36660 19984 36712
rect 20036 36660 20042 36712
rect 21542 36660 21548 36712
rect 21600 36700 21606 36712
rect 22281 36703 22339 36709
rect 22281 36700 22293 36703
rect 21600 36672 22293 36700
rect 21600 36660 21606 36672
rect 22281 36669 22293 36672
rect 22327 36669 22339 36703
rect 22281 36663 22339 36669
rect 22554 36660 22560 36712
rect 22612 36700 22618 36712
rect 24320 36700 24348 36796
rect 24780 36777 24808 36876
rect 25498 36796 25504 36848
rect 25556 36796 25562 36848
rect 27706 36836 27712 36848
rect 26436 36808 27712 36836
rect 24765 36771 24823 36777
rect 24765 36737 24777 36771
rect 24811 36737 24823 36771
rect 26436 36768 26464 36808
rect 27706 36796 27712 36808
rect 27764 36796 27770 36848
rect 27341 36771 27399 36777
rect 27341 36768 27353 36771
rect 24765 36731 24823 36737
rect 26252 36740 26464 36768
rect 26528 36740 27353 36768
rect 26252 36712 26280 36740
rect 22612 36672 24348 36700
rect 22612 36660 22618 36672
rect 24394 36660 24400 36712
rect 24452 36700 24458 36712
rect 25041 36703 25099 36709
rect 25041 36700 25053 36703
rect 24452 36672 25053 36700
rect 24452 36660 24458 36672
rect 25041 36669 25053 36672
rect 25087 36669 25099 36703
rect 25041 36663 25099 36669
rect 26234 36660 26240 36712
rect 26292 36660 26298 36712
rect 26528 36709 26556 36740
rect 27341 36737 27353 36740
rect 27387 36768 27399 36771
rect 28074 36768 28080 36780
rect 27387 36740 28080 36768
rect 27387 36737 27399 36740
rect 27341 36731 27399 36737
rect 28074 36728 28080 36740
rect 28132 36728 28138 36780
rect 28460 36777 28488 36876
rect 31846 36864 31852 36876
rect 31904 36904 31910 36916
rect 31904 36876 32352 36904
rect 31904 36864 31910 36876
rect 28718 36796 28724 36848
rect 28776 36796 28782 36848
rect 28994 36796 29000 36848
rect 29052 36836 29058 36848
rect 29052 36808 29210 36836
rect 29052 36796 29058 36808
rect 28445 36771 28503 36777
rect 28445 36737 28457 36771
rect 28491 36737 28503 36771
rect 28445 36731 28503 36737
rect 31113 36771 31171 36777
rect 31113 36737 31125 36771
rect 31159 36768 31171 36771
rect 32214 36768 32220 36780
rect 31159 36740 32220 36768
rect 31159 36737 31171 36740
rect 31113 36731 31171 36737
rect 32214 36728 32220 36740
rect 32272 36728 32278 36780
rect 32324 36777 32352 36876
rect 32416 36876 37964 36904
rect 32309 36771 32367 36777
rect 32309 36737 32321 36771
rect 32355 36737 32367 36771
rect 32309 36731 32367 36737
rect 26513 36703 26571 36709
rect 26513 36669 26525 36703
rect 26559 36669 26571 36703
rect 26513 36663 26571 36669
rect 27614 36660 27620 36712
rect 27672 36700 27678 36712
rect 30193 36703 30251 36709
rect 30193 36700 30205 36703
rect 27672 36672 30205 36700
rect 27672 36660 27678 36672
rect 30193 36669 30205 36672
rect 30239 36700 30251 36703
rect 31294 36700 31300 36712
rect 30239 36672 31300 36700
rect 30239 36669 30251 36672
rect 30193 36663 30251 36669
rect 31294 36660 31300 36672
rect 31352 36660 31358 36712
rect 31573 36703 31631 36709
rect 31573 36669 31585 36703
rect 31619 36700 31631 36703
rect 31662 36700 31668 36712
rect 31619 36672 31668 36700
rect 31619 36669 31631 36672
rect 31573 36663 31631 36669
rect 26142 36592 26148 36644
rect 26200 36632 26206 36644
rect 26602 36632 26608 36644
rect 26200 36604 26608 36632
rect 26200 36592 26206 36604
rect 26602 36592 26608 36604
rect 26660 36592 26666 36644
rect 31588 36632 31616 36663
rect 31662 36660 31668 36672
rect 31720 36700 31726 36712
rect 32416 36700 32444 36876
rect 35710 36845 35716 36848
rect 35704 36799 35716 36845
rect 35710 36796 35716 36799
rect 35768 36796 35774 36848
rect 35802 36796 35808 36848
rect 35860 36836 35866 36848
rect 37829 36839 37887 36845
rect 37829 36836 37841 36839
rect 35860 36808 37841 36836
rect 35860 36796 35866 36808
rect 37829 36805 37841 36808
rect 37875 36805 37887 36839
rect 37829 36799 37887 36805
rect 32576 36771 32634 36777
rect 32576 36737 32588 36771
rect 32622 36768 32634 36771
rect 33042 36768 33048 36780
rect 32622 36740 33048 36768
rect 32622 36737 32634 36740
rect 32576 36731 32634 36737
rect 33042 36728 33048 36740
rect 33100 36768 33106 36780
rect 33965 36771 34023 36777
rect 33965 36768 33977 36771
rect 33100 36740 33977 36768
rect 33100 36728 33106 36740
rect 33965 36737 33977 36740
rect 34011 36737 34023 36771
rect 33965 36731 34023 36737
rect 34514 36728 34520 36780
rect 34572 36728 34578 36780
rect 36078 36728 36084 36780
rect 36136 36768 36142 36780
rect 37936 36777 37964 36876
rect 37461 36771 37519 36777
rect 37461 36768 37473 36771
rect 36136 36740 37473 36768
rect 36136 36728 36142 36740
rect 37461 36737 37473 36740
rect 37507 36737 37519 36771
rect 37461 36731 37519 36737
rect 37645 36771 37703 36777
rect 37645 36737 37657 36771
rect 37691 36737 37703 36771
rect 37645 36731 37703 36737
rect 37921 36771 37979 36777
rect 37921 36737 37933 36771
rect 37967 36737 37979 36771
rect 37921 36731 37979 36737
rect 31720 36672 32444 36700
rect 31720 36660 31726 36672
rect 34606 36660 34612 36712
rect 34664 36660 34670 36712
rect 35437 36703 35495 36709
rect 35437 36669 35449 36703
rect 35483 36669 35495 36703
rect 37660 36700 37688 36731
rect 38010 36700 38016 36712
rect 37660 36672 38016 36700
rect 35437 36663 35495 36669
rect 29748 36604 31616 36632
rect 19300 36536 19748 36564
rect 19300 36524 19306 36536
rect 21450 36524 21456 36576
rect 21508 36524 21514 36576
rect 23658 36524 23664 36576
rect 23716 36564 23722 36576
rect 29086 36564 29092 36576
rect 23716 36536 29092 36564
rect 23716 36524 23722 36536
rect 29086 36524 29092 36536
rect 29144 36524 29150 36576
rect 29362 36524 29368 36576
rect 29420 36564 29426 36576
rect 29748 36564 29776 36604
rect 34146 36592 34152 36644
rect 34204 36632 34210 36644
rect 35452 36632 35480 36663
rect 38010 36660 38016 36672
rect 38068 36660 38074 36712
rect 34204 36604 35480 36632
rect 34204 36592 34210 36604
rect 29420 36536 29776 36564
rect 29420 36524 29426 36536
rect 29914 36524 29920 36576
rect 29972 36564 29978 36576
rect 32582 36564 32588 36576
rect 29972 36536 32588 36564
rect 29972 36524 29978 36536
rect 32582 36524 32588 36536
rect 32640 36524 32646 36576
rect 33226 36524 33232 36576
rect 33284 36564 33290 36576
rect 33689 36567 33747 36573
rect 33689 36564 33701 36567
rect 33284 36536 33701 36564
rect 33284 36524 33290 36536
rect 33689 36533 33701 36536
rect 33735 36533 33747 36567
rect 33689 36527 33747 36533
rect 34793 36567 34851 36573
rect 34793 36533 34805 36567
rect 34839 36564 34851 36567
rect 36170 36564 36176 36576
rect 34839 36536 36176 36564
rect 34839 36533 34851 36536
rect 34793 36527 34851 36533
rect 36170 36524 36176 36536
rect 36228 36524 36234 36576
rect 36446 36524 36452 36576
rect 36504 36564 36510 36576
rect 36817 36567 36875 36573
rect 36817 36564 36829 36567
rect 36504 36536 36829 36564
rect 36504 36524 36510 36536
rect 36817 36533 36829 36536
rect 36863 36533 36875 36567
rect 36817 36527 36875 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 2590 36320 2596 36372
rect 2648 36320 2654 36372
rect 3326 36320 3332 36372
rect 3384 36320 3390 36372
rect 5258 36320 5264 36372
rect 5316 36320 5322 36372
rect 6730 36320 6736 36372
rect 6788 36320 6794 36372
rect 7742 36320 7748 36372
rect 7800 36320 7806 36372
rect 7834 36320 7840 36372
rect 7892 36360 7898 36372
rect 9858 36360 9864 36372
rect 7892 36332 9864 36360
rect 7892 36320 7898 36332
rect 9858 36320 9864 36332
rect 9916 36320 9922 36372
rect 10502 36320 10508 36372
rect 10560 36320 10566 36372
rect 23339 36363 23397 36369
rect 10612 36332 23244 36360
rect 7190 36292 7196 36304
rect 2608 36264 7196 36292
rect 2608 36165 2636 36264
rect 7190 36252 7196 36264
rect 7248 36252 7254 36304
rect 8570 36252 8576 36304
rect 8628 36252 8634 36304
rect 9309 36295 9367 36301
rect 9309 36261 9321 36295
rect 9355 36292 9367 36295
rect 10410 36292 10416 36304
rect 9355 36264 10416 36292
rect 9355 36261 9367 36264
rect 9309 36255 9367 36261
rect 10410 36252 10416 36264
rect 10468 36252 10474 36304
rect 9214 36224 9220 36236
rect 2792 36196 6684 36224
rect 2792 36165 2820 36196
rect 2593 36159 2651 36165
rect 2593 36125 2605 36159
rect 2639 36125 2651 36159
rect 2593 36119 2651 36125
rect 2777 36159 2835 36165
rect 2777 36125 2789 36159
rect 2823 36125 2835 36159
rect 2777 36119 2835 36125
rect 3234 36116 3240 36168
rect 3292 36116 3298 36168
rect 4341 36159 4399 36165
rect 4341 36125 4353 36159
rect 4387 36156 4399 36159
rect 5074 36156 5080 36168
rect 4387 36128 5080 36156
rect 4387 36125 4399 36128
rect 4341 36119 4399 36125
rect 5074 36116 5080 36128
rect 5132 36116 5138 36168
rect 5169 36159 5227 36165
rect 5169 36125 5181 36159
rect 5215 36156 5227 36159
rect 5442 36156 5448 36168
rect 5215 36128 5448 36156
rect 5215 36125 5227 36128
rect 5169 36119 5227 36125
rect 5442 36116 5448 36128
rect 5500 36116 5506 36168
rect 5902 36116 5908 36168
rect 5960 36116 5966 36168
rect 6656 36165 6684 36196
rect 7576 36196 9220 36224
rect 6549 36159 6607 36165
rect 6549 36125 6561 36159
rect 6595 36125 6607 36159
rect 6549 36119 6607 36125
rect 6642 36159 6700 36165
rect 6642 36125 6654 36159
rect 6688 36156 6700 36159
rect 6688 36128 7420 36156
rect 6688 36125 6700 36128
rect 6642 36119 6700 36125
rect 4433 36091 4491 36097
rect 4433 36057 4445 36091
rect 4479 36088 4491 36091
rect 5810 36088 5816 36100
rect 4479 36060 5816 36088
rect 4479 36057 4491 36060
rect 4433 36051 4491 36057
rect 5810 36048 5816 36060
rect 5868 36048 5874 36100
rect 6086 36048 6092 36100
rect 6144 36048 6150 36100
rect 6564 36088 6592 36119
rect 7190 36088 7196 36100
rect 6564 36060 7196 36088
rect 7190 36048 7196 36060
rect 7248 36048 7254 36100
rect 7392 36088 7420 36128
rect 7466 36116 7472 36168
rect 7524 36116 7530 36168
rect 7576 36165 7604 36196
rect 9214 36184 9220 36196
rect 9272 36184 9278 36236
rect 9582 36184 9588 36236
rect 9640 36224 9646 36236
rect 9769 36227 9827 36233
rect 9769 36224 9781 36227
rect 9640 36196 9781 36224
rect 9640 36184 9646 36196
rect 9769 36193 9781 36196
rect 9815 36193 9827 36227
rect 9769 36187 9827 36193
rect 9858 36184 9864 36236
rect 9916 36184 9922 36236
rect 7561 36159 7619 36165
rect 7561 36125 7573 36159
rect 7607 36125 7619 36159
rect 10612 36156 10640 36332
rect 12710 36252 12716 36304
rect 12768 36292 12774 36304
rect 13081 36295 13139 36301
rect 13081 36292 13093 36295
rect 12768 36264 13093 36292
rect 12768 36252 12774 36264
rect 13081 36261 13093 36264
rect 13127 36261 13139 36295
rect 13081 36255 13139 36261
rect 14737 36295 14795 36301
rect 14737 36261 14749 36295
rect 14783 36292 14795 36295
rect 14918 36292 14924 36304
rect 14783 36264 14924 36292
rect 14783 36261 14795 36264
rect 14737 36255 14795 36261
rect 14918 36252 14924 36264
rect 14976 36252 14982 36304
rect 15838 36292 15844 36304
rect 15120 36264 15844 36292
rect 10962 36184 10968 36236
rect 11020 36224 11026 36236
rect 11057 36227 11115 36233
rect 11057 36224 11069 36227
rect 11020 36196 11069 36224
rect 11020 36184 11026 36196
rect 11057 36193 11069 36196
rect 11103 36193 11115 36227
rect 11057 36187 11115 36193
rect 11698 36184 11704 36236
rect 11756 36184 11762 36236
rect 15120 36224 15148 36264
rect 15838 36252 15844 36264
rect 15896 36252 15902 36304
rect 18414 36252 18420 36304
rect 18472 36292 18478 36304
rect 19429 36295 19487 36301
rect 19429 36292 19441 36295
rect 18472 36264 19441 36292
rect 18472 36252 18478 36264
rect 19429 36261 19441 36264
rect 19475 36261 19487 36295
rect 20438 36292 20444 36304
rect 19429 36255 19487 36261
rect 19996 36264 20444 36292
rect 13740 36196 15148 36224
rect 7561 36119 7619 36125
rect 7659 36128 10640 36156
rect 7659 36088 7687 36128
rect 11790 36116 11796 36168
rect 11848 36156 11854 36168
rect 13740 36165 13768 36196
rect 15194 36184 15200 36236
rect 15252 36184 15258 36236
rect 15289 36227 15347 36233
rect 15289 36193 15301 36227
rect 15335 36193 15347 36227
rect 18598 36224 18604 36236
rect 15289 36187 15347 36193
rect 18248 36196 18604 36224
rect 11957 36159 12015 36165
rect 11957 36156 11969 36159
rect 11848 36128 11969 36156
rect 11848 36116 11854 36128
rect 11957 36125 11969 36128
rect 12003 36125 12015 36159
rect 11957 36119 12015 36125
rect 13541 36159 13599 36165
rect 13541 36125 13553 36159
rect 13587 36125 13599 36159
rect 13541 36119 13599 36125
rect 13725 36159 13783 36165
rect 13725 36125 13737 36159
rect 13771 36125 13783 36159
rect 13725 36119 13783 36125
rect 7392 36060 7687 36088
rect 8110 36048 8116 36100
rect 8168 36088 8174 36100
rect 8205 36091 8263 36097
rect 8205 36088 8217 36091
rect 8168 36060 8217 36088
rect 8168 36048 8174 36060
rect 8205 36057 8217 36060
rect 8251 36057 8263 36091
rect 8205 36051 8263 36057
rect 8294 36048 8300 36100
rect 8352 36088 8358 36100
rect 8389 36091 8447 36097
rect 8389 36088 8401 36091
rect 8352 36060 8401 36088
rect 8352 36048 8358 36060
rect 8389 36057 8401 36060
rect 8435 36057 8447 36091
rect 8389 36051 8447 36057
rect 8478 36048 8484 36100
rect 8536 36088 8542 36100
rect 10873 36091 10931 36097
rect 10873 36088 10885 36091
rect 8536 36060 10885 36088
rect 8536 36048 8542 36060
rect 10873 36057 10885 36060
rect 10919 36088 10931 36091
rect 11698 36088 11704 36100
rect 10919 36060 11704 36088
rect 10919 36057 10931 36060
rect 10873 36051 10931 36057
rect 11698 36048 11704 36060
rect 11756 36048 11762 36100
rect 13556 36088 13584 36119
rect 14826 36116 14832 36168
rect 14884 36156 14890 36168
rect 15304 36156 15332 36187
rect 14884 36128 15332 36156
rect 15933 36159 15991 36165
rect 14884 36116 14890 36128
rect 15933 36125 15945 36159
rect 15979 36156 15991 36159
rect 17126 36156 17132 36168
rect 15979 36128 17132 36156
rect 15979 36125 15991 36128
rect 15933 36119 15991 36125
rect 17126 36116 17132 36128
rect 17184 36116 17190 36168
rect 18248 36165 18276 36196
rect 18598 36184 18604 36196
rect 18656 36224 18662 36236
rect 19996 36233 20024 36264
rect 20438 36252 20444 36264
rect 20496 36252 20502 36304
rect 23216 36292 23244 36332
rect 23339 36329 23351 36363
rect 23385 36360 23397 36363
rect 23566 36360 23572 36372
rect 23385 36332 23572 36360
rect 23385 36329 23397 36332
rect 23339 36323 23397 36329
rect 23566 36320 23572 36332
rect 23624 36320 23630 36372
rect 26234 36360 26240 36372
rect 25700 36332 26240 36360
rect 25700 36292 25728 36332
rect 26234 36320 26240 36332
rect 26292 36320 26298 36372
rect 27706 36320 27712 36372
rect 27764 36360 27770 36372
rect 29270 36360 29276 36372
rect 27764 36332 29276 36360
rect 27764 36320 27770 36332
rect 29270 36320 29276 36332
rect 29328 36320 29334 36372
rect 29822 36320 29828 36372
rect 29880 36360 29886 36372
rect 30837 36363 30895 36369
rect 30837 36360 30849 36363
rect 29880 36332 30849 36360
rect 29880 36320 29886 36332
rect 30837 36329 30849 36332
rect 30883 36329 30895 36363
rect 30837 36323 30895 36329
rect 32030 36320 32036 36372
rect 32088 36360 32094 36372
rect 32088 36332 34376 36360
rect 32088 36320 32094 36332
rect 29454 36292 29460 36304
rect 23216 36264 25728 36292
rect 25792 36264 29460 36292
rect 19889 36227 19947 36233
rect 19889 36224 19901 36227
rect 18656 36196 19901 36224
rect 18656 36184 18662 36196
rect 19889 36193 19901 36196
rect 19935 36193 19947 36227
rect 19889 36187 19947 36193
rect 19981 36227 20039 36233
rect 19981 36193 19993 36227
rect 20027 36193 20039 36227
rect 21542 36224 21548 36236
rect 19981 36187 20039 36193
rect 20088 36196 21548 36224
rect 18141 36159 18199 36165
rect 18141 36125 18153 36159
rect 18187 36125 18199 36159
rect 18141 36119 18199 36125
rect 18233 36159 18291 36165
rect 18233 36125 18245 36159
rect 18279 36125 18291 36159
rect 18233 36119 18291 36125
rect 16200 36091 16258 36097
rect 13556 36060 16160 36088
rect 3510 35980 3516 36032
rect 3568 36020 3574 36032
rect 7006 36020 7012 36032
rect 3568 35992 7012 36020
rect 3568 35980 3574 35992
rect 7006 35980 7012 35992
rect 7064 35980 7070 36032
rect 7558 35980 7564 36032
rect 7616 36020 7622 36032
rect 8128 36020 8156 36048
rect 7616 35992 8156 36020
rect 7616 35980 7622 35992
rect 9674 35980 9680 36032
rect 9732 35980 9738 36032
rect 10965 36023 11023 36029
rect 10965 35989 10977 36023
rect 11011 36020 11023 36023
rect 11146 36020 11152 36032
rect 11011 35992 11152 36020
rect 11011 35989 11023 35992
rect 10965 35983 11023 35989
rect 11146 35980 11152 35992
rect 11204 36020 11210 36032
rect 12066 36020 12072 36032
rect 11204 35992 12072 36020
rect 11204 35980 11210 35992
rect 12066 35980 12072 35992
rect 12124 35980 12130 36032
rect 13630 35980 13636 36032
rect 13688 35980 13694 36032
rect 15105 36023 15163 36029
rect 15105 35989 15117 36023
rect 15151 36020 15163 36023
rect 15746 36020 15752 36032
rect 15151 35992 15752 36020
rect 15151 35989 15163 35992
rect 15105 35983 15163 35989
rect 15746 35980 15752 35992
rect 15804 35980 15810 36032
rect 16132 36020 16160 36060
rect 16200 36057 16212 36091
rect 16246 36088 16258 36091
rect 16390 36088 16396 36100
rect 16246 36060 16396 36088
rect 16246 36057 16258 36060
rect 16200 36051 16258 36057
rect 16390 36048 16396 36060
rect 16448 36048 16454 36100
rect 17236 36060 18000 36088
rect 17236 36020 17264 36060
rect 16132 35992 17264 36020
rect 17310 35980 17316 36032
rect 17368 35980 17374 36032
rect 17972 36020 18000 36060
rect 18046 36020 18052 36032
rect 17972 35992 18052 36020
rect 18046 35980 18052 35992
rect 18104 35980 18110 36032
rect 18156 36020 18184 36119
rect 18414 36116 18420 36168
rect 18472 36116 18478 36168
rect 18506 36116 18512 36168
rect 18564 36156 18570 36168
rect 19242 36156 19248 36168
rect 18564 36128 19248 36156
rect 18564 36116 18570 36128
rect 19242 36116 19248 36128
rect 19300 36156 19306 36168
rect 20088 36156 20116 36196
rect 21542 36184 21548 36196
rect 21600 36184 21606 36236
rect 21913 36227 21971 36233
rect 21913 36193 21925 36227
rect 21959 36224 21971 36227
rect 22646 36224 22652 36236
rect 21959 36196 22652 36224
rect 21959 36193 21971 36196
rect 21913 36187 21971 36193
rect 22646 36184 22652 36196
rect 22704 36184 22710 36236
rect 24670 36184 24676 36236
rect 24728 36224 24734 36236
rect 24728 36196 25360 36224
rect 24728 36184 24734 36196
rect 19300 36128 20116 36156
rect 19300 36116 19306 36128
rect 20162 36116 20168 36168
rect 20220 36156 20226 36168
rect 20625 36159 20683 36165
rect 20625 36156 20637 36159
rect 20220 36128 20637 36156
rect 20220 36116 20226 36128
rect 20625 36125 20637 36128
rect 20671 36125 20683 36159
rect 20625 36119 20683 36125
rect 20898 36116 20904 36168
rect 20956 36116 20962 36168
rect 23842 36116 23848 36168
rect 23900 36116 23906 36168
rect 24029 36159 24087 36165
rect 24029 36125 24041 36159
rect 24075 36156 24087 36159
rect 24210 36156 24216 36168
rect 24075 36128 24216 36156
rect 24075 36125 24087 36128
rect 24029 36119 24087 36125
rect 24210 36116 24216 36128
rect 24268 36116 24274 36168
rect 24578 36116 24584 36168
rect 24636 36116 24642 36168
rect 24765 36159 24823 36165
rect 24765 36125 24777 36159
rect 24811 36125 24823 36159
rect 25332 36156 25360 36196
rect 25406 36184 25412 36236
rect 25464 36184 25470 36236
rect 25498 36184 25504 36236
rect 25556 36224 25562 36236
rect 25792 36233 25820 36264
rect 29454 36252 29460 36264
rect 29512 36292 29518 36304
rect 29914 36292 29920 36304
rect 29512 36264 29920 36292
rect 29512 36252 29518 36264
rect 29914 36252 29920 36264
rect 29972 36252 29978 36304
rect 32858 36252 32864 36304
rect 32916 36292 32922 36304
rect 34057 36295 34115 36301
rect 34057 36292 34069 36295
rect 32916 36264 34069 36292
rect 32916 36252 32922 36264
rect 34057 36261 34069 36264
rect 34103 36261 34115 36295
rect 34348 36292 34376 36332
rect 34422 36320 34428 36372
rect 34480 36360 34486 36372
rect 38013 36363 38071 36369
rect 38013 36360 38025 36363
rect 34480 36332 38025 36360
rect 34480 36320 34486 36332
rect 38013 36329 38025 36332
rect 38059 36329 38071 36363
rect 38013 36323 38071 36329
rect 36078 36292 36084 36304
rect 34348 36264 36084 36292
rect 34057 36255 34115 36261
rect 36078 36252 36084 36264
rect 36136 36252 36142 36304
rect 38102 36252 38108 36304
rect 38160 36252 38166 36304
rect 25777 36227 25835 36233
rect 25777 36224 25789 36227
rect 25556 36196 25789 36224
rect 25556 36184 25562 36196
rect 25777 36193 25789 36196
rect 25823 36193 25835 36227
rect 27614 36224 27620 36236
rect 25777 36187 25835 36193
rect 25884 36196 27620 36224
rect 25884 36156 25912 36196
rect 25332 36128 25912 36156
rect 24765 36119 24823 36125
rect 18598 36048 18604 36100
rect 18656 36088 18662 36100
rect 18877 36091 18935 36097
rect 18877 36088 18889 36091
rect 18656 36060 18889 36088
rect 18656 36048 18662 36060
rect 18877 36057 18889 36060
rect 18923 36057 18935 36091
rect 18877 36051 18935 36057
rect 18966 36048 18972 36100
rect 19024 36088 19030 36100
rect 21174 36088 21180 36100
rect 19024 36060 21180 36088
rect 19024 36048 19030 36060
rect 21174 36048 21180 36060
rect 21232 36048 21238 36100
rect 22278 36048 22284 36100
rect 22336 36048 22342 36100
rect 23860 36088 23888 36116
rect 24670 36088 24676 36100
rect 23860 36060 24676 36088
rect 24670 36048 24676 36060
rect 24728 36088 24734 36100
rect 24780 36088 24808 36119
rect 26050 36116 26056 36168
rect 26108 36156 26114 36168
rect 26602 36156 26608 36168
rect 26108 36128 26608 36156
rect 26108 36116 26114 36128
rect 26602 36116 26608 36128
rect 26660 36116 26666 36168
rect 26878 36116 26884 36168
rect 26936 36116 26942 36168
rect 26988 36142 27016 36196
rect 27614 36184 27620 36196
rect 27672 36184 27678 36236
rect 28534 36184 28540 36236
rect 28592 36224 28598 36236
rect 30009 36227 30067 36233
rect 28592 36196 28764 36224
rect 28592 36184 28598 36196
rect 27798 36116 27804 36168
rect 27856 36156 27862 36168
rect 28736 36165 28764 36196
rect 30009 36193 30021 36227
rect 30055 36224 30067 36227
rect 30098 36224 30104 36236
rect 30055 36196 30104 36224
rect 30055 36193 30067 36196
rect 30009 36187 30067 36193
rect 30098 36184 30104 36196
rect 30156 36224 30162 36236
rect 30374 36224 30380 36236
rect 30156 36196 30380 36224
rect 30156 36184 30162 36196
rect 30374 36184 30380 36196
rect 30432 36184 30438 36236
rect 31846 36184 31852 36236
rect 31904 36184 31910 36236
rect 32950 36184 32956 36236
rect 33008 36224 33014 36236
rect 38289 36227 38347 36233
rect 38289 36224 38301 36227
rect 33008 36196 35296 36224
rect 33008 36184 33014 36196
rect 28629 36159 28687 36165
rect 28629 36156 28641 36159
rect 27856 36128 28641 36156
rect 27856 36116 27862 36128
rect 28629 36125 28641 36128
rect 28675 36125 28687 36159
rect 28629 36119 28687 36125
rect 28721 36159 28779 36165
rect 28721 36125 28733 36159
rect 28767 36125 28779 36159
rect 28721 36119 28779 36125
rect 24728 36060 24808 36088
rect 24728 36048 24734 36060
rect 25038 36048 25044 36100
rect 25096 36088 25102 36100
rect 25894 36091 25952 36097
rect 25894 36088 25906 36091
rect 25096 36060 25906 36088
rect 25096 36048 25102 36060
rect 25894 36057 25906 36060
rect 25940 36088 25952 36091
rect 25940 36060 26188 36088
rect 25940 36057 25952 36060
rect 25894 36051 25952 36057
rect 19797 36023 19855 36029
rect 19797 36020 19809 36023
rect 18156 35992 19809 36020
rect 19797 35989 19809 35992
rect 19843 36020 19855 36023
rect 23106 36020 23112 36032
rect 19843 35992 23112 36020
rect 19843 35989 19855 35992
rect 19797 35983 19855 35989
rect 23106 35980 23112 35992
rect 23164 35980 23170 36032
rect 23566 35980 23572 36032
rect 23624 36020 23630 36032
rect 23937 36023 23995 36029
rect 23937 36020 23949 36023
rect 23624 35992 23949 36020
rect 23624 35980 23630 35992
rect 23937 35989 23949 35992
rect 23983 35989 23995 36023
rect 23937 35983 23995 35989
rect 24854 35980 24860 36032
rect 24912 35980 24918 36032
rect 25130 35980 25136 36032
rect 25188 36020 25194 36032
rect 25685 36023 25743 36029
rect 25685 36020 25697 36023
rect 25188 35992 25697 36020
rect 25188 35980 25194 35992
rect 25685 35989 25697 35992
rect 25731 35989 25743 36023
rect 25685 35983 25743 35989
rect 26050 35980 26056 36032
rect 26108 35980 26114 36032
rect 26160 36020 26188 36060
rect 26234 36048 26240 36100
rect 26292 36088 26298 36100
rect 27614 36088 27620 36100
rect 26292 36060 27620 36088
rect 26292 36048 26298 36060
rect 27614 36048 27620 36060
rect 27672 36048 27678 36100
rect 26970 36020 26976 36032
rect 26160 35992 26976 36020
rect 26970 35980 26976 35992
rect 27028 36020 27034 36032
rect 28074 36020 28080 36032
rect 27028 35992 28080 36020
rect 27028 35980 27034 35992
rect 28074 35980 28080 35992
rect 28132 35980 28138 36032
rect 28166 35980 28172 36032
rect 28224 36020 28230 36032
rect 28353 36023 28411 36029
rect 28353 36020 28365 36023
rect 28224 35992 28365 36020
rect 28224 35980 28230 35992
rect 28353 35989 28365 35992
rect 28399 35989 28411 36023
rect 28644 36020 28672 36119
rect 28810 36116 28816 36168
rect 28868 36116 28874 36168
rect 28902 36116 28908 36168
rect 28960 36156 28966 36168
rect 28997 36159 29055 36165
rect 28997 36156 29009 36159
rect 28960 36128 29009 36156
rect 28960 36116 28966 36128
rect 28997 36125 29009 36128
rect 29043 36125 29055 36159
rect 28997 36119 29055 36125
rect 29086 36116 29092 36168
rect 29144 36156 29150 36168
rect 29733 36159 29791 36165
rect 29733 36156 29745 36159
rect 29144 36128 29745 36156
rect 29144 36116 29150 36128
rect 29733 36125 29745 36128
rect 29779 36125 29791 36159
rect 29733 36119 29791 36125
rect 30834 36116 30840 36168
rect 30892 36156 30898 36168
rect 33873 36159 33931 36165
rect 33873 36156 33885 36159
rect 30892 36128 33885 36156
rect 30892 36116 30898 36128
rect 33873 36125 33885 36128
rect 33919 36125 33931 36159
rect 33873 36119 33931 36125
rect 34885 36159 34943 36165
rect 34885 36125 34897 36159
rect 34931 36125 34943 36159
rect 34885 36119 34943 36125
rect 30098 36048 30104 36100
rect 30156 36088 30162 36100
rect 30745 36091 30803 36097
rect 30745 36088 30757 36091
rect 30156 36060 30757 36088
rect 30156 36048 30162 36060
rect 30745 36057 30757 36060
rect 30791 36057 30803 36091
rect 30745 36051 30803 36057
rect 31938 36048 31944 36100
rect 31996 36088 32002 36100
rect 32094 36091 32152 36097
rect 32094 36088 32106 36091
rect 31996 36060 32106 36088
rect 31996 36048 32002 36060
rect 32094 36057 32106 36060
rect 32140 36057 32152 36091
rect 34900 36088 34928 36119
rect 32094 36051 32152 36057
rect 33152 36060 34928 36088
rect 35161 36091 35219 36097
rect 33152 36020 33180 36060
rect 35161 36057 35173 36091
rect 35207 36057 35219 36091
rect 35268 36088 35296 36196
rect 37099 36196 38301 36224
rect 36078 36116 36084 36168
rect 36136 36116 36142 36168
rect 36170 36116 36176 36168
rect 36228 36156 36234 36168
rect 36337 36159 36395 36165
rect 36337 36156 36349 36159
rect 36228 36128 36349 36156
rect 36228 36116 36234 36128
rect 36337 36125 36349 36128
rect 36383 36125 36395 36159
rect 37099 36156 37127 36196
rect 38289 36193 38301 36196
rect 38335 36193 38347 36227
rect 38289 36187 38347 36193
rect 36337 36119 36395 36125
rect 36464 36128 37127 36156
rect 38013 36159 38071 36165
rect 36464 36088 36492 36128
rect 38013 36125 38025 36159
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 35268 36060 36492 36088
rect 35161 36051 35219 36057
rect 28644 35992 33180 36020
rect 33229 36023 33287 36029
rect 28353 35983 28411 35989
rect 33229 35989 33241 36023
rect 33275 36020 33287 36023
rect 33318 36020 33324 36032
rect 33275 35992 33324 36020
rect 33275 35989 33287 35992
rect 33229 35983 33287 35989
rect 33318 35980 33324 35992
rect 33376 35980 33382 36032
rect 33410 35980 33416 36032
rect 33468 36020 33474 36032
rect 35176 36020 35204 36051
rect 36538 36048 36544 36100
rect 36596 36088 36602 36100
rect 38028 36088 38056 36119
rect 36596 36060 38056 36088
rect 36596 36048 36602 36060
rect 33468 35992 35204 36020
rect 33468 35980 33474 35992
rect 37182 35980 37188 36032
rect 37240 36020 37246 36032
rect 37461 36023 37519 36029
rect 37461 36020 37473 36023
rect 37240 35992 37473 36020
rect 37240 35980 37246 35992
rect 37461 35989 37473 35992
rect 37507 35989 37519 36023
rect 37461 35983 37519 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 4433 35819 4491 35825
rect 4433 35785 4445 35819
rect 4479 35816 4491 35819
rect 4798 35816 4804 35828
rect 4479 35788 4804 35816
rect 4479 35785 4491 35788
rect 4433 35779 4491 35785
rect 4798 35776 4804 35788
rect 4856 35776 4862 35828
rect 5997 35819 6055 35825
rect 5997 35785 6009 35819
rect 6043 35816 6055 35819
rect 6178 35816 6184 35828
rect 6043 35788 6184 35816
rect 6043 35785 6055 35788
rect 5997 35779 6055 35785
rect 6178 35776 6184 35788
rect 6236 35776 6242 35828
rect 6638 35776 6644 35828
rect 6696 35776 6702 35828
rect 9401 35819 9459 35825
rect 9401 35785 9413 35819
rect 9447 35816 9459 35819
rect 9582 35816 9588 35828
rect 9447 35788 9588 35816
rect 9447 35785 9459 35788
rect 9401 35779 9459 35785
rect 9582 35776 9588 35788
rect 9640 35816 9646 35828
rect 10321 35819 10379 35825
rect 10321 35816 10333 35819
rect 9640 35788 10333 35816
rect 9640 35776 9646 35788
rect 10321 35785 10333 35788
rect 10367 35785 10379 35819
rect 10321 35779 10379 35785
rect 14461 35819 14519 35825
rect 14461 35785 14473 35819
rect 14507 35816 14519 35819
rect 15930 35816 15936 35828
rect 14507 35788 15936 35816
rect 14507 35785 14519 35788
rect 14461 35779 14519 35785
rect 15930 35776 15936 35788
rect 15988 35776 15994 35828
rect 17310 35776 17316 35828
rect 17368 35816 17374 35828
rect 17405 35819 17463 35825
rect 17405 35816 17417 35819
rect 17368 35788 17417 35816
rect 17368 35776 17374 35788
rect 17405 35785 17417 35788
rect 17451 35785 17463 35819
rect 19150 35816 19156 35828
rect 17405 35779 17463 35785
rect 17512 35788 19156 35816
rect 3418 35708 3424 35760
rect 3476 35748 3482 35760
rect 5350 35748 5356 35760
rect 3476 35720 5356 35748
rect 3476 35708 3482 35720
rect 3896 35689 3924 35720
rect 5350 35708 5356 35720
rect 5408 35708 5414 35760
rect 5442 35708 5448 35760
rect 5500 35748 5506 35760
rect 5500 35720 6592 35748
rect 5500 35708 5506 35720
rect 3697 35683 3755 35689
rect 3697 35649 3709 35683
rect 3743 35649 3755 35683
rect 3697 35643 3755 35649
rect 3881 35683 3939 35689
rect 3881 35649 3893 35683
rect 3927 35649 3939 35683
rect 3881 35643 3939 35649
rect 3712 35612 3740 35643
rect 4338 35640 4344 35692
rect 4396 35640 4402 35692
rect 4522 35640 4528 35692
rect 4580 35640 4586 35692
rect 4798 35640 4804 35692
rect 4856 35640 4862 35692
rect 4982 35640 4988 35692
rect 5040 35640 5046 35692
rect 5077 35683 5135 35689
rect 5077 35649 5089 35683
rect 5123 35680 5135 35683
rect 5258 35680 5264 35692
rect 5123 35652 5264 35680
rect 5123 35649 5135 35652
rect 5077 35643 5135 35649
rect 5258 35640 5264 35652
rect 5316 35640 5322 35692
rect 5721 35683 5779 35689
rect 5721 35649 5733 35683
rect 5767 35680 5779 35683
rect 5810 35680 5816 35692
rect 5767 35652 5816 35680
rect 5767 35649 5779 35652
rect 5721 35643 5779 35649
rect 5810 35640 5816 35652
rect 5868 35640 5874 35692
rect 6564 35689 6592 35720
rect 6914 35708 6920 35760
rect 6972 35748 6978 35760
rect 9766 35748 9772 35760
rect 6972 35720 9772 35748
rect 6972 35708 6978 35720
rect 6549 35683 6607 35689
rect 6549 35649 6561 35683
rect 6595 35680 6607 35683
rect 7098 35680 7104 35692
rect 6595 35652 7104 35680
rect 6595 35649 6607 35652
rect 6549 35643 6607 35649
rect 7098 35640 7104 35652
rect 7156 35640 7162 35692
rect 7300 35689 7328 35720
rect 9766 35708 9772 35720
rect 9824 35708 9830 35760
rect 10226 35708 10232 35760
rect 10284 35708 10290 35760
rect 13633 35751 13691 35757
rect 13633 35717 13645 35751
rect 13679 35748 13691 35751
rect 17512 35748 17540 35788
rect 19150 35776 19156 35788
rect 19208 35776 19214 35828
rect 19242 35776 19248 35828
rect 19300 35816 19306 35828
rect 19300 35788 21036 35816
rect 19300 35776 19306 35788
rect 13679 35720 17540 35748
rect 13679 35717 13691 35720
rect 13633 35711 13691 35717
rect 7285 35683 7343 35689
rect 7285 35649 7297 35683
rect 7331 35649 7343 35683
rect 7285 35643 7343 35649
rect 7374 35640 7380 35692
rect 7432 35640 7438 35692
rect 8110 35680 8116 35692
rect 7484 35652 8116 35680
rect 5445 35615 5503 35621
rect 3712 35584 4844 35612
rect 4816 35553 4844 35584
rect 5445 35581 5457 35615
rect 5491 35612 5503 35615
rect 5997 35615 6055 35621
rect 5997 35612 6009 35615
rect 5491 35584 6009 35612
rect 5491 35581 5503 35584
rect 5445 35575 5503 35581
rect 5997 35581 6009 35584
rect 6043 35612 6055 35615
rect 6822 35612 6828 35624
rect 6043 35584 6828 35612
rect 6043 35581 6055 35584
rect 5997 35575 6055 35581
rect 6822 35572 6828 35584
rect 6880 35572 6886 35624
rect 4801 35547 4859 35553
rect 4801 35513 4813 35547
rect 4847 35513 4859 35547
rect 4801 35507 4859 35513
rect 5813 35547 5871 35553
rect 5813 35513 5825 35547
rect 5859 35544 5871 35547
rect 7484 35544 7512 35652
rect 8110 35640 8116 35652
rect 8168 35640 8174 35692
rect 8288 35683 8346 35689
rect 8288 35649 8300 35683
rect 8334 35680 8346 35683
rect 9122 35680 9128 35692
rect 8334 35652 9128 35680
rect 8334 35649 8346 35652
rect 8288 35643 8346 35649
rect 9122 35640 9128 35652
rect 9180 35640 9186 35692
rect 11698 35640 11704 35692
rect 11756 35680 11762 35692
rect 11977 35683 12035 35689
rect 11977 35680 11989 35683
rect 11756 35652 11989 35680
rect 11756 35640 11762 35652
rect 11977 35649 11989 35652
rect 12023 35649 12035 35683
rect 11977 35643 12035 35649
rect 12066 35640 12072 35692
rect 12124 35640 12130 35692
rect 12253 35683 12311 35689
rect 12253 35649 12265 35683
rect 12299 35680 12311 35683
rect 12434 35680 12440 35692
rect 12299 35652 12440 35680
rect 12299 35649 12311 35652
rect 12253 35643 12311 35649
rect 7650 35572 7656 35624
rect 7708 35612 7714 35624
rect 8021 35615 8079 35621
rect 8021 35612 8033 35615
rect 7708 35584 8033 35612
rect 7708 35572 7714 35584
rect 8021 35581 8033 35584
rect 8067 35581 8079 35615
rect 8021 35575 8079 35581
rect 9858 35572 9864 35624
rect 9916 35612 9922 35624
rect 10413 35615 10471 35621
rect 10413 35612 10425 35615
rect 9916 35584 10425 35612
rect 9916 35572 9922 35584
rect 10413 35581 10425 35584
rect 10459 35612 10471 35615
rect 12268 35612 12296 35643
rect 12434 35640 12440 35652
rect 12492 35640 12498 35692
rect 13078 35640 13084 35692
rect 13136 35680 13142 35692
rect 13265 35683 13323 35689
rect 13265 35680 13277 35683
rect 13136 35652 13277 35680
rect 13136 35640 13142 35652
rect 13265 35649 13277 35652
rect 13311 35649 13323 35683
rect 13265 35643 13323 35649
rect 13449 35683 13507 35689
rect 13449 35649 13461 35683
rect 13495 35680 13507 35683
rect 13495 35652 15148 35680
rect 13495 35649 13507 35652
rect 13449 35643 13507 35649
rect 10459 35584 12434 35612
rect 10459 35581 10471 35584
rect 10413 35575 10471 35581
rect 5859 35516 7512 35544
rect 7561 35547 7619 35553
rect 5859 35513 5871 35516
rect 5813 35507 5871 35513
rect 7561 35513 7573 35547
rect 7607 35544 7619 35547
rect 7926 35544 7932 35556
rect 7607 35516 7932 35544
rect 7607 35513 7619 35516
rect 7561 35507 7619 35513
rect 7926 35504 7932 35516
rect 7984 35504 7990 35556
rect 12406 35544 12434 35584
rect 12710 35572 12716 35624
rect 12768 35572 12774 35624
rect 14553 35615 14611 35621
rect 14553 35581 14565 35615
rect 14599 35581 14611 35615
rect 14553 35575 14611 35581
rect 14737 35615 14795 35621
rect 14737 35581 14749 35615
rect 14783 35581 14795 35615
rect 15120 35612 15148 35652
rect 15194 35640 15200 35692
rect 15252 35680 15258 35692
rect 15657 35683 15715 35689
rect 15657 35680 15669 35683
rect 15252 35652 15669 35680
rect 15252 35640 15258 35652
rect 15657 35649 15669 35652
rect 15703 35649 15715 35683
rect 15657 35643 15715 35649
rect 15746 35640 15752 35692
rect 15804 35640 15810 35692
rect 15841 35683 15899 35689
rect 15841 35649 15853 35683
rect 15887 35680 15899 35683
rect 17497 35683 17555 35689
rect 17497 35680 17509 35683
rect 15887 35652 17509 35680
rect 15887 35649 15899 35652
rect 15841 35643 15899 35649
rect 17497 35649 17509 35652
rect 17543 35680 17555 35683
rect 18322 35680 18328 35692
rect 17543 35652 18328 35680
rect 17543 35649 17555 35652
rect 17497 35643 17555 35649
rect 15470 35612 15476 35624
rect 15120 35584 15476 35612
rect 14737 35575 14795 35581
rect 12406 35516 14228 35544
rect 3694 35436 3700 35488
rect 3752 35436 3758 35488
rect 4522 35436 4528 35488
rect 4580 35476 4586 35488
rect 5442 35476 5448 35488
rect 4580 35448 5448 35476
rect 4580 35436 4586 35448
rect 5442 35436 5448 35448
rect 5500 35436 5506 35488
rect 5902 35436 5908 35488
rect 5960 35476 5966 35488
rect 9861 35479 9919 35485
rect 9861 35476 9873 35479
rect 5960 35448 9873 35476
rect 5960 35436 5966 35448
rect 9861 35445 9873 35448
rect 9907 35445 9919 35479
rect 9861 35439 9919 35445
rect 14090 35436 14096 35488
rect 14148 35436 14154 35488
rect 14200 35476 14228 35516
rect 14274 35504 14280 35556
rect 14332 35544 14338 35556
rect 14568 35544 14596 35575
rect 14332 35516 14596 35544
rect 14752 35544 14780 35575
rect 15470 35572 15476 35584
rect 15528 35572 15534 35624
rect 15565 35615 15623 35621
rect 15565 35581 15577 35615
rect 15611 35612 15623 35615
rect 15764 35612 15792 35640
rect 15611 35584 15792 35612
rect 15611 35581 15623 35584
rect 15565 35575 15623 35581
rect 15856 35544 15884 35643
rect 18322 35640 18328 35652
rect 18380 35640 18386 35692
rect 21008 35689 21036 35788
rect 21450 35776 21456 35828
rect 21508 35816 21514 35828
rect 21508 35788 23060 35816
rect 21508 35776 21514 35788
rect 21266 35708 21272 35760
rect 21324 35708 21330 35760
rect 22281 35751 22339 35757
rect 22281 35717 22293 35751
rect 22327 35748 22339 35751
rect 22370 35748 22376 35760
rect 22327 35720 22376 35748
rect 22327 35717 22339 35720
rect 22281 35711 22339 35717
rect 22370 35708 22376 35720
rect 22428 35708 22434 35760
rect 23032 35757 23060 35788
rect 23290 35776 23296 35828
rect 23348 35816 23354 35828
rect 23348 35788 26832 35816
rect 23348 35776 23354 35788
rect 23017 35751 23075 35757
rect 23017 35717 23029 35751
rect 23063 35717 23075 35751
rect 23017 35711 23075 35717
rect 23934 35708 23940 35760
rect 23992 35748 23998 35760
rect 23992 35720 24900 35748
rect 23992 35708 23998 35720
rect 20993 35683 21051 35689
rect 18432 35652 20760 35680
rect 16298 35572 16304 35624
rect 16356 35572 16362 35624
rect 17405 35615 17463 35621
rect 17405 35581 17417 35615
rect 17451 35612 17463 35615
rect 17954 35612 17960 35624
rect 17451 35584 17960 35612
rect 17451 35581 17463 35584
rect 17405 35575 17463 35581
rect 17954 35572 17960 35584
rect 18012 35572 18018 35624
rect 14752 35516 15884 35544
rect 14332 35504 14338 35516
rect 14752 35476 14780 35516
rect 17034 35504 17040 35556
rect 17092 35544 17098 35556
rect 18432 35544 18460 35652
rect 18506 35572 18512 35624
rect 18564 35572 18570 35624
rect 18785 35615 18843 35621
rect 18785 35581 18797 35615
rect 18831 35612 18843 35615
rect 20732 35612 20760 35652
rect 20993 35649 21005 35683
rect 21039 35649 21051 35683
rect 20993 35643 21051 35649
rect 22002 35640 22008 35692
rect 22060 35640 22066 35692
rect 23750 35640 23756 35692
rect 23808 35680 23814 35692
rect 23845 35683 23903 35689
rect 23845 35680 23857 35683
rect 23808 35652 23857 35680
rect 23808 35640 23814 35652
rect 23845 35649 23857 35652
rect 23891 35649 23903 35683
rect 23845 35643 23903 35649
rect 24026 35640 24032 35692
rect 24084 35680 24090 35692
rect 24872 35689 24900 35720
rect 25958 35708 25964 35760
rect 26016 35748 26022 35760
rect 26467 35751 26525 35757
rect 26016 35720 26280 35748
rect 26016 35708 26022 35720
rect 24397 35683 24455 35689
rect 24397 35680 24409 35683
rect 24084 35652 24409 35680
rect 24084 35640 24090 35652
rect 24397 35649 24409 35652
rect 24443 35649 24455 35683
rect 24397 35643 24455 35649
rect 24857 35683 24915 35689
rect 24857 35649 24869 35683
rect 24903 35680 24915 35683
rect 25130 35680 25136 35692
rect 24903 35652 25136 35680
rect 24903 35649 24915 35652
rect 24857 35643 24915 35649
rect 21450 35612 21456 35624
rect 18831 35584 20668 35612
rect 20732 35584 21456 35612
rect 18831 35581 18843 35584
rect 18785 35575 18843 35581
rect 17092 35516 18460 35544
rect 17092 35504 17098 35516
rect 19610 35504 19616 35556
rect 19668 35544 19674 35556
rect 20530 35544 20536 35556
rect 19668 35516 20536 35544
rect 19668 35504 19674 35516
rect 20530 35504 20536 35516
rect 20588 35504 20594 35556
rect 20640 35544 20668 35584
rect 21450 35572 21456 35584
rect 21508 35572 21514 35624
rect 22922 35572 22928 35624
rect 22980 35612 22986 35624
rect 24121 35615 24179 35621
rect 24121 35612 24133 35615
rect 22980 35584 24133 35612
rect 22980 35572 22986 35584
rect 24121 35581 24133 35584
rect 24167 35581 24179 35615
rect 24412 35612 24440 35643
rect 25130 35640 25136 35652
rect 25188 35640 25194 35692
rect 25498 35640 25504 35692
rect 25556 35640 25562 35692
rect 26252 35689 26280 35720
rect 26467 35717 26479 35751
rect 26513 35748 26525 35751
rect 26804 35748 26832 35788
rect 27338 35776 27344 35828
rect 27396 35816 27402 35828
rect 27798 35816 27804 35828
rect 27396 35788 27804 35816
rect 27396 35776 27402 35788
rect 27798 35776 27804 35788
rect 27856 35776 27862 35828
rect 28810 35776 28816 35828
rect 28868 35816 28874 35828
rect 32306 35816 32312 35828
rect 28868 35788 32312 35816
rect 28868 35776 28874 35788
rect 32306 35776 32312 35788
rect 32364 35776 32370 35828
rect 32766 35776 32772 35828
rect 32824 35816 32830 35828
rect 32861 35819 32919 35825
rect 32861 35816 32873 35819
rect 32824 35788 32873 35816
rect 32824 35776 32830 35788
rect 32861 35785 32873 35788
rect 32907 35785 32919 35819
rect 32861 35779 32919 35785
rect 32950 35776 32956 35828
rect 33008 35816 33014 35828
rect 33318 35816 33324 35828
rect 33008 35788 33324 35816
rect 33008 35776 33014 35788
rect 33318 35776 33324 35788
rect 33376 35776 33382 35828
rect 37550 35776 37556 35828
rect 37608 35776 37614 35828
rect 26513 35720 26740 35748
rect 26804 35720 31248 35748
rect 26513 35717 26525 35720
rect 26467 35711 26525 35717
rect 26145 35683 26203 35689
rect 26145 35649 26157 35683
rect 26191 35649 26203 35683
rect 26145 35643 26203 35649
rect 26237 35683 26295 35689
rect 26237 35649 26249 35683
rect 26283 35649 26295 35683
rect 26237 35643 26295 35649
rect 26329 35683 26387 35689
rect 26329 35649 26341 35683
rect 26375 35655 26464 35683
rect 26375 35649 26387 35655
rect 26329 35643 26387 35649
rect 24762 35612 24768 35624
rect 24412 35584 24768 35612
rect 24121 35575 24179 35581
rect 24762 35572 24768 35584
rect 24820 35612 24826 35624
rect 25222 35612 25228 35624
rect 24820 35584 25228 35612
rect 24820 35572 24826 35584
rect 25222 35572 25228 35584
rect 25280 35572 25286 35624
rect 25590 35572 25596 35624
rect 25648 35612 25654 35624
rect 26160 35612 26188 35643
rect 25648 35584 26280 35612
rect 25648 35572 25654 35584
rect 26252 35556 26280 35584
rect 25498 35544 25504 35556
rect 20640 35516 25504 35544
rect 25498 35504 25504 35516
rect 25556 35504 25562 35556
rect 26234 35504 26240 35556
rect 26292 35504 26298 35556
rect 14200 35448 14780 35476
rect 15286 35436 15292 35488
rect 15344 35476 15350 35488
rect 16945 35479 17003 35485
rect 16945 35476 16957 35479
rect 15344 35448 16957 35476
rect 15344 35436 15350 35448
rect 16945 35445 16957 35448
rect 16991 35445 17003 35479
rect 16945 35439 17003 35445
rect 18414 35436 18420 35488
rect 18472 35476 18478 35488
rect 19889 35479 19947 35485
rect 19889 35476 19901 35479
rect 18472 35448 19901 35476
rect 18472 35436 18478 35448
rect 19889 35445 19901 35448
rect 19935 35445 19947 35479
rect 19889 35439 19947 35445
rect 20346 35436 20352 35488
rect 20404 35476 20410 35488
rect 23109 35479 23167 35485
rect 23109 35476 23121 35479
rect 20404 35448 23121 35476
rect 20404 35436 20410 35448
rect 23109 35445 23121 35448
rect 23155 35476 23167 35479
rect 23750 35476 23756 35488
rect 23155 35448 23756 35476
rect 23155 35445 23167 35448
rect 23109 35439 23167 35445
rect 23750 35436 23756 35448
rect 23808 35436 23814 35488
rect 25958 35436 25964 35488
rect 26016 35436 26022 35488
rect 26436 35476 26464 35655
rect 26602 35572 26608 35624
rect 26660 35572 26666 35624
rect 26712 35612 26740 35720
rect 31220 35692 31248 35720
rect 31754 35708 31760 35760
rect 31812 35748 31818 35760
rect 31812 35720 32352 35748
rect 31812 35708 31818 35720
rect 27893 35683 27951 35689
rect 27893 35649 27905 35683
rect 27939 35680 27951 35683
rect 28626 35680 28632 35692
rect 27939 35652 28632 35680
rect 27939 35649 27951 35652
rect 27893 35643 27951 35649
rect 28626 35640 28632 35652
rect 28684 35640 28690 35692
rect 29822 35640 29828 35692
rect 29880 35640 29886 35692
rect 29914 35640 29920 35692
rect 29972 35640 29978 35692
rect 31202 35640 31208 35692
rect 31260 35640 31266 35692
rect 32324 35689 32352 35720
rect 32582 35708 32588 35760
rect 32640 35748 32646 35760
rect 33505 35751 33563 35757
rect 33505 35748 33517 35751
rect 32640 35720 33517 35748
rect 32640 35708 32646 35720
rect 33505 35717 33517 35720
rect 33551 35717 33563 35751
rect 33505 35711 33563 35717
rect 33962 35708 33968 35760
rect 34020 35748 34026 35760
rect 36538 35748 36544 35760
rect 34020 35720 36544 35748
rect 34020 35708 34026 35720
rect 36538 35708 36544 35720
rect 36596 35708 36602 35760
rect 36906 35708 36912 35760
rect 36964 35748 36970 35760
rect 38013 35751 38071 35757
rect 38013 35748 38025 35751
rect 36964 35720 38025 35748
rect 36964 35708 36970 35720
rect 38013 35717 38025 35720
rect 38059 35717 38071 35751
rect 38013 35711 38071 35717
rect 32309 35683 32367 35689
rect 32309 35649 32321 35683
rect 32355 35680 32367 35683
rect 33042 35680 33048 35692
rect 32355 35652 33048 35680
rect 32355 35649 32367 35652
rect 32309 35643 32367 35649
rect 33042 35640 33048 35652
rect 33100 35680 33106 35692
rect 33137 35683 33195 35689
rect 33137 35680 33149 35683
rect 33100 35652 33149 35680
rect 33100 35640 33106 35652
rect 33137 35649 33149 35652
rect 33183 35649 33195 35683
rect 33137 35643 33195 35649
rect 33318 35640 33324 35692
rect 33376 35640 33382 35692
rect 33778 35640 33784 35692
rect 33836 35680 33842 35692
rect 34405 35683 34463 35689
rect 34405 35680 34417 35683
rect 33836 35652 34417 35680
rect 33836 35640 33842 35652
rect 34405 35649 34417 35652
rect 34451 35649 34463 35683
rect 34405 35643 34463 35649
rect 36633 35683 36691 35689
rect 36633 35649 36645 35683
rect 36679 35680 36691 35683
rect 36998 35680 37004 35692
rect 36679 35652 37004 35680
rect 36679 35649 36691 35652
rect 36633 35643 36691 35649
rect 36998 35640 37004 35652
rect 37056 35640 37062 35692
rect 37366 35640 37372 35692
rect 37424 35680 37430 35692
rect 37921 35683 37979 35689
rect 37921 35680 37933 35683
rect 37424 35652 37933 35680
rect 37424 35640 37430 35652
rect 37921 35649 37933 35652
rect 37967 35649 37979 35683
rect 37921 35643 37979 35649
rect 26786 35612 26792 35624
rect 26712 35584 26792 35612
rect 26786 35572 26792 35584
rect 26844 35572 26850 35624
rect 27798 35572 27804 35624
rect 27856 35572 27862 35624
rect 28074 35572 28080 35624
rect 28132 35612 28138 35624
rect 28353 35615 28411 35621
rect 28353 35612 28365 35615
rect 28132 35584 28365 35612
rect 28132 35572 28138 35584
rect 28353 35581 28365 35584
rect 28399 35612 28411 35615
rect 28994 35612 29000 35624
rect 28399 35584 29000 35612
rect 28399 35581 28411 35584
rect 28353 35575 28411 35581
rect 28994 35572 29000 35584
rect 29052 35572 29058 35624
rect 30374 35572 30380 35624
rect 30432 35572 30438 35624
rect 30650 35572 30656 35624
rect 30708 35612 30714 35624
rect 31389 35615 31447 35621
rect 31389 35612 31401 35615
rect 30708 35584 31401 35612
rect 30708 35572 30714 35584
rect 31389 35581 31401 35584
rect 31435 35581 31447 35615
rect 31389 35575 31447 35581
rect 32122 35572 32128 35624
rect 32180 35612 32186 35624
rect 32585 35615 32643 35621
rect 32585 35612 32597 35615
rect 32180 35584 32597 35612
rect 32180 35572 32186 35584
rect 32585 35581 32597 35584
rect 32631 35581 32643 35615
rect 32585 35575 32643 35581
rect 32674 35572 32680 35624
rect 32732 35612 32738 35624
rect 33226 35612 33232 35624
rect 32732 35584 33232 35612
rect 32732 35572 32738 35584
rect 33226 35572 33232 35584
rect 33284 35572 33290 35624
rect 34146 35572 34152 35624
rect 34204 35572 34210 35624
rect 36354 35572 36360 35624
rect 36412 35612 36418 35624
rect 36909 35615 36967 35621
rect 36909 35612 36921 35615
rect 36412 35584 36921 35612
rect 36412 35572 36418 35584
rect 36909 35581 36921 35584
rect 36955 35581 36967 35615
rect 36909 35575 36967 35581
rect 38102 35572 38108 35624
rect 38160 35572 38166 35624
rect 26694 35504 26700 35556
rect 26752 35544 26758 35556
rect 33689 35547 33747 35553
rect 33689 35544 33701 35547
rect 26752 35516 33701 35544
rect 26752 35504 26758 35516
rect 33689 35513 33701 35516
rect 33735 35513 33747 35547
rect 36722 35544 36728 35556
rect 33689 35507 33747 35513
rect 35084 35516 36728 35544
rect 26878 35476 26884 35488
rect 26436 35448 26884 35476
rect 26878 35436 26884 35448
rect 26936 35436 26942 35488
rect 28258 35436 28264 35488
rect 28316 35436 28322 35488
rect 28629 35479 28687 35485
rect 28629 35445 28641 35479
rect 28675 35476 28687 35479
rect 28902 35476 28908 35488
rect 28675 35448 28908 35476
rect 28675 35445 28687 35448
rect 28629 35439 28687 35445
rect 28902 35436 28908 35448
rect 28960 35476 28966 35488
rect 29454 35476 29460 35488
rect 28960 35448 29460 35476
rect 28960 35436 28966 35448
rect 29454 35436 29460 35448
rect 29512 35436 29518 35488
rect 30282 35436 30288 35488
rect 30340 35436 30346 35488
rect 30466 35436 30472 35488
rect 30524 35436 30530 35488
rect 32674 35436 32680 35488
rect 32732 35436 32738 35488
rect 33594 35436 33600 35488
rect 33652 35476 33658 35488
rect 35084 35476 35112 35516
rect 36722 35504 36728 35516
rect 36780 35504 36786 35556
rect 33652 35448 35112 35476
rect 33652 35436 33658 35448
rect 35342 35436 35348 35488
rect 35400 35476 35406 35488
rect 35529 35479 35587 35485
rect 35529 35476 35541 35479
rect 35400 35448 35541 35476
rect 35400 35436 35406 35448
rect 35529 35445 35541 35448
rect 35575 35445 35587 35479
rect 35529 35439 35587 35445
rect 36449 35479 36507 35485
rect 36449 35445 36461 35479
rect 36495 35476 36507 35479
rect 36630 35476 36636 35488
rect 36495 35448 36636 35476
rect 36495 35445 36507 35448
rect 36449 35439 36507 35445
rect 36630 35436 36636 35448
rect 36688 35436 36694 35488
rect 36817 35479 36875 35485
rect 36817 35445 36829 35479
rect 36863 35476 36875 35479
rect 38930 35476 38936 35488
rect 36863 35448 38936 35476
rect 36863 35445 36875 35448
rect 36817 35439 36875 35445
rect 38930 35436 38936 35448
rect 38988 35436 38994 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 4338 35232 4344 35284
rect 4396 35272 4402 35284
rect 4982 35272 4988 35284
rect 4396 35244 4988 35272
rect 4396 35232 4402 35244
rect 4982 35232 4988 35244
rect 5040 35232 5046 35284
rect 5077 35275 5135 35281
rect 5077 35241 5089 35275
rect 5123 35272 5135 35275
rect 5258 35272 5264 35284
rect 5123 35244 5264 35272
rect 5123 35241 5135 35244
rect 5077 35235 5135 35241
rect 5258 35232 5264 35244
rect 5316 35232 5322 35284
rect 8389 35275 8447 35281
rect 8389 35241 8401 35275
rect 8435 35272 8447 35275
rect 8662 35272 8668 35284
rect 8435 35244 8668 35272
rect 8435 35241 8447 35244
rect 8389 35235 8447 35241
rect 8662 35232 8668 35244
rect 8720 35232 8726 35284
rect 9122 35232 9128 35284
rect 9180 35232 9186 35284
rect 11517 35275 11575 35281
rect 11517 35272 11529 35275
rect 9232 35244 11529 35272
rect 4801 35207 4859 35213
rect 4801 35173 4813 35207
rect 4847 35204 4859 35207
rect 5534 35204 5540 35216
rect 4847 35176 5540 35204
rect 4847 35173 4859 35176
rect 4801 35167 4859 35173
rect 4816 35136 4844 35167
rect 5534 35164 5540 35176
rect 5592 35164 5598 35216
rect 8018 35164 8024 35216
rect 8076 35204 8082 35216
rect 9232 35204 9260 35244
rect 11517 35241 11529 35244
rect 11563 35241 11575 35275
rect 11517 35235 11575 35241
rect 13630 35232 13636 35284
rect 13688 35272 13694 35284
rect 14461 35275 14519 35281
rect 14461 35272 14473 35275
rect 13688 35244 14473 35272
rect 13688 35232 13694 35244
rect 14461 35241 14473 35244
rect 14507 35241 14519 35275
rect 14461 35235 14519 35241
rect 16390 35232 16396 35284
rect 16448 35272 16454 35284
rect 16577 35275 16635 35281
rect 16577 35272 16589 35275
rect 16448 35244 16589 35272
rect 16448 35232 16454 35244
rect 16577 35241 16589 35244
rect 16623 35241 16635 35275
rect 16577 35235 16635 35241
rect 18138 35232 18144 35284
rect 18196 35272 18202 35284
rect 18509 35275 18567 35281
rect 18509 35272 18521 35275
rect 18196 35244 18521 35272
rect 18196 35232 18202 35244
rect 18509 35241 18521 35244
rect 18555 35241 18567 35275
rect 20346 35272 20352 35284
rect 18509 35235 18567 35241
rect 18616 35244 20352 35272
rect 8076 35176 9260 35204
rect 9416 35176 11560 35204
rect 8076 35164 8082 35176
rect 5721 35139 5779 35145
rect 5721 35136 5733 35139
rect 4264 35108 4844 35136
rect 5552 35108 5733 35136
rect 4264 35077 4292 35108
rect 5552 35080 5580 35108
rect 5721 35105 5733 35108
rect 5767 35136 5779 35139
rect 6914 35136 6920 35148
rect 5767 35108 6920 35136
rect 5767 35105 5779 35108
rect 5721 35099 5779 35105
rect 6914 35096 6920 35108
rect 6972 35096 6978 35148
rect 7374 35096 7380 35148
rect 7432 35136 7438 35148
rect 7432 35108 7972 35136
rect 7432 35096 7438 35108
rect 4249 35071 4307 35077
rect 4249 35037 4261 35071
rect 4295 35037 4307 35071
rect 4249 35031 4307 35037
rect 4338 35028 4344 35080
rect 4396 35028 4402 35080
rect 4433 35071 4491 35077
rect 4433 35037 4445 35071
rect 4479 35068 4491 35071
rect 4479 35040 5488 35068
rect 4479 35037 4491 35040
rect 4433 35031 4491 35037
rect 4356 35000 4384 35028
rect 4893 35003 4951 35009
rect 4893 35000 4905 35003
rect 4356 34972 4905 35000
rect 4893 34969 4905 34972
rect 4939 34969 4951 35003
rect 4893 34963 4951 34969
rect 4341 34935 4399 34941
rect 4341 34901 4353 34935
rect 4387 34932 4399 34935
rect 4614 34932 4620 34944
rect 4387 34904 4620 34932
rect 4387 34901 4399 34904
rect 4341 34895 4399 34901
rect 4614 34892 4620 34904
rect 4672 34892 4678 34944
rect 4798 34892 4804 34944
rect 4856 34932 4862 34944
rect 5074 34932 5080 34944
rect 5132 34941 5138 34944
rect 5132 34935 5151 34941
rect 4856 34904 5080 34932
rect 4856 34892 4862 34904
rect 5074 34892 5080 34904
rect 5139 34901 5151 34935
rect 5132 34895 5151 34901
rect 5261 34935 5319 34941
rect 5261 34901 5273 34935
rect 5307 34932 5319 34935
rect 5350 34932 5356 34944
rect 5307 34904 5356 34932
rect 5307 34901 5319 34904
rect 5261 34895 5319 34901
rect 5132 34892 5138 34895
rect 5350 34892 5356 34904
rect 5408 34892 5414 34944
rect 5460 34932 5488 35040
rect 5534 35028 5540 35080
rect 5592 35028 5598 35080
rect 5902 35028 5908 35080
rect 5960 35028 5966 35080
rect 6641 35071 6699 35077
rect 6641 35037 6653 35071
rect 6687 35068 6699 35071
rect 6730 35068 6736 35080
rect 6687 35040 6736 35068
rect 6687 35037 6699 35040
rect 6641 35031 6699 35037
rect 6730 35028 6736 35040
rect 6788 35028 6794 35080
rect 6822 35028 6828 35080
rect 6880 35028 6886 35080
rect 7466 35028 7472 35080
rect 7524 35028 7530 35080
rect 7653 35071 7711 35077
rect 7653 35037 7665 35071
rect 7699 35068 7711 35071
rect 7834 35068 7840 35080
rect 7699 35040 7840 35068
rect 7699 35037 7711 35040
rect 7653 35031 7711 35037
rect 7834 35028 7840 35040
rect 7892 35028 7898 35080
rect 6917 35003 6975 35009
rect 6917 34969 6929 35003
rect 6963 35000 6975 35003
rect 7282 35000 7288 35012
rect 6963 34972 7288 35000
rect 6963 34969 6975 34972
rect 6917 34963 6975 34969
rect 7282 34960 7288 34972
rect 7340 34960 7346 35012
rect 7742 34960 7748 35012
rect 7800 34960 7806 35012
rect 7944 35000 7972 35108
rect 8202 35028 8208 35080
rect 8260 35028 8266 35080
rect 8386 35028 8392 35080
rect 8444 35028 8450 35080
rect 9416 35068 9444 35176
rect 9582 35096 9588 35148
rect 9640 35096 9646 35148
rect 9677 35139 9735 35145
rect 9677 35105 9689 35139
rect 9723 35105 9735 35139
rect 9677 35099 9735 35105
rect 8496 35040 9444 35068
rect 8496 35000 8524 35040
rect 9490 35028 9496 35080
rect 9548 35068 9554 35080
rect 9692 35068 9720 35099
rect 10042 35096 10048 35148
rect 10100 35136 10106 35148
rect 10873 35139 10931 35145
rect 10873 35136 10885 35139
rect 10100 35108 10885 35136
rect 10100 35096 10106 35108
rect 10873 35105 10885 35108
rect 10919 35136 10931 35139
rect 11146 35136 11152 35148
rect 10919 35108 11152 35136
rect 10919 35105 10931 35108
rect 10873 35099 10931 35105
rect 11146 35096 11152 35108
rect 11204 35096 11210 35148
rect 11532 35136 11560 35176
rect 13078 35164 13084 35216
rect 13136 35204 13142 35216
rect 13136 35176 14596 35204
rect 13136 35164 13142 35176
rect 12710 35136 12716 35148
rect 11532 35108 12716 35136
rect 9548 35040 9720 35068
rect 9548 35028 9554 35040
rect 9766 35028 9772 35080
rect 9824 35068 9830 35080
rect 10318 35068 10324 35080
rect 9824 35040 10324 35068
rect 9824 35028 9830 35040
rect 10318 35028 10324 35040
rect 10376 35028 10382 35080
rect 10410 35028 10416 35080
rect 10468 35028 10474 35080
rect 11532 35077 11560 35108
rect 12710 35096 12716 35108
rect 12768 35096 12774 35148
rect 14568 35136 14596 35176
rect 14642 35164 14648 35216
rect 14700 35204 14706 35216
rect 18616 35204 18644 35244
rect 20346 35232 20352 35244
rect 20404 35232 20410 35284
rect 20530 35232 20536 35284
rect 20588 35272 20594 35284
rect 25866 35272 25872 35284
rect 20588 35244 25872 35272
rect 20588 35232 20594 35244
rect 25866 35232 25872 35244
rect 25924 35232 25930 35284
rect 26786 35232 26792 35284
rect 26844 35232 26850 35284
rect 27154 35232 27160 35284
rect 27212 35272 27218 35284
rect 27249 35275 27307 35281
rect 27249 35272 27261 35275
rect 27212 35244 27261 35272
rect 27212 35232 27218 35244
rect 27249 35241 27261 35244
rect 27295 35241 27307 35275
rect 27249 35235 27307 35241
rect 28442 35232 28448 35284
rect 28500 35272 28506 35284
rect 30239 35275 30297 35281
rect 30239 35272 30251 35275
rect 28500 35244 30251 35272
rect 28500 35232 28506 35244
rect 30239 35241 30251 35244
rect 30285 35241 30297 35275
rect 30239 35235 30297 35241
rect 32122 35232 32128 35284
rect 32180 35272 32186 35284
rect 32950 35272 32956 35284
rect 32180 35244 32956 35272
rect 32180 35232 32186 35244
rect 32950 35232 32956 35244
rect 33008 35232 33014 35284
rect 33045 35275 33103 35281
rect 33045 35241 33057 35275
rect 33091 35241 33103 35275
rect 33045 35235 33103 35241
rect 33229 35275 33287 35281
rect 33229 35241 33241 35275
rect 33275 35272 33287 35275
rect 34514 35272 34520 35284
rect 33275 35244 34520 35272
rect 33275 35241 33287 35244
rect 33229 35235 33287 35241
rect 14700 35176 18644 35204
rect 18877 35207 18935 35213
rect 14700 35164 14706 35176
rect 18877 35173 18889 35207
rect 18923 35204 18935 35207
rect 19978 35204 19984 35216
rect 18923 35176 19984 35204
rect 18923 35173 18935 35176
rect 18877 35167 18935 35173
rect 19978 35164 19984 35176
rect 20036 35204 20042 35216
rect 20898 35204 20904 35216
rect 20036 35176 20904 35204
rect 20036 35164 20042 35176
rect 20898 35164 20904 35176
rect 20956 35164 20962 35216
rect 21450 35164 21456 35216
rect 21508 35204 21514 35216
rect 23842 35204 23848 35216
rect 21508 35176 23848 35204
rect 21508 35164 21514 35176
rect 23842 35164 23848 35176
rect 23900 35164 23906 35216
rect 25130 35164 25136 35216
rect 25188 35164 25194 35216
rect 26053 35207 26111 35213
rect 26053 35173 26065 35207
rect 26099 35173 26111 35207
rect 26053 35167 26111 35173
rect 28077 35207 28135 35213
rect 28077 35173 28089 35207
rect 28123 35204 28135 35207
rect 28258 35204 28264 35216
rect 28123 35176 28264 35204
rect 28123 35173 28135 35176
rect 28077 35167 28135 35173
rect 14568 35108 14688 35136
rect 11517 35071 11575 35077
rect 11517 35037 11529 35071
rect 11563 35037 11575 35071
rect 11517 35031 11575 35037
rect 12158 35028 12164 35080
rect 12216 35068 12222 35080
rect 12345 35071 12403 35077
rect 12345 35068 12357 35071
rect 12216 35040 12357 35068
rect 12216 35028 12222 35040
rect 12345 35037 12357 35040
rect 12391 35037 12403 35071
rect 12345 35031 12403 35037
rect 13262 35028 13268 35080
rect 13320 35028 13326 35080
rect 13541 35071 13599 35077
rect 13541 35037 13553 35071
rect 13587 35068 13599 35071
rect 14550 35068 14556 35080
rect 13587 35040 14556 35068
rect 13587 35037 13599 35040
rect 13541 35031 13599 35037
rect 14550 35028 14556 35040
rect 14608 35028 14614 35080
rect 14660 35068 14688 35108
rect 14826 35096 14832 35148
rect 14884 35136 14890 35148
rect 17126 35136 17132 35148
rect 14884 35108 17132 35136
rect 14884 35096 14890 35108
rect 17126 35096 17132 35108
rect 17184 35096 17190 35148
rect 17402 35096 17408 35148
rect 17460 35136 17466 35148
rect 17865 35139 17923 35145
rect 17865 35136 17877 35139
rect 17460 35108 17877 35136
rect 17460 35096 17466 35108
rect 17865 35105 17877 35108
rect 17911 35105 17923 35139
rect 17865 35099 17923 35105
rect 18049 35139 18107 35145
rect 18049 35105 18061 35139
rect 18095 35136 18107 35139
rect 18690 35136 18696 35148
rect 18095 35108 18696 35136
rect 18095 35105 18107 35108
rect 18049 35099 18107 35105
rect 18690 35096 18696 35108
rect 18748 35096 18754 35148
rect 21266 35136 21272 35148
rect 19306 35108 21272 35136
rect 15473 35071 15531 35077
rect 15473 35068 15485 35071
rect 14660 35040 15485 35068
rect 15473 35037 15485 35040
rect 15519 35037 15531 35071
rect 15473 35031 15531 35037
rect 9674 35000 9680 35012
rect 7944 34972 8524 35000
rect 8588 34972 9680 35000
rect 5994 34932 6000 34944
rect 5460 34904 6000 34932
rect 5994 34892 6000 34904
rect 6052 34892 6058 34944
rect 6086 34892 6092 34944
rect 6144 34892 6150 34944
rect 6546 34892 6552 34944
rect 6604 34932 6610 34944
rect 7190 34932 7196 34944
rect 6604 34904 7196 34932
rect 6604 34892 6610 34904
rect 7190 34892 7196 34904
rect 7248 34892 7254 34944
rect 8588 34941 8616 34972
rect 9674 34960 9680 34972
rect 9732 34960 9738 35012
rect 12618 35000 12624 35012
rect 10980 34972 12624 35000
rect 8573 34935 8631 34941
rect 8573 34901 8585 34935
rect 8619 34901 8631 34935
rect 8573 34895 8631 34901
rect 9398 34892 9404 34944
rect 9456 34932 9462 34944
rect 9493 34935 9551 34941
rect 9493 34932 9505 34935
rect 9456 34904 9505 34932
rect 9456 34892 9462 34904
rect 9493 34901 9505 34904
rect 9539 34901 9551 34935
rect 9493 34895 9551 34901
rect 9582 34892 9588 34944
rect 9640 34932 9646 34944
rect 10980 34932 11008 34972
rect 12618 34960 12624 34972
rect 12676 34960 12682 35012
rect 14369 35003 14427 35009
rect 14369 34969 14381 35003
rect 14415 34969 14427 35003
rect 15488 35000 15516 35031
rect 15562 35028 15568 35080
rect 15620 35068 15626 35080
rect 15657 35071 15715 35077
rect 15657 35068 15669 35071
rect 15620 35040 15669 35068
rect 15620 35028 15626 35040
rect 15657 35037 15669 35040
rect 15703 35037 15715 35071
rect 15657 35031 15715 35037
rect 15749 35071 15807 35077
rect 15749 35037 15761 35071
rect 15795 35068 15807 35071
rect 16114 35068 16120 35080
rect 15795 35040 16120 35068
rect 15795 35037 15807 35040
rect 15749 35031 15807 35037
rect 16114 35028 16120 35040
rect 16172 35028 16178 35080
rect 17037 35071 17095 35077
rect 17037 35037 17049 35071
rect 17083 35068 17095 35071
rect 17310 35068 17316 35080
rect 17083 35040 17316 35068
rect 17083 35037 17095 35040
rect 17037 35031 17095 35037
rect 17310 35028 17316 35040
rect 17368 35028 17374 35080
rect 17773 35071 17831 35077
rect 17773 35037 17785 35071
rect 17819 35068 17831 35071
rect 18322 35068 18328 35080
rect 17819 35040 18328 35068
rect 17819 35037 17831 35040
rect 17773 35031 17831 35037
rect 18322 35028 18328 35040
rect 18380 35028 18386 35080
rect 18509 35071 18567 35077
rect 18509 35037 18521 35071
rect 18555 35037 18567 35071
rect 18509 35031 18567 35037
rect 18601 35071 18659 35077
rect 18601 35037 18613 35071
rect 18647 35068 18659 35071
rect 19306 35068 19334 35108
rect 21266 35096 21272 35108
rect 21324 35096 21330 35148
rect 23382 35096 23388 35148
rect 23440 35136 23446 35148
rect 23661 35139 23719 35145
rect 23661 35136 23673 35139
rect 23440 35108 23673 35136
rect 23440 35096 23446 35108
rect 23661 35105 23673 35108
rect 23707 35136 23719 35139
rect 24673 35139 24731 35145
rect 24673 35136 24685 35139
rect 23707 35108 24685 35136
rect 23707 35105 23719 35108
rect 23661 35099 23719 35105
rect 24673 35105 24685 35108
rect 24719 35136 24731 35139
rect 24719 35108 25176 35136
rect 24719 35105 24731 35108
rect 24673 35099 24731 35105
rect 18647 35040 19334 35068
rect 18647 35037 18659 35040
rect 18601 35031 18659 35037
rect 16850 35000 16856 35012
rect 15488 34972 16856 35000
rect 14369 34963 14427 34969
rect 9640 34904 11008 34932
rect 9640 34892 9646 34904
rect 11606 34892 11612 34944
rect 11664 34932 11670 34944
rect 14090 34932 14096 34944
rect 11664 34904 14096 34932
rect 11664 34892 11670 34904
rect 14090 34892 14096 34904
rect 14148 34932 14154 34944
rect 14384 34932 14412 34963
rect 16850 34960 16856 34972
rect 16908 34960 16914 35012
rect 16945 35003 17003 35009
rect 16945 34969 16957 35003
rect 16991 35000 17003 35003
rect 17954 35000 17960 35012
rect 16991 34972 17960 35000
rect 16991 34969 17003 34972
rect 16945 34963 17003 34969
rect 17954 34960 17960 34972
rect 18012 34960 18018 35012
rect 18524 35000 18552 35031
rect 19610 35028 19616 35080
rect 19668 35028 19674 35080
rect 19978 35028 19984 35080
rect 20036 35068 20042 35080
rect 20438 35068 20444 35080
rect 20036 35040 20444 35068
rect 20036 35028 20042 35040
rect 20438 35028 20444 35040
rect 20496 35028 20502 35080
rect 20622 35028 20628 35080
rect 20680 35028 20686 35080
rect 20714 35028 20720 35080
rect 20772 35028 20778 35080
rect 20806 35028 20812 35080
rect 20864 35028 20870 35080
rect 21361 35071 21419 35077
rect 21361 35037 21373 35071
rect 21407 35068 21419 35071
rect 21634 35068 21640 35080
rect 21407 35040 21640 35068
rect 21407 35037 21419 35040
rect 21361 35031 21419 35037
rect 21634 35028 21640 35040
rect 21692 35028 21698 35080
rect 22554 35028 22560 35080
rect 22612 35028 22618 35080
rect 23474 35028 23480 35080
rect 23532 35028 23538 35080
rect 23750 35028 23756 35080
rect 23808 35068 23814 35080
rect 24765 35071 24823 35077
rect 24765 35068 24777 35071
rect 23808 35040 24777 35068
rect 23808 35028 23814 35040
rect 24765 35037 24777 35040
rect 24811 35068 24823 35071
rect 25038 35068 25044 35080
rect 24811 35040 25044 35068
rect 24811 35037 24823 35040
rect 24765 35031 24823 35037
rect 25038 35028 25044 35040
rect 25096 35028 25102 35080
rect 25148 35068 25176 35108
rect 25222 35096 25228 35148
rect 25280 35096 25286 35148
rect 25498 35096 25504 35148
rect 25556 35136 25562 35148
rect 26068 35136 26096 35167
rect 28258 35164 28264 35176
rect 28316 35164 28322 35216
rect 28537 35207 28595 35213
rect 28537 35173 28549 35207
rect 28583 35204 28595 35207
rect 28994 35204 29000 35216
rect 28583 35176 29000 35204
rect 28583 35173 28595 35176
rect 28537 35167 28595 35173
rect 28994 35164 29000 35176
rect 29052 35204 29058 35216
rect 30377 35207 30435 35213
rect 30377 35204 30389 35207
rect 29052 35176 30389 35204
rect 29052 35164 29058 35176
rect 30377 35173 30389 35176
rect 30423 35173 30435 35207
rect 33060 35204 33088 35235
rect 34514 35232 34520 35244
rect 34572 35232 34578 35284
rect 34790 35232 34796 35284
rect 34848 35272 34854 35284
rect 37274 35272 37280 35284
rect 34848 35244 37280 35272
rect 34848 35232 34854 35244
rect 37274 35232 37280 35244
rect 37332 35232 37338 35284
rect 34054 35204 34060 35216
rect 33060 35176 34060 35204
rect 30377 35167 30435 35173
rect 34054 35164 34060 35176
rect 34112 35164 34118 35216
rect 36630 35164 36636 35216
rect 36688 35204 36694 35216
rect 37734 35204 37740 35216
rect 36688 35176 37740 35204
rect 36688 35164 36694 35176
rect 37734 35164 37740 35176
rect 37792 35164 37798 35216
rect 27246 35136 27252 35148
rect 25556 35108 26096 35136
rect 26252 35108 27252 35136
rect 25556 35096 25562 35108
rect 26252 35068 26280 35108
rect 27246 35096 27252 35108
rect 27304 35136 27310 35148
rect 28626 35136 28632 35148
rect 27304 35108 28632 35136
rect 27304 35096 27310 35108
rect 28626 35096 28632 35108
rect 28684 35096 28690 35148
rect 29178 35136 29184 35148
rect 28966 35108 29184 35136
rect 25148 35040 26280 35068
rect 26326 35028 26332 35080
rect 26384 35028 26390 35080
rect 26878 35028 26884 35080
rect 26936 35068 26942 35080
rect 26973 35071 27031 35077
rect 26973 35068 26985 35071
rect 26936 35040 26985 35068
rect 26936 35028 26942 35040
rect 26973 35037 26985 35040
rect 27019 35037 27031 35071
rect 26973 35031 27031 35037
rect 27062 35028 27068 35080
rect 27120 35028 27126 35080
rect 28966 35068 28994 35108
rect 29178 35096 29184 35108
rect 29236 35096 29242 35148
rect 29914 35096 29920 35148
rect 29972 35136 29978 35148
rect 30469 35139 30527 35145
rect 30469 35136 30481 35139
rect 29972 35108 30481 35136
rect 29972 35096 29978 35108
rect 30469 35105 30481 35108
rect 30515 35105 30527 35139
rect 30469 35099 30527 35105
rect 31846 35096 31852 35148
rect 31904 35136 31910 35148
rect 32398 35136 32404 35148
rect 31904 35108 32404 35136
rect 31904 35096 31910 35108
rect 32398 35096 32404 35108
rect 32456 35096 32462 35148
rect 33870 35096 33876 35148
rect 33928 35096 33934 35148
rect 34333 35139 34391 35145
rect 34333 35105 34345 35139
rect 34379 35105 34391 35139
rect 34333 35099 34391 35105
rect 27172 35040 28994 35068
rect 19334 35000 19340 35012
rect 18524 34972 19340 35000
rect 19334 34960 19340 34972
rect 19392 34960 19398 35012
rect 19426 34960 19432 35012
rect 19484 34960 19490 35012
rect 21082 35000 21088 35012
rect 20364 34972 21088 35000
rect 14148 34904 14412 34932
rect 15289 34935 15347 34941
rect 14148 34892 14154 34904
rect 15289 34901 15301 34935
rect 15335 34932 15347 34935
rect 15654 34932 15660 34944
rect 15335 34904 15660 34932
rect 15335 34901 15347 34904
rect 15289 34895 15347 34901
rect 15654 34892 15660 34904
rect 15712 34892 15718 34944
rect 18049 34935 18107 34941
rect 18049 34901 18061 34935
rect 18095 34932 18107 34935
rect 20364 34932 20392 34972
rect 21082 34960 21088 34972
rect 21140 34960 21146 35012
rect 21913 35003 21971 35009
rect 21913 34969 21925 35003
rect 21959 34969 21971 35003
rect 21913 34963 21971 34969
rect 18095 34904 20392 34932
rect 18095 34901 18107 34904
rect 18049 34895 18107 34901
rect 20438 34892 20444 34944
rect 20496 34892 20502 34944
rect 20714 34892 20720 34944
rect 20772 34932 20778 34944
rect 21726 34932 21732 34944
rect 20772 34904 21732 34932
rect 20772 34892 20778 34904
rect 21726 34892 21732 34904
rect 21784 34892 21790 34944
rect 21928 34932 21956 34963
rect 22462 34960 22468 35012
rect 22520 35000 22526 35012
rect 22833 35003 22891 35009
rect 22833 35000 22845 35003
rect 22520 34972 22845 35000
rect 22520 34960 22526 34972
rect 22833 34969 22845 34972
rect 22879 35000 22891 35003
rect 24026 35000 24032 35012
rect 22879 34972 24032 35000
rect 22879 34969 22891 34972
rect 22833 34963 22891 34969
rect 24026 34960 24032 34972
rect 24084 34960 24090 35012
rect 24670 34960 24676 35012
rect 24728 35000 24734 35012
rect 25406 35000 25412 35012
rect 24728 34972 25412 35000
rect 24728 34960 24734 34972
rect 25406 34960 25412 34972
rect 25464 35000 25470 35012
rect 25593 35003 25651 35009
rect 25593 35000 25605 35003
rect 25464 34972 25605 35000
rect 25464 34960 25470 34972
rect 25593 34969 25605 34972
rect 25639 34969 25651 35003
rect 25593 34963 25651 34969
rect 25866 34960 25872 35012
rect 25924 35000 25930 35012
rect 26053 35003 26111 35009
rect 26053 35000 26065 35003
rect 25924 34972 26065 35000
rect 25924 34960 25930 34972
rect 26053 34969 26065 34972
rect 26099 34969 26111 35003
rect 27172 35000 27200 35040
rect 29270 35028 29276 35080
rect 29328 35068 29334 35080
rect 31478 35068 31484 35080
rect 29328 35040 31484 35068
rect 29328 35028 29334 35040
rect 31478 35028 31484 35040
rect 31536 35028 31542 35080
rect 32766 35028 32772 35080
rect 32824 35068 32830 35080
rect 33965 35071 34023 35077
rect 33965 35068 33977 35071
rect 32824 35040 33977 35068
rect 32824 35028 32830 35040
rect 33965 35037 33977 35040
rect 34011 35037 34023 35071
rect 33965 35031 34023 35037
rect 26053 34963 26111 34969
rect 26160 34972 27200 35000
rect 22554 34932 22560 34944
rect 21928 34904 22560 34932
rect 22554 34892 22560 34904
rect 22612 34892 22618 34944
rect 25130 34892 25136 34944
rect 25188 34932 25194 34944
rect 25682 34932 25688 34944
rect 25188 34904 25688 34932
rect 25188 34892 25194 34904
rect 25682 34892 25688 34904
rect 25740 34932 25746 34944
rect 26160 34932 26188 34972
rect 27246 34960 27252 35012
rect 27304 35000 27310 35012
rect 27304 34972 29040 35000
rect 27304 34960 27310 34972
rect 25740 34904 26188 34932
rect 26237 34935 26295 34941
rect 25740 34892 25746 34904
rect 26237 34901 26249 34935
rect 26283 34932 26295 34935
rect 26326 34932 26332 34944
rect 26283 34904 26332 34932
rect 26283 34901 26295 34904
rect 26237 34895 26295 34901
rect 26326 34892 26332 34904
rect 26384 34892 26390 34944
rect 27798 34892 27804 34944
rect 27856 34932 27862 34944
rect 28810 34932 28816 34944
rect 27856 34904 28816 34932
rect 27856 34892 27862 34904
rect 28810 34892 28816 34904
rect 28868 34932 28874 34944
rect 28905 34935 28963 34941
rect 28905 34932 28917 34935
rect 28868 34904 28917 34932
rect 28868 34892 28874 34904
rect 28905 34901 28917 34904
rect 28951 34901 28963 34935
rect 29012 34932 29040 34972
rect 29178 34960 29184 35012
rect 29236 35000 29242 35012
rect 30098 35000 30104 35012
rect 29236 34972 30104 35000
rect 29236 34960 29242 34972
rect 30098 34960 30104 34972
rect 30156 34960 30162 35012
rect 30668 34972 30880 35000
rect 30668 34932 30696 34972
rect 29012 34904 30696 34932
rect 28905 34895 28963 34901
rect 30742 34892 30748 34944
rect 30800 34892 30806 34944
rect 30852 34932 30880 34972
rect 31294 34960 31300 35012
rect 31352 34960 31358 35012
rect 32674 34960 32680 35012
rect 32732 35000 32738 35012
rect 32861 35003 32919 35009
rect 32861 35000 32873 35003
rect 32732 34972 32873 35000
rect 32732 34960 32738 34972
rect 32861 34969 32873 34972
rect 32907 34969 32919 35003
rect 34348 35000 34376 35099
rect 34698 35096 34704 35148
rect 34756 35136 34762 35148
rect 34756 35108 35112 35136
rect 34756 35096 34762 35108
rect 34422 35028 34428 35080
rect 34480 35068 34486 35080
rect 35084 35077 35112 35108
rect 36538 35096 36544 35148
rect 36596 35136 36602 35148
rect 38378 35136 38384 35148
rect 36596 35108 38384 35136
rect 36596 35096 36602 35108
rect 38378 35096 38384 35108
rect 38436 35096 38442 35148
rect 34885 35071 34943 35077
rect 34885 35068 34897 35071
rect 34480 35040 34897 35068
rect 34480 35028 34486 35040
rect 34885 35037 34897 35040
rect 34931 35037 34943 35071
rect 34885 35031 34943 35037
rect 35069 35071 35127 35077
rect 35069 35037 35081 35071
rect 35115 35037 35127 35071
rect 35069 35031 35127 35037
rect 35250 35028 35256 35080
rect 35308 35068 35314 35080
rect 35434 35068 35440 35080
rect 35308 35040 35440 35068
rect 35308 35028 35314 35040
rect 35434 35028 35440 35040
rect 35492 35028 35498 35080
rect 35529 35071 35587 35077
rect 35529 35037 35541 35071
rect 35575 35068 35587 35071
rect 36078 35068 36084 35080
rect 35575 35040 36084 35068
rect 35575 35037 35587 35040
rect 35529 35031 35587 35037
rect 36078 35028 36084 35040
rect 36136 35028 36142 35080
rect 36170 35028 36176 35080
rect 36228 35068 36234 35080
rect 37366 35068 37372 35080
rect 36228 35040 37372 35068
rect 36228 35028 36234 35040
rect 37366 35028 37372 35040
rect 37424 35028 37430 35080
rect 37458 35028 37464 35080
rect 37516 35028 37522 35080
rect 37737 35071 37795 35077
rect 37737 35068 37749 35071
rect 37568 35040 37749 35068
rect 35774 35003 35832 35009
rect 35774 35000 35786 35003
rect 32861 34963 32919 34969
rect 32968 34972 34284 35000
rect 34348 34972 35786 35000
rect 32968 34932 32996 34972
rect 30852 34904 32996 34932
rect 33042 34892 33048 34944
rect 33100 34892 33106 34944
rect 34256 34932 34284 34972
rect 35774 34969 35786 34972
rect 35820 34969 35832 35003
rect 35774 34963 35832 34969
rect 36722 34960 36728 35012
rect 36780 35000 36786 35012
rect 37568 35000 37596 35040
rect 37737 35037 37749 35040
rect 37783 35037 37795 35071
rect 37737 35031 37795 35037
rect 37829 35071 37887 35077
rect 37829 35037 37841 35071
rect 37875 35068 37887 35071
rect 37918 35068 37924 35080
rect 37875 35040 37924 35068
rect 37875 35037 37887 35040
rect 37829 35031 37887 35037
rect 37918 35028 37924 35040
rect 37976 35028 37982 35080
rect 36780 34972 37596 35000
rect 36780 34960 36786 34972
rect 37642 34960 37648 35012
rect 37700 34960 37706 35012
rect 34974 34932 34980 34944
rect 34256 34904 34980 34932
rect 34974 34892 34980 34904
rect 35032 34892 35038 34944
rect 35066 34892 35072 34944
rect 35124 34892 35130 34944
rect 36814 34892 36820 34944
rect 36872 34932 36878 34944
rect 36909 34935 36967 34941
rect 36909 34932 36921 34935
rect 36872 34904 36921 34932
rect 36872 34892 36878 34904
rect 36909 34901 36921 34904
rect 36955 34901 36967 34935
rect 36909 34895 36967 34901
rect 37366 34892 37372 34944
rect 37424 34932 37430 34944
rect 38013 34935 38071 34941
rect 38013 34932 38025 34935
rect 37424 34904 38025 34932
rect 37424 34892 37430 34904
rect 38013 34901 38025 34904
rect 38059 34901 38071 34935
rect 38013 34895 38071 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 3602 34688 3608 34740
rect 3660 34688 3666 34740
rect 4341 34731 4399 34737
rect 4341 34697 4353 34731
rect 4387 34728 4399 34731
rect 4890 34728 4896 34740
rect 4387 34700 4896 34728
rect 4387 34697 4399 34700
rect 4341 34691 4399 34697
rect 4890 34688 4896 34700
rect 4948 34688 4954 34740
rect 5166 34688 5172 34740
rect 5224 34728 5230 34740
rect 6546 34728 6552 34740
rect 5224 34700 6552 34728
rect 5224 34688 5230 34700
rect 6546 34688 6552 34700
rect 6604 34688 6610 34740
rect 11974 34728 11980 34740
rect 6656 34700 11980 34728
rect 5902 34660 5908 34672
rect 5000 34632 5908 34660
rect 3237 34595 3295 34601
rect 3237 34561 3249 34595
rect 3283 34592 3295 34595
rect 3510 34592 3516 34604
rect 3283 34564 3516 34592
rect 3283 34561 3295 34564
rect 3237 34555 3295 34561
rect 3510 34552 3516 34564
rect 3568 34552 3574 34604
rect 4154 34552 4160 34604
rect 4212 34552 4218 34604
rect 4341 34595 4399 34601
rect 4341 34561 4353 34595
rect 4387 34592 4399 34595
rect 4893 34598 4951 34601
rect 5000 34598 5028 34632
rect 5902 34620 5908 34632
rect 5960 34620 5966 34672
rect 4893 34595 5028 34598
rect 4387 34564 4568 34592
rect 4387 34561 4399 34564
rect 4341 34555 4399 34561
rect 4540 34456 4568 34564
rect 4893 34561 4905 34595
rect 4939 34570 5028 34595
rect 5077 34595 5135 34601
rect 4939 34561 4951 34570
rect 4893 34555 4951 34561
rect 5077 34561 5089 34595
rect 5123 34592 5135 34595
rect 5534 34592 5540 34604
rect 5123 34564 5540 34592
rect 5123 34561 5135 34564
rect 5077 34555 5135 34561
rect 5092 34456 5120 34555
rect 5534 34552 5540 34564
rect 5592 34552 5598 34604
rect 5718 34552 5724 34604
rect 5776 34552 5782 34604
rect 6656 34601 6684 34700
rect 11974 34688 11980 34700
rect 12032 34728 12038 34740
rect 14645 34731 14703 34737
rect 12032 34700 14412 34728
rect 12032 34688 12038 34700
rect 7190 34620 7196 34672
rect 7248 34660 7254 34672
rect 11701 34663 11759 34669
rect 7248 34632 10180 34660
rect 7248 34620 7254 34632
rect 5813 34595 5871 34601
rect 5813 34561 5825 34595
rect 5859 34592 5871 34595
rect 6641 34595 6699 34601
rect 5859 34564 6592 34592
rect 5859 34561 5871 34564
rect 5813 34555 5871 34561
rect 5169 34527 5227 34533
rect 5169 34493 5181 34527
rect 5215 34524 5227 34527
rect 5828 34524 5856 34555
rect 5215 34496 5856 34524
rect 5215 34493 5227 34496
rect 5169 34487 5227 34493
rect 5902 34484 5908 34536
rect 5960 34484 5966 34536
rect 6564 34524 6592 34564
rect 6641 34561 6653 34595
rect 6687 34561 6699 34595
rect 6641 34555 6699 34561
rect 6825 34595 6883 34601
rect 6825 34561 6837 34595
rect 6871 34592 6883 34595
rect 6914 34592 6920 34604
rect 6871 34564 6920 34592
rect 6871 34561 6883 34564
rect 6825 34555 6883 34561
rect 6914 34552 6920 34564
rect 6972 34552 6978 34604
rect 7006 34552 7012 34604
rect 7064 34592 7070 34604
rect 7377 34595 7435 34601
rect 7377 34592 7389 34595
rect 7064 34564 7389 34592
rect 7064 34552 7070 34564
rect 7377 34561 7389 34564
rect 7423 34561 7435 34595
rect 7561 34595 7619 34601
rect 7561 34592 7573 34595
rect 7377 34555 7435 34561
rect 7475 34564 7573 34592
rect 7190 34524 7196 34536
rect 6564 34496 7196 34524
rect 7190 34484 7196 34496
rect 7248 34484 7254 34536
rect 7475 34524 7503 34564
rect 7561 34561 7573 34564
rect 7607 34561 7619 34595
rect 7561 34555 7619 34561
rect 7834 34552 7840 34604
rect 7892 34592 7898 34604
rect 8018 34592 8024 34604
rect 7892 34564 8024 34592
rect 7892 34552 7898 34564
rect 8018 34552 8024 34564
rect 8076 34592 8082 34604
rect 8205 34595 8263 34601
rect 8205 34592 8217 34595
rect 8076 34564 8217 34592
rect 8076 34552 8082 34564
rect 8205 34561 8217 34564
rect 8251 34561 8263 34595
rect 8205 34555 8263 34561
rect 8389 34595 8447 34601
rect 8389 34561 8401 34595
rect 8435 34561 8447 34595
rect 8389 34555 8447 34561
rect 8404 34524 8432 34555
rect 9030 34552 9036 34604
rect 9088 34592 9094 34604
rect 9309 34595 9367 34601
rect 9309 34592 9321 34595
rect 9088 34564 9321 34592
rect 9088 34552 9094 34564
rect 9309 34561 9321 34564
rect 9355 34561 9367 34595
rect 9309 34555 9367 34561
rect 9398 34552 9404 34604
rect 9456 34592 9462 34604
rect 9493 34595 9551 34601
rect 9493 34592 9505 34595
rect 9456 34564 9505 34592
rect 9456 34552 9462 34564
rect 9493 34561 9505 34564
rect 9539 34592 9551 34595
rect 9539 34564 9996 34592
rect 9539 34561 9551 34564
rect 9493 34555 9551 34561
rect 9125 34527 9183 34533
rect 7300 34496 8984 34524
rect 4540 34428 5120 34456
rect 5534 34416 5540 34468
rect 5592 34456 5598 34468
rect 6641 34459 6699 34465
rect 6641 34456 6653 34459
rect 5592 34428 6653 34456
rect 5592 34416 5598 34428
rect 6641 34425 6653 34428
rect 6687 34456 6699 34459
rect 7300 34456 7328 34496
rect 6687 34428 7328 34456
rect 6687 34425 6699 34428
rect 6641 34419 6699 34425
rect 7374 34416 7380 34468
rect 7432 34456 7438 34468
rect 7558 34456 7564 34468
rect 7432 34428 7564 34456
rect 7432 34416 7438 34428
rect 7558 34416 7564 34428
rect 7616 34416 7622 34468
rect 8570 34416 8576 34468
rect 8628 34416 8634 34468
rect 8956 34456 8984 34496
rect 9125 34493 9137 34527
rect 9171 34524 9183 34527
rect 9766 34524 9772 34536
rect 9171 34496 9772 34524
rect 9171 34493 9183 34496
rect 9125 34487 9183 34493
rect 9766 34484 9772 34496
rect 9824 34484 9830 34536
rect 9968 34524 9996 34564
rect 10042 34552 10048 34604
rect 10100 34552 10106 34604
rect 10152 34601 10180 34632
rect 11701 34629 11713 34663
rect 11747 34660 11759 34663
rect 14274 34660 14280 34672
rect 11747 34632 14280 34660
rect 11747 34629 11759 34632
rect 11701 34623 11759 34629
rect 14274 34620 14280 34632
rect 14332 34620 14338 34672
rect 14384 34604 14412 34700
rect 14645 34697 14657 34731
rect 14691 34728 14703 34731
rect 15194 34728 15200 34740
rect 14691 34700 15200 34728
rect 14691 34697 14703 34700
rect 14645 34691 14703 34697
rect 15194 34688 15200 34700
rect 15252 34688 15258 34740
rect 15470 34688 15476 34740
rect 15528 34688 15534 34740
rect 17126 34688 17132 34740
rect 17184 34728 17190 34740
rect 19886 34728 19892 34740
rect 17184 34700 19892 34728
rect 17184 34688 17190 34700
rect 19886 34688 19892 34700
rect 19944 34688 19950 34740
rect 19981 34731 20039 34737
rect 19981 34697 19993 34731
rect 20027 34728 20039 34731
rect 20070 34728 20076 34740
rect 20027 34700 20076 34728
rect 20027 34697 20039 34700
rect 19981 34691 20039 34697
rect 20070 34688 20076 34700
rect 20128 34688 20134 34740
rect 20898 34688 20904 34740
rect 20956 34688 20962 34740
rect 21085 34731 21143 34737
rect 21085 34697 21097 34731
rect 21131 34728 21143 34731
rect 21174 34728 21180 34740
rect 21131 34700 21180 34728
rect 21131 34697 21143 34700
rect 21085 34691 21143 34697
rect 21174 34688 21180 34700
rect 21232 34688 21238 34740
rect 22646 34688 22652 34740
rect 22704 34688 22710 34740
rect 23842 34688 23848 34740
rect 23900 34728 23906 34740
rect 31846 34728 31852 34740
rect 23900 34700 31852 34728
rect 23900 34688 23906 34700
rect 20438 34660 20444 34672
rect 14752 34632 17356 34660
rect 10137 34595 10195 34601
rect 10137 34561 10149 34595
rect 10183 34592 10195 34595
rect 10318 34592 10324 34604
rect 10183 34564 10324 34592
rect 10183 34561 10195 34564
rect 10137 34555 10195 34561
rect 10318 34552 10324 34564
rect 10376 34552 10382 34604
rect 11885 34595 11943 34601
rect 11885 34561 11897 34595
rect 11931 34592 11943 34595
rect 11974 34592 11980 34604
rect 11931 34564 11980 34592
rect 11931 34561 11943 34564
rect 11885 34555 11943 34561
rect 11900 34524 11928 34555
rect 11974 34552 11980 34564
rect 12032 34552 12038 34604
rect 12158 34552 12164 34604
rect 12216 34552 12222 34604
rect 13449 34595 13507 34601
rect 13449 34561 13461 34595
rect 13495 34592 13507 34595
rect 13998 34592 14004 34604
rect 13495 34564 14004 34592
rect 13495 34561 13507 34564
rect 13449 34555 13507 34561
rect 13998 34552 14004 34564
rect 14056 34592 14062 34604
rect 14056 34564 14136 34592
rect 14056 34552 14062 34564
rect 9968 34496 11928 34524
rect 12434 34484 12440 34536
rect 12492 34524 12498 34536
rect 13725 34527 13783 34533
rect 13725 34524 13737 34527
rect 12492 34496 13737 34524
rect 12492 34484 12498 34496
rect 13725 34493 13737 34496
rect 13771 34493 13783 34527
rect 14108 34524 14136 34564
rect 14182 34552 14188 34604
rect 14240 34552 14246 34604
rect 14366 34552 14372 34604
rect 14424 34552 14430 34604
rect 14461 34595 14519 34601
rect 14461 34561 14473 34595
rect 14507 34592 14519 34595
rect 14642 34592 14648 34604
rect 14507 34564 14648 34592
rect 14507 34561 14519 34564
rect 14461 34555 14519 34561
rect 14642 34552 14648 34564
rect 14700 34552 14706 34604
rect 14752 34524 14780 34632
rect 15010 34552 15016 34604
rect 15068 34592 15074 34604
rect 15197 34595 15255 34601
rect 15197 34592 15209 34595
rect 15068 34564 15209 34592
rect 15068 34552 15074 34564
rect 15197 34561 15209 34564
rect 15243 34561 15255 34595
rect 15197 34555 15255 34561
rect 15381 34595 15439 34601
rect 15381 34561 15393 34595
rect 15427 34561 15439 34595
rect 15381 34555 15439 34561
rect 14108 34496 14780 34524
rect 13725 34487 13783 34493
rect 15102 34484 15108 34536
rect 15160 34524 15166 34536
rect 15396 34524 15424 34555
rect 16850 34552 16856 34604
rect 16908 34592 16914 34604
rect 17328 34601 17356 34632
rect 19812 34632 20444 34660
rect 17221 34595 17279 34601
rect 17221 34592 17233 34595
rect 16908 34564 17233 34592
rect 16908 34552 16914 34564
rect 17221 34561 17233 34564
rect 17267 34561 17279 34595
rect 17221 34555 17279 34561
rect 17313 34595 17371 34601
rect 17313 34561 17325 34595
rect 17359 34561 17371 34595
rect 17313 34555 17371 34561
rect 15160 34496 15424 34524
rect 17328 34524 17356 34555
rect 17494 34552 17500 34604
rect 17552 34552 17558 34604
rect 17589 34595 17647 34601
rect 17589 34561 17601 34595
rect 17635 34592 17647 34595
rect 17678 34592 17684 34604
rect 17635 34564 17684 34592
rect 17635 34561 17647 34564
rect 17589 34555 17647 34561
rect 17678 34552 17684 34564
rect 17736 34552 17742 34604
rect 17954 34552 17960 34604
rect 18012 34592 18018 34604
rect 18233 34595 18291 34601
rect 18233 34592 18245 34595
rect 18012 34564 18245 34592
rect 18012 34552 18018 34564
rect 18233 34561 18245 34564
rect 18279 34561 18291 34595
rect 18233 34555 18291 34561
rect 19610 34552 19616 34604
rect 19668 34552 19674 34604
rect 19702 34552 19708 34604
rect 19760 34552 19766 34604
rect 19812 34601 19840 34632
rect 20438 34620 20444 34632
rect 20496 34620 20502 34672
rect 20916 34601 20944 34688
rect 23201 34663 23259 34669
rect 23201 34629 23213 34663
rect 23247 34660 23259 34663
rect 23382 34660 23388 34672
rect 23247 34632 23388 34660
rect 23247 34629 23259 34632
rect 23201 34623 23259 34629
rect 23382 34620 23388 34632
rect 23440 34620 23446 34672
rect 19797 34595 19855 34601
rect 19797 34561 19809 34595
rect 19843 34561 19855 34595
rect 19797 34555 19855 34561
rect 20901 34595 20959 34601
rect 20901 34561 20913 34595
rect 20947 34561 20959 34595
rect 20901 34555 20959 34561
rect 20990 34552 20996 34604
rect 21048 34592 21054 34604
rect 22005 34595 22063 34601
rect 22005 34592 22017 34595
rect 21048 34564 22017 34592
rect 21048 34552 21054 34564
rect 22005 34561 22017 34564
rect 22051 34561 22063 34595
rect 22005 34555 22063 34561
rect 22465 34595 22523 34601
rect 22465 34561 22477 34595
rect 22511 34561 22523 34595
rect 22465 34555 22523 34561
rect 17770 34524 17776 34536
rect 17328 34496 17776 34524
rect 15160 34484 15166 34496
rect 17770 34484 17776 34496
rect 17828 34484 17834 34536
rect 20809 34527 20867 34533
rect 20809 34493 20821 34527
rect 20855 34524 20867 34527
rect 21358 34524 21364 34536
rect 20855 34496 21364 34524
rect 20855 34493 20867 34496
rect 20809 34487 20867 34493
rect 21358 34484 21364 34496
rect 21416 34484 21422 34536
rect 21450 34484 21456 34536
rect 21508 34524 21514 34536
rect 22281 34527 22339 34533
rect 22281 34524 22293 34527
rect 21508 34496 22293 34524
rect 21508 34484 21514 34496
rect 22281 34493 22293 34496
rect 22327 34493 22339 34527
rect 22480 34524 22508 34555
rect 23014 34552 23020 34604
rect 23072 34592 23078 34604
rect 23109 34595 23167 34601
rect 23109 34592 23121 34595
rect 23072 34564 23121 34592
rect 23072 34552 23078 34564
rect 23109 34561 23121 34564
rect 23155 34561 23167 34595
rect 23109 34555 23167 34561
rect 23290 34552 23296 34604
rect 23348 34552 23354 34604
rect 23860 34601 23888 34688
rect 25590 34620 25596 34672
rect 25648 34620 25654 34672
rect 26602 34660 26608 34672
rect 25792 34632 26608 34660
rect 23845 34595 23903 34601
rect 23845 34561 23857 34595
rect 23891 34561 23903 34595
rect 23845 34555 23903 34561
rect 24210 34552 24216 34604
rect 24268 34552 24274 34604
rect 25608 34592 25636 34620
rect 25792 34601 25820 34632
rect 26602 34620 26608 34632
rect 26660 34660 26666 34672
rect 27154 34660 27160 34672
rect 26660 34632 27160 34660
rect 26660 34620 26666 34632
rect 27154 34620 27160 34632
rect 27212 34620 27218 34672
rect 27798 34660 27804 34672
rect 27448 34632 27804 34660
rect 25685 34595 25743 34601
rect 25685 34592 25697 34595
rect 25608 34564 25697 34592
rect 25685 34561 25697 34564
rect 25731 34561 25743 34595
rect 25685 34555 25743 34561
rect 25777 34595 25835 34601
rect 25777 34561 25789 34595
rect 25823 34561 25835 34595
rect 25777 34555 25835 34561
rect 25961 34595 26019 34601
rect 25961 34561 25973 34595
rect 26007 34561 26019 34595
rect 25961 34555 26019 34561
rect 26053 34595 26111 34601
rect 26053 34561 26065 34595
rect 26099 34593 26111 34595
rect 26099 34592 26168 34593
rect 26418 34592 26424 34604
rect 26099 34565 26424 34592
rect 26099 34561 26111 34565
rect 26140 34564 26424 34565
rect 26053 34555 26111 34561
rect 25976 34524 26004 34555
rect 26418 34552 26424 34564
rect 26476 34552 26482 34604
rect 26786 34552 26792 34604
rect 26844 34592 26850 34604
rect 27448 34601 27476 34632
rect 27798 34620 27804 34632
rect 27856 34620 27862 34672
rect 27890 34620 27896 34672
rect 27948 34620 27954 34672
rect 27433 34595 27491 34601
rect 27433 34592 27445 34595
rect 26844 34564 27445 34592
rect 26844 34552 26850 34564
rect 27433 34561 27445 34564
rect 27479 34561 27491 34595
rect 27433 34555 27491 34561
rect 27522 34552 27528 34604
rect 27580 34552 27586 34604
rect 28258 34592 28264 34604
rect 27724 34564 28264 34592
rect 22480 34496 26004 34524
rect 26436 34524 26464 34552
rect 27724 34524 27752 34564
rect 28258 34552 28264 34564
rect 28316 34552 28322 34604
rect 28537 34595 28595 34601
rect 28537 34561 28549 34595
rect 28583 34592 28595 34595
rect 28644 34592 28672 34700
rect 31846 34688 31852 34700
rect 31904 34688 31910 34740
rect 33870 34688 33876 34740
rect 33928 34728 33934 34740
rect 34149 34731 34207 34737
rect 34149 34728 34161 34731
rect 33928 34700 34161 34728
rect 33928 34688 33934 34700
rect 34149 34697 34161 34700
rect 34195 34697 34207 34731
rect 34149 34691 34207 34697
rect 34606 34688 34612 34740
rect 34664 34728 34670 34740
rect 35345 34731 35403 34737
rect 35345 34728 35357 34731
rect 34664 34700 35357 34728
rect 34664 34688 34670 34700
rect 35345 34697 35357 34700
rect 35391 34697 35403 34731
rect 35345 34691 35403 34697
rect 36906 34688 36912 34740
rect 36964 34688 36970 34740
rect 37090 34688 37096 34740
rect 37148 34728 37154 34740
rect 37461 34731 37519 34737
rect 37461 34728 37473 34731
rect 37148 34700 37473 34728
rect 37148 34688 37154 34700
rect 37461 34697 37473 34700
rect 37507 34697 37519 34731
rect 37461 34691 37519 34697
rect 28994 34620 29000 34672
rect 29052 34660 29058 34672
rect 33686 34660 33692 34672
rect 29052 34632 32536 34660
rect 29052 34620 29058 34632
rect 30098 34592 30104 34604
rect 28583 34564 28672 34592
rect 29472 34564 30104 34592
rect 28583 34561 28595 34564
rect 28537 34555 28595 34561
rect 26436 34496 27752 34524
rect 22281 34487 22339 34493
rect 25608 34468 25636 34496
rect 27798 34484 27804 34536
rect 27856 34524 27862 34536
rect 29472 34524 29500 34564
rect 30098 34552 30104 34564
rect 30156 34552 30162 34604
rect 30374 34552 30380 34604
rect 30432 34592 30438 34604
rect 30650 34592 30656 34604
rect 30432 34564 30656 34592
rect 30432 34552 30438 34564
rect 30650 34552 30656 34564
rect 30708 34552 30714 34604
rect 30742 34552 30748 34604
rect 30800 34552 30806 34604
rect 32508 34601 32536 34632
rect 32968 34632 33692 34660
rect 32493 34595 32551 34601
rect 30944 34564 31754 34592
rect 27856 34496 29500 34524
rect 27856 34484 27862 34496
rect 29546 34484 29552 34536
rect 29604 34484 29610 34536
rect 30116 34524 30144 34552
rect 30944 34524 30972 34564
rect 30116 34496 30972 34524
rect 31018 34484 31024 34536
rect 31076 34524 31082 34536
rect 31294 34524 31300 34536
rect 31076 34496 31300 34524
rect 31076 34484 31082 34496
rect 31294 34484 31300 34496
rect 31352 34484 31358 34536
rect 31726 34524 31754 34564
rect 32493 34561 32505 34595
rect 32539 34561 32551 34595
rect 32858 34592 32864 34604
rect 32493 34555 32551 34561
rect 32600 34564 32864 34592
rect 32600 34524 32628 34564
rect 32858 34552 32864 34564
rect 32916 34552 32922 34604
rect 31726 34496 32628 34524
rect 32674 34484 32680 34536
rect 32732 34484 32738 34536
rect 32769 34527 32827 34533
rect 32769 34493 32781 34527
rect 32815 34524 32827 34527
rect 32968 34524 32996 34632
rect 33686 34620 33692 34632
rect 33744 34620 33750 34672
rect 33781 34663 33839 34669
rect 33781 34629 33793 34663
rect 33827 34660 33839 34663
rect 34330 34660 34336 34672
rect 33827 34632 34336 34660
rect 33827 34629 33839 34632
rect 33781 34623 33839 34629
rect 34330 34620 34336 34632
rect 34388 34660 34394 34672
rect 34977 34663 35035 34669
rect 34977 34660 34989 34663
rect 34388 34632 34989 34660
rect 34388 34620 34394 34632
rect 34977 34629 34989 34632
rect 35023 34629 35035 34663
rect 37182 34660 37188 34672
rect 34977 34623 35035 34629
rect 36648 34632 37188 34660
rect 33502 34552 33508 34604
rect 33560 34552 33566 34604
rect 33594 34552 33600 34604
rect 33652 34592 33658 34604
rect 33873 34595 33931 34601
rect 33652 34564 33697 34592
rect 33652 34552 33658 34564
rect 33873 34561 33885 34595
rect 33919 34561 33931 34595
rect 33873 34555 33931 34561
rect 33970 34595 34028 34601
rect 33970 34561 33982 34595
rect 34016 34561 34028 34595
rect 33970 34555 34028 34561
rect 32815 34496 32996 34524
rect 32815 34493 32827 34496
rect 32769 34487 32827 34493
rect 32876 34468 32904 34496
rect 33410 34484 33416 34536
rect 33468 34524 33474 34536
rect 33888 34524 33916 34555
rect 33468 34496 33916 34524
rect 33985 34524 34013 34555
rect 34146 34552 34152 34604
rect 34204 34592 34210 34604
rect 34701 34595 34759 34601
rect 34701 34592 34713 34595
rect 34204 34564 34713 34592
rect 34204 34552 34210 34564
rect 34701 34561 34713 34564
rect 34747 34561 34759 34595
rect 34701 34555 34759 34561
rect 34794 34595 34852 34601
rect 34794 34561 34806 34595
rect 34840 34561 34852 34595
rect 34794 34555 34852 34561
rect 34809 34524 34837 34555
rect 35066 34552 35072 34604
rect 35124 34552 35130 34604
rect 35158 34552 35164 34604
rect 35216 34601 35222 34604
rect 35216 34592 35224 34601
rect 35216 34564 35261 34592
rect 35216 34555 35224 34564
rect 35216 34552 35222 34555
rect 35618 34552 35624 34604
rect 35676 34592 35682 34604
rect 36265 34595 36323 34601
rect 36265 34592 36277 34595
rect 35676 34564 36277 34592
rect 35676 34552 35682 34564
rect 36265 34561 36277 34564
rect 36311 34561 36323 34595
rect 36265 34555 36323 34561
rect 36358 34595 36416 34601
rect 36358 34561 36370 34595
rect 36404 34561 36416 34595
rect 36358 34555 36416 34561
rect 35434 34524 35440 34536
rect 33985 34496 34744 34524
rect 34809 34496 35440 34524
rect 33468 34484 33474 34496
rect 34716 34468 34744 34496
rect 35434 34484 35440 34496
rect 35492 34484 35498 34536
rect 36170 34484 36176 34536
rect 36228 34524 36234 34536
rect 36373 34524 36401 34555
rect 36538 34552 36544 34604
rect 36596 34552 36602 34604
rect 36648 34601 36676 34632
rect 37182 34620 37188 34632
rect 37240 34620 37246 34672
rect 36633 34595 36691 34601
rect 36633 34561 36645 34595
rect 36679 34561 36691 34595
rect 36633 34555 36691 34561
rect 36228 34496 36401 34524
rect 36228 34484 36234 34496
rect 9490 34456 9496 34468
rect 8956 34428 9496 34456
rect 9490 34416 9496 34428
rect 9548 34416 9554 34468
rect 10870 34416 10876 34468
rect 10928 34456 10934 34468
rect 11977 34459 12035 34465
rect 11977 34456 11989 34459
rect 10928 34428 11989 34456
rect 10928 34416 10934 34428
rect 11977 34425 11989 34428
rect 12023 34425 12035 34459
rect 11977 34419 12035 34425
rect 12069 34459 12127 34465
rect 12069 34425 12081 34459
rect 12115 34456 12127 34459
rect 12802 34456 12808 34468
rect 12115 34428 12808 34456
rect 12115 34425 12127 34428
rect 12069 34419 12127 34425
rect 12802 34416 12808 34428
rect 12860 34416 12866 34468
rect 12894 34416 12900 34468
rect 12952 34456 12958 34468
rect 12952 34428 13400 34456
rect 12952 34416 12958 34428
rect 4154 34348 4160 34400
rect 4212 34388 4218 34400
rect 7098 34388 7104 34400
rect 4212 34360 7104 34388
rect 4212 34348 4218 34360
rect 7098 34348 7104 34360
rect 7156 34348 7162 34400
rect 7469 34391 7527 34397
rect 7469 34357 7481 34391
rect 7515 34388 7527 34391
rect 9582 34388 9588 34400
rect 7515 34360 9588 34388
rect 7515 34357 7527 34360
rect 7469 34351 7527 34357
rect 9582 34348 9588 34360
rect 9640 34348 9646 34400
rect 10134 34348 10140 34400
rect 10192 34388 10198 34400
rect 10321 34391 10379 34397
rect 10321 34388 10333 34391
rect 10192 34360 10333 34388
rect 10192 34348 10198 34360
rect 10321 34357 10333 34360
rect 10367 34357 10379 34391
rect 10321 34351 10379 34357
rect 13262 34348 13268 34400
rect 13320 34348 13326 34400
rect 13372 34388 13400 34428
rect 13538 34416 13544 34468
rect 13596 34456 13602 34468
rect 16022 34456 16028 34468
rect 13596 34428 16028 34456
rect 13596 34416 13602 34428
rect 16022 34416 16028 34428
rect 16080 34416 16086 34468
rect 17037 34459 17095 34465
rect 17037 34425 17049 34459
rect 17083 34456 17095 34459
rect 17083 34428 18184 34456
rect 17083 34425 17095 34428
rect 17037 34419 17095 34425
rect 13630 34388 13636 34400
rect 13372 34360 13636 34388
rect 13630 34348 13636 34360
rect 13688 34348 13694 34400
rect 13814 34348 13820 34400
rect 13872 34388 13878 34400
rect 14185 34391 14243 34397
rect 14185 34388 14197 34391
rect 13872 34360 14197 34388
rect 13872 34348 13878 34360
rect 14185 34357 14197 34360
rect 14231 34388 14243 34391
rect 14458 34388 14464 34400
rect 14231 34360 14464 34388
rect 14231 34357 14243 34360
rect 14185 34351 14243 34357
rect 14458 34348 14464 34360
rect 14516 34348 14522 34400
rect 14642 34348 14648 34400
rect 14700 34388 14706 34400
rect 17954 34388 17960 34400
rect 14700 34360 17960 34388
rect 14700 34348 14706 34360
rect 17954 34348 17960 34360
rect 18012 34348 18018 34400
rect 18156 34388 18184 34428
rect 18322 34416 18328 34468
rect 18380 34456 18386 34468
rect 18417 34459 18475 34465
rect 18417 34456 18429 34459
rect 18380 34428 18429 34456
rect 18380 34416 18386 34428
rect 18417 34425 18429 34428
rect 18463 34425 18475 34459
rect 18417 34419 18475 34425
rect 19334 34416 19340 34468
rect 19392 34456 19398 34468
rect 25222 34456 25228 34468
rect 19392 34428 25228 34456
rect 19392 34416 19398 34428
rect 25222 34416 25228 34428
rect 25280 34416 25286 34468
rect 25590 34416 25596 34468
rect 25648 34416 25654 34468
rect 25866 34416 25872 34468
rect 25924 34456 25930 34468
rect 32398 34456 32404 34468
rect 25924 34428 32404 34456
rect 25924 34416 25930 34428
rect 32398 34416 32404 34428
rect 32456 34416 32462 34468
rect 32858 34416 32864 34468
rect 32916 34416 32922 34468
rect 33134 34416 33140 34468
rect 33192 34456 33198 34468
rect 34422 34456 34428 34468
rect 33192 34428 34428 34456
rect 33192 34416 33198 34428
rect 34422 34416 34428 34428
rect 34480 34416 34486 34468
rect 34698 34416 34704 34468
rect 34756 34456 34762 34468
rect 35158 34456 35164 34468
rect 34756 34428 35164 34456
rect 34756 34416 34762 34428
rect 35158 34416 35164 34428
rect 35216 34416 35222 34468
rect 35452 34456 35480 34484
rect 36648 34456 36676 34555
rect 36722 34552 36728 34604
rect 36780 34601 36786 34604
rect 36780 34592 36788 34601
rect 36780 34564 36825 34592
rect 36780 34555 36788 34564
rect 36780 34552 36786 34555
rect 37826 34552 37832 34604
rect 37884 34552 37890 34604
rect 37921 34527 37979 34533
rect 37921 34524 37933 34527
rect 36740 34496 37933 34524
rect 36740 34468 36768 34496
rect 37921 34493 37933 34496
rect 37967 34493 37979 34527
rect 37921 34487 37979 34493
rect 38102 34484 38108 34536
rect 38160 34484 38166 34536
rect 35452 34428 36676 34456
rect 36722 34416 36728 34468
rect 36780 34416 36786 34468
rect 36814 34416 36820 34468
rect 36872 34456 36878 34468
rect 37182 34456 37188 34468
rect 36872 34428 37188 34456
rect 36872 34416 36878 34428
rect 37182 34416 37188 34428
rect 37240 34416 37246 34468
rect 20714 34388 20720 34400
rect 18156 34360 20720 34388
rect 20714 34348 20720 34360
rect 20772 34348 20778 34400
rect 20806 34348 20812 34400
rect 20864 34348 20870 34400
rect 21082 34348 21088 34400
rect 21140 34388 21146 34400
rect 21818 34388 21824 34400
rect 21140 34360 21824 34388
rect 21140 34348 21146 34360
rect 21818 34348 21824 34360
rect 21876 34348 21882 34400
rect 22094 34348 22100 34400
rect 22152 34348 22158 34400
rect 22646 34348 22652 34400
rect 22704 34388 22710 34400
rect 24210 34388 24216 34400
rect 22704 34360 24216 34388
rect 22704 34348 22710 34360
rect 24210 34348 24216 34360
rect 24268 34348 24274 34400
rect 25498 34348 25504 34400
rect 25556 34348 25562 34400
rect 27246 34348 27252 34400
rect 27304 34348 27310 34400
rect 27890 34348 27896 34400
rect 27948 34388 27954 34400
rect 28810 34388 28816 34400
rect 27948 34360 28816 34388
rect 27948 34348 27954 34360
rect 28810 34348 28816 34360
rect 28868 34348 28874 34400
rect 30834 34348 30840 34400
rect 30892 34348 30898 34400
rect 32309 34391 32367 34397
rect 32309 34357 32321 34391
rect 32355 34388 32367 34391
rect 32490 34388 32496 34400
rect 32355 34360 32496 34388
rect 32355 34357 32367 34360
rect 32309 34351 32367 34357
rect 32490 34348 32496 34360
rect 32548 34348 32554 34400
rect 33870 34348 33876 34400
rect 33928 34388 33934 34400
rect 37458 34388 37464 34400
rect 33928 34360 37464 34388
rect 33928 34348 33934 34360
rect 37458 34348 37464 34360
rect 37516 34348 37522 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 4982 34144 4988 34196
rect 5040 34184 5046 34196
rect 5169 34187 5227 34193
rect 5169 34184 5181 34187
rect 5040 34156 5181 34184
rect 5040 34144 5046 34156
rect 5169 34153 5181 34156
rect 5215 34153 5227 34187
rect 5169 34147 5227 34153
rect 5905 34187 5963 34193
rect 5905 34153 5917 34187
rect 5951 34184 5963 34187
rect 6822 34184 6828 34196
rect 5951 34156 6828 34184
rect 5951 34153 5963 34156
rect 5905 34147 5963 34153
rect 6822 34144 6828 34156
rect 6880 34144 6886 34196
rect 7558 34144 7564 34196
rect 7616 34184 7622 34196
rect 8202 34184 8208 34196
rect 7616 34156 8208 34184
rect 7616 34144 7622 34156
rect 8202 34144 8208 34156
rect 8260 34144 8266 34196
rect 8570 34144 8576 34196
rect 8628 34184 8634 34196
rect 9585 34187 9643 34193
rect 9585 34184 9597 34187
rect 8628 34156 9597 34184
rect 8628 34144 8634 34156
rect 9585 34153 9597 34156
rect 9631 34184 9643 34187
rect 9674 34184 9680 34196
rect 9631 34156 9680 34184
rect 9631 34153 9643 34156
rect 9585 34147 9643 34153
rect 9674 34144 9680 34156
rect 9732 34144 9738 34196
rect 13078 34184 13084 34196
rect 9784 34156 13084 34184
rect 5077 34119 5135 34125
rect 5077 34085 5089 34119
rect 5123 34116 5135 34119
rect 7926 34116 7932 34128
rect 5123 34088 7932 34116
rect 5123 34085 5135 34088
rect 5077 34079 5135 34085
rect 7926 34076 7932 34088
rect 7984 34076 7990 34128
rect 8018 34076 8024 34128
rect 8076 34116 8082 34128
rect 9784 34116 9812 34156
rect 13078 34144 13084 34156
rect 13136 34144 13142 34196
rect 13354 34184 13360 34196
rect 13280 34156 13360 34184
rect 8076 34088 9168 34116
rect 8076 34076 8082 34088
rect 5166 34048 5172 34060
rect 4356 34020 5172 34048
rect 4062 33940 4068 33992
rect 4120 33940 4126 33992
rect 4356 33989 4384 34020
rect 5166 34008 5172 34020
rect 5224 34008 5230 34060
rect 5261 34051 5319 34057
rect 5261 34017 5273 34051
rect 5307 34048 5319 34051
rect 5534 34048 5540 34060
rect 5307 34020 5540 34048
rect 5307 34017 5319 34020
rect 5261 34011 5319 34017
rect 4341 33983 4399 33989
rect 4341 33949 4353 33983
rect 4387 33949 4399 33983
rect 4341 33943 4399 33949
rect 4525 33983 4583 33989
rect 4525 33949 4537 33983
rect 4571 33949 4583 33983
rect 4525 33943 4583 33949
rect 4080 33912 4108 33940
rect 4540 33912 4568 33943
rect 4982 33940 4988 33992
rect 5040 33940 5046 33992
rect 4080 33884 4568 33912
rect 4890 33872 4896 33924
rect 4948 33912 4954 33924
rect 5276 33912 5304 34011
rect 5534 34008 5540 34020
rect 5592 34008 5598 34060
rect 6086 34008 6092 34060
rect 6144 34048 6150 34060
rect 6546 34048 6552 34060
rect 6144 34020 6552 34048
rect 6144 34008 6150 34020
rect 6546 34008 6552 34020
rect 6604 34008 6610 34060
rect 8303 34048 8432 34056
rect 8573 34051 8631 34057
rect 8573 34048 8585 34051
rect 8303 34028 8585 34048
rect 5721 33983 5779 33989
rect 5721 33949 5733 33983
rect 5767 33949 5779 33983
rect 5721 33943 5779 33949
rect 5905 33983 5963 33989
rect 5905 33949 5917 33983
rect 5951 33980 5963 33983
rect 6178 33980 6184 33992
rect 5951 33952 6184 33980
rect 5951 33949 5963 33952
rect 5905 33943 5963 33949
rect 4948 33884 5304 33912
rect 5736 33912 5764 33943
rect 6178 33940 6184 33952
rect 6236 33940 6242 33992
rect 6638 33980 6644 33992
rect 6288 33952 6644 33980
rect 6288 33912 6316 33952
rect 6638 33940 6644 33952
rect 6696 33940 6702 33992
rect 7282 33940 7288 33992
rect 7340 33980 7346 33992
rect 7377 33983 7435 33989
rect 7377 33980 7389 33983
rect 7340 33952 7389 33980
rect 7340 33940 7346 33952
rect 7377 33949 7389 33952
rect 7423 33949 7435 33983
rect 7377 33943 7435 33949
rect 7466 33940 7472 33992
rect 7524 33940 7530 33992
rect 7834 33940 7840 33992
rect 7892 33980 7898 33992
rect 8303 33980 8331 34028
rect 8404 34020 8585 34028
rect 8573 34017 8585 34020
rect 8619 34048 8631 34051
rect 8938 34048 8944 34060
rect 8619 34020 8944 34048
rect 8619 34017 8631 34020
rect 8573 34011 8631 34017
rect 8938 34008 8944 34020
rect 8996 34008 9002 34060
rect 7892 33952 8331 33980
rect 7892 33940 7898 33952
rect 8386 33940 8392 33992
rect 8444 33940 8450 33992
rect 5736 33884 6316 33912
rect 4948 33872 4954 33884
rect 6546 33872 6552 33924
rect 6604 33872 6610 33924
rect 6730 33872 6736 33924
rect 6788 33872 6794 33924
rect 6914 33872 6920 33924
rect 6972 33872 6978 33924
rect 7098 33872 7104 33924
rect 7156 33912 7162 33924
rect 8205 33915 8263 33921
rect 8205 33912 8217 33915
rect 7156 33884 8217 33912
rect 7156 33872 7162 33884
rect 8205 33881 8217 33884
rect 8251 33912 8263 33915
rect 9030 33912 9036 33924
rect 8251 33884 9036 33912
rect 8251 33881 8263 33884
rect 8205 33875 8263 33881
rect 9030 33872 9036 33884
rect 9088 33872 9094 33924
rect 9140 33912 9168 34088
rect 9508 34088 9812 34116
rect 9861 34119 9919 34125
rect 9508 33989 9536 34088
rect 9861 34085 9873 34119
rect 9907 34116 9919 34119
rect 13170 34116 13176 34128
rect 9907 34088 13176 34116
rect 9907 34085 9919 34088
rect 9861 34079 9919 34085
rect 13170 34076 13176 34088
rect 13228 34076 13234 34128
rect 9674 34008 9680 34060
rect 9732 34048 9738 34060
rect 13280 34048 13308 34156
rect 13354 34144 13360 34156
rect 13412 34144 13418 34196
rect 14550 34144 14556 34196
rect 14608 34144 14614 34196
rect 14734 34144 14740 34196
rect 14792 34144 14798 34196
rect 15838 34144 15844 34196
rect 15896 34184 15902 34196
rect 15896 34156 19840 34184
rect 15896 34144 15902 34156
rect 17405 34119 17463 34125
rect 17405 34116 17417 34119
rect 14936 34088 17417 34116
rect 9732 34020 13308 34048
rect 9732 34008 9738 34020
rect 14366 34008 14372 34060
rect 14424 34008 14430 34060
rect 14936 33992 14964 34088
rect 17405 34085 17417 34088
rect 17451 34085 17463 34119
rect 17405 34079 17463 34085
rect 17494 34076 17500 34128
rect 17552 34116 17558 34128
rect 18874 34116 18880 34128
rect 17552 34088 18880 34116
rect 17552 34076 17558 34088
rect 18874 34076 18880 34088
rect 18932 34076 18938 34128
rect 19702 34116 19708 34128
rect 19444 34088 19708 34116
rect 15562 34008 15568 34060
rect 15620 34048 15626 34060
rect 15746 34048 15752 34060
rect 15620 34020 15752 34048
rect 15620 34008 15626 34020
rect 15746 34008 15752 34020
rect 15804 34008 15810 34060
rect 15838 34008 15844 34060
rect 15896 34008 15902 34060
rect 16209 34051 16267 34057
rect 16209 34017 16221 34051
rect 16255 34048 16267 34051
rect 16255 34020 17816 34048
rect 16255 34017 16267 34020
rect 16209 34011 16267 34017
rect 9493 33983 9551 33989
rect 9493 33949 9505 33983
rect 9539 33949 9551 33983
rect 9493 33943 9551 33949
rect 9585 33983 9643 33989
rect 9585 33949 9597 33983
rect 9631 33980 9643 33983
rect 9766 33980 9772 33992
rect 9631 33952 9772 33980
rect 9631 33949 9643 33952
rect 9585 33943 9643 33949
rect 9766 33940 9772 33952
rect 9824 33940 9830 33992
rect 10318 33940 10324 33992
rect 10376 33940 10382 33992
rect 10689 33983 10747 33989
rect 10689 33949 10701 33983
rect 10735 33980 10747 33983
rect 10870 33980 10876 33992
rect 10735 33952 10876 33980
rect 10735 33949 10747 33952
rect 10689 33943 10747 33949
rect 10870 33940 10876 33952
rect 10928 33940 10934 33992
rect 11057 33983 11115 33989
rect 11057 33949 11069 33983
rect 11103 33980 11115 33983
rect 11146 33980 11152 33992
rect 11103 33952 11152 33980
rect 11103 33949 11115 33952
rect 11057 33943 11115 33949
rect 11146 33940 11152 33952
rect 11204 33940 11210 33992
rect 11514 33940 11520 33992
rect 11572 33980 11578 33992
rect 11977 33983 12035 33989
rect 11977 33980 11989 33983
rect 11572 33952 11989 33980
rect 11572 33940 11578 33952
rect 11977 33949 11989 33952
rect 12023 33949 12035 33983
rect 11977 33943 12035 33949
rect 12345 33983 12403 33989
rect 12345 33949 12357 33983
rect 12391 33980 12403 33983
rect 12434 33980 12440 33992
rect 12391 33952 12440 33980
rect 12391 33949 12403 33952
rect 12345 33943 12403 33949
rect 12434 33940 12440 33952
rect 12492 33940 12498 33992
rect 12526 33940 12532 33992
rect 12584 33940 12590 33992
rect 13004 33982 13288 33990
rect 13357 33983 13415 33989
rect 13357 33982 13369 33983
rect 13004 33962 13369 33982
rect 13004 33912 13032 33962
rect 13260 33954 13369 33962
rect 13357 33949 13369 33954
rect 13403 33949 13415 33983
rect 13357 33943 13415 33949
rect 13449 33983 13507 33989
rect 13449 33949 13461 33983
rect 13495 33949 13507 33983
rect 13449 33943 13507 33949
rect 9140 33884 13032 33912
rect 13170 33872 13176 33924
rect 13228 33872 13234 33924
rect 13464 33912 13492 33943
rect 13630 33940 13636 33992
rect 13688 33940 13694 33992
rect 13725 33983 13783 33989
rect 13725 33949 13737 33983
rect 13771 33980 13783 33983
rect 13814 33980 13820 33992
rect 13771 33952 13820 33980
rect 13771 33949 13783 33952
rect 13725 33943 13783 33949
rect 13814 33940 13820 33952
rect 13872 33940 13878 33992
rect 14553 33983 14611 33989
rect 14553 33949 14565 33983
rect 14599 33980 14611 33983
rect 14642 33980 14648 33992
rect 14599 33952 14648 33980
rect 14599 33949 14611 33952
rect 14553 33943 14611 33949
rect 14642 33940 14648 33952
rect 14700 33980 14706 33992
rect 14826 33980 14832 33992
rect 14700 33952 14832 33980
rect 14700 33940 14706 33952
rect 14826 33940 14832 33952
rect 14884 33940 14890 33992
rect 14918 33940 14924 33992
rect 14976 33940 14982 33992
rect 15102 33940 15108 33992
rect 15160 33980 15166 33992
rect 15473 33983 15531 33989
rect 15473 33980 15485 33983
rect 15160 33952 15485 33980
rect 15160 33940 15166 33952
rect 15473 33949 15485 33952
rect 15519 33949 15531 33983
rect 15473 33943 15531 33949
rect 15654 33940 15660 33992
rect 15712 33940 15718 33992
rect 16022 33940 16028 33992
rect 16080 33940 16086 33992
rect 16666 33940 16672 33992
rect 16724 33940 16730 33992
rect 17788 33989 17816 34020
rect 18230 34008 18236 34060
rect 18288 34048 18294 34060
rect 19444 34057 19472 34088
rect 19702 34076 19708 34088
rect 19760 34076 19766 34128
rect 19812 34125 19840 34156
rect 20622 34144 20628 34196
rect 20680 34184 20686 34196
rect 21269 34187 21327 34193
rect 21269 34184 21281 34187
rect 20680 34156 21281 34184
rect 20680 34144 20686 34156
rect 21269 34153 21281 34156
rect 21315 34184 21327 34187
rect 21634 34184 21640 34196
rect 21315 34156 21640 34184
rect 21315 34153 21327 34156
rect 21269 34147 21327 34153
rect 21634 34144 21640 34156
rect 21692 34144 21698 34196
rect 21818 34144 21824 34196
rect 21876 34184 21882 34196
rect 21913 34187 21971 34193
rect 21913 34184 21925 34187
rect 21876 34156 21925 34184
rect 21876 34144 21882 34156
rect 21913 34153 21925 34156
rect 21959 34153 21971 34187
rect 22094 34184 22100 34196
rect 21913 34147 21971 34153
rect 22066 34144 22100 34184
rect 22152 34144 22158 34196
rect 23014 34184 23020 34196
rect 22204 34156 23020 34184
rect 19797 34119 19855 34125
rect 19797 34085 19809 34119
rect 19843 34085 19855 34119
rect 19797 34079 19855 34085
rect 21358 34076 21364 34128
rect 21416 34116 21422 34128
rect 22066 34116 22094 34144
rect 21416 34088 22094 34116
rect 21416 34076 21422 34088
rect 19429 34051 19487 34057
rect 19429 34048 19441 34051
rect 18288 34020 19441 34048
rect 18288 34008 18294 34020
rect 19429 34017 19441 34020
rect 19475 34017 19487 34051
rect 19429 34011 19487 34017
rect 19518 34008 19524 34060
rect 19576 34048 19582 34060
rect 19576 34020 19748 34048
rect 19576 34008 19582 34020
rect 17773 33983 17831 33989
rect 17773 33949 17785 33983
rect 17819 33949 17831 33983
rect 17773 33943 17831 33949
rect 17954 33940 17960 33992
rect 18012 33980 18018 33992
rect 18509 33983 18567 33989
rect 18509 33980 18521 33983
rect 18012 33952 18521 33980
rect 18012 33940 18018 33952
rect 18509 33949 18521 33952
rect 18555 33949 18567 33983
rect 18509 33943 18567 33949
rect 18693 33983 18751 33989
rect 18693 33949 18705 33983
rect 18739 33949 18751 33983
rect 18693 33943 18751 33949
rect 13372 33884 13492 33912
rect 13648 33912 13676 33940
rect 13648 33884 14136 33912
rect 4062 33804 4068 33856
rect 4120 33844 4126 33856
rect 4433 33847 4491 33853
rect 4433 33844 4445 33847
rect 4120 33816 4445 33844
rect 4120 33804 4126 33816
rect 4433 33813 4445 33816
rect 4479 33813 4491 33847
rect 4433 33807 4491 33813
rect 6086 33804 6092 33856
rect 6144 33804 6150 33856
rect 6178 33804 6184 33856
rect 6236 33844 6242 33856
rect 7466 33844 7472 33856
rect 6236 33816 7472 33844
rect 6236 33804 6242 33816
rect 7466 33804 7472 33816
rect 7524 33804 7530 33856
rect 7742 33804 7748 33856
rect 7800 33804 7806 33856
rect 7926 33804 7932 33856
rect 7984 33844 7990 33856
rect 12342 33844 12348 33856
rect 7984 33816 12348 33844
rect 7984 33804 7990 33816
rect 12342 33804 12348 33816
rect 12400 33804 12406 33856
rect 12986 33804 12992 33856
rect 13044 33844 13050 33856
rect 13372 33844 13400 33884
rect 13044 33816 13400 33844
rect 13044 33804 13050 33816
rect 13446 33804 13452 33856
rect 13504 33844 13510 33856
rect 13998 33844 14004 33856
rect 13504 33816 14004 33844
rect 13504 33804 13510 33816
rect 13998 33804 14004 33816
rect 14056 33804 14062 33856
rect 14108 33844 14136 33884
rect 14182 33872 14188 33924
rect 14240 33912 14246 33924
rect 14277 33915 14335 33921
rect 14277 33912 14289 33915
rect 14240 33884 14289 33912
rect 14240 33872 14246 33884
rect 14277 33881 14289 33884
rect 14323 33881 14335 33915
rect 14277 33875 14335 33881
rect 17586 33872 17592 33924
rect 17644 33872 17650 33924
rect 18708 33912 18736 33943
rect 18874 33940 18880 33992
rect 18932 33980 18938 33992
rect 19720 33989 19748 34020
rect 20346 34008 20352 34060
rect 20404 34048 20410 34060
rect 21085 34051 21143 34057
rect 21085 34048 21097 34051
rect 20404 34020 21097 34048
rect 20404 34008 20410 34020
rect 21085 34017 21097 34020
rect 21131 34048 21143 34051
rect 21131 34020 22048 34048
rect 21131 34017 21143 34020
rect 21085 34011 21143 34017
rect 19613 33983 19671 33989
rect 19613 33980 19625 33983
rect 18932 33952 19625 33980
rect 18932 33940 18938 33952
rect 19613 33949 19625 33952
rect 19659 33949 19671 33983
rect 19613 33943 19671 33949
rect 19705 33983 19763 33989
rect 19705 33949 19717 33983
rect 19751 33949 19763 33983
rect 19705 33943 19763 33949
rect 19889 33983 19947 33989
rect 19889 33949 19901 33983
rect 19935 33980 19947 33983
rect 20622 33980 20628 33992
rect 19935 33952 20628 33980
rect 19935 33949 19947 33952
rect 19889 33943 19947 33949
rect 20622 33940 20628 33952
rect 20680 33940 20686 33992
rect 21266 33940 21272 33992
rect 21324 33940 21330 33992
rect 21542 33940 21548 33992
rect 21600 33980 21606 33992
rect 21913 33983 21971 33989
rect 21913 33980 21925 33983
rect 21600 33952 21925 33980
rect 21600 33940 21606 33952
rect 21913 33949 21925 33952
rect 21959 33949 21971 33983
rect 22020 33980 22048 34020
rect 22094 34008 22100 34060
rect 22152 34048 22158 34060
rect 22204 34048 22232 34156
rect 23014 34144 23020 34156
rect 23072 34144 23078 34196
rect 23845 34187 23903 34193
rect 23845 34153 23857 34187
rect 23891 34184 23903 34187
rect 23934 34184 23940 34196
rect 23891 34156 23940 34184
rect 23891 34153 23903 34156
rect 23845 34147 23903 34153
rect 23934 34144 23940 34156
rect 23992 34144 23998 34196
rect 24029 34187 24087 34193
rect 24029 34153 24041 34187
rect 24075 34184 24087 34187
rect 24394 34184 24400 34196
rect 24075 34156 24400 34184
rect 24075 34153 24087 34156
rect 24029 34147 24087 34153
rect 24394 34144 24400 34156
rect 24452 34144 24458 34196
rect 24854 34144 24860 34196
rect 24912 34144 24918 34196
rect 24946 34144 24952 34196
rect 25004 34184 25010 34196
rect 25774 34184 25780 34196
rect 25004 34156 25780 34184
rect 25004 34144 25010 34156
rect 25774 34144 25780 34156
rect 25832 34144 25838 34196
rect 27706 34144 27712 34196
rect 27764 34184 27770 34196
rect 31570 34184 31576 34196
rect 27764 34156 31576 34184
rect 27764 34144 27770 34156
rect 31570 34144 31576 34156
rect 31628 34144 31634 34196
rect 31846 34144 31852 34196
rect 31904 34184 31910 34196
rect 33134 34184 33140 34196
rect 31904 34156 33140 34184
rect 31904 34144 31910 34156
rect 33134 34144 33140 34156
rect 33192 34144 33198 34196
rect 33689 34187 33747 34193
rect 33689 34153 33701 34187
rect 33735 34184 33747 34187
rect 34146 34184 34152 34196
rect 33735 34156 34152 34184
rect 33735 34153 33747 34156
rect 33689 34147 33747 34153
rect 34146 34144 34152 34156
rect 34204 34144 34210 34196
rect 34238 34144 34244 34196
rect 34296 34184 34302 34196
rect 34422 34184 34428 34196
rect 34296 34156 34428 34184
rect 34296 34144 34302 34156
rect 34422 34144 34428 34156
rect 34480 34144 34486 34196
rect 34606 34144 34612 34196
rect 34664 34144 34670 34196
rect 34698 34144 34704 34196
rect 34756 34184 34762 34196
rect 34756 34156 34928 34184
rect 34756 34144 34762 34156
rect 25225 34119 25283 34125
rect 25225 34116 25237 34119
rect 22152 34020 22232 34048
rect 22572 34088 25237 34116
rect 22152 34008 22158 34020
rect 22189 33983 22247 33989
rect 22020 33952 22094 33980
rect 21913 33943 21971 33949
rect 20714 33912 20720 33924
rect 18708 33884 20720 33912
rect 20714 33872 20720 33884
rect 20772 33872 20778 33924
rect 20993 33915 21051 33921
rect 20993 33881 21005 33915
rect 21039 33912 21051 33915
rect 22066 33912 22094 33952
rect 22189 33949 22201 33983
rect 22235 33949 22247 33983
rect 22189 33943 22247 33949
rect 22204 33912 22232 33943
rect 22572 33912 22600 34088
rect 25225 34085 25237 34088
rect 25271 34085 25283 34119
rect 25225 34079 25283 34085
rect 25314 34076 25320 34128
rect 25372 34116 25378 34128
rect 27430 34116 27436 34128
rect 25372 34088 27436 34116
rect 25372 34076 25378 34088
rect 27430 34076 27436 34088
rect 27488 34076 27494 34128
rect 27893 34119 27951 34125
rect 27893 34085 27905 34119
rect 27939 34085 27951 34119
rect 27893 34079 27951 34085
rect 22922 34008 22928 34060
rect 22980 34008 22986 34060
rect 23106 34008 23112 34060
rect 23164 34008 23170 34060
rect 23750 34008 23756 34060
rect 23808 34008 23814 34060
rect 23934 34008 23940 34060
rect 23992 34048 23998 34060
rect 27908 34048 27936 34079
rect 28074 34076 28080 34128
rect 28132 34116 28138 34128
rect 30561 34119 30619 34125
rect 30561 34116 30573 34119
rect 28132 34088 30573 34116
rect 28132 34076 28138 34088
rect 30561 34085 30573 34088
rect 30607 34116 30619 34119
rect 31018 34116 31024 34128
rect 30607 34088 31024 34116
rect 30607 34085 30619 34088
rect 30561 34079 30619 34085
rect 31018 34076 31024 34088
rect 31076 34076 31082 34128
rect 31202 34076 31208 34128
rect 31260 34116 31266 34128
rect 31260 34088 31984 34116
rect 31260 34076 31266 34088
rect 31846 34048 31852 34060
rect 23992 34020 27936 34048
rect 28000 34020 31852 34048
rect 23992 34008 23998 34020
rect 22646 33940 22652 33992
rect 22704 33980 22710 33992
rect 22833 33983 22891 33989
rect 22833 33980 22845 33983
rect 22704 33952 22845 33980
rect 22704 33940 22710 33952
rect 22833 33949 22845 33952
rect 22879 33949 22891 33983
rect 22833 33943 22891 33949
rect 23014 33940 23020 33992
rect 23072 33980 23078 33992
rect 23845 33983 23903 33989
rect 23845 33980 23857 33983
rect 23072 33952 23857 33980
rect 23072 33940 23078 33952
rect 23845 33949 23857 33952
rect 23891 33949 23903 33983
rect 23845 33943 23903 33949
rect 24946 33940 24952 33992
rect 25004 33940 25010 33992
rect 25041 33983 25099 33989
rect 25041 33949 25053 33983
rect 25087 33980 25099 33983
rect 25314 33980 25320 33992
rect 25087 33952 25320 33980
rect 25087 33949 25099 33952
rect 25041 33943 25099 33949
rect 25314 33940 25320 33952
rect 25372 33940 25378 33992
rect 26053 33983 26111 33989
rect 26053 33949 26065 33983
rect 26099 33949 26111 33983
rect 26053 33943 26111 33949
rect 21039 33884 21864 33912
rect 22066 33884 22232 33912
rect 22296 33884 22600 33912
rect 21039 33881 21051 33884
rect 20993 33875 21051 33881
rect 15470 33844 15476 33856
rect 14108 33816 15476 33844
rect 15470 33804 15476 33816
rect 15528 33804 15534 33856
rect 16850 33804 16856 33856
rect 16908 33804 16914 33856
rect 16942 33804 16948 33856
rect 17000 33844 17006 33856
rect 17681 33847 17739 33853
rect 17681 33844 17693 33847
rect 17000 33816 17693 33844
rect 17000 33804 17006 33816
rect 17681 33813 17693 33816
rect 17727 33813 17739 33847
rect 17681 33807 17739 33813
rect 17957 33847 18015 33853
rect 17957 33813 17969 33847
rect 18003 33844 18015 33847
rect 18782 33844 18788 33856
rect 18003 33816 18788 33844
rect 18003 33813 18015 33816
rect 17957 33807 18015 33813
rect 18782 33804 18788 33816
rect 18840 33804 18846 33856
rect 18874 33804 18880 33856
rect 18932 33804 18938 33856
rect 20898 33804 20904 33856
rect 20956 33844 20962 33856
rect 21453 33847 21511 33853
rect 21453 33844 21465 33847
rect 20956 33816 21465 33844
rect 20956 33804 20962 33816
rect 21453 33813 21465 33816
rect 21499 33813 21511 33847
rect 21836 33844 21864 33884
rect 22296 33844 22324 33884
rect 22738 33872 22744 33924
rect 22796 33912 22802 33924
rect 23569 33915 23627 33921
rect 23569 33912 23581 33915
rect 22796 33884 23581 33912
rect 22796 33872 22802 33884
rect 23569 33881 23581 33884
rect 23615 33881 23627 33915
rect 23569 33875 23627 33881
rect 24118 33872 24124 33924
rect 24176 33912 24182 33924
rect 24394 33912 24400 33924
rect 24176 33884 24400 33912
rect 24176 33872 24182 33884
rect 24394 33872 24400 33884
rect 24452 33872 24458 33924
rect 24578 33872 24584 33924
rect 24636 33872 24642 33924
rect 25406 33872 25412 33924
rect 25464 33912 25470 33924
rect 26068 33912 26096 33943
rect 26142 33940 26148 33992
rect 26200 33940 26206 33992
rect 26234 33940 26240 33992
rect 26292 33940 26298 33992
rect 26329 33983 26387 33989
rect 26329 33949 26341 33983
rect 26375 33949 26387 33983
rect 26329 33943 26387 33949
rect 25464 33884 26096 33912
rect 26344 33912 26372 33943
rect 26418 33940 26424 33992
rect 26476 33980 26482 33992
rect 27065 33983 27123 33989
rect 27065 33980 27077 33983
rect 26476 33952 27077 33980
rect 26476 33940 26482 33952
rect 27065 33949 27077 33952
rect 27111 33949 27123 33983
rect 27065 33943 27123 33949
rect 27154 33940 27160 33992
rect 27212 33980 27218 33992
rect 27249 33983 27307 33989
rect 27249 33980 27261 33983
rect 27212 33952 27261 33980
rect 27212 33940 27218 33952
rect 27249 33949 27261 33952
rect 27295 33949 27307 33983
rect 27249 33943 27307 33949
rect 27341 33983 27399 33989
rect 27341 33949 27353 33983
rect 27387 33980 27399 33983
rect 27522 33980 27528 33992
rect 27387 33952 27528 33980
rect 27387 33949 27399 33952
rect 27341 33943 27399 33949
rect 27522 33940 27528 33952
rect 27580 33940 27586 33992
rect 27614 33940 27620 33992
rect 27672 33980 27678 33992
rect 28000 33980 28028 34020
rect 31846 34008 31852 34020
rect 31904 34008 31910 34060
rect 31956 34057 31984 34088
rect 32122 34076 32128 34128
rect 32180 34116 32186 34128
rect 32180 34088 33553 34116
rect 32180 34076 32186 34088
rect 31941 34051 31999 34057
rect 31941 34017 31953 34051
rect 31987 34017 31999 34051
rect 31941 34011 31999 34017
rect 32490 34008 32496 34060
rect 32548 34048 32554 34060
rect 32548 34020 33364 34048
rect 32548 34008 32554 34020
rect 27672 33952 28028 33980
rect 28077 33983 28135 33989
rect 27672 33940 27678 33952
rect 28077 33949 28089 33983
rect 28123 33949 28135 33983
rect 28077 33943 28135 33949
rect 26510 33912 26516 33924
rect 26344 33884 26516 33912
rect 25464 33872 25470 33884
rect 26510 33872 26516 33884
rect 26568 33912 26574 33924
rect 27798 33912 27804 33924
rect 26568 33884 27804 33912
rect 26568 33872 26574 33884
rect 27798 33872 27804 33884
rect 27856 33872 27862 33924
rect 27890 33872 27896 33924
rect 27948 33912 27954 33924
rect 28092 33912 28120 33943
rect 28166 33940 28172 33992
rect 28224 33940 28230 33992
rect 28537 33983 28595 33989
rect 28537 33949 28549 33983
rect 28583 33980 28595 33983
rect 28810 33980 28816 33992
rect 28583 33952 28816 33980
rect 28583 33949 28595 33952
rect 28537 33943 28595 33949
rect 28810 33940 28816 33952
rect 28868 33940 28874 33992
rect 28997 33983 29055 33989
rect 28997 33949 29009 33983
rect 29043 33980 29055 33983
rect 29086 33980 29092 33992
rect 29043 33952 29092 33980
rect 29043 33949 29055 33952
rect 28997 33943 29055 33949
rect 29086 33940 29092 33952
rect 29144 33940 29150 33992
rect 29181 33983 29239 33989
rect 29181 33949 29193 33983
rect 29227 33980 29239 33983
rect 29270 33980 29276 33992
rect 29227 33952 29276 33980
rect 29227 33949 29239 33952
rect 29181 33943 29239 33949
rect 29270 33940 29276 33952
rect 29328 33940 29334 33992
rect 29825 33983 29883 33989
rect 29825 33949 29837 33983
rect 29871 33949 29883 33983
rect 29825 33943 29883 33949
rect 27948 33884 28120 33912
rect 27948 33872 27954 33884
rect 28350 33872 28356 33924
rect 28408 33912 28414 33924
rect 28445 33915 28503 33921
rect 28445 33912 28457 33915
rect 28408 33884 28457 33912
rect 28408 33872 28414 33884
rect 28445 33881 28457 33884
rect 28491 33881 28503 33915
rect 28445 33875 28503 33881
rect 28626 33872 28632 33924
rect 28684 33912 28690 33924
rect 29840 33912 29868 33943
rect 30282 33940 30288 33992
rect 30340 33940 30346 33992
rect 31202 33980 31208 33992
rect 30392 33952 31208 33980
rect 28684 33884 29868 33912
rect 28684 33872 28690 33884
rect 30006 33872 30012 33924
rect 30064 33872 30070 33924
rect 21836 33816 22324 33844
rect 21453 33807 21511 33813
rect 22370 33804 22376 33856
rect 22428 33804 22434 33856
rect 22554 33804 22560 33856
rect 22612 33844 22618 33856
rect 23014 33844 23020 33856
rect 22612 33816 23020 33844
rect 22612 33804 22618 33816
rect 23014 33804 23020 33816
rect 23072 33804 23078 33856
rect 23109 33847 23167 33853
rect 23109 33813 23121 33847
rect 23155 33844 23167 33847
rect 25590 33844 25596 33856
rect 23155 33816 25596 33844
rect 23155 33813 23167 33816
rect 23109 33807 23167 33813
rect 25590 33804 25596 33816
rect 25648 33804 25654 33856
rect 25682 33804 25688 33856
rect 25740 33844 25746 33856
rect 25869 33847 25927 33853
rect 25869 33844 25881 33847
rect 25740 33816 25881 33844
rect 25740 33804 25746 33816
rect 25869 33813 25881 33816
rect 25915 33813 25927 33847
rect 25869 33807 25927 33813
rect 26881 33847 26939 33853
rect 26881 33813 26893 33847
rect 26927 33844 26939 33847
rect 27154 33844 27160 33856
rect 26927 33816 27160 33844
rect 26927 33813 26939 33816
rect 26881 33807 26939 33813
rect 27154 33804 27160 33816
rect 27212 33804 27218 33856
rect 28166 33804 28172 33856
rect 28224 33844 28230 33856
rect 28718 33844 28724 33856
rect 28224 33816 28724 33844
rect 28224 33804 28230 33816
rect 28718 33804 28724 33816
rect 28776 33804 28782 33856
rect 29086 33804 29092 33856
rect 29144 33804 29150 33856
rect 29454 33804 29460 33856
rect 29512 33844 29518 33856
rect 30392 33844 30420 33952
rect 31202 33940 31208 33952
rect 31260 33940 31266 33992
rect 31386 33940 31392 33992
rect 31444 33940 31450 33992
rect 32858 33940 32864 33992
rect 32916 33980 32922 33992
rect 33226 33989 33232 33992
rect 33045 33983 33103 33989
rect 33045 33980 33057 33983
rect 32916 33952 33057 33980
rect 32916 33940 32922 33952
rect 33045 33949 33057 33952
rect 33091 33949 33103 33983
rect 33045 33943 33103 33949
rect 33183 33983 33232 33989
rect 33183 33949 33195 33983
rect 33229 33949 33232 33983
rect 33183 33943 33232 33949
rect 33198 33940 33232 33943
rect 33284 33940 33290 33992
rect 33336 33989 33364 34020
rect 33321 33983 33379 33989
rect 33321 33949 33333 33983
rect 33367 33949 33379 33983
rect 33321 33943 33379 33949
rect 33410 33940 33416 33992
rect 33468 33940 33474 33992
rect 33525 33989 33553 34088
rect 33686 34008 33692 34060
rect 33744 34048 33750 34060
rect 34241 34051 34299 34057
rect 34241 34048 34253 34051
rect 33744 34020 34253 34048
rect 33744 34008 33750 34020
rect 34241 34017 34253 34020
rect 34287 34017 34299 34051
rect 34624 34048 34652 34144
rect 34900 34128 34928 34156
rect 35710 34144 35716 34196
rect 35768 34184 35774 34196
rect 38286 34184 38292 34196
rect 35768 34156 38292 34184
rect 35768 34144 35774 34156
rect 38286 34144 38292 34156
rect 38344 34144 38350 34196
rect 34882 34076 34888 34128
rect 34940 34116 34946 34128
rect 34940 34088 35393 34116
rect 34940 34076 34946 34088
rect 34241 34011 34299 34017
rect 34348 34020 34652 34048
rect 33510 33983 33568 33989
rect 33510 33949 33522 33983
rect 33556 33949 33568 33983
rect 33510 33943 33568 33949
rect 30742 33872 30748 33924
rect 30800 33912 30806 33924
rect 33198 33912 33226 33940
rect 30800 33884 33226 33912
rect 33525 33912 33553 33943
rect 34054 33940 34060 33992
rect 34112 33980 34118 33992
rect 34348 33989 34376 34020
rect 35250 34008 35256 34060
rect 35308 34008 35314 34060
rect 34149 33983 34207 33989
rect 34149 33980 34161 33983
rect 34112 33952 34161 33980
rect 34112 33940 34118 33952
rect 34149 33949 34161 33952
rect 34195 33949 34207 33983
rect 34149 33943 34207 33949
rect 34333 33983 34391 33989
rect 34333 33949 34345 33983
rect 34379 33949 34391 33983
rect 34333 33943 34391 33949
rect 34514 33940 34520 33992
rect 34572 33980 34578 33992
rect 34885 33983 34943 33989
rect 34885 33980 34897 33983
rect 34572 33952 34897 33980
rect 34572 33940 34578 33952
rect 34885 33949 34897 33952
rect 34931 33949 34943 33983
rect 34885 33943 34943 33949
rect 35033 33983 35091 33989
rect 35033 33949 35045 33983
rect 35079 33980 35091 33983
rect 35268 33980 35296 34008
rect 35365 33989 35393 34088
rect 35710 34008 35716 34060
rect 35768 34008 35774 34060
rect 36078 34008 36084 34060
rect 36136 34048 36142 34060
rect 36814 34048 36820 34060
rect 36136 34020 36820 34048
rect 36136 34008 36142 34020
rect 36814 34008 36820 34020
rect 36872 34008 36878 34060
rect 35079 33952 35296 33980
rect 35350 33983 35408 33989
rect 35079 33949 35091 33952
rect 35033 33943 35091 33949
rect 35350 33949 35362 33983
rect 35396 33949 35408 33983
rect 35728 33980 35756 34008
rect 35350 33943 35408 33949
rect 35452 33952 35756 33980
rect 33686 33912 33692 33924
rect 33525 33884 33692 33912
rect 30800 33872 30806 33884
rect 33686 33872 33692 33884
rect 33744 33872 33750 33924
rect 35161 33915 35219 33921
rect 35161 33912 35173 33915
rect 34348 33884 35173 33912
rect 34348 33856 34376 33884
rect 35161 33881 35173 33884
rect 35207 33881 35219 33915
rect 35161 33875 35219 33881
rect 35253 33915 35311 33921
rect 35253 33881 35265 33915
rect 35299 33912 35311 33915
rect 35452 33912 35480 33952
rect 35986 33940 35992 33992
rect 36044 33940 36050 33992
rect 37090 33989 37096 33992
rect 36173 33983 36231 33989
rect 36173 33949 36185 33983
rect 36219 33949 36231 33983
rect 37084 33980 37096 33989
rect 37051 33952 37096 33980
rect 36173 33943 36231 33949
rect 37084 33943 37096 33952
rect 35299 33884 35480 33912
rect 35299 33881 35311 33884
rect 35253 33875 35311 33881
rect 35710 33872 35716 33924
rect 35768 33912 35774 33924
rect 36188 33912 36216 33943
rect 37090 33940 37096 33943
rect 37148 33940 37154 33992
rect 35768 33884 36216 33912
rect 35768 33872 35774 33884
rect 36262 33872 36268 33924
rect 36320 33912 36326 33924
rect 37826 33912 37832 33924
rect 36320 33884 37832 33912
rect 36320 33872 36326 33884
rect 37826 33872 37832 33884
rect 37884 33912 37890 33924
rect 37884 33884 38240 33912
rect 37884 33872 37890 33884
rect 29512 33816 30420 33844
rect 29512 33804 29518 33816
rect 30466 33804 30472 33856
rect 30524 33844 30530 33856
rect 33594 33844 33600 33856
rect 30524 33816 33600 33844
rect 30524 33804 30530 33816
rect 33594 33804 33600 33816
rect 33652 33804 33658 33856
rect 34330 33804 34336 33856
rect 34388 33804 34394 33856
rect 34606 33804 34612 33856
rect 34664 33844 34670 33856
rect 35529 33847 35587 33853
rect 35529 33844 35541 33847
rect 34664 33816 35541 33844
rect 34664 33804 34670 33816
rect 35529 33813 35541 33816
rect 35575 33813 35587 33847
rect 35529 33807 35587 33813
rect 35802 33804 35808 33856
rect 35860 33844 35866 33856
rect 36081 33847 36139 33853
rect 36081 33844 36093 33847
rect 35860 33816 36093 33844
rect 35860 33804 35866 33816
rect 36081 33813 36093 33816
rect 36127 33813 36139 33847
rect 36081 33807 36139 33813
rect 36170 33804 36176 33856
rect 36228 33844 36234 33856
rect 36446 33844 36452 33856
rect 36228 33816 36452 33844
rect 36228 33804 36234 33816
rect 36446 33804 36452 33816
rect 36504 33804 36510 33856
rect 38212 33853 38240 33884
rect 38197 33847 38255 33853
rect 38197 33813 38209 33847
rect 38243 33813 38255 33847
rect 38197 33807 38255 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 4525 33643 4583 33649
rect 4525 33609 4537 33643
rect 4571 33640 4583 33643
rect 4798 33640 4804 33652
rect 4571 33612 4804 33640
rect 4571 33609 4583 33612
rect 4525 33603 4583 33609
rect 4798 33600 4804 33612
rect 4856 33600 4862 33652
rect 4982 33600 4988 33652
rect 5040 33640 5046 33652
rect 8570 33640 8576 33652
rect 5040 33612 8576 33640
rect 5040 33600 5046 33612
rect 8570 33600 8576 33612
rect 8628 33600 8634 33652
rect 9585 33643 9643 33649
rect 9585 33640 9597 33643
rect 8772 33612 9597 33640
rect 3970 33532 3976 33584
rect 4028 33572 4034 33584
rect 7742 33572 7748 33584
rect 4028 33544 4108 33572
rect 4028 33532 4034 33544
rect 4080 33513 4108 33544
rect 4540 33544 7748 33572
rect 4540 33513 4568 33544
rect 7742 33532 7748 33544
rect 7800 33532 7806 33584
rect 7920 33575 7978 33581
rect 7920 33541 7932 33575
rect 7966 33572 7978 33575
rect 8772 33572 8800 33612
rect 9585 33609 9597 33612
rect 9631 33609 9643 33643
rect 9585 33603 9643 33609
rect 9950 33600 9956 33652
rect 10008 33600 10014 33652
rect 13446 33640 13452 33652
rect 11164 33612 13452 33640
rect 7966 33544 8800 33572
rect 7966 33541 7978 33544
rect 7920 33535 7978 33541
rect 8938 33532 8944 33584
rect 8996 33572 9002 33584
rect 10781 33575 10839 33581
rect 8996 33544 10732 33572
rect 8996 33532 9002 33544
rect 3881 33507 3939 33513
rect 3881 33473 3893 33507
rect 3927 33473 3939 33507
rect 3881 33467 3939 33473
rect 4065 33507 4123 33513
rect 4065 33473 4077 33507
rect 4111 33473 4123 33507
rect 4065 33467 4123 33473
rect 4341 33507 4399 33513
rect 4341 33473 4353 33507
rect 4387 33473 4399 33507
rect 4341 33467 4399 33473
rect 4525 33507 4583 33513
rect 4525 33473 4537 33507
rect 4571 33473 4583 33507
rect 4525 33467 4583 33473
rect 3896 33368 3924 33467
rect 4356 33436 4384 33467
rect 4798 33464 4804 33516
rect 4856 33504 4862 33516
rect 5169 33507 5227 33513
rect 5169 33504 5181 33507
rect 4856 33476 5181 33504
rect 4856 33464 4862 33476
rect 5169 33473 5181 33476
rect 5215 33473 5227 33507
rect 5169 33467 5227 33473
rect 5350 33464 5356 33516
rect 5408 33464 5414 33516
rect 5810 33464 5816 33516
rect 5868 33464 5874 33516
rect 5997 33507 6055 33513
rect 5997 33473 6009 33507
rect 6043 33473 6055 33507
rect 5997 33467 6055 33473
rect 6825 33507 6883 33513
rect 6825 33473 6837 33507
rect 6871 33502 6883 33507
rect 7009 33507 7067 33513
rect 6871 33474 6960 33502
rect 6871 33473 6883 33474
rect 6825 33467 6883 33473
rect 4890 33436 4896 33448
rect 4356 33408 4896 33436
rect 4890 33396 4896 33408
rect 4948 33396 4954 33448
rect 5626 33396 5632 33448
rect 5684 33436 5690 33448
rect 6012 33436 6040 33467
rect 6546 33436 6552 33448
rect 5684 33408 6552 33436
rect 5684 33396 5690 33408
rect 6546 33396 6552 33408
rect 6604 33396 6610 33448
rect 6932 33436 6960 33474
rect 7009 33473 7021 33507
rect 7055 33504 7067 33507
rect 7098 33504 7104 33516
rect 7055 33476 7104 33504
rect 7055 33473 7067 33476
rect 7009 33467 7067 33473
rect 7098 33464 7104 33476
rect 7156 33464 7162 33516
rect 7561 33507 7619 33513
rect 7561 33473 7573 33507
rect 7607 33504 7619 33507
rect 8754 33504 8760 33516
rect 7607 33476 8760 33504
rect 7607 33473 7619 33476
rect 7561 33467 7619 33473
rect 7576 33436 7604 33467
rect 8754 33464 8760 33476
rect 8812 33464 8818 33516
rect 9490 33464 9496 33516
rect 9548 33504 9554 33516
rect 10704 33504 10732 33544
rect 10781 33541 10793 33575
rect 10827 33572 10839 33575
rect 11054 33572 11060 33584
rect 10827 33544 11060 33572
rect 10827 33541 10839 33544
rect 10781 33535 10839 33541
rect 11054 33532 11060 33544
rect 11112 33532 11118 33584
rect 11164 33581 11192 33612
rect 13446 33600 13452 33612
rect 13504 33600 13510 33652
rect 13538 33600 13544 33652
rect 13596 33640 13602 33652
rect 14918 33640 14924 33652
rect 13596 33612 14924 33640
rect 13596 33600 13602 33612
rect 14918 33600 14924 33612
rect 14976 33600 14982 33652
rect 15102 33600 15108 33652
rect 15160 33600 15166 33652
rect 15746 33640 15752 33652
rect 15203 33612 15752 33640
rect 11149 33575 11207 33581
rect 11149 33541 11161 33575
rect 11195 33541 11207 33575
rect 11149 33535 11207 33541
rect 12342 33532 12348 33584
rect 12400 33572 12406 33584
rect 12437 33575 12495 33581
rect 12437 33572 12449 33575
rect 12400 33544 12449 33572
rect 12400 33532 12406 33544
rect 12437 33541 12449 33544
rect 12483 33541 12495 33575
rect 12437 33535 12495 33541
rect 13262 33532 13268 33584
rect 13320 33572 13326 33584
rect 13320 33544 13932 33572
rect 13320 33532 13326 33544
rect 10962 33504 10968 33516
rect 9548 33476 10180 33504
rect 10704 33476 10968 33504
rect 9548 33464 9554 33476
rect 6932 33408 7604 33436
rect 7650 33396 7656 33448
rect 7708 33396 7714 33448
rect 8662 33396 8668 33448
rect 8720 33436 8726 33448
rect 9858 33436 9864 33448
rect 8720 33408 9864 33436
rect 8720 33396 8726 33408
rect 9858 33396 9864 33408
rect 9916 33396 9922 33448
rect 10042 33396 10048 33448
rect 10100 33396 10106 33448
rect 10152 33445 10180 33476
rect 10962 33464 10968 33476
rect 11020 33464 11026 33516
rect 11698 33464 11704 33516
rect 11756 33464 11762 33516
rect 11882 33464 11888 33516
rect 11940 33504 11946 33516
rect 11977 33507 12035 33513
rect 11977 33504 11989 33507
rect 11940 33476 11989 33504
rect 11940 33464 11946 33476
rect 11977 33473 11989 33476
rect 12023 33473 12035 33507
rect 11977 33467 12035 33473
rect 12618 33464 12624 33516
rect 12676 33464 12682 33516
rect 13630 33504 13636 33516
rect 12728 33476 13636 33504
rect 10137 33439 10195 33445
rect 10137 33405 10149 33439
rect 10183 33405 10195 33439
rect 10137 33399 10195 33405
rect 10686 33396 10692 33448
rect 10744 33436 10750 33448
rect 12728 33436 12756 33476
rect 13630 33464 13636 33476
rect 13688 33504 13694 33516
rect 13904 33513 13932 33544
rect 14642 33532 14648 33584
rect 14700 33572 14706 33584
rect 15203 33572 15231 33612
rect 15746 33600 15752 33612
rect 15804 33600 15810 33652
rect 16942 33600 16948 33652
rect 17000 33600 17006 33652
rect 17402 33600 17408 33652
rect 17460 33600 17466 33652
rect 17586 33600 17592 33652
rect 17644 33640 17650 33652
rect 17862 33640 17868 33652
rect 17644 33612 17868 33640
rect 17644 33600 17650 33612
rect 17862 33600 17868 33612
rect 17920 33600 17926 33652
rect 18874 33600 18880 33652
rect 18932 33640 18938 33652
rect 21266 33640 21272 33652
rect 18932 33612 21272 33640
rect 18932 33600 18938 33612
rect 21266 33600 21272 33612
rect 21324 33600 21330 33652
rect 21450 33600 21456 33652
rect 21508 33600 21514 33652
rect 22186 33600 22192 33652
rect 22244 33640 22250 33652
rect 24118 33640 24124 33652
rect 22244 33612 24124 33640
rect 22244 33600 22250 33612
rect 24118 33600 24124 33612
rect 24176 33600 24182 33652
rect 27246 33640 27252 33652
rect 25056 33612 27252 33640
rect 15473 33575 15531 33581
rect 15473 33572 15485 33575
rect 14700 33544 15231 33572
rect 15304 33544 15485 33572
rect 14700 33532 14706 33544
rect 13725 33507 13783 33513
rect 13725 33504 13737 33507
rect 13688 33476 13737 33504
rect 13688 33464 13694 33476
rect 13725 33473 13737 33476
rect 13771 33473 13783 33507
rect 13904 33507 13967 33513
rect 13904 33482 13921 33507
rect 13725 33467 13783 33473
rect 13909 33473 13921 33482
rect 13955 33473 13967 33507
rect 13909 33467 13967 33473
rect 13998 33464 14004 33516
rect 14056 33464 14062 33516
rect 14550 33464 14556 33516
rect 14608 33504 14614 33516
rect 15102 33504 15108 33516
rect 14608 33476 15108 33504
rect 14608 33464 14614 33476
rect 15102 33464 15108 33476
rect 15160 33464 15166 33516
rect 10744 33408 12756 33436
rect 10744 33396 10750 33408
rect 13170 33396 13176 33448
rect 13228 33436 13234 33448
rect 13538 33436 13544 33448
rect 13228 33408 13544 33436
rect 13228 33396 13234 33408
rect 13538 33396 13544 33408
rect 13596 33396 13602 33448
rect 13814 33396 13820 33448
rect 13872 33396 13878 33448
rect 7193 33371 7251 33377
rect 7193 33368 7205 33371
rect 3896 33340 7205 33368
rect 7193 33337 7205 33340
rect 7239 33368 7251 33371
rect 7282 33368 7288 33380
rect 7239 33340 7288 33368
rect 7239 33337 7251 33340
rect 7193 33331 7251 33337
rect 7282 33328 7288 33340
rect 7340 33328 7346 33380
rect 7374 33328 7380 33380
rect 7432 33368 7438 33380
rect 7668 33368 7696 33396
rect 7432 33340 7696 33368
rect 9033 33371 9091 33377
rect 7432 33328 7438 33340
rect 9033 33337 9045 33371
rect 9079 33368 9091 33371
rect 9950 33368 9956 33380
rect 9079 33340 9956 33368
rect 9079 33337 9091 33340
rect 9033 33331 9091 33337
rect 9950 33328 9956 33340
rect 10008 33328 10014 33380
rect 11793 33371 11851 33377
rect 11793 33337 11805 33371
rect 11839 33368 11851 33371
rect 12066 33368 12072 33380
rect 11839 33340 12072 33368
rect 11839 33337 11851 33340
rect 11793 33331 11851 33337
rect 12066 33328 12072 33340
rect 12124 33328 12130 33380
rect 14274 33328 14280 33380
rect 14332 33368 14338 33380
rect 15304 33368 15332 33544
rect 15473 33541 15485 33544
rect 15519 33541 15531 33575
rect 15473 33535 15531 33541
rect 15562 33532 15568 33584
rect 15620 33532 15626 33584
rect 15654 33532 15660 33584
rect 15712 33572 15718 33584
rect 17313 33575 17371 33581
rect 17313 33572 17325 33575
rect 15712 33544 17325 33572
rect 15712 33532 15718 33544
rect 17313 33541 17325 33544
rect 17359 33541 17371 33575
rect 20070 33572 20076 33584
rect 17313 33535 17371 33541
rect 18708 33544 20076 33572
rect 15381 33507 15439 33513
rect 15381 33473 15393 33507
rect 15427 33473 15439 33507
rect 15381 33467 15439 33473
rect 14332 33340 15332 33368
rect 15396 33368 15424 33467
rect 15746 33464 15752 33516
rect 15804 33464 15810 33516
rect 15841 33507 15899 33513
rect 15841 33473 15853 33507
rect 15887 33504 15899 33507
rect 15930 33504 15936 33516
rect 15887 33476 15936 33504
rect 15887 33473 15899 33476
rect 15841 33467 15899 33473
rect 15930 33464 15936 33476
rect 15988 33464 15994 33516
rect 16482 33464 16488 33516
rect 16540 33504 16546 33516
rect 17221 33507 17279 33513
rect 17221 33504 17233 33507
rect 16540 33476 17233 33504
rect 16540 33464 16546 33476
rect 17221 33473 17233 33476
rect 17267 33473 17279 33507
rect 17221 33467 17279 33473
rect 17586 33464 17592 33516
rect 17644 33504 17650 33516
rect 17644 33476 17816 33504
rect 17644 33464 17650 33476
rect 15764 33436 15792 33464
rect 16942 33436 16948 33448
rect 15764 33408 16948 33436
rect 16942 33396 16948 33408
rect 17000 33436 17006 33448
rect 17678 33436 17684 33448
rect 17000 33408 17684 33436
rect 17000 33396 17006 33408
rect 17678 33396 17684 33408
rect 17736 33396 17742 33448
rect 17788 33436 17816 33476
rect 18414 33464 18420 33516
rect 18472 33504 18478 33516
rect 18509 33507 18567 33513
rect 18509 33504 18521 33507
rect 18472 33476 18521 33504
rect 18472 33464 18478 33476
rect 18509 33473 18521 33476
rect 18555 33473 18567 33507
rect 18509 33467 18567 33473
rect 18601 33439 18659 33445
rect 18601 33436 18613 33439
rect 17788 33408 18613 33436
rect 18601 33405 18613 33408
rect 18647 33405 18659 33439
rect 18601 33399 18659 33405
rect 17402 33368 17408 33380
rect 15396 33340 17408 33368
rect 14332 33328 14338 33340
rect 3878 33260 3884 33312
rect 3936 33260 3942 33312
rect 4798 33260 4804 33312
rect 4856 33260 4862 33312
rect 4890 33260 4896 33312
rect 4948 33300 4954 33312
rect 5261 33303 5319 33309
rect 5261 33300 5273 33303
rect 4948 33272 5273 33300
rect 4948 33260 4954 33272
rect 5261 33269 5273 33272
rect 5307 33269 5319 33303
rect 5261 33263 5319 33269
rect 5810 33260 5816 33312
rect 5868 33260 5874 33312
rect 6546 33260 6552 33312
rect 6604 33300 6610 33312
rect 6822 33300 6828 33312
rect 6604 33272 6828 33300
rect 6604 33260 6610 33272
rect 6822 33260 6828 33272
rect 6880 33260 6886 33312
rect 8570 33260 8576 33312
rect 8628 33300 8634 33312
rect 10134 33300 10140 33312
rect 8628 33272 10140 33300
rect 8628 33260 8634 33272
rect 10134 33260 10140 33272
rect 10192 33260 10198 33312
rect 11698 33260 11704 33312
rect 11756 33260 11762 33312
rect 12713 33303 12771 33309
rect 12713 33269 12725 33303
rect 12759 33300 12771 33303
rect 12802 33300 12808 33312
rect 12759 33272 12808 33300
rect 12759 33269 12771 33272
rect 12713 33263 12771 33269
rect 12802 33260 12808 33272
rect 12860 33260 12866 33312
rect 13722 33260 13728 33312
rect 13780 33300 13786 33312
rect 13814 33300 13820 33312
rect 13780 33272 13820 33300
rect 13780 33260 13786 33272
rect 13814 33260 13820 33272
rect 13872 33300 13878 33312
rect 15010 33300 15016 33312
rect 13872 33272 15016 33300
rect 13872 33260 13878 33272
rect 15010 33260 15016 33272
rect 15068 33260 15074 33312
rect 15304 33300 15332 33340
rect 17402 33328 17408 33340
rect 17460 33328 17466 33380
rect 18708 33368 18736 33544
rect 20070 33532 20076 33544
rect 20128 33532 20134 33584
rect 23661 33575 23719 33581
rect 23661 33541 23673 33575
rect 23707 33572 23719 33575
rect 24854 33572 24860 33584
rect 23707 33544 24860 33572
rect 23707 33541 23719 33544
rect 23661 33535 23719 33541
rect 22005 33529 22063 33535
rect 24854 33532 24860 33544
rect 24912 33532 24918 33584
rect 25056 33572 25084 33612
rect 27246 33600 27252 33612
rect 27304 33600 27310 33652
rect 27338 33600 27344 33652
rect 27396 33640 27402 33652
rect 28537 33643 28595 33649
rect 28537 33640 28549 33643
rect 27396 33612 28549 33640
rect 27396 33600 27402 33612
rect 28537 33609 28549 33612
rect 28583 33609 28595 33643
rect 28537 33603 28595 33609
rect 30190 33600 30196 33652
rect 30248 33600 30254 33652
rect 30558 33600 30564 33652
rect 30616 33600 30622 33652
rect 32858 33600 32864 33652
rect 32916 33640 32922 33652
rect 32916 33612 35480 33640
rect 32916 33600 32922 33612
rect 24964 33544 25084 33572
rect 22005 33526 22017 33529
rect 21940 33516 22017 33526
rect 19797 33507 19855 33513
rect 19797 33473 19809 33507
rect 19843 33504 19855 33507
rect 20438 33504 20444 33516
rect 19843 33476 20444 33504
rect 19843 33473 19855 33476
rect 19797 33467 19855 33473
rect 20438 33464 20444 33476
rect 20496 33464 20502 33516
rect 20993 33507 21051 33513
rect 20993 33473 21005 33507
rect 21039 33473 21051 33507
rect 20993 33467 21051 33473
rect 21269 33507 21327 33513
rect 21269 33473 21281 33507
rect 21315 33504 21327 33507
rect 21450 33504 21456 33516
rect 21315 33476 21456 33504
rect 21315 33473 21327 33476
rect 21269 33467 21327 33473
rect 19426 33396 19432 33448
rect 19484 33436 19490 33448
rect 19981 33439 20039 33445
rect 19981 33436 19993 33439
rect 19484 33408 19993 33436
rect 19484 33396 19490 33408
rect 19981 33405 19993 33408
rect 20027 33405 20039 33439
rect 19981 33399 20039 33405
rect 20254 33368 20260 33380
rect 17512 33340 18736 33368
rect 18800 33340 20260 33368
rect 17512 33300 17540 33340
rect 15304 33272 17540 33300
rect 17589 33303 17647 33309
rect 17589 33269 17601 33303
rect 17635 33300 17647 33303
rect 17770 33300 17776 33312
rect 17635 33272 17776 33300
rect 17635 33269 17647 33272
rect 17589 33263 17647 33269
rect 17770 33260 17776 33272
rect 17828 33260 17834 33312
rect 17954 33260 17960 33312
rect 18012 33300 18018 33312
rect 18693 33303 18751 33309
rect 18693 33300 18705 33303
rect 18012 33272 18705 33300
rect 18012 33260 18018 33272
rect 18693 33269 18705 33272
rect 18739 33300 18751 33303
rect 18800 33300 18828 33340
rect 20254 33328 20260 33340
rect 20312 33328 20318 33380
rect 21008 33368 21036 33467
rect 21450 33464 21456 33476
rect 21508 33464 21514 33516
rect 21910 33464 21916 33516
rect 21968 33498 22017 33516
rect 21968 33464 21974 33498
rect 22005 33495 22017 33498
rect 22051 33495 22063 33529
rect 22005 33489 22063 33495
rect 22189 33507 22247 33513
rect 22189 33473 22201 33507
rect 22235 33473 22247 33507
rect 22189 33467 22247 33473
rect 21082 33396 21088 33448
rect 21140 33396 21146 33448
rect 22204 33436 22232 33467
rect 22278 33464 22284 33516
rect 22336 33464 22342 33516
rect 22373 33507 22431 33513
rect 22373 33473 22385 33507
rect 22419 33504 22431 33507
rect 22419 33476 22508 33504
rect 22419 33473 22431 33476
rect 22373 33467 22431 33473
rect 22480 33436 22508 33476
rect 22554 33464 22560 33516
rect 22612 33464 22618 33516
rect 22738 33464 22744 33516
rect 22796 33504 22802 33516
rect 23290 33504 23296 33516
rect 22796 33476 23296 33504
rect 22796 33464 22802 33476
rect 23290 33464 23296 33476
rect 23348 33464 23354 33516
rect 23937 33507 23995 33513
rect 23937 33504 23949 33507
rect 23584 33476 23949 33504
rect 23584 33448 23612 33476
rect 23937 33473 23949 33476
rect 23983 33473 23995 33507
rect 23937 33467 23995 33473
rect 24026 33464 24032 33516
rect 24084 33504 24090 33516
rect 24578 33504 24584 33516
rect 24084 33476 24584 33504
rect 24084 33464 24090 33476
rect 24578 33464 24584 33476
rect 24636 33464 24642 33516
rect 24964 33513 24992 33544
rect 25682 33532 25688 33584
rect 25740 33532 25746 33584
rect 27157 33575 27215 33581
rect 27157 33541 27169 33575
rect 27203 33572 27215 33575
rect 28902 33572 28908 33584
rect 27203 33544 28908 33572
rect 27203 33541 27215 33544
rect 27157 33535 27215 33541
rect 28902 33532 28908 33544
rect 28960 33532 28966 33584
rect 29365 33575 29423 33581
rect 29365 33541 29377 33575
rect 29411 33572 29423 33575
rect 29638 33572 29644 33584
rect 29411 33544 29644 33572
rect 29411 33541 29423 33544
rect 29365 33535 29423 33541
rect 24949 33507 25007 33513
rect 24949 33473 24961 33507
rect 24995 33473 25007 33507
rect 24949 33467 25007 33473
rect 25038 33464 25044 33516
rect 25096 33464 25102 33516
rect 25590 33464 25596 33516
rect 25648 33504 25654 33516
rect 25648 33476 26096 33504
rect 25648 33464 25654 33476
rect 23198 33436 23204 33448
rect 22204 33408 22324 33436
rect 22480 33408 23204 33436
rect 22296 33380 22324 33408
rect 23198 33396 23204 33408
rect 23256 33396 23262 33448
rect 23566 33396 23572 33448
rect 23624 33396 23630 33448
rect 23753 33439 23811 33445
rect 23753 33405 23765 33439
rect 23799 33436 23811 33439
rect 23842 33436 23848 33448
rect 23799 33408 23848 33436
rect 23799 33405 23811 33408
rect 23753 33399 23811 33405
rect 23842 33396 23848 33408
rect 23900 33396 23906 33448
rect 24118 33396 24124 33448
rect 24176 33436 24182 33448
rect 25682 33436 25688 33448
rect 24176 33408 25688 33436
rect 24176 33396 24182 33408
rect 25682 33396 25688 33408
rect 25740 33396 25746 33448
rect 25866 33396 25872 33448
rect 25924 33436 25930 33448
rect 25961 33439 26019 33445
rect 25961 33436 25973 33439
rect 25924 33408 25973 33436
rect 25924 33396 25930 33408
rect 25961 33405 25973 33408
rect 26007 33405 26019 33439
rect 26068 33436 26096 33476
rect 26142 33464 26148 33516
rect 26200 33464 26206 33516
rect 26786 33464 26792 33516
rect 26844 33504 26850 33516
rect 27430 33504 27436 33516
rect 26844 33476 27436 33504
rect 26844 33464 26850 33476
rect 27430 33464 27436 33476
rect 27488 33464 27494 33516
rect 27522 33464 27528 33516
rect 27580 33504 27586 33516
rect 28169 33507 28227 33513
rect 28169 33504 28181 33507
rect 27580 33476 28181 33504
rect 27580 33464 27586 33476
rect 28169 33473 28181 33476
rect 28215 33504 28227 33507
rect 29380 33504 29408 33535
rect 29638 33532 29644 33544
rect 29696 33532 29702 33584
rect 29822 33532 29828 33584
rect 29880 33572 29886 33584
rect 29880 33544 30972 33572
rect 29880 33532 29886 33544
rect 28215 33476 29408 33504
rect 29549 33507 29607 33513
rect 28215 33473 28227 33476
rect 28169 33467 28227 33473
rect 29549 33473 29561 33507
rect 29595 33504 29607 33507
rect 30006 33504 30012 33516
rect 29595 33476 30012 33504
rect 29595 33473 29607 33476
rect 29549 33467 29607 33473
rect 30006 33464 30012 33476
rect 30064 33464 30070 33516
rect 30374 33504 30380 33516
rect 30116 33476 30380 33504
rect 27249 33439 27307 33445
rect 27249 33436 27261 33439
rect 26068 33408 27261 33436
rect 25961 33399 26019 33405
rect 27249 33405 27261 33408
rect 27295 33436 27307 33439
rect 27295 33408 27752 33436
rect 27295 33405 27307 33408
rect 27249 33399 27307 33405
rect 22002 33368 22008 33380
rect 21008 33340 22008 33368
rect 22002 33328 22008 33340
rect 22060 33328 22066 33380
rect 22278 33328 22284 33380
rect 22336 33368 22342 33380
rect 22462 33368 22468 33380
rect 22336 33340 22468 33368
rect 22336 33328 22342 33340
rect 22462 33328 22468 33340
rect 22520 33328 22526 33380
rect 23474 33328 23480 33380
rect 23532 33368 23538 33380
rect 27617 33371 27675 33377
rect 27617 33368 27629 33371
rect 23532 33340 27629 33368
rect 23532 33328 23538 33340
rect 27617 33337 27629 33340
rect 27663 33337 27675 33371
rect 27724 33368 27752 33408
rect 27890 33396 27896 33448
rect 27948 33436 27954 33448
rect 28261 33439 28319 33445
rect 28261 33436 28273 33439
rect 27948 33408 28273 33436
rect 27948 33396 27954 33408
rect 28261 33405 28273 33408
rect 28307 33436 28319 33439
rect 30116 33436 30144 33476
rect 30374 33464 30380 33476
rect 30432 33504 30438 33516
rect 30944 33513 30972 33544
rect 32490 33532 32496 33584
rect 32548 33572 32554 33584
rect 33134 33572 33140 33584
rect 32548 33544 33140 33572
rect 32548 33532 32554 33544
rect 33134 33532 33140 33544
rect 33192 33532 33198 33584
rect 33686 33572 33692 33584
rect 33520 33544 33692 33572
rect 30837 33507 30895 33513
rect 30837 33504 30849 33507
rect 30432 33476 30849 33504
rect 30432 33464 30438 33476
rect 30837 33473 30849 33476
rect 30883 33473 30895 33507
rect 30837 33467 30895 33473
rect 30929 33507 30987 33513
rect 30929 33473 30941 33507
rect 30975 33473 30987 33507
rect 30929 33467 30987 33473
rect 31018 33464 31024 33516
rect 31076 33464 31082 33516
rect 31205 33507 31263 33513
rect 31205 33473 31217 33507
rect 31251 33473 31263 33507
rect 31205 33467 31263 33473
rect 28307 33408 30144 33436
rect 28307 33405 28319 33408
rect 28261 33399 28319 33405
rect 30190 33396 30196 33448
rect 30248 33436 30254 33448
rect 31220 33436 31248 33467
rect 32858 33464 32864 33516
rect 32916 33464 32922 33516
rect 33009 33507 33067 33513
rect 33009 33473 33021 33507
rect 33055 33504 33067 33507
rect 33237 33507 33295 33513
rect 33055 33473 33088 33504
rect 33009 33467 33088 33473
rect 33237 33473 33249 33507
rect 33283 33473 33295 33507
rect 33237 33467 33295 33473
rect 33326 33507 33384 33513
rect 33326 33473 33338 33507
rect 33372 33504 33384 33507
rect 33520 33504 33548 33544
rect 33686 33532 33692 33544
rect 33744 33532 33750 33584
rect 34164 33544 34652 33572
rect 33870 33504 33876 33516
rect 33372 33476 33548 33504
rect 33704 33476 33876 33504
rect 33372 33473 33384 33476
rect 33326 33467 33384 33473
rect 33060 33436 33088 33467
rect 30248 33408 31248 33436
rect 32969 33408 33088 33436
rect 33249 33436 33277 33467
rect 33704 33448 33732 33476
rect 33870 33464 33876 33476
rect 33928 33464 33934 33516
rect 34164 33513 34192 33544
rect 33965 33507 34023 33513
rect 33965 33473 33977 33507
rect 34011 33473 34023 33507
rect 33965 33467 34023 33473
rect 34113 33507 34192 33513
rect 34113 33473 34125 33507
rect 34159 33476 34192 33507
rect 34159 33473 34171 33476
rect 34113 33467 34171 33473
rect 33686 33436 33692 33448
rect 33249 33408 33692 33436
rect 30248 33396 30254 33408
rect 32582 33368 32588 33380
rect 27724 33340 32588 33368
rect 27617 33331 27675 33337
rect 32582 33328 32588 33340
rect 32640 33328 32646 33380
rect 18739 33272 18828 33300
rect 18739 33269 18751 33272
rect 18693 33263 18751 33269
rect 18874 33260 18880 33312
rect 18932 33260 18938 33312
rect 21174 33260 21180 33312
rect 21232 33260 21238 33312
rect 21266 33260 21272 33312
rect 21324 33300 21330 33312
rect 22094 33300 22100 33312
rect 21324 33272 22100 33300
rect 21324 33260 21330 33272
rect 22094 33260 22100 33272
rect 22152 33260 22158 33312
rect 22741 33303 22799 33309
rect 22741 33269 22753 33303
rect 22787 33300 22799 33303
rect 22922 33300 22928 33312
rect 22787 33272 22928 33300
rect 22787 33269 22799 33272
rect 22741 33263 22799 33269
rect 22922 33260 22928 33272
rect 22980 33260 22986 33312
rect 23937 33303 23995 33309
rect 23937 33269 23949 33303
rect 23983 33300 23995 33303
rect 24026 33300 24032 33312
rect 23983 33272 24032 33300
rect 23983 33269 23995 33272
rect 23937 33263 23995 33269
rect 24026 33260 24032 33272
rect 24084 33260 24090 33312
rect 24121 33303 24179 33309
rect 24121 33269 24133 33303
rect 24167 33300 24179 33303
rect 24394 33300 24400 33312
rect 24167 33272 24400 33300
rect 24167 33269 24179 33272
rect 24121 33263 24179 33269
rect 24394 33260 24400 33272
rect 24452 33260 24458 33312
rect 25041 33303 25099 33309
rect 25041 33269 25053 33303
rect 25087 33300 25099 33303
rect 25130 33300 25136 33312
rect 25087 33272 25136 33300
rect 25087 33269 25099 33272
rect 25041 33263 25099 33269
rect 25130 33260 25136 33272
rect 25188 33260 25194 33312
rect 25222 33260 25228 33312
rect 25280 33260 25286 33312
rect 25682 33260 25688 33312
rect 25740 33300 25746 33312
rect 25777 33303 25835 33309
rect 25777 33300 25789 33303
rect 25740 33272 25789 33300
rect 25740 33260 25746 33272
rect 25777 33269 25789 33272
rect 25823 33300 25835 33303
rect 26050 33300 26056 33312
rect 25823 33272 26056 33300
rect 25823 33269 25835 33272
rect 25777 33263 25835 33269
rect 26050 33260 26056 33272
rect 26108 33260 26114 33312
rect 26326 33260 26332 33312
rect 26384 33260 26390 33312
rect 27154 33260 27160 33312
rect 27212 33260 27218 33312
rect 27338 33260 27344 33312
rect 27396 33300 27402 33312
rect 27890 33300 27896 33312
rect 27396 33272 27896 33300
rect 27396 33260 27402 33272
rect 27890 33260 27896 33272
rect 27948 33260 27954 33312
rect 28166 33260 28172 33312
rect 28224 33260 28230 33312
rect 28626 33260 28632 33312
rect 28684 33300 28690 33312
rect 29270 33300 29276 33312
rect 28684 33272 29276 33300
rect 28684 33260 28690 33272
rect 29270 33260 29276 33272
rect 29328 33260 29334 33312
rect 29638 33260 29644 33312
rect 29696 33260 29702 33312
rect 30650 33260 30656 33312
rect 30708 33300 30714 33312
rect 32766 33300 32772 33312
rect 30708 33272 32772 33300
rect 30708 33260 30714 33272
rect 32766 33260 32772 33272
rect 32824 33260 32830 33312
rect 32969 33300 32997 33408
rect 33686 33396 33692 33408
rect 33744 33396 33750 33448
rect 33505 33371 33563 33377
rect 33505 33337 33517 33371
rect 33551 33368 33563 33371
rect 33980 33368 34008 33467
rect 34238 33464 34244 33516
rect 34296 33464 34302 33516
rect 34330 33464 34336 33516
rect 34388 33464 34394 33516
rect 34430 33507 34488 33513
rect 34430 33473 34442 33507
rect 34476 33473 34488 33507
rect 34624 33504 34652 33544
rect 34790 33532 34796 33584
rect 34848 33572 34854 33584
rect 35345 33575 35403 33581
rect 35345 33572 35357 33575
rect 34848 33544 35357 33572
rect 34848 33532 34854 33544
rect 35345 33541 35357 33544
rect 35391 33541 35403 33575
rect 35452 33572 35480 33612
rect 35618 33600 35624 33652
rect 35676 33600 35682 33652
rect 38286 33640 38292 33652
rect 37752 33612 38292 33640
rect 35802 33572 35808 33584
rect 35452 33544 35808 33572
rect 35345 33535 35403 33541
rect 35802 33532 35808 33544
rect 35860 33532 35866 33584
rect 37366 33572 37372 33584
rect 36096 33544 37372 33572
rect 34624 33476 35020 33504
rect 34430 33467 34488 33473
rect 34445 33436 34473 33467
rect 34882 33436 34888 33448
rect 33551 33340 34008 33368
rect 34072 33408 34888 33436
rect 33551 33337 33563 33340
rect 33505 33331 33563 33337
rect 34072 33312 34100 33408
rect 34882 33396 34888 33408
rect 34940 33396 34946 33448
rect 34422 33328 34428 33380
rect 34480 33368 34486 33380
rect 34992 33368 35020 33476
rect 35066 33464 35072 33516
rect 35124 33464 35130 33516
rect 35250 33464 35256 33516
rect 35308 33464 35314 33516
rect 36096 33513 36124 33544
rect 37366 33532 37372 33544
rect 37424 33532 37430 33584
rect 36262 33513 36268 33516
rect 35437 33507 35495 33513
rect 35437 33473 35449 33507
rect 35483 33473 35495 33507
rect 35437 33467 35495 33473
rect 36081 33507 36139 33513
rect 36081 33473 36093 33507
rect 36127 33473 36139 33507
rect 36081 33467 36139 33473
rect 36229 33507 36268 33513
rect 36229 33473 36241 33507
rect 36229 33467 36268 33473
rect 35452 33436 35480 33467
rect 36262 33464 36268 33467
rect 36320 33464 36326 33516
rect 36357 33507 36415 33513
rect 36357 33473 36369 33507
rect 36403 33473 36415 33507
rect 36357 33467 36415 33473
rect 35710 33436 35716 33448
rect 35452 33408 35716 33436
rect 35710 33396 35716 33408
rect 35768 33396 35774 33448
rect 35894 33396 35900 33448
rect 35952 33436 35958 33448
rect 36372 33436 36400 33467
rect 36446 33464 36452 33516
rect 36504 33464 36510 33516
rect 36630 33513 36636 33516
rect 36587 33507 36636 33513
rect 36587 33473 36599 33507
rect 36633 33473 36636 33507
rect 36587 33467 36636 33473
rect 36630 33464 36636 33467
rect 36688 33464 36694 33516
rect 37461 33507 37519 33513
rect 37461 33473 37473 33507
rect 37507 33473 37519 33507
rect 37461 33467 37519 33473
rect 35952 33408 36584 33436
rect 35952 33396 35958 33408
rect 36280 33380 36308 33408
rect 36556 33380 36584 33408
rect 36906 33396 36912 33448
rect 36964 33436 36970 33448
rect 37476 33436 37504 33467
rect 37642 33464 37648 33516
rect 37700 33464 37706 33516
rect 37752 33513 37780 33612
rect 38286 33600 38292 33612
rect 38344 33600 38350 33652
rect 37737 33507 37795 33513
rect 37737 33473 37749 33507
rect 37783 33473 37795 33507
rect 37737 33467 37795 33473
rect 37829 33507 37887 33513
rect 37829 33473 37841 33507
rect 37875 33504 37887 33507
rect 37918 33504 37924 33516
rect 37875 33476 37924 33504
rect 37875 33473 37887 33476
rect 37829 33467 37887 33473
rect 37918 33464 37924 33476
rect 37976 33464 37982 33516
rect 39390 33436 39396 33448
rect 36964 33408 39396 33436
rect 36964 33396 36970 33408
rect 39390 33396 39396 33408
rect 39448 33396 39454 33448
rect 36170 33368 36176 33380
rect 34480 33340 36176 33368
rect 34480 33328 34486 33340
rect 36170 33328 36176 33340
rect 36228 33328 36234 33380
rect 36262 33328 36268 33380
rect 36320 33328 36326 33380
rect 36538 33328 36544 33380
rect 36596 33328 36602 33380
rect 36648 33340 37412 33368
rect 33594 33300 33600 33312
rect 32969 33272 33600 33300
rect 33594 33260 33600 33272
rect 33652 33260 33658 33312
rect 34054 33260 34060 33312
rect 34112 33260 34118 33312
rect 34609 33303 34667 33309
rect 34609 33269 34621 33303
rect 34655 33300 34667 33303
rect 36648 33300 36676 33340
rect 37384 33312 37412 33340
rect 34655 33272 36676 33300
rect 34655 33269 34667 33272
rect 34609 33263 34667 33269
rect 36722 33260 36728 33312
rect 36780 33260 36786 33312
rect 37366 33260 37372 33312
rect 37424 33260 37430 33312
rect 38010 33260 38016 33312
rect 38068 33260 38074 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 7834 33096 7840 33108
rect 4540 33068 7840 33096
rect 4540 32901 4568 33068
rect 7834 33056 7840 33068
rect 7892 33056 7898 33108
rect 8113 33099 8171 33105
rect 8113 33065 8125 33099
rect 8159 33096 8171 33099
rect 10042 33096 10048 33108
rect 8159 33068 10048 33096
rect 8159 33065 8171 33068
rect 8113 33059 8171 33065
rect 10042 33056 10048 33068
rect 10100 33056 10106 33108
rect 10962 33056 10968 33108
rect 11020 33096 11026 33108
rect 11882 33096 11888 33108
rect 11020 33068 11888 33096
rect 11020 33056 11026 33068
rect 11882 33056 11888 33068
rect 11940 33056 11946 33108
rect 12618 33056 12624 33108
rect 12676 33096 12682 33108
rect 12894 33096 12900 33108
rect 12676 33068 12900 33096
rect 12676 33056 12682 33068
rect 12894 33056 12900 33068
rect 12952 33056 12958 33108
rect 13262 33056 13268 33108
rect 13320 33056 13326 33108
rect 13538 33056 13544 33108
rect 13596 33096 13602 33108
rect 13998 33096 14004 33108
rect 13596 33068 14004 33096
rect 13596 33056 13602 33068
rect 13998 33056 14004 33068
rect 14056 33056 14062 33108
rect 14369 33099 14427 33105
rect 14369 33065 14381 33099
rect 14415 33065 14427 33099
rect 14369 33059 14427 33065
rect 4614 32988 4620 33040
rect 4672 33028 4678 33040
rect 5813 33031 5871 33037
rect 5813 33028 5825 33031
rect 4672 33000 5825 33028
rect 4672 32988 4678 33000
rect 5813 32997 5825 33000
rect 5859 32997 5871 33031
rect 5813 32991 5871 32997
rect 6178 32988 6184 33040
rect 6236 33028 6242 33040
rect 6454 33028 6460 33040
rect 6236 33000 6460 33028
rect 6236 32988 6242 33000
rect 6454 32988 6460 33000
rect 6512 32988 6518 33040
rect 7653 33031 7711 33037
rect 7653 32997 7665 33031
rect 7699 33028 7711 33031
rect 8018 33028 8024 33040
rect 7699 33000 8024 33028
rect 7699 32997 7711 33000
rect 7653 32991 7711 32997
rect 8018 32988 8024 33000
rect 8076 32988 8082 33040
rect 8478 32988 8484 33040
rect 8536 33028 8542 33040
rect 11701 33031 11759 33037
rect 11701 33028 11713 33031
rect 8536 33000 11713 33028
rect 8536 32988 8542 33000
rect 11701 32997 11713 33000
rect 11747 32997 11759 33031
rect 11701 32991 11759 32997
rect 12158 32988 12164 33040
rect 12216 33028 12222 33040
rect 12805 33031 12863 33037
rect 12805 33028 12817 33031
rect 12216 33000 12817 33028
rect 12216 32988 12222 33000
rect 12805 32997 12817 33000
rect 12851 32997 12863 33031
rect 12805 32991 12863 32997
rect 13354 32988 13360 33040
rect 13412 33028 13418 33040
rect 14384 33028 14412 33059
rect 15286 33056 15292 33108
rect 15344 33056 15350 33108
rect 15565 33099 15623 33105
rect 15565 33065 15577 33099
rect 15611 33096 15623 33099
rect 15654 33096 15660 33108
rect 15611 33068 15660 33096
rect 15611 33065 15623 33068
rect 15565 33059 15623 33065
rect 15654 33056 15660 33068
rect 15712 33056 15718 33108
rect 15838 33056 15844 33108
rect 15896 33096 15902 33108
rect 16025 33099 16083 33105
rect 16025 33096 16037 33099
rect 15896 33068 16037 33096
rect 15896 33056 15902 33068
rect 16025 33065 16037 33068
rect 16071 33096 16083 33099
rect 16114 33096 16120 33108
rect 16071 33068 16120 33096
rect 16071 33065 16083 33068
rect 16025 33059 16083 33065
rect 16114 33056 16120 33068
rect 16172 33056 16178 33108
rect 16482 33056 16488 33108
rect 16540 33056 16546 33108
rect 17218 33056 17224 33108
rect 17276 33096 17282 33108
rect 17405 33099 17463 33105
rect 17405 33096 17417 33099
rect 17276 33068 17417 33096
rect 17276 33056 17282 33068
rect 17405 33065 17417 33068
rect 17451 33065 17463 33099
rect 17405 33059 17463 33065
rect 17589 33099 17647 33105
rect 17589 33065 17601 33099
rect 17635 33096 17647 33099
rect 17862 33096 17868 33108
rect 17635 33068 17868 33096
rect 17635 33065 17647 33068
rect 17589 33059 17647 33065
rect 17862 33056 17868 33068
rect 17920 33056 17926 33108
rect 18966 33056 18972 33108
rect 19024 33096 19030 33108
rect 19978 33096 19984 33108
rect 19024 33068 19984 33096
rect 19024 33056 19030 33068
rect 19978 33056 19984 33068
rect 20036 33056 20042 33108
rect 20346 33056 20352 33108
rect 20404 33056 20410 33108
rect 20622 33056 20628 33108
rect 20680 33096 20686 33108
rect 20680 33068 22324 33096
rect 20680 33056 20686 33068
rect 13412 33000 14412 33028
rect 15212 33000 16243 33028
rect 13412 32988 13418 33000
rect 5261 32963 5319 32969
rect 5261 32929 5273 32963
rect 5307 32960 5319 32963
rect 8202 32960 8208 32972
rect 5307 32932 8208 32960
rect 5307 32929 5319 32932
rect 5261 32923 5319 32929
rect 8202 32920 8208 32932
rect 8260 32920 8266 32972
rect 8570 32920 8576 32972
rect 8628 32920 8634 32972
rect 8662 32920 8668 32972
rect 8720 32920 8726 32972
rect 9214 32920 9220 32972
rect 9272 32960 9278 32972
rect 9401 32963 9459 32969
rect 9401 32960 9413 32963
rect 9272 32932 9413 32960
rect 9272 32920 9278 32932
rect 9401 32929 9413 32932
rect 9447 32929 9459 32963
rect 9401 32923 9459 32929
rect 9674 32920 9680 32972
rect 9732 32960 9738 32972
rect 11333 32963 11391 32969
rect 9732 32932 10824 32960
rect 9732 32920 9738 32932
rect 4525 32895 4583 32901
rect 4525 32861 4537 32895
rect 4571 32861 4583 32895
rect 4525 32855 4583 32861
rect 4709 32895 4767 32901
rect 4709 32861 4721 32895
rect 4755 32892 4767 32895
rect 4982 32892 4988 32904
rect 4755 32864 4988 32892
rect 4755 32861 4767 32864
rect 4709 32855 4767 32861
rect 4982 32852 4988 32864
rect 5040 32852 5046 32904
rect 5169 32895 5227 32901
rect 5169 32861 5181 32895
rect 5215 32892 5227 32895
rect 5353 32895 5411 32901
rect 5215 32864 5304 32892
rect 5215 32861 5227 32864
rect 5169 32855 5227 32861
rect 4617 32759 4675 32765
rect 4617 32725 4629 32759
rect 4663 32756 4675 32759
rect 5166 32756 5172 32768
rect 4663 32728 5172 32756
rect 4663 32725 4675 32728
rect 4617 32719 4675 32725
rect 5166 32716 5172 32728
rect 5224 32716 5230 32768
rect 5276 32756 5304 32864
rect 5353 32861 5365 32895
rect 5399 32861 5411 32895
rect 5353 32855 5411 32861
rect 5368 32824 5396 32855
rect 5626 32852 5632 32904
rect 5684 32852 5690 32904
rect 5718 32852 5724 32904
rect 5776 32892 5782 32904
rect 5813 32895 5871 32901
rect 5813 32892 5825 32895
rect 5776 32864 5825 32892
rect 5776 32852 5782 32864
rect 5813 32861 5825 32864
rect 5859 32861 5871 32895
rect 5813 32855 5871 32861
rect 5997 32895 6055 32901
rect 5997 32861 6009 32895
rect 6043 32892 6055 32895
rect 6362 32892 6368 32904
rect 6043 32864 6368 32892
rect 6043 32861 6055 32864
rect 5997 32855 6055 32861
rect 6362 32852 6368 32864
rect 6420 32852 6426 32904
rect 6454 32852 6460 32904
rect 6512 32892 6518 32904
rect 6549 32895 6607 32901
rect 6549 32892 6561 32895
rect 6512 32864 6561 32892
rect 6512 32852 6518 32864
rect 6549 32861 6561 32864
rect 6595 32861 6607 32895
rect 6549 32855 6607 32861
rect 6730 32852 6736 32904
rect 6788 32892 6794 32904
rect 6788 32864 6960 32892
rect 6788 32852 6794 32864
rect 5644 32824 5672 32852
rect 6932 32836 6960 32864
rect 7190 32852 7196 32904
rect 7248 32892 7254 32904
rect 7285 32895 7343 32901
rect 7285 32892 7297 32895
rect 7248 32864 7297 32892
rect 7248 32852 7254 32864
rect 7285 32861 7297 32864
rect 7331 32861 7343 32895
rect 7285 32855 7343 32861
rect 7834 32852 7840 32904
rect 7892 32892 7898 32904
rect 8297 32895 8355 32901
rect 8297 32892 8309 32895
rect 7892 32864 8309 32892
rect 7892 32852 7898 32864
rect 8297 32861 8309 32864
rect 8343 32861 8355 32895
rect 8297 32855 8355 32861
rect 8478 32852 8484 32904
rect 8536 32852 8542 32904
rect 8680 32892 8708 32920
rect 8588 32864 8708 32892
rect 6914 32824 6920 32836
rect 5368 32796 6920 32824
rect 6914 32784 6920 32796
rect 6972 32824 6978 32836
rect 7469 32827 7527 32833
rect 7469 32824 7481 32827
rect 6972 32796 7481 32824
rect 6972 32784 6978 32796
rect 7469 32793 7481 32796
rect 7515 32824 7527 32827
rect 7926 32824 7932 32836
rect 7515 32796 7932 32824
rect 7515 32793 7527 32796
rect 7469 32787 7527 32793
rect 7926 32784 7932 32796
rect 7984 32824 7990 32836
rect 8588 32824 8616 32864
rect 8846 32852 8852 32904
rect 8904 32892 8910 32904
rect 9309 32895 9367 32901
rect 9309 32892 9321 32895
rect 8904 32864 9321 32892
rect 8904 32852 8910 32864
rect 9309 32861 9321 32864
rect 9355 32861 9367 32895
rect 9309 32855 9367 32861
rect 9490 32852 9496 32904
rect 9548 32852 9554 32904
rect 9582 32852 9588 32904
rect 9640 32852 9646 32904
rect 10410 32852 10416 32904
rect 10468 32852 10474 32904
rect 10686 32852 10692 32904
rect 10744 32852 10750 32904
rect 9508 32824 9536 32852
rect 7984 32796 8616 32824
rect 9048 32796 9536 32824
rect 10796 32824 10824 32932
rect 11333 32929 11345 32963
rect 11379 32960 11391 32963
rect 11379 32932 12020 32960
rect 11379 32929 11391 32932
rect 11333 32923 11391 32929
rect 11422 32852 11428 32904
rect 11480 32892 11486 32904
rect 11517 32895 11575 32901
rect 11517 32892 11529 32895
rect 11480 32864 11529 32892
rect 11480 32852 11486 32864
rect 11517 32861 11529 32864
rect 11563 32861 11575 32895
rect 11517 32855 11575 32861
rect 11606 32852 11612 32904
rect 11664 32852 11670 32904
rect 11790 32852 11796 32904
rect 11848 32852 11854 32904
rect 11992 32892 12020 32932
rect 12066 32920 12072 32972
rect 12124 32960 12130 32972
rect 12437 32963 12495 32969
rect 12437 32960 12449 32963
rect 12124 32932 12449 32960
rect 12124 32920 12130 32932
rect 12437 32929 12449 32932
rect 12483 32929 12495 32963
rect 14090 32960 14096 32972
rect 12437 32923 12495 32929
rect 12544 32932 14096 32960
rect 12544 32892 12572 32932
rect 14090 32920 14096 32932
rect 14148 32920 14154 32972
rect 14369 32963 14427 32969
rect 14369 32929 14381 32963
rect 14415 32960 14427 32963
rect 14642 32960 14648 32972
rect 14415 32932 14648 32960
rect 14415 32929 14427 32932
rect 14369 32923 14427 32929
rect 14642 32920 14648 32932
rect 14700 32920 14706 32972
rect 15010 32920 15016 32972
rect 15068 32960 15074 32972
rect 15212 32969 15240 33000
rect 15197 32963 15255 32969
rect 15197 32960 15209 32963
rect 15068 32932 15209 32960
rect 15068 32920 15074 32932
rect 15197 32929 15209 32932
rect 15243 32929 15255 32963
rect 15746 32960 15752 32972
rect 15197 32923 15255 32929
rect 15304 32932 15752 32960
rect 11992 32864 12572 32892
rect 12621 32895 12679 32901
rect 12621 32861 12633 32895
rect 12667 32861 12679 32895
rect 12621 32855 12679 32861
rect 12342 32824 12348 32836
rect 10796 32796 12348 32824
rect 7984 32784 7990 32796
rect 5442 32756 5448 32768
rect 5276 32728 5448 32756
rect 5442 32716 5448 32728
rect 5500 32716 5506 32768
rect 6733 32759 6791 32765
rect 6733 32725 6745 32759
rect 6779 32756 6791 32759
rect 9048 32756 9076 32796
rect 9324 32768 9352 32796
rect 12342 32784 12348 32796
rect 12400 32784 12406 32836
rect 12434 32784 12440 32836
rect 12492 32824 12498 32836
rect 12636 32824 12664 32855
rect 12710 32852 12716 32904
rect 12768 32892 12774 32904
rect 13449 32895 13507 32901
rect 13449 32892 13461 32895
rect 12768 32864 13461 32892
rect 12768 32852 12774 32864
rect 13449 32861 13461 32864
rect 13495 32861 13507 32895
rect 13449 32855 13507 32861
rect 13538 32852 13544 32904
rect 13596 32892 13602 32904
rect 13725 32895 13783 32901
rect 13725 32892 13737 32895
rect 13596 32864 13737 32892
rect 13596 32852 13602 32864
rect 13725 32861 13737 32864
rect 13771 32892 13783 32895
rect 14182 32892 14188 32904
rect 13771 32864 14188 32892
rect 13771 32861 13783 32864
rect 13725 32855 13783 32861
rect 14182 32852 14188 32864
rect 14240 32852 14246 32904
rect 14277 32895 14335 32901
rect 14277 32861 14289 32895
rect 14323 32892 14335 32895
rect 15304 32892 15332 32932
rect 15746 32920 15752 32932
rect 15804 32960 15810 32972
rect 16117 32963 16175 32969
rect 16117 32960 16129 32963
rect 15804 32932 16129 32960
rect 15804 32920 15810 32932
rect 16117 32929 16129 32932
rect 16163 32929 16175 32963
rect 16117 32923 16175 32929
rect 14323 32864 15332 32892
rect 14323 32861 14335 32864
rect 14277 32855 14335 32861
rect 15378 32852 15384 32904
rect 15436 32852 15442 32904
rect 15470 32852 15476 32904
rect 15528 32892 15534 32904
rect 16025 32895 16083 32901
rect 16025 32892 16037 32895
rect 15528 32864 16037 32892
rect 15528 32852 15534 32864
rect 16025 32861 16037 32864
rect 16071 32861 16083 32895
rect 16215 32892 16243 33000
rect 17310 32988 17316 33040
rect 17368 33028 17374 33040
rect 17678 33028 17684 33040
rect 17368 33000 17684 33028
rect 17368 32988 17374 33000
rect 17678 32988 17684 33000
rect 17736 32988 17742 33040
rect 18414 32988 18420 33040
rect 18472 33028 18478 33040
rect 21591 33031 21649 33037
rect 21591 33028 21603 33031
rect 18472 33000 21603 33028
rect 18472 32988 18478 33000
rect 21591 32997 21603 33000
rect 21637 33028 21649 33031
rect 21818 33028 21824 33040
rect 21637 33000 21824 33028
rect 21637 32997 21649 33000
rect 21591 32991 21649 32997
rect 21818 32988 21824 33000
rect 21876 32988 21882 33040
rect 22094 33028 22100 33040
rect 22020 33000 22100 33028
rect 18874 32920 18880 32972
rect 18932 32960 18938 32972
rect 22020 32960 22048 33000
rect 22094 32988 22100 33000
rect 22152 32988 22158 33040
rect 22296 33028 22324 33068
rect 22370 33056 22376 33108
rect 22428 33096 22434 33108
rect 23569 33099 23627 33105
rect 23569 33096 23581 33099
rect 22428 33068 23581 33096
rect 22428 33056 22434 33068
rect 23569 33065 23581 33068
rect 23615 33065 23627 33099
rect 23569 33059 23627 33065
rect 23750 33056 23756 33108
rect 23808 33096 23814 33108
rect 24029 33099 24087 33105
rect 24029 33096 24041 33099
rect 23808 33068 24041 33096
rect 23808 33056 23814 33068
rect 24029 33065 24041 33068
rect 24075 33065 24087 33099
rect 24029 33059 24087 33065
rect 24486 33056 24492 33108
rect 24544 33096 24550 33108
rect 24544 33068 24993 33096
rect 24544 33056 24550 33068
rect 24581 33031 24639 33037
rect 24581 33028 24593 33031
rect 22296 33000 24593 33028
rect 24581 32997 24593 33000
rect 24627 32997 24639 33031
rect 24965 33028 24993 33068
rect 25038 33056 25044 33108
rect 25096 33096 25102 33108
rect 26421 33099 26479 33105
rect 26421 33096 26433 33099
rect 25096 33068 26433 33096
rect 25096 33056 25102 33068
rect 26421 33065 26433 33068
rect 26467 33096 26479 33099
rect 26694 33096 26700 33108
rect 26467 33068 26700 33096
rect 26467 33065 26479 33068
rect 26421 33059 26479 33065
rect 26694 33056 26700 33068
rect 26752 33056 26758 33108
rect 27617 33099 27675 33105
rect 27617 33065 27629 33099
rect 27663 33096 27675 33099
rect 27663 33068 28304 33096
rect 27663 33065 27675 33068
rect 27617 33059 27675 33065
rect 25222 33028 25228 33040
rect 24965 33000 25228 33028
rect 24581 32991 24639 32997
rect 25222 32988 25228 33000
rect 25280 32988 25286 33040
rect 25314 32988 25320 33040
rect 25372 33028 25378 33040
rect 25866 33028 25872 33040
rect 25372 33000 25872 33028
rect 25372 32988 25378 33000
rect 25866 32988 25872 33000
rect 25924 32988 25930 33040
rect 26329 33031 26387 33037
rect 26329 32997 26341 33031
rect 26375 33028 26387 33031
rect 26786 33028 26792 33040
rect 26375 33000 26792 33028
rect 26375 32997 26387 33000
rect 26329 32991 26387 32997
rect 26786 32988 26792 33000
rect 26844 32988 26850 33040
rect 27801 33031 27859 33037
rect 27801 32997 27813 33031
rect 27847 33028 27859 33031
rect 27890 33028 27896 33040
rect 27847 33000 27896 33028
rect 27847 32997 27859 33000
rect 27801 32991 27859 32997
rect 27890 32988 27896 33000
rect 27948 32988 27954 33040
rect 18932 32932 20208 32960
rect 18932 32920 18938 32932
rect 16301 32895 16359 32901
rect 16301 32892 16313 32895
rect 16215 32864 16313 32892
rect 16025 32855 16083 32861
rect 16301 32861 16313 32864
rect 16347 32861 16359 32895
rect 16301 32855 16359 32861
rect 16850 32852 16856 32904
rect 16908 32892 16914 32904
rect 17037 32895 17095 32901
rect 17037 32892 17049 32895
rect 16908 32864 17049 32892
rect 16908 32852 16914 32864
rect 17037 32861 17049 32864
rect 17083 32861 17095 32895
rect 17037 32855 17095 32861
rect 18049 32895 18107 32901
rect 18049 32861 18061 32895
rect 18095 32861 18107 32895
rect 18049 32855 18107 32861
rect 15105 32827 15163 32833
rect 15105 32824 15117 32827
rect 12492 32796 12664 32824
rect 12728 32796 15117 32824
rect 12492 32784 12498 32796
rect 6779 32728 9076 32756
rect 6779 32725 6791 32728
rect 6733 32719 6791 32725
rect 9122 32716 9128 32768
rect 9180 32716 9186 32768
rect 9306 32716 9312 32768
rect 9364 32716 9370 32768
rect 10410 32716 10416 32768
rect 10468 32756 10474 32768
rect 11790 32756 11796 32768
rect 10468 32728 11796 32756
rect 10468 32716 10474 32728
rect 11790 32716 11796 32728
rect 11848 32716 11854 32768
rect 11882 32716 11888 32768
rect 11940 32756 11946 32768
rect 12728 32756 12756 32796
rect 15105 32793 15117 32796
rect 15151 32793 15163 32827
rect 15105 32787 15163 32793
rect 15488 32796 15700 32824
rect 11940 32728 12756 32756
rect 11940 32716 11946 32728
rect 12894 32716 12900 32768
rect 12952 32756 12958 32768
rect 13633 32759 13691 32765
rect 13633 32756 13645 32759
rect 12952 32728 13645 32756
rect 12952 32716 12958 32728
rect 13633 32725 13645 32728
rect 13679 32756 13691 32759
rect 14182 32756 14188 32768
rect 13679 32728 14188 32756
rect 13679 32725 13691 32728
rect 13633 32719 13691 32725
rect 14182 32716 14188 32728
rect 14240 32716 14246 32768
rect 14274 32716 14280 32768
rect 14332 32756 14338 32768
rect 14645 32759 14703 32765
rect 14645 32756 14657 32759
rect 14332 32728 14657 32756
rect 14332 32716 14338 32728
rect 14645 32725 14657 32728
rect 14691 32756 14703 32759
rect 15488 32756 15516 32796
rect 14691 32728 15516 32756
rect 15672 32756 15700 32796
rect 17405 32759 17463 32765
rect 17405 32756 17417 32759
rect 15672 32728 17417 32756
rect 14691 32725 14703 32728
rect 14645 32719 14703 32725
rect 17405 32725 17417 32728
rect 17451 32725 17463 32759
rect 18064 32756 18092 32855
rect 19426 32852 19432 32904
rect 19484 32892 19490 32904
rect 20180 32901 20208 32932
rect 21744 32932 22048 32960
rect 22299 32932 22692 32960
rect 19797 32895 19855 32901
rect 19797 32892 19809 32895
rect 19484 32864 19809 32892
rect 19484 32852 19490 32864
rect 19797 32861 19809 32864
rect 19843 32861 19855 32895
rect 19797 32855 19855 32861
rect 20165 32895 20223 32901
rect 20165 32861 20177 32895
rect 20211 32861 20223 32895
rect 20165 32855 20223 32861
rect 20622 32852 20628 32904
rect 20680 32892 20686 32904
rect 20809 32895 20867 32901
rect 20809 32892 20821 32895
rect 20680 32864 20821 32892
rect 20680 32852 20686 32864
rect 20809 32861 20821 32864
rect 20855 32861 20867 32895
rect 20809 32855 20867 32861
rect 20993 32895 21051 32901
rect 20993 32861 21005 32895
rect 21039 32892 21051 32895
rect 21082 32892 21088 32904
rect 21039 32864 21088 32892
rect 21039 32861 21051 32864
rect 20993 32855 21051 32861
rect 21082 32852 21088 32864
rect 21140 32852 21146 32904
rect 21174 32852 21180 32904
rect 21232 32892 21238 32904
rect 21744 32901 21772 32932
rect 21442 32895 21500 32901
rect 21442 32892 21454 32895
rect 21232 32864 21454 32892
rect 21232 32852 21238 32864
rect 21442 32861 21454 32864
rect 21488 32861 21500 32895
rect 21442 32855 21500 32861
rect 21729 32895 21787 32901
rect 21729 32861 21741 32895
rect 21775 32861 21787 32895
rect 21729 32855 21787 32861
rect 21925 32892 21983 32895
rect 22299 32892 22327 32932
rect 21925 32889 22327 32892
rect 21925 32855 21937 32889
rect 21971 32864 22327 32889
rect 22557 32895 22615 32901
rect 21971 32855 21983 32864
rect 22557 32861 22569 32895
rect 22603 32861 22615 32895
rect 22557 32855 22615 32861
rect 21925 32849 21983 32855
rect 18322 32784 18328 32836
rect 18380 32784 18386 32836
rect 18414 32784 18420 32836
rect 18472 32824 18478 32836
rect 19981 32827 20039 32833
rect 19981 32824 19993 32827
rect 18472 32796 19993 32824
rect 18472 32784 18478 32796
rect 19981 32793 19993 32796
rect 20027 32793 20039 32827
rect 19981 32787 20039 32793
rect 20073 32827 20131 32833
rect 20073 32793 20085 32827
rect 20119 32824 20131 32827
rect 21266 32824 21272 32836
rect 20119 32796 21272 32824
rect 20119 32793 20131 32796
rect 20073 32787 20131 32793
rect 21266 32784 21272 32796
rect 21324 32784 21330 32836
rect 22572 32768 22600 32855
rect 22664 32824 22692 32932
rect 22738 32920 22744 32972
rect 22796 32920 22802 32972
rect 23750 32920 23756 32972
rect 23808 32960 23814 32972
rect 26878 32960 26884 32972
rect 23808 32932 26884 32960
rect 23808 32920 23814 32932
rect 26878 32920 26884 32932
rect 26936 32920 26942 32972
rect 28276 32960 28304 33068
rect 28350 33056 28356 33108
rect 28408 33096 28414 33108
rect 30466 33096 30472 33108
rect 28408 33068 30472 33096
rect 28408 33056 28414 33068
rect 30466 33056 30472 33068
rect 30524 33056 30530 33108
rect 30650 33056 30656 33108
rect 30708 33096 30714 33108
rect 30926 33096 30932 33108
rect 30708 33068 30932 33096
rect 30708 33056 30714 33068
rect 30926 33056 30932 33068
rect 30984 33056 30990 33108
rect 31389 33099 31447 33105
rect 31389 33065 31401 33099
rect 31435 33096 31447 33099
rect 32490 33096 32496 33108
rect 31435 33068 32496 33096
rect 31435 33065 31447 33068
rect 31389 33059 31447 33065
rect 32490 33056 32496 33068
rect 32548 33056 32554 33108
rect 33318 33056 33324 33108
rect 33376 33096 33382 33108
rect 33597 33099 33655 33105
rect 33376 33068 33548 33096
rect 33376 33056 33382 33068
rect 28442 32988 28448 33040
rect 28500 33028 28506 33040
rect 31754 33028 31760 33040
rect 28500 33000 31760 33028
rect 28500 32988 28506 33000
rect 31754 32988 31760 33000
rect 31812 32988 31818 33040
rect 32122 32988 32128 33040
rect 32180 33028 32186 33040
rect 32180 33000 33456 33028
rect 32180 32988 32186 33000
rect 28828 32960 28948 32968
rect 29362 32960 29368 32972
rect 28276 32949 28948 32960
rect 29006 32949 29368 32960
rect 28276 32940 29368 32949
rect 28276 32932 28856 32940
rect 28920 32932 29368 32940
rect 28920 32921 29034 32932
rect 29362 32920 29368 32932
rect 29420 32960 29426 32972
rect 29546 32960 29552 32972
rect 29420 32932 29552 32960
rect 29420 32920 29426 32932
rect 29546 32920 29552 32932
rect 29604 32920 29610 32972
rect 29730 32920 29736 32972
rect 29788 32960 29794 32972
rect 30009 32963 30067 32969
rect 30009 32960 30021 32963
rect 29788 32932 30021 32960
rect 29788 32920 29794 32932
rect 30009 32929 30021 32932
rect 30055 32929 30067 32963
rect 30009 32923 30067 32929
rect 30374 32920 30380 32972
rect 30432 32960 30438 32972
rect 31018 32960 31024 32972
rect 30432 32932 31024 32960
rect 30432 32920 30438 32932
rect 31018 32920 31024 32932
rect 31076 32920 31082 32972
rect 31478 32920 31484 32972
rect 31536 32960 31542 32972
rect 31536 32932 32444 32960
rect 31536 32920 31542 32932
rect 22833 32895 22891 32901
rect 22833 32861 22845 32895
rect 22879 32892 22891 32895
rect 23290 32892 23296 32904
rect 22879 32864 23296 32892
rect 22879 32861 22891 32864
rect 22833 32855 22891 32861
rect 23290 32852 23296 32864
rect 23348 32852 23354 32904
rect 23569 32895 23627 32901
rect 23569 32861 23581 32895
rect 23615 32892 23627 32895
rect 23658 32892 23664 32904
rect 23615 32864 23664 32892
rect 23615 32861 23627 32864
rect 23569 32855 23627 32861
rect 23658 32852 23664 32864
rect 23716 32852 23722 32904
rect 23842 32852 23848 32904
rect 23900 32892 23906 32904
rect 24394 32892 24400 32904
rect 23900 32864 24400 32892
rect 23900 32852 23906 32864
rect 24394 32852 24400 32864
rect 24452 32852 24458 32904
rect 24762 32852 24768 32904
rect 24820 32892 24826 32904
rect 24857 32895 24915 32901
rect 24857 32892 24869 32895
rect 24820 32864 24869 32892
rect 24820 32852 24826 32864
rect 24857 32861 24869 32864
rect 24903 32861 24915 32895
rect 24857 32855 24915 32861
rect 24946 32852 24952 32904
rect 25004 32852 25010 32904
rect 25038 32852 25044 32904
rect 25096 32852 25102 32904
rect 25222 32852 25228 32904
rect 25280 32852 25286 32904
rect 25961 32895 26019 32901
rect 25961 32861 25973 32895
rect 26007 32892 26019 32895
rect 26050 32892 26056 32904
rect 26007 32864 26056 32892
rect 26007 32861 26019 32864
rect 25961 32855 26019 32861
rect 26050 32852 26056 32864
rect 26108 32852 26114 32904
rect 27430 32852 27436 32904
rect 27488 32852 27494 32904
rect 27522 32852 27528 32904
rect 27580 32892 27586 32904
rect 28166 32892 28172 32904
rect 27580 32864 28172 32892
rect 27580 32852 27586 32864
rect 28166 32852 28172 32864
rect 28224 32852 28230 32904
rect 28350 32852 28356 32904
rect 28408 32852 28414 32904
rect 28810 32852 28816 32904
rect 28868 32852 28874 32904
rect 29917 32895 29975 32901
rect 29917 32861 29929 32895
rect 29963 32861 29975 32895
rect 29917 32855 29975 32861
rect 22922 32824 22928 32836
rect 22664 32796 22928 32824
rect 22922 32784 22928 32796
rect 22980 32784 22986 32836
rect 23474 32784 23480 32836
rect 23532 32824 23538 32836
rect 24670 32824 24676 32836
rect 23532 32796 24676 32824
rect 23532 32784 23538 32796
rect 24670 32784 24676 32796
rect 24728 32784 24734 32836
rect 25314 32784 25320 32836
rect 25372 32824 25378 32836
rect 29270 32824 29276 32836
rect 25372 32796 29276 32824
rect 25372 32784 25378 32796
rect 29270 32784 29276 32796
rect 29328 32784 29334 32836
rect 29730 32784 29736 32836
rect 29788 32824 29794 32836
rect 29932 32824 29960 32855
rect 30190 32852 30196 32904
rect 30248 32852 30254 32904
rect 31941 32895 31999 32901
rect 31941 32892 31953 32895
rect 30300 32864 31953 32892
rect 29788 32796 29960 32824
rect 29788 32784 29794 32796
rect 19058 32756 19064 32768
rect 18064 32728 19064 32756
rect 17405 32719 17463 32725
rect 19058 32716 19064 32728
rect 19116 32716 19122 32768
rect 19150 32716 19156 32768
rect 19208 32756 19214 32768
rect 20806 32756 20812 32768
rect 19208 32728 20812 32756
rect 19208 32716 19214 32728
rect 20806 32716 20812 32728
rect 20864 32716 20870 32768
rect 20898 32716 20904 32768
rect 20956 32716 20962 32768
rect 21450 32716 21456 32768
rect 21508 32756 21514 32768
rect 21821 32759 21879 32765
rect 21821 32756 21833 32759
rect 21508 32728 21833 32756
rect 21508 32716 21514 32728
rect 21821 32725 21833 32728
rect 21867 32725 21879 32759
rect 21821 32719 21879 32725
rect 22094 32716 22100 32768
rect 22152 32756 22158 32768
rect 22554 32756 22560 32768
rect 22152 32728 22560 32756
rect 22152 32716 22158 32728
rect 22554 32716 22560 32728
rect 22612 32716 22618 32768
rect 23198 32716 23204 32768
rect 23256 32756 23262 32768
rect 26142 32756 26148 32768
rect 23256 32728 26148 32756
rect 23256 32716 23262 32728
rect 26142 32716 26148 32728
rect 26200 32756 26206 32768
rect 28445 32759 28503 32765
rect 28445 32756 28457 32759
rect 26200 32728 28457 32756
rect 26200 32716 26206 32728
rect 28445 32725 28457 32728
rect 28491 32725 28503 32759
rect 28445 32719 28503 32725
rect 28902 32716 28908 32768
rect 28960 32756 28966 32768
rect 30300 32756 30328 32864
rect 31941 32861 31953 32864
rect 31987 32861 31999 32895
rect 31941 32855 31999 32861
rect 32033 32895 32091 32901
rect 32033 32861 32045 32895
rect 32079 32892 32091 32895
rect 32122 32892 32128 32904
rect 32079 32864 32128 32892
rect 32079 32861 32091 32864
rect 32033 32855 32091 32861
rect 32122 32852 32128 32864
rect 32180 32852 32186 32904
rect 32306 32852 32312 32904
rect 32364 32852 32370 32904
rect 32416 32824 32444 32932
rect 32784 32932 33089 32960
rect 32493 32895 32551 32901
rect 32493 32861 32505 32895
rect 32539 32892 32551 32895
rect 32582 32892 32588 32904
rect 32539 32864 32588 32892
rect 32539 32861 32551 32864
rect 32493 32855 32551 32861
rect 32582 32852 32588 32864
rect 32640 32852 32646 32904
rect 32674 32852 32680 32904
rect 32732 32892 32738 32904
rect 32784 32892 32812 32932
rect 32732 32864 32812 32892
rect 32732 32852 32738 32864
rect 32858 32852 32864 32904
rect 32916 32892 32922 32904
rect 33061 32901 33089 32932
rect 33428 32904 33456 33000
rect 33520 32960 33548 33068
rect 33597 33065 33609 33099
rect 33643 33096 33655 33099
rect 34514 33096 34520 33108
rect 33643 33068 34520 33096
rect 33643 33065 33655 33068
rect 33597 33059 33655 33065
rect 34514 33056 34520 33068
rect 34572 33056 34578 33108
rect 38010 33096 38016 33108
rect 35544 33068 38016 33096
rect 34146 32988 34152 33040
rect 34204 33028 34210 33040
rect 34241 33031 34299 33037
rect 34241 33028 34253 33031
rect 34204 33000 34253 33028
rect 34204 32988 34210 33000
rect 34241 32997 34253 33000
rect 34287 32997 34299 33031
rect 34241 32991 34299 32997
rect 33520 32932 34192 32960
rect 32953 32895 33011 32901
rect 32953 32892 32965 32895
rect 32916 32864 32965 32892
rect 32916 32852 32922 32864
rect 32953 32861 32965 32864
rect 32999 32861 33011 32895
rect 32953 32855 33011 32861
rect 33046 32895 33104 32901
rect 33046 32861 33058 32895
rect 33092 32861 33104 32895
rect 33046 32855 33104 32861
rect 33134 32852 33140 32904
rect 33192 32892 33198 32904
rect 33229 32895 33287 32901
rect 33229 32892 33241 32895
rect 33192 32864 33241 32892
rect 33192 32852 33198 32864
rect 33229 32861 33241 32864
rect 33275 32861 33287 32895
rect 33229 32855 33287 32861
rect 33318 32852 33324 32904
rect 33376 32852 33382 32904
rect 33410 32852 33416 32904
rect 33468 32901 33474 32904
rect 34164 32901 34192 32932
rect 34330 32920 34336 32972
rect 34388 32920 34394 32972
rect 33468 32892 33476 32901
rect 34057 32895 34115 32901
rect 33468 32864 33513 32892
rect 33468 32855 33476 32864
rect 34057 32861 34069 32895
rect 34103 32861 34115 32895
rect 34057 32855 34115 32861
rect 34149 32895 34207 32901
rect 34149 32861 34161 32895
rect 34195 32861 34207 32895
rect 34149 32855 34207 32861
rect 33468 32852 33474 32855
rect 34072 32824 34100 32855
rect 34514 32852 34520 32904
rect 34572 32892 34578 32904
rect 34885 32895 34943 32901
rect 34885 32892 34897 32895
rect 34572 32864 34897 32892
rect 34572 32852 34578 32864
rect 34885 32861 34897 32864
rect 34931 32861 34943 32895
rect 34885 32855 34943 32861
rect 35066 32852 35072 32904
rect 35124 32852 35130 32904
rect 35544 32901 35572 33068
rect 38010 33056 38016 33068
rect 38068 33056 38074 33108
rect 35710 32960 35716 32972
rect 35637 32932 35716 32960
rect 35637 32901 35665 32932
rect 35710 32920 35716 32932
rect 35768 32920 35774 32972
rect 36722 32960 36728 32972
rect 35912 32932 36728 32960
rect 35529 32895 35587 32901
rect 35529 32861 35541 32895
rect 35575 32861 35587 32895
rect 35529 32855 35587 32861
rect 35622 32895 35680 32901
rect 35622 32861 35634 32895
rect 35668 32861 35680 32895
rect 35912 32892 35940 32932
rect 36722 32920 36728 32932
rect 36780 32920 36786 32972
rect 35622 32855 35680 32861
rect 35728 32864 35940 32892
rect 36035 32895 36093 32901
rect 35728 32824 35756 32864
rect 36035 32861 36047 32895
rect 36081 32892 36093 32895
rect 36630 32892 36636 32904
rect 36081 32864 36636 32892
rect 36081 32861 36093 32864
rect 36035 32855 36093 32861
rect 36630 32852 36636 32864
rect 36688 32852 36694 32904
rect 36817 32895 36875 32901
rect 36817 32861 36829 32895
rect 36863 32861 36875 32895
rect 36817 32855 36875 32861
rect 32416 32796 34100 32824
rect 34624 32796 35756 32824
rect 28960 32728 30328 32756
rect 28960 32716 28966 32728
rect 31754 32716 31760 32768
rect 31812 32756 31818 32768
rect 34624 32756 34652 32796
rect 35802 32784 35808 32836
rect 35860 32784 35866 32836
rect 35897 32827 35955 32833
rect 35897 32793 35909 32827
rect 35943 32793 35955 32827
rect 35897 32787 35955 32793
rect 31812 32728 34652 32756
rect 31812 32716 31818 32728
rect 34698 32716 34704 32768
rect 34756 32756 34762 32768
rect 34977 32759 35035 32765
rect 34977 32756 34989 32759
rect 34756 32728 34989 32756
rect 34756 32716 34762 32728
rect 34977 32725 34989 32728
rect 35023 32725 35035 32759
rect 34977 32719 35035 32725
rect 35342 32716 35348 32768
rect 35400 32756 35406 32768
rect 35710 32756 35716 32768
rect 35400 32728 35716 32756
rect 35400 32716 35406 32728
rect 35710 32716 35716 32728
rect 35768 32756 35774 32768
rect 35912 32756 35940 32787
rect 36538 32784 36544 32836
rect 36596 32824 36602 32836
rect 36832 32824 36860 32855
rect 36596 32796 36860 32824
rect 37084 32827 37142 32833
rect 36596 32784 36602 32796
rect 37084 32793 37096 32827
rect 37130 32824 37142 32827
rect 37458 32824 37464 32836
rect 37130 32796 37464 32824
rect 37130 32793 37142 32796
rect 37084 32787 37142 32793
rect 37458 32784 37464 32796
rect 37516 32784 37522 32836
rect 35768 32728 35940 32756
rect 35768 32716 35774 32728
rect 36170 32716 36176 32768
rect 36228 32716 36234 32768
rect 37826 32716 37832 32768
rect 37884 32756 37890 32768
rect 38197 32759 38255 32765
rect 38197 32756 38209 32759
rect 37884 32728 38209 32756
rect 37884 32716 37890 32728
rect 38197 32725 38209 32728
rect 38243 32725 38255 32759
rect 38197 32719 38255 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 4157 32555 4215 32561
rect 4157 32521 4169 32555
rect 4203 32552 4215 32555
rect 8478 32552 8484 32564
rect 4203 32524 8484 32552
rect 4203 32521 4215 32524
rect 4157 32515 4215 32521
rect 8478 32512 8484 32524
rect 8536 32552 8542 32564
rect 13814 32552 13820 32564
rect 8536 32524 10088 32552
rect 8536 32512 8542 32524
rect 7098 32484 7104 32496
rect 4080 32456 7104 32484
rect 4080 32425 4108 32456
rect 7098 32444 7104 32456
rect 7156 32444 7162 32496
rect 7828 32487 7886 32493
rect 7828 32453 7840 32487
rect 7874 32484 7886 32487
rect 9122 32484 9128 32496
rect 7874 32456 9128 32484
rect 7874 32453 7886 32456
rect 7828 32447 7886 32453
rect 9122 32444 9128 32456
rect 9180 32444 9186 32496
rect 10060 32493 10088 32524
rect 11072 32524 13820 32552
rect 10045 32487 10103 32493
rect 10045 32453 10057 32487
rect 10091 32453 10103 32487
rect 10045 32447 10103 32453
rect 10965 32429 11023 32435
rect 4065 32419 4123 32425
rect 4065 32385 4077 32419
rect 4111 32385 4123 32419
rect 4065 32379 4123 32385
rect 4522 32376 4528 32428
rect 4580 32416 4586 32428
rect 4709 32419 4767 32425
rect 4709 32416 4721 32419
rect 4580 32388 4721 32416
rect 4580 32376 4586 32388
rect 4709 32385 4721 32388
rect 4755 32385 4767 32419
rect 4709 32379 4767 32385
rect 4893 32419 4951 32425
rect 4893 32385 4905 32419
rect 4939 32385 4951 32419
rect 4893 32379 4951 32385
rect 2682 32308 2688 32360
rect 2740 32348 2746 32360
rect 4908 32348 4936 32379
rect 5810 32376 5816 32428
rect 5868 32376 5874 32428
rect 5905 32419 5963 32425
rect 5905 32385 5917 32419
rect 5951 32385 5963 32419
rect 5905 32379 5963 32385
rect 2740 32320 4936 32348
rect 5920 32348 5948 32379
rect 5994 32376 6000 32428
rect 6052 32376 6058 32428
rect 6730 32376 6736 32428
rect 6788 32376 6794 32428
rect 6914 32376 6920 32428
rect 6972 32376 6978 32428
rect 8294 32376 8300 32428
rect 8352 32416 8358 32428
rect 9030 32416 9036 32428
rect 8352 32388 9036 32416
rect 8352 32376 8358 32388
rect 9030 32376 9036 32388
rect 9088 32376 9094 32428
rect 9769 32419 9827 32425
rect 9769 32385 9781 32419
rect 9815 32385 9827 32419
rect 9769 32379 9827 32385
rect 6362 32348 6368 32360
rect 5920 32320 6368 32348
rect 2740 32308 2746 32320
rect 6362 32308 6368 32320
rect 6420 32308 6426 32360
rect 6748 32348 6776 32376
rect 7006 32348 7012 32360
rect 6748 32320 7012 32348
rect 7006 32308 7012 32320
rect 7064 32308 7070 32360
rect 7374 32308 7380 32360
rect 7432 32348 7438 32360
rect 7561 32351 7619 32357
rect 7561 32348 7573 32351
rect 7432 32320 7573 32348
rect 7432 32308 7438 32320
rect 7561 32317 7573 32320
rect 7607 32317 7619 32351
rect 7561 32311 7619 32317
rect 8754 32308 8760 32360
rect 8812 32348 8818 32360
rect 9398 32348 9404 32360
rect 8812 32320 9404 32348
rect 8812 32308 8818 32320
rect 9398 32308 9404 32320
rect 9456 32308 9462 32360
rect 9784 32348 9812 32379
rect 9950 32376 9956 32428
rect 10008 32376 10014 32428
rect 10134 32376 10140 32428
rect 10192 32376 10198 32428
rect 10965 32395 10977 32429
rect 11011 32426 11023 32429
rect 11072 32426 11100 32524
rect 13814 32512 13820 32524
rect 13872 32512 13878 32564
rect 13998 32512 14004 32564
rect 14056 32552 14062 32564
rect 15838 32552 15844 32564
rect 14056 32524 15844 32552
rect 14056 32512 14062 32524
rect 15838 32512 15844 32524
rect 15896 32512 15902 32564
rect 16114 32512 16120 32564
rect 16172 32552 16178 32564
rect 19150 32552 19156 32564
rect 16172 32524 19156 32552
rect 16172 32512 16178 32524
rect 19150 32512 19156 32524
rect 19208 32512 19214 32564
rect 19426 32512 19432 32564
rect 19484 32552 19490 32564
rect 19613 32555 19671 32561
rect 19613 32552 19625 32555
rect 19484 32524 19625 32552
rect 19484 32512 19490 32524
rect 19613 32521 19625 32524
rect 19659 32521 19671 32555
rect 19613 32515 19671 32521
rect 20257 32555 20315 32561
rect 20257 32521 20269 32555
rect 20303 32552 20315 32555
rect 22094 32552 22100 32564
rect 20303 32524 22100 32552
rect 20303 32521 20315 32524
rect 20257 32515 20315 32521
rect 22094 32512 22100 32524
rect 22152 32512 22158 32564
rect 22186 32512 22192 32564
rect 22244 32552 22250 32564
rect 22281 32555 22339 32561
rect 22281 32552 22293 32555
rect 22244 32524 22293 32552
rect 22244 32512 22250 32524
rect 22281 32521 22293 32524
rect 22327 32521 22339 32555
rect 23750 32552 23756 32564
rect 22281 32515 22339 32521
rect 22388 32524 23756 32552
rect 11790 32444 11796 32496
rect 11848 32444 11854 32496
rect 11977 32487 12035 32493
rect 11977 32453 11989 32487
rect 12023 32484 12035 32487
rect 12023 32456 12756 32484
rect 12023 32453 12035 32456
rect 11977 32447 12035 32453
rect 11011 32398 11100 32426
rect 11149 32419 11207 32425
rect 11011 32395 11023 32398
rect 10965 32389 11023 32395
rect 11149 32385 11161 32419
rect 11195 32416 11207 32419
rect 11238 32416 11244 32428
rect 11195 32388 11244 32416
rect 11195 32385 11207 32388
rect 11149 32379 11207 32385
rect 11238 32376 11244 32388
rect 11296 32376 11302 32428
rect 11330 32376 11336 32428
rect 11388 32416 11394 32428
rect 12253 32419 12311 32425
rect 12253 32416 12265 32419
rect 11388 32388 12265 32416
rect 11388 32376 11394 32388
rect 12253 32385 12265 32388
rect 12299 32385 12311 32419
rect 12253 32379 12311 32385
rect 10502 32348 10508 32360
rect 9784 32320 10508 32348
rect 10502 32308 10508 32320
rect 10560 32348 10566 32360
rect 11348 32348 11376 32376
rect 10560 32320 11376 32348
rect 10560 32308 10566 32320
rect 11790 32308 11796 32360
rect 11848 32348 11854 32360
rect 12526 32348 12532 32360
rect 11848 32320 12532 32348
rect 11848 32308 11854 32320
rect 12526 32308 12532 32320
rect 12584 32308 12590 32360
rect 12728 32348 12756 32456
rect 12986 32444 12992 32496
rect 13044 32484 13050 32496
rect 14826 32484 14832 32496
rect 13044 32456 14832 32484
rect 13044 32444 13050 32456
rect 14826 32444 14832 32456
rect 14884 32484 14890 32496
rect 15194 32484 15200 32496
rect 14884 32456 15200 32484
rect 14884 32444 14890 32456
rect 15194 32444 15200 32456
rect 15252 32444 15258 32496
rect 17954 32444 17960 32496
rect 18012 32444 18018 32496
rect 18049 32487 18107 32493
rect 18049 32453 18061 32487
rect 18095 32484 18107 32487
rect 18322 32484 18328 32496
rect 18095 32456 18328 32484
rect 18095 32453 18107 32456
rect 18049 32447 18107 32453
rect 18322 32444 18328 32456
rect 18380 32444 18386 32496
rect 20714 32484 20720 32496
rect 19444 32456 20720 32484
rect 12802 32376 12808 32428
rect 12860 32416 12866 32428
rect 12897 32419 12955 32425
rect 12897 32416 12909 32419
rect 12860 32388 12909 32416
rect 12860 32376 12866 32388
rect 12897 32385 12909 32388
rect 12943 32385 12955 32419
rect 12897 32379 12955 32385
rect 13909 32419 13967 32425
rect 13909 32385 13921 32419
rect 13955 32416 13967 32419
rect 14090 32416 14096 32428
rect 13955 32388 14096 32416
rect 13955 32385 13967 32388
rect 13909 32379 13967 32385
rect 14090 32376 14096 32388
rect 14148 32376 14154 32428
rect 15470 32376 15476 32428
rect 15528 32376 15534 32428
rect 16942 32376 16948 32428
rect 17000 32376 17006 32428
rect 17126 32376 17132 32428
rect 17184 32416 17190 32428
rect 17494 32416 17500 32428
rect 17184 32388 17500 32416
rect 17184 32376 17190 32388
rect 17494 32376 17500 32388
rect 17552 32376 17558 32428
rect 17770 32376 17776 32428
rect 17828 32376 17834 32428
rect 18141 32419 18199 32425
rect 18141 32385 18153 32419
rect 18187 32416 18199 32419
rect 18230 32416 18236 32428
rect 18187 32388 18236 32416
rect 18187 32385 18199 32388
rect 18141 32379 18199 32385
rect 18230 32376 18236 32388
rect 18288 32376 18294 32428
rect 19444 32425 19472 32456
rect 20714 32444 20720 32456
rect 20772 32444 20778 32496
rect 20806 32444 20812 32496
rect 20864 32444 20870 32496
rect 22388 32484 22416 32524
rect 23750 32512 23756 32524
rect 23808 32512 23814 32564
rect 24762 32512 24768 32564
rect 24820 32552 24826 32564
rect 25406 32552 25412 32564
rect 24820 32524 25412 32552
rect 24820 32512 24826 32524
rect 25406 32512 25412 32524
rect 25464 32512 25470 32564
rect 25498 32512 25504 32564
rect 25556 32512 25562 32564
rect 36170 32552 36176 32564
rect 27632 32524 36176 32552
rect 23474 32484 23480 32496
rect 21008 32456 22416 32484
rect 22756 32456 23480 32484
rect 19429 32419 19487 32425
rect 19429 32385 19441 32419
rect 19475 32385 19487 32419
rect 19429 32379 19487 32385
rect 19705 32419 19763 32425
rect 19705 32385 19717 32419
rect 19751 32416 19763 32419
rect 19978 32416 19984 32428
rect 19751 32388 19984 32416
rect 19751 32385 19763 32388
rect 19705 32379 19763 32385
rect 19978 32376 19984 32388
rect 20036 32376 20042 32428
rect 20165 32419 20223 32425
rect 20165 32385 20177 32419
rect 20211 32385 20223 32419
rect 20165 32379 20223 32385
rect 12986 32348 12992 32360
rect 12728 32320 12992 32348
rect 12986 32308 12992 32320
rect 13044 32308 13050 32360
rect 13078 32308 13084 32360
rect 13136 32308 13142 32360
rect 14185 32351 14243 32357
rect 14185 32348 14197 32351
rect 13188 32320 14197 32348
rect 5166 32240 5172 32292
rect 5224 32280 5230 32292
rect 5626 32280 5632 32292
rect 5224 32252 5632 32280
rect 5224 32240 5230 32252
rect 5626 32240 5632 32252
rect 5684 32240 5690 32292
rect 7098 32240 7104 32292
rect 7156 32240 7162 32292
rect 9674 32280 9680 32292
rect 8496 32252 9680 32280
rect 4062 32172 4068 32224
rect 4120 32212 4126 32224
rect 4614 32212 4620 32224
rect 4120 32184 4620 32212
rect 4120 32172 4126 32184
rect 4614 32172 4620 32184
rect 4672 32172 4678 32224
rect 4706 32172 4712 32224
rect 4764 32172 4770 32224
rect 5810 32172 5816 32224
rect 5868 32212 5874 32224
rect 8496 32212 8524 32252
rect 9674 32240 9680 32252
rect 9732 32240 9738 32292
rect 10689 32283 10747 32289
rect 10689 32249 10701 32283
rect 10735 32280 10747 32283
rect 11238 32280 11244 32292
rect 10735 32252 11244 32280
rect 10735 32249 10747 32252
rect 10689 32243 10747 32249
rect 11238 32240 11244 32252
rect 11296 32240 11302 32292
rect 12544 32280 12572 32308
rect 13188 32280 13216 32320
rect 14185 32317 14197 32320
rect 14231 32317 14243 32351
rect 14185 32311 14243 32317
rect 15010 32308 15016 32360
rect 15068 32348 15074 32360
rect 15289 32351 15347 32357
rect 15289 32348 15301 32351
rect 15068 32320 15301 32348
rect 15068 32308 15074 32320
rect 15289 32317 15301 32320
rect 15335 32317 15347 32351
rect 19334 32348 19340 32360
rect 15289 32311 15347 32317
rect 16960 32320 19340 32348
rect 12544 32252 13216 32280
rect 13262 32240 13268 32292
rect 13320 32280 13326 32292
rect 15378 32280 15384 32292
rect 13320 32252 15384 32280
rect 13320 32240 13326 32252
rect 15378 32240 15384 32252
rect 15436 32240 15442 32292
rect 16960 32280 16988 32320
rect 19334 32308 19340 32320
rect 19392 32308 19398 32360
rect 20180 32348 20208 32379
rect 20346 32376 20352 32428
rect 20404 32376 20410 32428
rect 21008 32425 21036 32456
rect 20993 32419 21051 32425
rect 20993 32385 21005 32419
rect 21039 32385 21051 32419
rect 20993 32379 21051 32385
rect 21085 32419 21143 32425
rect 21085 32385 21097 32419
rect 21131 32416 21143 32419
rect 21634 32416 21640 32428
rect 21131 32388 21640 32416
rect 21131 32385 21143 32388
rect 21085 32379 21143 32385
rect 21634 32376 21640 32388
rect 21692 32376 21698 32428
rect 22186 32376 22192 32428
rect 22244 32416 22250 32428
rect 22462 32416 22468 32428
rect 22244 32388 22468 32416
rect 22244 32376 22250 32388
rect 22462 32376 22468 32388
rect 22520 32376 22526 32428
rect 22649 32422 22707 32425
rect 22756 32422 22784 32456
rect 23474 32444 23480 32456
rect 23532 32444 23538 32496
rect 27338 32484 27344 32496
rect 23768 32456 27344 32484
rect 22649 32419 22784 32422
rect 22649 32385 22661 32419
rect 22695 32394 22784 32419
rect 22695 32385 22707 32394
rect 22649 32379 22707 32385
rect 22830 32376 22836 32428
rect 22888 32416 22894 32428
rect 22925 32419 22983 32425
rect 22925 32416 22937 32419
rect 22888 32388 22937 32416
rect 22888 32376 22894 32388
rect 22925 32385 22937 32388
rect 22971 32385 22983 32419
rect 22925 32379 22983 32385
rect 20180 32320 22692 32348
rect 15580 32252 16988 32280
rect 5868 32184 8524 32212
rect 5868 32172 5874 32184
rect 8570 32172 8576 32224
rect 8628 32212 8634 32224
rect 8754 32212 8760 32224
rect 8628 32184 8760 32212
rect 8628 32172 8634 32184
rect 8754 32172 8760 32184
rect 8812 32172 8818 32224
rect 8938 32172 8944 32224
rect 8996 32172 9002 32224
rect 9030 32172 9036 32224
rect 9088 32212 9094 32224
rect 9766 32212 9772 32224
rect 9088 32184 9772 32212
rect 9088 32172 9094 32184
rect 9766 32172 9772 32184
rect 9824 32172 9830 32224
rect 9858 32172 9864 32224
rect 9916 32212 9922 32224
rect 10321 32215 10379 32221
rect 10321 32212 10333 32215
rect 9916 32184 10333 32212
rect 9916 32172 9922 32184
rect 10321 32181 10333 32184
rect 10367 32181 10379 32215
rect 10321 32175 10379 32181
rect 11054 32172 11060 32224
rect 11112 32172 11118 32224
rect 11606 32172 11612 32224
rect 11664 32212 11670 32224
rect 11943 32215 12001 32221
rect 11943 32212 11955 32215
rect 11664 32184 11955 32212
rect 11664 32172 11670 32184
rect 11943 32181 11955 32184
rect 11989 32181 12001 32215
rect 11943 32175 12001 32181
rect 15102 32172 15108 32224
rect 15160 32212 15166 32224
rect 15197 32215 15255 32221
rect 15197 32212 15209 32215
rect 15160 32184 15209 32212
rect 15160 32172 15166 32184
rect 15197 32181 15209 32184
rect 15243 32212 15255 32215
rect 15580 32212 15608 32252
rect 15243 32184 15608 32212
rect 15243 32181 15255 32184
rect 15197 32175 15255 32181
rect 15654 32172 15660 32224
rect 15712 32172 15718 32224
rect 16960 32221 16988 32252
rect 18046 32240 18052 32292
rect 18104 32280 18110 32292
rect 18874 32280 18880 32292
rect 18104 32252 18880 32280
rect 18104 32240 18110 32252
rect 18874 32240 18880 32252
rect 18932 32240 18938 32292
rect 21269 32283 21327 32289
rect 19168 32252 21220 32280
rect 16945 32215 17003 32221
rect 16945 32181 16957 32215
rect 16991 32181 17003 32215
rect 16945 32175 17003 32181
rect 17313 32215 17371 32221
rect 17313 32181 17325 32215
rect 17359 32212 17371 32215
rect 17862 32212 17868 32224
rect 17359 32184 17868 32212
rect 17359 32181 17371 32184
rect 17313 32175 17371 32181
rect 17862 32172 17868 32184
rect 17920 32172 17926 32224
rect 18230 32172 18236 32224
rect 18288 32212 18294 32224
rect 18325 32215 18383 32221
rect 18325 32212 18337 32215
rect 18288 32184 18337 32212
rect 18288 32172 18294 32184
rect 18325 32181 18337 32184
rect 18371 32181 18383 32215
rect 18325 32175 18383 32181
rect 18782 32172 18788 32224
rect 18840 32212 18846 32224
rect 19168 32212 19196 32252
rect 18840 32184 19196 32212
rect 18840 32172 18846 32184
rect 19242 32172 19248 32224
rect 19300 32172 19306 32224
rect 19334 32172 19340 32224
rect 19392 32212 19398 32224
rect 20530 32212 20536 32224
rect 19392 32184 20536 32212
rect 19392 32172 19398 32184
rect 20530 32172 20536 32184
rect 20588 32172 20594 32224
rect 20990 32172 20996 32224
rect 21048 32172 21054 32224
rect 21192 32212 21220 32252
rect 21269 32249 21281 32283
rect 21315 32280 21327 32283
rect 21726 32280 21732 32292
rect 21315 32252 21732 32280
rect 21315 32249 21327 32252
rect 21269 32243 21327 32249
rect 21726 32240 21732 32252
rect 21784 32240 21790 32292
rect 22462 32240 22468 32292
rect 22520 32280 22526 32292
rect 22557 32283 22615 32289
rect 22557 32280 22569 32283
rect 22520 32252 22569 32280
rect 22520 32240 22526 32252
rect 22557 32249 22569 32252
rect 22603 32249 22615 32283
rect 22664 32280 22692 32320
rect 22738 32308 22744 32360
rect 22796 32348 22802 32360
rect 23768 32348 23796 32456
rect 27338 32444 27344 32456
rect 27396 32444 27402 32496
rect 23845 32419 23903 32425
rect 23845 32385 23857 32419
rect 23891 32416 23903 32419
rect 24026 32416 24032 32428
rect 23891 32388 24032 32416
rect 23891 32385 23903 32388
rect 23845 32379 23903 32385
rect 24026 32376 24032 32388
rect 24084 32376 24090 32428
rect 24949 32419 25007 32425
rect 24949 32385 24961 32419
rect 24995 32416 25007 32419
rect 25130 32416 25136 32428
rect 24995 32388 25136 32416
rect 24995 32385 25007 32388
rect 24949 32379 25007 32385
rect 25130 32376 25136 32388
rect 25188 32376 25194 32428
rect 25314 32376 25320 32428
rect 25372 32376 25378 32428
rect 26145 32419 26203 32425
rect 26145 32385 26157 32419
rect 26191 32416 26203 32419
rect 27522 32416 27528 32428
rect 26191 32388 27528 32416
rect 26191 32385 26203 32388
rect 26145 32379 26203 32385
rect 27522 32376 27528 32388
rect 27580 32376 27586 32428
rect 27632 32425 27660 32524
rect 36170 32512 36176 32524
rect 36228 32512 36234 32564
rect 37458 32512 37464 32564
rect 37516 32512 37522 32564
rect 37826 32512 37832 32564
rect 37884 32512 37890 32564
rect 27893 32487 27951 32493
rect 27893 32453 27905 32487
rect 27939 32484 27951 32487
rect 27939 32456 29224 32484
rect 27939 32453 27951 32456
rect 27893 32447 27951 32453
rect 27617 32419 27675 32425
rect 27617 32385 27629 32419
rect 27663 32385 27675 32419
rect 27617 32379 27675 32385
rect 27798 32376 27804 32428
rect 27856 32416 27862 32428
rect 27856 32388 28212 32416
rect 27856 32376 27862 32388
rect 22796 32320 23796 32348
rect 22796 32308 22802 32320
rect 24118 32308 24124 32360
rect 24176 32308 24182 32360
rect 24762 32308 24768 32360
rect 24820 32348 24826 32360
rect 24857 32351 24915 32357
rect 24857 32348 24869 32351
rect 24820 32320 24869 32348
rect 24820 32308 24826 32320
rect 24857 32317 24869 32320
rect 24903 32317 24915 32351
rect 24857 32311 24915 32317
rect 25406 32308 25412 32360
rect 25464 32348 25470 32360
rect 25774 32348 25780 32360
rect 25464 32320 25780 32348
rect 25464 32308 25470 32320
rect 25774 32308 25780 32320
rect 25832 32308 25838 32360
rect 26421 32351 26479 32357
rect 26421 32317 26433 32351
rect 26467 32348 26479 32351
rect 28184 32348 28212 32388
rect 28258 32376 28264 32428
rect 28316 32416 28322 32428
rect 28718 32425 28724 32428
rect 28537 32419 28595 32425
rect 28537 32416 28549 32419
rect 28316 32388 28549 32416
rect 28316 32376 28322 32388
rect 28537 32385 28549 32388
rect 28583 32385 28595 32419
rect 28537 32379 28595 32385
rect 28684 32419 28724 32425
rect 28684 32385 28696 32419
rect 28684 32379 28724 32385
rect 28718 32376 28724 32379
rect 28776 32376 28782 32428
rect 28902 32348 28908 32360
rect 26467 32320 27936 32348
rect 28184 32320 28908 32348
rect 26467 32317 26479 32320
rect 26421 32311 26479 32317
rect 22830 32280 22836 32292
rect 22664 32252 22836 32280
rect 22557 32243 22615 32249
rect 22830 32240 22836 32252
rect 22888 32280 22894 32292
rect 23842 32280 23848 32292
rect 22888 32252 23848 32280
rect 22888 32240 22894 32252
rect 23842 32240 23848 32252
rect 23900 32280 23906 32292
rect 24578 32280 24584 32292
rect 23900 32252 24584 32280
rect 23900 32240 23906 32252
rect 24578 32240 24584 32252
rect 24636 32240 24642 32292
rect 24670 32240 24676 32292
rect 24728 32280 24734 32292
rect 25038 32280 25044 32292
rect 24728 32252 25044 32280
rect 24728 32240 24734 32252
rect 25038 32240 25044 32252
rect 25096 32240 25102 32292
rect 25317 32215 25375 32221
rect 25317 32212 25329 32215
rect 21192 32184 25329 32212
rect 25317 32181 25329 32184
rect 25363 32181 25375 32215
rect 25317 32175 25375 32181
rect 25406 32172 25412 32224
rect 25464 32212 25470 32224
rect 26510 32212 26516 32224
rect 25464 32184 26516 32212
rect 25464 32172 25470 32184
rect 26510 32172 26516 32184
rect 26568 32172 26574 32224
rect 27908 32212 27936 32320
rect 28902 32308 28908 32320
rect 28960 32308 28966 32360
rect 28994 32308 29000 32360
rect 29052 32308 29058 32360
rect 28166 32240 28172 32292
rect 28224 32280 28230 32292
rect 28813 32283 28871 32289
rect 28813 32280 28825 32283
rect 28224 32252 28825 32280
rect 28224 32240 28230 32252
rect 28813 32249 28825 32252
rect 28859 32249 28871 32283
rect 29196 32280 29224 32456
rect 29822 32444 29828 32496
rect 29880 32484 29886 32496
rect 30282 32484 30288 32496
rect 29880 32456 30288 32484
rect 29880 32444 29886 32456
rect 30282 32444 30288 32456
rect 30340 32444 30346 32496
rect 31202 32444 31208 32496
rect 31260 32484 31266 32496
rect 31260 32456 32536 32484
rect 31260 32444 31266 32456
rect 29454 32376 29460 32428
rect 29512 32416 29518 32428
rect 29733 32419 29791 32425
rect 29733 32416 29745 32419
rect 29512 32388 29745 32416
rect 29512 32376 29518 32388
rect 29733 32385 29745 32388
rect 29779 32385 29791 32419
rect 29733 32379 29791 32385
rect 29917 32419 29975 32425
rect 29917 32385 29929 32419
rect 29963 32416 29975 32419
rect 30098 32416 30104 32428
rect 29963 32388 30104 32416
rect 29963 32385 29975 32388
rect 29917 32379 29975 32385
rect 30098 32376 30104 32388
rect 30156 32376 30162 32428
rect 30650 32376 30656 32428
rect 30708 32376 30714 32428
rect 31018 32376 31024 32428
rect 31076 32376 31082 32428
rect 31570 32376 31576 32428
rect 31628 32376 31634 32428
rect 31757 32419 31815 32425
rect 31757 32385 31769 32419
rect 31803 32416 31815 32419
rect 31938 32416 31944 32428
rect 31803 32388 31944 32416
rect 31803 32385 31815 32388
rect 31757 32379 31815 32385
rect 31938 32376 31944 32388
rect 31996 32376 32002 32428
rect 32306 32376 32312 32428
rect 32364 32376 32370 32428
rect 32508 32425 32536 32456
rect 33226 32444 33232 32496
rect 33284 32484 33290 32496
rect 34149 32487 34207 32493
rect 34149 32484 34161 32487
rect 33284 32456 34161 32484
rect 33284 32444 33290 32456
rect 34149 32453 34161 32456
rect 34195 32453 34207 32487
rect 34149 32447 34207 32453
rect 34422 32444 34428 32496
rect 34480 32484 34486 32496
rect 36188 32484 36216 32512
rect 37921 32487 37979 32493
rect 37921 32484 37933 32487
rect 34480 32456 35940 32484
rect 36188 32456 37933 32484
rect 34480 32444 34486 32456
rect 32493 32419 32551 32425
rect 32493 32385 32505 32419
rect 32539 32385 32551 32419
rect 32493 32379 32551 32385
rect 32582 32376 32588 32428
rect 32640 32416 32646 32428
rect 32640 32388 32997 32416
rect 32640 32376 32646 32388
rect 29270 32308 29276 32360
rect 29328 32348 29334 32360
rect 30926 32348 30932 32360
rect 29328 32320 30932 32348
rect 29328 32308 29334 32320
rect 30926 32308 30932 32320
rect 30984 32308 30990 32360
rect 32324 32348 32352 32376
rect 32769 32351 32827 32357
rect 32769 32348 32781 32351
rect 32324 32320 32781 32348
rect 32769 32317 32781 32320
rect 32815 32317 32827 32351
rect 32969 32348 32997 32388
rect 33042 32376 33048 32428
rect 33100 32376 33106 32428
rect 33318 32376 33324 32428
rect 33376 32416 33382 32428
rect 33873 32419 33931 32425
rect 33873 32416 33885 32419
rect 33376 32388 33885 32416
rect 33376 32376 33382 32388
rect 33873 32385 33885 32388
rect 33919 32385 33931 32419
rect 33873 32379 33931 32385
rect 34057 32419 34115 32425
rect 34057 32385 34069 32419
rect 34103 32385 34115 32419
rect 34057 32379 34115 32385
rect 34241 32419 34299 32425
rect 34241 32385 34253 32419
rect 34287 32416 34299 32419
rect 34606 32416 34612 32428
rect 34287 32388 34612 32416
rect 34287 32385 34299 32388
rect 34241 32379 34299 32385
rect 34072 32348 34100 32379
rect 34606 32376 34612 32388
rect 34664 32376 34670 32428
rect 34882 32376 34888 32428
rect 34940 32416 34946 32428
rect 35912 32425 35940 32456
rect 37921 32453 37933 32456
rect 37967 32453 37979 32487
rect 37921 32447 37979 32453
rect 35069 32419 35127 32425
rect 35069 32416 35081 32419
rect 34940 32388 35081 32416
rect 34940 32376 34946 32388
rect 35069 32385 35081 32388
rect 35115 32385 35127 32419
rect 35069 32379 35127 32385
rect 35897 32419 35955 32425
rect 35897 32385 35909 32419
rect 35943 32385 35955 32419
rect 35897 32379 35955 32385
rect 36081 32419 36139 32425
rect 36081 32385 36093 32419
rect 36127 32385 36139 32419
rect 36081 32379 36139 32385
rect 32969 32320 34100 32348
rect 32769 32311 32827 32317
rect 33888 32292 33916 32320
rect 34790 32308 34796 32360
rect 34848 32348 34854 32360
rect 34977 32351 35035 32357
rect 34977 32348 34989 32351
rect 34848 32320 34989 32348
rect 34848 32308 34854 32320
rect 34977 32317 34989 32320
rect 35023 32317 35035 32351
rect 34977 32311 35035 32317
rect 35618 32308 35624 32360
rect 35676 32348 35682 32360
rect 35802 32348 35808 32360
rect 35676 32320 35808 32348
rect 35676 32308 35682 32320
rect 35802 32308 35808 32320
rect 35860 32348 35866 32360
rect 36096 32348 36124 32379
rect 36170 32376 36176 32428
rect 36228 32376 36234 32428
rect 36265 32419 36323 32425
rect 36265 32385 36277 32419
rect 36311 32385 36323 32419
rect 36265 32379 36323 32385
rect 35860 32320 36124 32348
rect 35860 32308 35866 32320
rect 29196 32252 33269 32280
rect 28813 32243 28871 32249
rect 29270 32212 29276 32224
rect 27908 32184 29276 32212
rect 29270 32172 29276 32184
rect 29328 32172 29334 32224
rect 29822 32172 29828 32224
rect 29880 32212 29886 32224
rect 30101 32215 30159 32221
rect 30101 32212 30113 32215
rect 29880 32184 30113 32212
rect 29880 32172 29886 32184
rect 30101 32181 30113 32184
rect 30147 32181 30159 32215
rect 30101 32175 30159 32181
rect 32398 32172 32404 32224
rect 32456 32172 32462 32224
rect 32950 32172 32956 32224
rect 33008 32212 33014 32224
rect 33137 32215 33195 32221
rect 33137 32212 33149 32215
rect 33008 32184 33149 32212
rect 33008 32172 33014 32184
rect 33137 32181 33149 32184
rect 33183 32181 33195 32215
rect 33241 32212 33269 32252
rect 33870 32240 33876 32292
rect 33928 32240 33934 32292
rect 34425 32283 34483 32289
rect 34425 32249 34437 32283
rect 34471 32280 34483 32283
rect 36078 32280 36084 32292
rect 34471 32252 36084 32280
rect 34471 32249 34483 32252
rect 34425 32243 34483 32249
rect 36078 32240 36084 32252
rect 36136 32240 36142 32292
rect 36280 32280 36308 32379
rect 38010 32308 38016 32360
rect 38068 32308 38074 32360
rect 36722 32280 36728 32292
rect 36280 32252 36728 32280
rect 36722 32240 36728 32252
rect 36780 32280 36786 32292
rect 37918 32280 37924 32292
rect 36780 32252 37924 32280
rect 36780 32240 36786 32252
rect 37918 32240 37924 32252
rect 37976 32240 37982 32292
rect 34974 32212 34980 32224
rect 33241 32184 34980 32212
rect 33137 32175 33195 32181
rect 34974 32172 34980 32184
rect 35032 32172 35038 32224
rect 35342 32172 35348 32224
rect 35400 32212 35406 32224
rect 35437 32215 35495 32221
rect 35437 32212 35449 32215
rect 35400 32184 35449 32212
rect 35400 32172 35406 32184
rect 35437 32181 35449 32184
rect 35483 32181 35495 32215
rect 35437 32175 35495 32181
rect 35894 32172 35900 32224
rect 35952 32212 35958 32224
rect 36449 32215 36507 32221
rect 36449 32212 36461 32215
rect 35952 32184 36461 32212
rect 35952 32172 35958 32184
rect 36449 32181 36461 32184
rect 36495 32181 36507 32215
rect 36449 32175 36507 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 6362 32008 6368 32020
rect 4356 31980 6368 32008
rect 4356 31813 4384 31980
rect 6362 31968 6368 31980
rect 6420 32008 6426 32020
rect 7006 32008 7012 32020
rect 6420 31980 7012 32008
rect 6420 31968 6426 31980
rect 7006 31968 7012 31980
rect 7064 32008 7070 32020
rect 7653 32011 7711 32017
rect 7653 32008 7665 32011
rect 7064 31980 7665 32008
rect 7064 31968 7070 31980
rect 7653 31977 7665 31980
rect 7699 31977 7711 32011
rect 7653 31971 7711 31977
rect 8389 32011 8447 32017
rect 8389 31977 8401 32011
rect 8435 32008 8447 32011
rect 8478 32008 8484 32020
rect 8435 31980 8484 32008
rect 8435 31977 8447 31980
rect 8389 31971 8447 31977
rect 8478 31968 8484 31980
rect 8536 31968 8542 32020
rect 8588 31980 9168 32008
rect 5810 31940 5816 31952
rect 4540 31912 5816 31940
rect 4430 31832 4436 31884
rect 4488 31832 4494 31884
rect 4540 31813 4568 31912
rect 5810 31900 5816 31912
rect 5868 31900 5874 31952
rect 6825 31943 6883 31949
rect 6825 31909 6837 31943
rect 6871 31940 6883 31943
rect 8588 31940 8616 31980
rect 6871 31912 8616 31940
rect 9140 31940 9168 31980
rect 9398 31968 9404 32020
rect 9456 32008 9462 32020
rect 10134 32008 10140 32020
rect 9456 31980 10140 32008
rect 9456 31968 9462 31980
rect 10134 31968 10140 31980
rect 10192 31968 10198 32020
rect 11793 32011 11851 32017
rect 11793 31977 11805 32011
rect 11839 32008 11851 32011
rect 12250 32008 12256 32020
rect 11839 31980 12256 32008
rect 11839 31977 11851 31980
rect 11793 31971 11851 31977
rect 12250 31968 12256 31980
rect 12308 31968 12314 32020
rect 13078 32008 13084 32020
rect 12360 31980 13084 32008
rect 9582 31940 9588 31952
rect 9140 31912 9588 31940
rect 6871 31909 6883 31912
rect 6825 31903 6883 31909
rect 9582 31900 9588 31912
rect 9640 31900 9646 31952
rect 9766 31900 9772 31952
rect 9824 31940 9830 31952
rect 12360 31940 12388 31980
rect 13078 31968 13084 31980
rect 13136 31968 13142 32020
rect 13906 32008 13912 32020
rect 13188 31980 13912 32008
rect 12986 31940 12992 31952
rect 9824 31912 12388 31940
rect 12452 31912 12992 31940
rect 9824 31900 9830 31912
rect 5442 31832 5448 31884
rect 5500 31872 5506 31884
rect 5500 31844 6776 31872
rect 5500 31832 5506 31844
rect 4341 31807 4399 31813
rect 4341 31773 4353 31807
rect 4387 31773 4399 31807
rect 4341 31767 4399 31773
rect 4525 31807 4583 31813
rect 4525 31773 4537 31807
rect 4571 31773 4583 31807
rect 4525 31767 4583 31773
rect 4893 31807 4951 31813
rect 4893 31773 4905 31807
rect 4939 31804 4951 31807
rect 4982 31804 4988 31816
rect 4939 31776 4988 31804
rect 4939 31773 4951 31776
rect 4893 31767 4951 31773
rect 4982 31764 4988 31776
rect 5040 31804 5046 31816
rect 5169 31807 5227 31813
rect 5169 31804 5181 31807
rect 5040 31776 5181 31804
rect 5040 31764 5046 31776
rect 5169 31773 5181 31776
rect 5215 31773 5227 31807
rect 5169 31767 5227 31773
rect 5350 31764 5356 31816
rect 5408 31764 5414 31816
rect 5810 31764 5816 31816
rect 5868 31764 5874 31816
rect 5994 31764 6000 31816
rect 6052 31764 6058 31816
rect 6362 31764 6368 31816
rect 6420 31804 6426 31816
rect 6420 31776 6500 31804
rect 6420 31764 6426 31776
rect 5261 31739 5319 31745
rect 5261 31705 5273 31739
rect 5307 31736 5319 31739
rect 6178 31736 6184 31748
rect 5307 31708 6184 31736
rect 5307 31705 5319 31708
rect 5261 31699 5319 31705
rect 6178 31696 6184 31708
rect 6236 31696 6242 31748
rect 4614 31628 4620 31680
rect 4672 31668 4678 31680
rect 4890 31668 4896 31680
rect 4672 31640 4896 31668
rect 4672 31628 4678 31640
rect 4890 31628 4896 31640
rect 4948 31628 4954 31680
rect 5534 31628 5540 31680
rect 5592 31668 5598 31680
rect 5905 31671 5963 31677
rect 5905 31668 5917 31671
rect 5592 31640 5917 31668
rect 5592 31628 5598 31640
rect 5905 31637 5917 31640
rect 5951 31637 5963 31671
rect 6472 31668 6500 31776
rect 6546 31764 6552 31816
rect 6604 31764 6610 31816
rect 6638 31764 6644 31816
rect 6696 31764 6702 31816
rect 6748 31736 6776 31844
rect 7926 31832 7932 31884
rect 7984 31872 7990 31884
rect 8205 31875 8263 31881
rect 8205 31872 8217 31875
rect 7984 31844 8217 31872
rect 7984 31832 7990 31844
rect 8205 31841 8217 31844
rect 8251 31841 8263 31875
rect 8205 31835 8263 31841
rect 9398 31832 9404 31884
rect 9456 31832 9462 31884
rect 9490 31832 9496 31884
rect 9548 31832 9554 31884
rect 10134 31832 10140 31884
rect 10192 31872 10198 31884
rect 11330 31872 11336 31884
rect 10192 31844 10548 31872
rect 10192 31832 10198 31844
rect 10520 31816 10548 31844
rect 10704 31844 11336 31872
rect 7285 31807 7343 31813
rect 7285 31773 7297 31807
rect 7331 31804 7343 31807
rect 8018 31804 8024 31816
rect 7331 31776 8024 31804
rect 7331 31773 7343 31776
rect 7285 31767 7343 31773
rect 8018 31764 8024 31776
rect 8076 31764 8082 31816
rect 8294 31764 8300 31816
rect 8352 31804 8358 31816
rect 8389 31807 8447 31813
rect 8389 31804 8401 31807
rect 8352 31776 8401 31804
rect 8352 31764 8358 31776
rect 8389 31773 8401 31776
rect 8435 31773 8447 31807
rect 8570 31804 8576 31816
rect 8389 31767 8447 31773
rect 8496 31776 8576 31804
rect 7469 31739 7527 31745
rect 7469 31736 7481 31739
rect 6748 31708 7481 31736
rect 7469 31705 7481 31708
rect 7515 31736 7527 31739
rect 7558 31736 7564 31748
rect 7515 31708 7564 31736
rect 7515 31705 7527 31708
rect 7469 31699 7527 31705
rect 7558 31696 7564 31708
rect 7616 31696 7622 31748
rect 7650 31696 7656 31748
rect 7708 31736 7714 31748
rect 8113 31739 8171 31745
rect 8113 31736 8125 31739
rect 7708 31708 8125 31736
rect 7708 31696 7714 31708
rect 8113 31705 8125 31708
rect 8159 31736 8171 31739
rect 8496 31736 8524 31776
rect 8570 31764 8576 31776
rect 8628 31804 8634 31816
rect 9214 31804 9220 31816
rect 8628 31776 9220 31804
rect 8628 31764 8634 31776
rect 9214 31764 9220 31776
rect 9272 31764 9278 31816
rect 9585 31807 9643 31813
rect 9585 31773 9597 31807
rect 9631 31773 9643 31807
rect 9585 31767 9643 31773
rect 9677 31807 9735 31813
rect 9677 31773 9689 31807
rect 9723 31804 9735 31807
rect 9766 31804 9772 31816
rect 9723 31776 9772 31804
rect 9723 31773 9735 31776
rect 9677 31767 9735 31773
rect 8159 31708 8524 31736
rect 8159 31705 8171 31708
rect 8113 31699 8171 31705
rect 8662 31696 8668 31748
rect 8720 31736 8726 31748
rect 9600 31736 9628 31767
rect 9766 31764 9772 31776
rect 9824 31764 9830 31816
rect 10410 31764 10416 31816
rect 10468 31764 10474 31816
rect 10502 31764 10508 31816
rect 10560 31804 10566 31816
rect 10704 31813 10732 31844
rect 11330 31832 11336 31844
rect 11388 31832 11394 31884
rect 11716 31844 12388 31872
rect 10597 31807 10655 31813
rect 10597 31804 10609 31807
rect 10560 31776 10609 31804
rect 10560 31764 10566 31776
rect 10597 31773 10609 31776
rect 10643 31773 10655 31807
rect 10597 31767 10655 31773
rect 10689 31807 10747 31813
rect 10689 31773 10701 31807
rect 10735 31773 10747 31807
rect 10689 31767 10747 31773
rect 10778 31764 10784 31816
rect 10836 31764 10842 31816
rect 11514 31764 11520 31816
rect 11572 31764 11578 31816
rect 11716 31813 11744 31844
rect 11701 31807 11759 31813
rect 11701 31773 11713 31807
rect 11747 31773 11759 31807
rect 11701 31767 11759 31773
rect 8720 31708 9628 31736
rect 12360 31736 12388 31844
rect 12452 31813 12480 31912
rect 12986 31900 12992 31912
rect 13044 31940 13050 31952
rect 13188 31940 13216 31980
rect 13906 31968 13912 31980
rect 13964 31968 13970 32020
rect 14458 31968 14464 32020
rect 14516 32008 14522 32020
rect 14918 32008 14924 32020
rect 14516 31980 14924 32008
rect 14516 31968 14522 31980
rect 14918 31968 14924 31980
rect 14976 31968 14982 32020
rect 16206 31968 16212 32020
rect 16264 31968 16270 32020
rect 16850 31968 16856 32020
rect 16908 32008 16914 32020
rect 17129 32011 17187 32017
rect 17129 32008 17141 32011
rect 16908 31980 17141 32008
rect 16908 31968 16914 31980
rect 17129 31977 17141 31980
rect 17175 31977 17187 32011
rect 17129 31971 17187 31977
rect 17494 31968 17500 32020
rect 17552 32008 17558 32020
rect 17552 31980 18368 32008
rect 17552 31968 17558 31980
rect 13044 31912 13216 31940
rect 13044 31900 13050 31912
rect 13446 31900 13452 31952
rect 13504 31940 13510 31952
rect 15286 31940 15292 31952
rect 13504 31912 15292 31940
rect 13504 31900 13510 31912
rect 15286 31900 15292 31912
rect 15344 31900 15350 31952
rect 15381 31943 15439 31949
rect 15381 31909 15393 31943
rect 15427 31909 15439 31943
rect 15381 31903 15439 31909
rect 16485 31943 16543 31949
rect 16485 31909 16497 31943
rect 16531 31940 16543 31943
rect 16574 31940 16580 31952
rect 16531 31912 16580 31940
rect 16531 31909 16543 31912
rect 16485 31903 16543 31909
rect 12526 31832 12532 31884
rect 12584 31872 12590 31884
rect 12584 31844 13308 31872
rect 12584 31832 12590 31844
rect 12437 31807 12495 31813
rect 12437 31773 12449 31807
rect 12483 31773 12495 31807
rect 12437 31767 12495 31773
rect 12986 31764 12992 31816
rect 13044 31804 13050 31816
rect 13170 31804 13176 31816
rect 13044 31776 13176 31804
rect 13044 31764 13050 31776
rect 13170 31764 13176 31776
rect 13228 31764 13234 31816
rect 13280 31813 13308 31844
rect 14182 31832 14188 31884
rect 14240 31872 14246 31884
rect 15010 31872 15016 31884
rect 14240 31844 15016 31872
rect 14240 31832 14246 31844
rect 15010 31832 15016 31844
rect 15068 31832 15074 31884
rect 15396 31872 15424 31903
rect 16574 31900 16580 31912
rect 16632 31900 16638 31952
rect 17954 31900 17960 31952
rect 18012 31900 18018 31952
rect 17494 31872 17500 31884
rect 15396 31844 17500 31872
rect 17494 31832 17500 31844
rect 17552 31832 17558 31884
rect 17972 31872 18000 31900
rect 18340 31872 18368 31980
rect 18782 31968 18788 32020
rect 18840 32008 18846 32020
rect 19886 32008 19892 32020
rect 18840 31980 19892 32008
rect 18840 31968 18846 31980
rect 19886 31968 19892 31980
rect 19944 31968 19950 32020
rect 19981 32011 20039 32017
rect 19981 31977 19993 32011
rect 20027 31977 20039 32011
rect 19981 31971 20039 31977
rect 20349 32011 20407 32017
rect 20349 31977 20361 32011
rect 20395 32008 20407 32011
rect 20990 32008 20996 32020
rect 20395 31980 20996 32008
rect 20395 31977 20407 31980
rect 20349 31971 20407 31977
rect 18414 31900 18420 31952
rect 18472 31940 18478 31952
rect 18509 31943 18567 31949
rect 18509 31940 18521 31943
rect 18472 31912 18521 31940
rect 18472 31900 18478 31912
rect 18509 31909 18521 31912
rect 18555 31909 18567 31943
rect 18509 31903 18567 31909
rect 18874 31900 18880 31952
rect 18932 31940 18938 31952
rect 19996 31940 20024 31971
rect 20990 31968 20996 31980
rect 21048 31968 21054 32020
rect 21177 32011 21235 32017
rect 21177 31977 21189 32011
rect 21223 32008 21235 32011
rect 22370 32008 22376 32020
rect 21223 31980 22376 32008
rect 21223 31977 21235 31980
rect 21177 31971 21235 31977
rect 22370 31968 22376 31980
rect 22428 31968 22434 32020
rect 22462 31968 22468 32020
rect 22520 32008 22526 32020
rect 22646 32008 22652 32020
rect 22520 31980 22652 32008
rect 22520 31968 22526 31980
rect 22646 31968 22652 31980
rect 22704 31968 22710 32020
rect 24762 31968 24768 32020
rect 24820 31968 24826 32020
rect 26510 32008 26516 32020
rect 24965 31980 26516 32008
rect 18932 31912 20024 31940
rect 18932 31900 18938 31912
rect 20622 31900 20628 31952
rect 20680 31940 20686 31952
rect 21266 31940 21272 31952
rect 20680 31912 21272 31940
rect 20680 31900 20686 31912
rect 21266 31900 21272 31912
rect 21324 31900 21330 31952
rect 21358 31900 21364 31952
rect 21416 31900 21422 31952
rect 24965 31940 24993 31980
rect 26510 31968 26516 31980
rect 26568 31968 26574 32020
rect 26878 31968 26884 32020
rect 26936 32008 26942 32020
rect 27614 32008 27620 32020
rect 26936 31980 27620 32008
rect 26936 31968 26942 31980
rect 27614 31968 27620 31980
rect 27672 31968 27678 32020
rect 28350 31968 28356 32020
rect 28408 32008 28414 32020
rect 28445 32011 28503 32017
rect 28445 32008 28457 32011
rect 28408 31980 28457 32008
rect 28408 31968 28414 31980
rect 28445 31977 28457 31980
rect 28491 31977 28503 32011
rect 31754 32008 31760 32020
rect 28445 31971 28503 31977
rect 28920 31980 31760 32008
rect 25314 31940 25320 31952
rect 23308 31912 24993 31940
rect 25148 31912 25320 31940
rect 20073 31875 20131 31881
rect 17972 31844 18276 31872
rect 18340 31844 19840 31872
rect 13265 31807 13323 31813
rect 13265 31773 13277 31807
rect 13311 31773 13323 31807
rect 13265 31767 13323 31773
rect 13354 31764 13360 31816
rect 13412 31804 13418 31816
rect 13630 31804 13636 31816
rect 13412 31776 13636 31804
rect 13412 31764 13418 31776
rect 13630 31764 13636 31776
rect 13688 31764 13694 31816
rect 14274 31764 14280 31816
rect 14332 31764 14338 31816
rect 14458 31764 14464 31816
rect 14516 31804 14522 31816
rect 15197 31807 15255 31813
rect 15197 31804 15209 31807
rect 14516 31776 15209 31804
rect 14516 31764 14522 31776
rect 15197 31773 15209 31776
rect 15243 31804 15255 31807
rect 15470 31804 15476 31816
rect 15243 31776 15476 31804
rect 15243 31773 15255 31776
rect 15197 31767 15255 31773
rect 15470 31764 15476 31776
rect 15528 31764 15534 31816
rect 16114 31764 16120 31816
rect 16172 31764 16178 31816
rect 16298 31764 16304 31816
rect 16356 31764 16362 31816
rect 17770 31804 17776 31816
rect 16399 31776 17776 31804
rect 12360 31708 14780 31736
rect 8720 31696 8726 31708
rect 6638 31668 6644 31680
rect 6472 31640 6644 31668
rect 5905 31631 5963 31637
rect 6638 31628 6644 31640
rect 6696 31628 6702 31680
rect 6730 31628 6736 31680
rect 6788 31668 6794 31680
rect 7926 31668 7932 31680
rect 6788 31640 7932 31668
rect 6788 31628 6794 31640
rect 7926 31628 7932 31640
rect 7984 31628 7990 31680
rect 8202 31628 8208 31680
rect 8260 31668 8266 31680
rect 8573 31671 8631 31677
rect 8573 31668 8585 31671
rect 8260 31640 8585 31668
rect 8260 31628 8266 31640
rect 8573 31637 8585 31640
rect 8619 31637 8631 31671
rect 8573 31631 8631 31637
rect 9030 31628 9036 31680
rect 9088 31668 9094 31680
rect 9217 31671 9275 31677
rect 9217 31668 9229 31671
rect 9088 31640 9229 31668
rect 9088 31628 9094 31640
rect 9217 31637 9229 31640
rect 9263 31637 9275 31671
rect 9217 31631 9275 31637
rect 10686 31628 10692 31680
rect 10744 31668 10750 31680
rect 10965 31671 11023 31677
rect 10965 31668 10977 31671
rect 10744 31640 10977 31668
rect 10744 31628 10750 31640
rect 10965 31637 10977 31640
rect 11011 31637 11023 31671
rect 10965 31631 11023 31637
rect 12342 31628 12348 31680
rect 12400 31668 12406 31680
rect 13446 31668 13452 31680
rect 12400 31640 13452 31668
rect 12400 31628 12406 31640
rect 13446 31628 13452 31640
rect 13504 31628 13510 31680
rect 14366 31628 14372 31680
rect 14424 31628 14430 31680
rect 14752 31668 14780 31708
rect 14826 31696 14832 31748
rect 14884 31736 14890 31748
rect 14921 31739 14979 31745
rect 14921 31736 14933 31739
rect 14884 31708 14933 31736
rect 14884 31696 14890 31708
rect 14921 31705 14933 31708
rect 14967 31705 14979 31739
rect 14921 31699 14979 31705
rect 15286 31696 15292 31748
rect 15344 31736 15350 31748
rect 16399 31736 16427 31776
rect 17770 31764 17776 31776
rect 17828 31804 17834 31816
rect 17957 31807 18015 31813
rect 17957 31804 17969 31807
rect 17828 31776 17969 31804
rect 17828 31764 17834 31776
rect 17957 31773 17969 31776
rect 18003 31773 18015 31807
rect 18248 31804 18276 31844
rect 18325 31807 18383 31813
rect 18325 31804 18337 31807
rect 18248 31776 18337 31804
rect 17957 31767 18015 31773
rect 18325 31773 18337 31776
rect 18371 31773 18383 31807
rect 18598 31804 18604 31816
rect 18325 31767 18383 31773
rect 18432 31776 18604 31804
rect 15344 31708 16427 31736
rect 16945 31739 17003 31745
rect 15344 31696 15350 31708
rect 16945 31705 16957 31739
rect 16991 31736 17003 31739
rect 17402 31736 17408 31748
rect 16991 31708 17408 31736
rect 16991 31705 17003 31708
rect 16945 31699 17003 31705
rect 17402 31696 17408 31708
rect 17460 31696 17466 31748
rect 18141 31739 18199 31745
rect 18141 31705 18153 31739
rect 18187 31705 18199 31739
rect 18141 31699 18199 31705
rect 18233 31739 18291 31745
rect 18233 31705 18245 31739
rect 18279 31736 18291 31739
rect 18432 31736 18460 31776
rect 18598 31764 18604 31776
rect 18656 31764 18662 31816
rect 19812 31813 19840 31844
rect 20073 31841 20085 31875
rect 20119 31872 20131 31875
rect 20806 31872 20812 31884
rect 20119 31844 20812 31872
rect 20119 31841 20131 31844
rect 20073 31835 20131 31841
rect 20806 31832 20812 31844
rect 20864 31832 20870 31884
rect 21726 31872 21732 31884
rect 20916 31844 21732 31872
rect 19797 31807 19855 31813
rect 19797 31773 19809 31807
rect 19843 31773 19855 31807
rect 19797 31767 19855 31773
rect 19886 31764 19892 31816
rect 19944 31804 19950 31816
rect 20916 31804 20944 31844
rect 21726 31832 21732 31844
rect 21784 31832 21790 31884
rect 23014 31832 23020 31884
rect 23072 31872 23078 31884
rect 23308 31881 23336 31912
rect 23293 31875 23351 31881
rect 23293 31872 23305 31875
rect 23072 31844 23305 31872
rect 23072 31832 23078 31844
rect 23293 31841 23305 31844
rect 23339 31841 23351 31875
rect 23293 31835 23351 31841
rect 24946 31832 24952 31884
rect 25004 31832 25010 31884
rect 25038 31832 25044 31884
rect 25096 31832 25102 31884
rect 25148 31881 25176 31912
rect 25314 31900 25320 31912
rect 25372 31900 25378 31952
rect 25682 31900 25688 31952
rect 25740 31940 25746 31952
rect 26145 31943 26203 31949
rect 26145 31940 26157 31943
rect 25740 31912 26157 31940
rect 25740 31900 25746 31912
rect 26145 31909 26157 31912
rect 26191 31909 26203 31943
rect 26145 31903 26203 31909
rect 26237 31943 26295 31949
rect 26237 31909 26249 31943
rect 26283 31940 26295 31943
rect 26970 31940 26976 31952
rect 26283 31912 26976 31940
rect 26283 31909 26295 31912
rect 26237 31903 26295 31909
rect 26970 31900 26976 31912
rect 27028 31900 27034 31952
rect 27522 31900 27528 31952
rect 27580 31940 27586 31952
rect 28920 31940 28948 31980
rect 31754 31968 31760 31980
rect 31812 31968 31818 32020
rect 31938 31968 31944 32020
rect 31996 32008 32002 32020
rect 31996 31980 33180 32008
rect 31996 31968 32002 31980
rect 27580 31912 28948 31940
rect 27580 31900 27586 31912
rect 28994 31900 29000 31952
rect 29052 31900 29058 31952
rect 29196 31912 29684 31940
rect 25133 31875 25191 31881
rect 25133 31841 25145 31875
rect 25179 31841 25191 31875
rect 25133 31835 25191 31841
rect 25225 31875 25283 31881
rect 25225 31841 25237 31875
rect 25271 31872 25283 31875
rect 25406 31872 25412 31884
rect 25271 31844 25412 31872
rect 25271 31841 25283 31844
rect 25225 31835 25283 31841
rect 25406 31832 25412 31844
rect 25464 31832 25470 31884
rect 19944 31776 20944 31804
rect 19944 31764 19950 31776
rect 20990 31764 20996 31816
rect 21048 31764 21054 31816
rect 21085 31807 21143 31813
rect 21085 31773 21097 31807
rect 21131 31773 21143 31807
rect 21085 31767 21143 31773
rect 18279 31708 18460 31736
rect 18279 31705 18291 31708
rect 18233 31699 18291 31705
rect 17034 31668 17040 31680
rect 14752 31640 17040 31668
rect 17034 31628 17040 31640
rect 17092 31628 17098 31680
rect 17126 31628 17132 31680
rect 17184 31677 17190 31680
rect 17184 31671 17203 31677
rect 17191 31637 17203 31671
rect 17184 31631 17203 31637
rect 17313 31671 17371 31677
rect 17313 31637 17325 31671
rect 17359 31668 17371 31671
rect 17770 31668 17776 31680
rect 17359 31640 17776 31668
rect 17359 31637 17371 31640
rect 17313 31631 17371 31637
rect 17184 31628 17190 31631
rect 17770 31628 17776 31640
rect 17828 31668 17834 31680
rect 18046 31668 18052 31680
rect 17828 31640 18052 31668
rect 17828 31628 17834 31640
rect 18046 31628 18052 31640
rect 18104 31668 18110 31680
rect 18156 31668 18184 31699
rect 20070 31696 20076 31748
rect 20128 31736 20134 31748
rect 20530 31736 20536 31748
rect 20128 31708 20536 31736
rect 20128 31696 20134 31708
rect 20530 31696 20536 31708
rect 20588 31696 20594 31748
rect 21100 31736 21128 31767
rect 21910 31764 21916 31816
rect 21968 31764 21974 31816
rect 22094 31764 22100 31816
rect 22152 31764 22158 31816
rect 22554 31764 22560 31816
rect 22612 31804 22618 31816
rect 22741 31807 22799 31813
rect 22741 31804 22753 31807
rect 22612 31776 22753 31804
rect 22612 31764 22618 31776
rect 22741 31773 22753 31776
rect 22787 31773 22799 31807
rect 22741 31767 22799 31773
rect 22925 31807 22983 31813
rect 22925 31773 22937 31807
rect 22971 31804 22983 31807
rect 23382 31804 23388 31816
rect 22971 31776 23388 31804
rect 22971 31773 22983 31776
rect 22925 31767 22983 31773
rect 23382 31764 23388 31776
rect 23440 31764 23446 31816
rect 23937 31807 23995 31813
rect 23937 31773 23949 31807
rect 23983 31804 23995 31807
rect 25700 31804 25728 31900
rect 25774 31832 25780 31884
rect 25832 31832 25838 31884
rect 26050 31832 26056 31884
rect 26108 31872 26114 31884
rect 26329 31875 26387 31881
rect 26329 31872 26341 31875
rect 26108 31844 26341 31872
rect 26108 31832 26114 31844
rect 26329 31841 26341 31844
rect 26375 31872 26387 31875
rect 26418 31872 26424 31884
rect 26375 31844 26424 31872
rect 26375 31841 26387 31844
rect 26329 31835 26387 31841
rect 26418 31832 26424 31844
rect 26476 31832 26482 31884
rect 26510 31832 26516 31884
rect 26568 31872 26574 31884
rect 29196 31872 29224 31912
rect 26568 31844 29224 31872
rect 26568 31832 26574 31844
rect 23983 31776 25728 31804
rect 27433 31807 27491 31813
rect 23983 31773 23995 31776
rect 23937 31767 23995 31773
rect 27433 31773 27445 31807
rect 27479 31804 27491 31807
rect 28442 31804 28448 31816
rect 27479 31776 28448 31804
rect 27479 31773 27491 31776
rect 27433 31767 27491 31773
rect 28442 31764 28448 31776
rect 28500 31764 28506 31816
rect 28626 31764 28632 31816
rect 28684 31764 28690 31816
rect 28813 31807 28871 31813
rect 28813 31773 28825 31807
rect 28859 31773 28871 31807
rect 28813 31767 28871 31773
rect 21450 31736 21456 31748
rect 21100 31708 21456 31736
rect 21450 31696 21456 31708
rect 21508 31696 21514 31748
rect 24026 31736 24032 31748
rect 22066 31708 24032 31736
rect 18104 31640 18184 31668
rect 18104 31628 18110 31640
rect 18874 31628 18880 31680
rect 18932 31668 18938 31680
rect 22066 31668 22094 31708
rect 24026 31696 24032 31708
rect 24084 31696 24090 31748
rect 24578 31696 24584 31748
rect 24636 31736 24642 31748
rect 25038 31736 25044 31748
rect 24636 31708 25044 31736
rect 24636 31696 24642 31708
rect 25038 31696 25044 31708
rect 25096 31736 25102 31748
rect 25096 31708 26648 31736
rect 25096 31696 25102 31708
rect 18932 31640 22094 31668
rect 22281 31671 22339 31677
rect 18932 31628 18938 31640
rect 22281 31637 22293 31671
rect 22327 31668 22339 31671
rect 23382 31668 23388 31680
rect 22327 31640 23388 31668
rect 22327 31637 22339 31640
rect 22281 31631 22339 31637
rect 23382 31628 23388 31640
rect 23440 31628 23446 31680
rect 23934 31628 23940 31680
rect 23992 31628 23998 31680
rect 24486 31628 24492 31680
rect 24544 31668 24550 31680
rect 26050 31668 26056 31680
rect 24544 31640 26056 31668
rect 24544 31628 24550 31640
rect 26050 31628 26056 31640
rect 26108 31628 26114 31680
rect 26620 31677 26648 31708
rect 27706 31696 27712 31748
rect 27764 31696 27770 31748
rect 27890 31696 27896 31748
rect 27948 31736 27954 31748
rect 28353 31739 28411 31745
rect 28353 31736 28365 31739
rect 27948 31708 28365 31736
rect 27948 31696 27954 31708
rect 28353 31705 28365 31708
rect 28399 31705 28411 31739
rect 28353 31699 28411 31705
rect 28534 31696 28540 31748
rect 28592 31736 28598 31748
rect 28828 31736 28856 31767
rect 29546 31764 29552 31816
rect 29604 31764 29610 31816
rect 29564 31736 29592 31764
rect 28592 31708 28856 31736
rect 28920 31708 29592 31736
rect 29656 31736 29684 31912
rect 30006 31900 30012 31952
rect 30064 31900 30070 31952
rect 32490 31900 32496 31952
rect 32548 31940 32554 31952
rect 32858 31940 32864 31952
rect 32548 31912 32864 31940
rect 32548 31900 32554 31912
rect 32858 31900 32864 31912
rect 32916 31900 32922 31952
rect 33152 31940 33180 31980
rect 33502 31968 33508 32020
rect 33560 32008 33566 32020
rect 33597 32011 33655 32017
rect 33597 32008 33609 32011
rect 33560 31980 33609 32008
rect 33560 31968 33566 31980
rect 33597 31977 33609 31980
rect 33643 31977 33655 32011
rect 34606 32008 34612 32020
rect 33597 31971 33655 31977
rect 33693 31980 34612 32008
rect 33693 31940 33721 31980
rect 34606 31968 34612 31980
rect 34664 31968 34670 32020
rect 35526 32008 35532 32020
rect 34900 31980 35532 32008
rect 33152 31912 33721 31940
rect 34054 31900 34060 31952
rect 34112 31900 34118 31952
rect 29822 31832 29828 31884
rect 29880 31832 29886 31884
rect 30024 31872 30052 31900
rect 31852 31884 31904 31890
rect 29932 31844 30052 31872
rect 29733 31807 29791 31813
rect 29733 31773 29745 31807
rect 29779 31804 29791 31807
rect 29932 31804 29960 31844
rect 30098 31832 30104 31884
rect 30156 31872 30162 31884
rect 30282 31872 30288 31884
rect 30156 31844 30288 31872
rect 30156 31832 30162 31844
rect 30282 31832 30288 31844
rect 30340 31832 30346 31884
rect 30377 31875 30435 31881
rect 30377 31841 30389 31875
rect 30423 31872 30435 31875
rect 30466 31872 30472 31884
rect 30423 31844 30472 31872
rect 30423 31841 30435 31844
rect 30377 31835 30435 31841
rect 30466 31832 30472 31844
rect 30524 31832 30530 31884
rect 30926 31832 30932 31884
rect 30984 31872 30990 31884
rect 31113 31875 31171 31881
rect 31113 31872 31125 31875
rect 30984 31844 31125 31872
rect 30984 31832 30990 31844
rect 31113 31841 31125 31844
rect 31159 31872 31171 31875
rect 31202 31872 31208 31884
rect 31159 31844 31208 31872
rect 31159 31841 31171 31844
rect 31113 31835 31171 31841
rect 31202 31832 31208 31844
rect 31260 31832 31266 31884
rect 34900 31881 34928 31980
rect 35526 31968 35532 31980
rect 35584 32008 35590 32020
rect 36538 32008 36544 32020
rect 35584 31980 36544 32008
rect 35584 31968 35590 31980
rect 36538 31968 36544 31980
rect 36596 32008 36602 32020
rect 36998 32008 37004 32020
rect 36596 31980 37004 32008
rect 36596 31968 36602 31980
rect 36998 31968 37004 31980
rect 37056 31968 37062 32020
rect 36265 31943 36323 31949
rect 36265 31909 36277 31943
rect 36311 31909 36323 31943
rect 36265 31903 36323 31909
rect 34885 31875 34943 31881
rect 31852 31826 31904 31832
rect 33061 31844 34837 31872
rect 29779 31776 29960 31804
rect 29779 31773 29791 31776
rect 29733 31767 29791 31773
rect 30006 31764 30012 31816
rect 30064 31804 30070 31816
rect 30190 31804 30196 31816
rect 30064 31776 30196 31804
rect 30064 31764 30070 31776
rect 30190 31764 30196 31776
rect 30248 31764 30254 31816
rect 31478 31764 31484 31816
rect 31536 31764 31542 31816
rect 32125 31807 32183 31813
rect 32125 31773 32137 31807
rect 32171 31773 32183 31807
rect 32125 31767 32183 31773
rect 32140 31736 32168 31767
rect 32950 31764 32956 31816
rect 33008 31764 33014 31816
rect 33061 31813 33089 31844
rect 33046 31807 33104 31813
rect 33046 31773 33058 31807
rect 33092 31773 33104 31807
rect 33046 31767 33104 31773
rect 29656 31708 32168 31736
rect 28592 31696 28598 31708
rect 26605 31671 26663 31677
rect 26605 31637 26617 31671
rect 26651 31668 26663 31671
rect 27246 31668 27252 31680
rect 26651 31640 27252 31668
rect 26651 31637 26663 31640
rect 26605 31631 26663 31637
rect 27246 31628 27252 31640
rect 27304 31628 27310 31680
rect 28258 31628 28264 31680
rect 28316 31668 28322 31680
rect 28920 31668 28948 31708
rect 32214 31696 32220 31748
rect 32272 31736 32278 31748
rect 33061 31736 33089 31767
rect 33410 31764 33416 31816
rect 33468 31813 33474 31816
rect 33468 31804 33476 31813
rect 33468 31776 33513 31804
rect 33468 31767 33476 31776
rect 33468 31764 33474 31767
rect 33594 31764 33600 31816
rect 33652 31804 33658 31816
rect 33652 31776 33916 31804
rect 33652 31764 33658 31776
rect 32272 31708 33089 31736
rect 32272 31696 32278 31708
rect 33226 31696 33232 31748
rect 33284 31696 33290 31748
rect 33318 31696 33324 31748
rect 33376 31696 33382 31748
rect 33888 31736 33916 31776
rect 33962 31764 33968 31816
rect 34020 31804 34026 31816
rect 34333 31807 34391 31813
rect 34333 31804 34345 31807
rect 34020 31776 34345 31804
rect 34020 31764 34026 31776
rect 34333 31773 34345 31776
rect 34379 31773 34391 31807
rect 34809 31804 34837 31844
rect 34885 31841 34897 31875
rect 34931 31841 34943 31875
rect 36280 31872 36308 31903
rect 36446 31900 36452 31952
rect 36504 31940 36510 31952
rect 36633 31943 36691 31949
rect 36633 31940 36645 31943
rect 36504 31912 36645 31940
rect 36504 31900 36510 31912
rect 36633 31909 36645 31912
rect 36679 31909 36691 31943
rect 36633 31903 36691 31909
rect 36280 31844 36492 31872
rect 34885 31835 34943 31841
rect 35158 31813 35164 31816
rect 34809 31776 35112 31804
rect 34333 31767 34391 31773
rect 34057 31739 34115 31745
rect 34057 31736 34069 31739
rect 33888 31708 34069 31736
rect 34057 31705 34069 31708
rect 34103 31705 34115 31739
rect 34057 31699 34115 31705
rect 34241 31739 34299 31745
rect 34241 31705 34253 31739
rect 34287 31736 34299 31739
rect 34514 31736 34520 31748
rect 34287 31708 34520 31736
rect 34287 31705 34299 31708
rect 34241 31699 34299 31705
rect 34514 31696 34520 31708
rect 34572 31696 34578 31748
rect 34698 31696 34704 31748
rect 34756 31736 34762 31748
rect 34882 31736 34888 31748
rect 34756 31708 34888 31736
rect 34756 31696 34762 31708
rect 34882 31696 34888 31708
rect 34940 31696 34946 31748
rect 35084 31736 35112 31776
rect 35152 31767 35164 31813
rect 35216 31804 35222 31816
rect 35216 31776 35252 31804
rect 35158 31764 35164 31767
rect 35216 31764 35222 31776
rect 36464 31736 36492 31844
rect 36814 31832 36820 31884
rect 36872 31832 36878 31884
rect 37084 31807 37142 31813
rect 37084 31773 37096 31807
rect 37130 31804 37142 31807
rect 37458 31804 37464 31816
rect 37130 31776 37464 31804
rect 37130 31773 37142 31776
rect 37084 31767 37142 31773
rect 37458 31764 37464 31776
rect 37516 31764 37522 31816
rect 38010 31736 38016 31748
rect 35084 31708 36400 31736
rect 36464 31708 38016 31736
rect 28316 31640 28948 31668
rect 28316 31628 28322 31640
rect 29546 31628 29552 31680
rect 29604 31668 29610 31680
rect 30190 31668 30196 31680
rect 29604 31640 30196 31668
rect 29604 31628 29610 31640
rect 30190 31628 30196 31640
rect 30248 31628 30254 31680
rect 31570 31628 31576 31680
rect 31628 31668 31634 31680
rect 31874 31671 31932 31677
rect 31874 31668 31886 31671
rect 31628 31640 31886 31668
rect 31628 31628 31634 31640
rect 31874 31637 31886 31640
rect 31920 31637 31932 31671
rect 31874 31631 31932 31637
rect 32950 31628 32956 31680
rect 33008 31668 33014 31680
rect 33336 31668 33364 31696
rect 36372 31680 36400 31708
rect 38010 31696 38016 31708
rect 38068 31696 38074 31748
rect 33008 31640 33364 31668
rect 33008 31628 33014 31640
rect 33502 31628 33508 31680
rect 33560 31668 33566 31680
rect 34422 31668 34428 31680
rect 33560 31640 34428 31668
rect 33560 31628 33566 31640
rect 34422 31628 34428 31640
rect 34480 31628 34486 31680
rect 34606 31628 34612 31680
rect 34664 31668 34670 31680
rect 35250 31668 35256 31680
rect 34664 31640 35256 31668
rect 34664 31628 34670 31640
rect 35250 31628 35256 31640
rect 35308 31668 35314 31680
rect 35802 31668 35808 31680
rect 35308 31640 35808 31668
rect 35308 31628 35314 31640
rect 35802 31628 35808 31640
rect 35860 31628 35866 31680
rect 36354 31628 36360 31680
rect 36412 31628 36418 31680
rect 36814 31628 36820 31680
rect 36872 31668 36878 31680
rect 37182 31668 37188 31680
rect 36872 31640 37188 31668
rect 36872 31628 36878 31640
rect 37182 31628 37188 31640
rect 37240 31628 37246 31680
rect 37826 31628 37832 31680
rect 37884 31668 37890 31680
rect 38197 31671 38255 31677
rect 38197 31668 38209 31671
rect 37884 31640 38209 31668
rect 37884 31628 37890 31640
rect 38197 31637 38209 31640
rect 38243 31637 38255 31671
rect 38197 31631 38255 31637
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 10870 31464 10876 31476
rect 7116 31436 10876 31464
rect 5166 31288 5172 31340
rect 5224 31288 5230 31340
rect 5353 31331 5411 31337
rect 5353 31297 5365 31331
rect 5399 31297 5411 31331
rect 5353 31291 5411 31297
rect 5074 31220 5080 31272
rect 5132 31260 5138 31272
rect 5368 31260 5396 31291
rect 5718 31288 5724 31340
rect 5776 31328 5782 31340
rect 5813 31331 5871 31337
rect 5813 31328 5825 31331
rect 5776 31300 5825 31328
rect 5776 31288 5782 31300
rect 5813 31297 5825 31300
rect 5859 31297 5871 31331
rect 5813 31291 5871 31297
rect 5997 31331 6055 31337
rect 5997 31297 6009 31331
rect 6043 31328 6055 31331
rect 6730 31328 6736 31340
rect 6043 31300 6736 31328
rect 6043 31297 6055 31300
rect 5997 31291 6055 31297
rect 6730 31288 6736 31300
rect 6788 31288 6794 31340
rect 7116 31337 7144 31436
rect 10870 31424 10876 31436
rect 10928 31424 10934 31476
rect 10962 31424 10968 31476
rect 11020 31464 11026 31476
rect 12710 31464 12716 31476
rect 11020 31436 12716 31464
rect 11020 31424 11026 31436
rect 12710 31424 12716 31436
rect 12768 31424 12774 31476
rect 13630 31424 13636 31476
rect 13688 31424 13694 31476
rect 14366 31424 14372 31476
rect 14424 31464 14430 31476
rect 20990 31464 20996 31476
rect 14424 31436 20996 31464
rect 14424 31424 14430 31436
rect 20990 31424 20996 31436
rect 21048 31424 21054 31476
rect 21174 31424 21180 31476
rect 21232 31464 21238 31476
rect 22186 31464 22192 31476
rect 21232 31436 22192 31464
rect 21232 31424 21238 31436
rect 22186 31424 22192 31436
rect 22244 31424 22250 31476
rect 23106 31424 23112 31476
rect 23164 31464 23170 31476
rect 32030 31464 32036 31476
rect 23164 31436 25912 31464
rect 23164 31424 23170 31436
rect 7377 31399 7435 31405
rect 7377 31365 7389 31399
rect 7423 31396 7435 31399
rect 7834 31396 7840 31408
rect 7423 31368 7840 31396
rect 7423 31365 7435 31368
rect 7377 31359 7435 31365
rect 7834 31356 7840 31368
rect 7892 31356 7898 31408
rect 8938 31396 8944 31408
rect 8220 31368 8944 31396
rect 7101 31331 7159 31337
rect 7101 31297 7113 31331
rect 7147 31297 7159 31331
rect 7101 31291 7159 31297
rect 7190 31288 7196 31340
rect 7248 31328 7254 31340
rect 7285 31331 7343 31337
rect 7285 31328 7297 31331
rect 7248 31300 7297 31328
rect 7248 31288 7254 31300
rect 7285 31297 7297 31300
rect 7331 31328 7343 31331
rect 7650 31328 7656 31340
rect 7331 31300 7656 31328
rect 7331 31297 7343 31300
rect 7285 31291 7343 31297
rect 7650 31288 7656 31300
rect 7708 31288 7714 31340
rect 7926 31288 7932 31340
rect 7984 31288 7990 31340
rect 8018 31288 8024 31340
rect 8076 31288 8082 31340
rect 8220 31337 8248 31368
rect 8938 31356 8944 31368
rect 8996 31356 9002 31408
rect 9214 31356 9220 31408
rect 9272 31396 9278 31408
rect 9490 31396 9496 31408
rect 9272 31368 9496 31396
rect 9272 31356 9278 31368
rect 9490 31356 9496 31368
rect 9548 31356 9554 31408
rect 10686 31396 10692 31408
rect 9692 31368 10692 31396
rect 8205 31331 8263 31337
rect 8205 31297 8217 31331
rect 8251 31297 8263 31331
rect 8205 31291 8263 31297
rect 8849 31331 8907 31337
rect 8849 31297 8861 31331
rect 8895 31297 8907 31331
rect 8849 31291 8907 31297
rect 9033 31331 9091 31337
rect 9033 31297 9045 31331
rect 9079 31328 9091 31331
rect 9398 31328 9404 31340
rect 9079 31300 9404 31328
rect 9079 31297 9091 31300
rect 9033 31291 9091 31297
rect 5132 31232 5396 31260
rect 5132 31220 5138 31232
rect 5368 31192 5396 31232
rect 5902 31220 5908 31272
rect 5960 31220 5966 31272
rect 7742 31220 7748 31272
rect 7800 31260 7806 31272
rect 8665 31263 8723 31269
rect 8665 31260 8677 31263
rect 7800 31232 8677 31260
rect 7800 31220 7806 31232
rect 8665 31229 8677 31232
rect 8711 31260 8723 31263
rect 8754 31260 8760 31272
rect 8711 31232 8760 31260
rect 8711 31229 8723 31232
rect 8665 31223 8723 31229
rect 8754 31220 8760 31232
rect 8812 31220 8818 31272
rect 7650 31192 7656 31204
rect 5368 31164 7656 31192
rect 7650 31152 7656 31164
rect 7708 31152 7714 31204
rect 7834 31152 7840 31204
rect 7892 31192 7898 31204
rect 8864 31192 8892 31291
rect 9398 31288 9404 31300
rect 9456 31288 9462 31340
rect 9692 31337 9720 31368
rect 10686 31356 10692 31368
rect 10744 31356 10750 31408
rect 11330 31356 11336 31408
rect 11388 31396 11394 31408
rect 13648 31396 13676 31424
rect 11388 31368 13676 31396
rect 11388 31356 11394 31368
rect 9677 31331 9735 31337
rect 9677 31297 9689 31331
rect 9723 31297 9735 31331
rect 10137 31331 10195 31337
rect 10137 31328 10149 31331
rect 9677 31291 9735 31297
rect 9784 31300 10149 31328
rect 9306 31220 9312 31272
rect 9364 31260 9370 31272
rect 9784 31260 9812 31300
rect 10137 31297 10149 31300
rect 10183 31297 10195 31331
rect 10137 31291 10195 31297
rect 10870 31288 10876 31340
rect 10928 31288 10934 31340
rect 11054 31288 11060 31340
rect 11112 31288 11118 31340
rect 12342 31288 12348 31340
rect 12400 31288 12406 31340
rect 12434 31288 12440 31340
rect 12492 31328 12498 31340
rect 12912 31337 12940 31368
rect 13722 31356 13728 31408
rect 13780 31396 13786 31408
rect 15194 31396 15200 31408
rect 13780 31368 14044 31396
rect 13780 31356 13786 31368
rect 12529 31331 12587 31337
rect 12529 31328 12541 31331
rect 12492 31300 12541 31328
rect 12492 31288 12498 31300
rect 12529 31297 12541 31300
rect 12575 31297 12587 31331
rect 12529 31291 12587 31297
rect 12897 31331 12955 31337
rect 12897 31297 12909 31331
rect 12943 31297 12955 31331
rect 12897 31291 12955 31297
rect 13078 31288 13084 31340
rect 13136 31328 13142 31340
rect 13357 31331 13415 31337
rect 13357 31328 13369 31331
rect 13136 31300 13369 31328
rect 13136 31288 13142 31300
rect 13357 31297 13369 31300
rect 13403 31328 13415 31331
rect 13403 31300 13492 31328
rect 13403 31297 13415 31300
rect 13357 31291 13415 31297
rect 9364 31232 9812 31260
rect 9364 31220 9370 31232
rect 9858 31220 9864 31272
rect 9916 31220 9922 31272
rect 9953 31263 10011 31269
rect 9953 31229 9965 31263
rect 9999 31260 10011 31263
rect 11149 31263 11207 31269
rect 9999 31232 11100 31260
rect 9999 31229 10011 31232
rect 9953 31223 10011 31229
rect 11072 31204 11100 31232
rect 11149 31229 11161 31263
rect 11195 31229 11207 31263
rect 11149 31223 11207 31229
rect 7892 31164 8892 31192
rect 7892 31152 7898 31164
rect 8938 31152 8944 31204
rect 8996 31192 9002 31204
rect 8996 31164 9674 31192
rect 8996 31152 9002 31164
rect 5169 31127 5227 31133
rect 5169 31093 5181 31127
rect 5215 31124 5227 31127
rect 5442 31124 5448 31136
rect 5215 31096 5448 31124
rect 5215 31093 5227 31096
rect 5169 31087 5227 31093
rect 5442 31084 5448 31096
rect 5500 31084 5506 31136
rect 8294 31084 8300 31136
rect 8352 31124 8358 31136
rect 9030 31124 9036 31136
rect 8352 31096 9036 31124
rect 8352 31084 8358 31096
rect 9030 31084 9036 31096
rect 9088 31084 9094 31136
rect 9122 31084 9128 31136
rect 9180 31124 9186 31136
rect 9493 31127 9551 31133
rect 9493 31124 9505 31127
rect 9180 31096 9505 31124
rect 9180 31084 9186 31096
rect 9493 31093 9505 31096
rect 9539 31093 9551 31127
rect 9646 31124 9674 31164
rect 9766 31152 9772 31204
rect 9824 31192 9830 31204
rect 10410 31192 10416 31204
rect 9824 31164 10416 31192
rect 9824 31152 9830 31164
rect 10410 31152 10416 31164
rect 10468 31152 10474 31204
rect 11054 31152 11060 31204
rect 11112 31152 11118 31204
rect 11164 31192 11192 31223
rect 11514 31220 11520 31272
rect 11572 31260 11578 31272
rect 12618 31260 12624 31272
rect 11572 31232 12624 31260
rect 11572 31220 11578 31232
rect 12618 31220 12624 31232
rect 12676 31260 12682 31272
rect 13262 31260 13268 31272
rect 12676 31232 13268 31260
rect 12676 31220 12682 31232
rect 13262 31220 13268 31232
rect 13320 31220 13326 31272
rect 13464 31260 13492 31300
rect 13538 31288 13544 31340
rect 13596 31328 13602 31340
rect 13633 31331 13691 31337
rect 13633 31328 13645 31331
rect 13596 31300 13645 31328
rect 13596 31288 13602 31300
rect 13633 31297 13645 31300
rect 13679 31328 13691 31331
rect 13814 31328 13820 31340
rect 13679 31300 13820 31328
rect 13679 31297 13691 31300
rect 13633 31291 13691 31297
rect 13814 31288 13820 31300
rect 13872 31288 13878 31340
rect 13906 31288 13912 31340
rect 13964 31288 13970 31340
rect 14016 31337 14044 31368
rect 14844 31368 15200 31396
rect 14844 31337 14872 31368
rect 15194 31356 15200 31368
rect 15252 31356 15258 31408
rect 15930 31356 15936 31408
rect 15988 31396 15994 31408
rect 16117 31399 16175 31405
rect 16117 31396 16129 31399
rect 15988 31368 16129 31396
rect 15988 31356 15994 31368
rect 16117 31365 16129 31368
rect 16163 31396 16175 31399
rect 17586 31396 17592 31408
rect 16163 31368 17592 31396
rect 16163 31365 16175 31368
rect 16117 31359 16175 31365
rect 17586 31356 17592 31368
rect 17644 31356 17650 31408
rect 18230 31356 18236 31408
rect 18288 31396 18294 31408
rect 18386 31399 18444 31405
rect 18386 31396 18398 31399
rect 18288 31368 18398 31396
rect 18288 31356 18294 31368
rect 18386 31365 18398 31368
rect 18432 31365 18444 31399
rect 18386 31359 18444 31365
rect 20438 31356 20444 31408
rect 20496 31356 20502 31408
rect 23658 31396 23664 31408
rect 20916 31368 23664 31396
rect 14001 31331 14059 31337
rect 14001 31297 14013 31331
rect 14047 31297 14059 31331
rect 14001 31291 14059 31297
rect 14829 31331 14887 31337
rect 14829 31297 14841 31331
rect 14875 31297 14887 31331
rect 14829 31291 14887 31297
rect 13722 31260 13728 31272
rect 13464 31232 13728 31260
rect 13722 31220 13728 31232
rect 13780 31220 13786 31272
rect 14185 31263 14243 31269
rect 14185 31229 14197 31263
rect 14231 31260 14243 31263
rect 14366 31260 14372 31272
rect 14231 31232 14372 31260
rect 14231 31229 14243 31232
rect 14185 31223 14243 31229
rect 14366 31220 14372 31232
rect 14424 31220 14430 31272
rect 11974 31192 11980 31204
rect 11164 31164 11980 31192
rect 11974 31152 11980 31164
rect 12032 31192 12038 31204
rect 12802 31192 12808 31204
rect 12032 31164 12808 31192
rect 12032 31152 12038 31164
rect 12802 31152 12808 31164
rect 12860 31152 12866 31204
rect 14844 31192 14872 31291
rect 14918 31288 14924 31340
rect 14976 31328 14982 31340
rect 15289 31331 15347 31337
rect 15289 31328 15301 31331
rect 14976 31300 15301 31328
rect 14976 31288 14982 31300
rect 15289 31297 15301 31300
rect 15335 31297 15347 31331
rect 15289 31291 15347 31297
rect 16850 31288 16856 31340
rect 16908 31288 16914 31340
rect 17126 31328 17132 31340
rect 16960 31300 17132 31328
rect 15010 31220 15016 31272
rect 15068 31260 15074 31272
rect 15381 31263 15439 31269
rect 15381 31260 15393 31263
rect 15068 31232 15393 31260
rect 15068 31220 15074 31232
rect 15381 31229 15393 31232
rect 15427 31260 15439 31263
rect 16960 31260 16988 31300
rect 17126 31288 17132 31300
rect 17184 31288 17190 31340
rect 17402 31288 17408 31340
rect 17460 31328 17466 31340
rect 19426 31328 19432 31340
rect 17460 31300 19432 31328
rect 17460 31288 17466 31300
rect 19426 31288 19432 31300
rect 19484 31288 19490 31340
rect 20254 31337 20260 31340
rect 20248 31291 20260 31337
rect 20254 31288 20260 31291
rect 20312 31288 20318 31340
rect 20456 31328 20484 31356
rect 20916 31328 20944 31368
rect 20456 31300 20944 31328
rect 22462 31288 22468 31340
rect 22520 31328 22526 31340
rect 22520 31300 22600 31328
rect 22520 31288 22526 31300
rect 15427 31232 16988 31260
rect 17037 31263 17095 31269
rect 15427 31229 15439 31232
rect 15381 31223 15439 31229
rect 17037 31229 17049 31263
rect 17083 31229 17095 31263
rect 17037 31223 17095 31229
rect 18141 31263 18199 31269
rect 18141 31229 18153 31263
rect 18187 31229 18199 31263
rect 18141 31223 18199 31229
rect 13924 31164 14872 31192
rect 9950 31124 9956 31136
rect 9646 31096 9956 31124
rect 9493 31087 9551 31093
rect 9950 31084 9956 31096
rect 10008 31124 10014 31136
rect 10870 31124 10876 31136
rect 10008 31096 10876 31124
rect 10008 31084 10014 31096
rect 10870 31084 10876 31096
rect 10928 31084 10934 31136
rect 12250 31084 12256 31136
rect 12308 31124 12314 31136
rect 12618 31124 12624 31136
rect 12308 31096 12624 31124
rect 12308 31084 12314 31096
rect 12618 31084 12624 31096
rect 12676 31084 12682 31136
rect 12710 31084 12716 31136
rect 12768 31124 12774 31136
rect 13924 31124 13952 31164
rect 15194 31152 15200 31204
rect 15252 31192 15258 31204
rect 16574 31192 16580 31204
rect 15252 31164 16580 31192
rect 15252 31152 15258 31164
rect 16574 31152 16580 31164
rect 16632 31152 16638 31204
rect 16850 31152 16856 31204
rect 16908 31192 16914 31204
rect 17052 31192 17080 31223
rect 16908 31164 17080 31192
rect 16908 31152 16914 31164
rect 18156 31136 18184 31223
rect 19334 31220 19340 31272
rect 19392 31260 19398 31272
rect 19981 31263 20039 31269
rect 19981 31260 19993 31263
rect 19392 31232 19993 31260
rect 19392 31220 19398 31232
rect 19981 31229 19993 31232
rect 20027 31229 20039 31263
rect 22572 31260 22600 31300
rect 22646 31288 22652 31340
rect 22704 31288 22710 31340
rect 23198 31328 23204 31340
rect 22756 31300 23204 31328
rect 22756 31260 22784 31300
rect 23198 31288 23204 31300
rect 23256 31288 23262 31340
rect 23308 31337 23336 31368
rect 23658 31356 23664 31368
rect 23716 31356 23722 31408
rect 23293 31331 23351 31337
rect 23293 31297 23305 31331
rect 23339 31297 23351 31331
rect 23293 31291 23351 31297
rect 23382 31288 23388 31340
rect 23440 31328 23446 31340
rect 25498 31328 25504 31340
rect 23440 31300 25504 31328
rect 23440 31288 23446 31300
rect 25498 31288 25504 31300
rect 25556 31288 25562 31340
rect 25590 31288 25596 31340
rect 25648 31288 25654 31340
rect 22572 31232 22784 31260
rect 19981 31223 20039 31229
rect 23106 31220 23112 31272
rect 23164 31260 23170 31272
rect 23753 31263 23811 31269
rect 23753 31260 23765 31263
rect 23164 31232 23765 31260
rect 23164 31220 23170 31232
rect 23753 31229 23765 31232
rect 23799 31229 23811 31263
rect 25884 31260 25912 31436
rect 26896 31436 32036 31464
rect 25961 31331 26019 31337
rect 25961 31297 25973 31331
rect 26007 31328 26019 31331
rect 26896 31328 26924 31436
rect 32030 31424 32036 31436
rect 32088 31424 32094 31476
rect 32490 31424 32496 31476
rect 32548 31424 32554 31476
rect 33318 31464 33324 31476
rect 33152 31436 33324 31464
rect 27614 31356 27620 31408
rect 27672 31396 27678 31408
rect 29086 31396 29092 31408
rect 27672 31368 29092 31396
rect 27672 31356 27678 31368
rect 29086 31356 29092 31368
rect 29144 31356 29150 31408
rect 29196 31368 29684 31396
rect 26007 31300 26924 31328
rect 26007 31297 26019 31300
rect 25961 31291 26019 31297
rect 26970 31288 26976 31340
rect 27028 31328 27034 31340
rect 27249 31331 27307 31337
rect 27249 31328 27261 31331
rect 27028 31300 27261 31328
rect 27028 31288 27034 31300
rect 27249 31297 27261 31300
rect 27295 31297 27307 31331
rect 27249 31291 27307 31297
rect 28077 31331 28135 31337
rect 28077 31297 28089 31331
rect 28123 31297 28135 31331
rect 28077 31291 28135 31297
rect 25884 31232 27292 31260
rect 23753 31223 23811 31229
rect 21266 31152 21272 31204
rect 21324 31192 21330 31204
rect 24946 31192 24952 31204
rect 21324 31164 24952 31192
rect 21324 31152 21330 31164
rect 24946 31152 24952 31164
rect 25004 31152 25010 31204
rect 27154 31192 27160 31204
rect 25976 31164 27160 31192
rect 12768 31096 13952 31124
rect 12768 31084 12774 31096
rect 16114 31084 16120 31136
rect 16172 31124 16178 31136
rect 16209 31127 16267 31133
rect 16209 31124 16221 31127
rect 16172 31096 16221 31124
rect 16172 31084 16178 31096
rect 16209 31093 16221 31096
rect 16255 31124 16267 31127
rect 17218 31124 17224 31136
rect 16255 31096 17224 31124
rect 16255 31093 16267 31096
rect 16209 31087 16267 31093
rect 17218 31084 17224 31096
rect 17276 31084 17282 31136
rect 18138 31084 18144 31136
rect 18196 31124 18202 31136
rect 18506 31124 18512 31136
rect 18196 31096 18512 31124
rect 18196 31084 18202 31096
rect 18506 31084 18512 31096
rect 18564 31084 18570 31136
rect 19058 31084 19064 31136
rect 19116 31124 19122 31136
rect 19521 31127 19579 31133
rect 19521 31124 19533 31127
rect 19116 31096 19533 31124
rect 19116 31084 19122 31096
rect 19521 31093 19533 31096
rect 19567 31124 19579 31127
rect 19978 31124 19984 31136
rect 19567 31096 19984 31124
rect 19567 31093 19579 31096
rect 19521 31087 19579 31093
rect 19978 31084 19984 31096
rect 20036 31084 20042 31136
rect 20622 31084 20628 31136
rect 20680 31124 20686 31136
rect 21361 31127 21419 31133
rect 21361 31124 21373 31127
rect 20680 31096 21373 31124
rect 20680 31084 20686 31096
rect 21361 31093 21373 31096
rect 21407 31124 21419 31127
rect 21818 31124 21824 31136
rect 21407 31096 21824 31124
rect 21407 31093 21419 31096
rect 21361 31087 21419 31093
rect 21818 31084 21824 31096
rect 21876 31084 21882 31136
rect 21910 31084 21916 31136
rect 21968 31124 21974 31136
rect 22554 31124 22560 31136
rect 21968 31096 22560 31124
rect 21968 31084 21974 31096
rect 22554 31084 22560 31096
rect 22612 31084 22618 31136
rect 22738 31084 22744 31136
rect 22796 31084 22802 31136
rect 25976 31133 26004 31164
rect 27154 31152 27160 31164
rect 27212 31152 27218 31204
rect 25961 31127 26019 31133
rect 25961 31093 25973 31127
rect 26007 31093 26019 31127
rect 25961 31087 26019 31093
rect 26142 31084 26148 31136
rect 26200 31084 26206 31136
rect 27264 31124 27292 31232
rect 27522 31220 27528 31272
rect 27580 31220 27586 31272
rect 28092 31192 28120 31291
rect 28626 31288 28632 31340
rect 28684 31328 28690 31340
rect 29196 31328 29224 31368
rect 28684 31300 29224 31328
rect 28684 31288 28690 31300
rect 29270 31288 29276 31340
rect 29328 31288 29334 31340
rect 29656 31328 29684 31368
rect 29730 31356 29736 31408
rect 29788 31396 29794 31408
rect 30101 31399 30159 31405
rect 30101 31396 30113 31399
rect 29788 31368 30113 31396
rect 29788 31356 29794 31368
rect 30101 31365 30113 31368
rect 30147 31365 30159 31399
rect 30101 31359 30159 31365
rect 30190 31356 30196 31408
rect 30248 31396 30254 31408
rect 30285 31399 30343 31405
rect 30285 31396 30297 31399
rect 30248 31368 30297 31396
rect 30248 31356 30254 31368
rect 30285 31365 30297 31368
rect 30331 31365 30343 31399
rect 32508 31396 32536 31424
rect 33152 31405 33180 31436
rect 33318 31424 33324 31436
rect 33376 31424 33382 31476
rect 34054 31424 34060 31476
rect 34112 31464 34118 31476
rect 34514 31464 34520 31476
rect 34112 31436 34520 31464
rect 34112 31424 34118 31436
rect 34514 31424 34520 31436
rect 34572 31424 34578 31476
rect 37458 31424 37464 31476
rect 37516 31424 37522 31476
rect 33137 31399 33195 31405
rect 30285 31359 30343 31365
rect 30576 31368 32536 31396
rect 32784 31368 32997 31396
rect 30576 31328 30604 31368
rect 29656 31300 30604 31328
rect 30650 31288 30656 31340
rect 30708 31328 30714 31340
rect 31021 31331 31079 31337
rect 31021 31328 31033 31331
rect 30708 31300 31033 31328
rect 30708 31288 30714 31300
rect 31021 31297 31033 31300
rect 31067 31297 31079 31331
rect 31021 31291 31079 31297
rect 31386 31288 31392 31340
rect 31444 31328 31450 31340
rect 31481 31331 31539 31337
rect 31481 31328 31493 31331
rect 31444 31300 31493 31328
rect 31444 31288 31450 31300
rect 31481 31297 31493 31300
rect 31527 31297 31539 31331
rect 32306 31328 32312 31340
rect 31481 31291 31539 31297
rect 31588 31300 32312 31328
rect 28534 31220 28540 31272
rect 28592 31220 28598 31272
rect 29288 31260 29316 31288
rect 29288 31232 30972 31260
rect 30834 31192 30840 31204
rect 28092 31164 30840 31192
rect 30834 31152 30840 31164
rect 30892 31152 30898 31204
rect 30944 31192 30972 31232
rect 31202 31220 31208 31272
rect 31260 31260 31266 31272
rect 31588 31269 31616 31300
rect 32306 31288 32312 31300
rect 32364 31288 32370 31340
rect 32490 31288 32496 31340
rect 32548 31328 32554 31340
rect 32784 31328 32812 31368
rect 32548 31300 32812 31328
rect 32548 31288 32554 31300
rect 32858 31288 32864 31340
rect 32916 31288 32922 31340
rect 32969 31337 32997 31368
rect 33137 31365 33149 31399
rect 33183 31365 33195 31399
rect 33137 31359 33195 31365
rect 33229 31399 33287 31405
rect 33229 31365 33241 31399
rect 33275 31396 33287 31399
rect 33502 31396 33508 31408
rect 33275 31368 33508 31396
rect 33275 31365 33287 31368
rect 33229 31359 33287 31365
rect 33502 31356 33508 31368
rect 33560 31356 33566 31408
rect 34238 31356 34244 31408
rect 34296 31356 34302 31408
rect 34698 31356 34704 31408
rect 34756 31396 34762 31408
rect 35345 31399 35403 31405
rect 35345 31396 35357 31399
rect 34756 31368 35357 31396
rect 34756 31356 34762 31368
rect 35345 31365 35357 31368
rect 35391 31365 35403 31399
rect 37826 31396 37832 31408
rect 35345 31359 35403 31365
rect 36372 31368 37832 31396
rect 36372 31340 36400 31368
rect 37826 31356 37832 31368
rect 37884 31356 37890 31408
rect 32954 31331 33012 31337
rect 32954 31297 32966 31331
rect 33000 31297 33012 31331
rect 32954 31291 33012 31297
rect 33326 31331 33384 31337
rect 33326 31297 33338 31331
rect 33372 31328 33384 31331
rect 33965 31331 34023 31337
rect 33372 31300 33406 31328
rect 33372 31297 33384 31300
rect 33326 31291 33384 31297
rect 33965 31297 33977 31331
rect 34011 31297 34023 31331
rect 33965 31291 34023 31297
rect 34113 31331 34171 31337
rect 34113 31297 34125 31331
rect 34159 31328 34171 31331
rect 34333 31331 34391 31337
rect 34159 31300 34284 31328
rect 34159 31297 34171 31300
rect 34113 31291 34171 31297
rect 31573 31263 31631 31269
rect 31573 31260 31585 31263
rect 31260 31232 31585 31260
rect 31260 31220 31266 31232
rect 31573 31229 31585 31232
rect 31619 31229 31631 31263
rect 31573 31223 31631 31229
rect 31754 31220 31760 31272
rect 31812 31260 31818 31272
rect 33134 31260 33140 31272
rect 31812 31232 33140 31260
rect 31812 31220 31818 31232
rect 33134 31220 33140 31232
rect 33192 31220 33198 31272
rect 33226 31220 33232 31272
rect 33284 31260 33290 31272
rect 33341 31260 33369 31291
rect 33410 31260 33416 31272
rect 33284 31232 33416 31260
rect 33284 31220 33290 31232
rect 33410 31220 33416 31232
rect 33468 31220 33474 31272
rect 32122 31192 32128 31204
rect 30944 31164 32128 31192
rect 32122 31152 32128 31164
rect 32180 31152 32186 31204
rect 33505 31195 33563 31201
rect 33505 31161 33517 31195
rect 33551 31192 33563 31195
rect 33980 31192 34008 31291
rect 33551 31164 34008 31192
rect 34256 31192 34284 31300
rect 34333 31297 34345 31331
rect 34379 31297 34391 31331
rect 34333 31291 34391 31297
rect 34348 31260 34376 31291
rect 34422 31288 34428 31340
rect 34480 31337 34486 31340
rect 34480 31328 34488 31337
rect 34480 31300 34525 31328
rect 34480 31291 34488 31300
rect 34480 31288 34486 31291
rect 34790 31288 34796 31340
rect 34848 31288 34854 31340
rect 35069 31331 35127 31337
rect 35069 31297 35081 31331
rect 35115 31297 35127 31331
rect 35069 31291 35127 31297
rect 34808 31260 34836 31288
rect 34348 31232 34836 31260
rect 35084 31260 35112 31291
rect 35250 31288 35256 31340
rect 35308 31288 35314 31340
rect 35434 31288 35440 31340
rect 35492 31288 35498 31340
rect 36078 31288 36084 31340
rect 36136 31328 36142 31340
rect 36354 31337 36360 31340
rect 36173 31331 36231 31337
rect 36173 31328 36185 31331
rect 36136 31300 36185 31328
rect 36136 31288 36142 31300
rect 36173 31297 36185 31300
rect 36219 31297 36231 31331
rect 36173 31291 36231 31297
rect 36321 31331 36360 31337
rect 36321 31297 36333 31331
rect 36321 31291 36360 31297
rect 36354 31288 36360 31291
rect 36412 31288 36418 31340
rect 36449 31331 36507 31337
rect 36449 31297 36461 31331
rect 36495 31297 36507 31331
rect 36449 31291 36507 31297
rect 36541 31331 36599 31337
rect 36541 31297 36553 31331
rect 36587 31297 36599 31331
rect 36541 31291 36599 31297
rect 35802 31260 35808 31272
rect 35084 31232 35808 31260
rect 35802 31220 35808 31232
rect 35860 31220 35866 31272
rect 36464 31260 36492 31291
rect 36188 31232 36492 31260
rect 36556 31260 36584 31291
rect 36630 31288 36636 31340
rect 36688 31337 36694 31340
rect 36688 31328 36696 31337
rect 36688 31300 36733 31328
rect 36688 31291 36696 31300
rect 36688 31288 36694 31291
rect 36814 31288 36820 31340
rect 36872 31288 36878 31340
rect 37921 31331 37979 31337
rect 37921 31328 37933 31331
rect 37246 31300 37933 31328
rect 36832 31260 36860 31288
rect 36556 31232 36860 31260
rect 36188 31204 36216 31232
rect 36648 31204 36676 31232
rect 34256 31164 35848 31192
rect 33551 31161 33563 31164
rect 33505 31155 33563 31161
rect 29270 31124 29276 31136
rect 27264 31096 29276 31124
rect 29270 31084 29276 31096
rect 29328 31084 29334 31136
rect 29730 31084 29736 31136
rect 29788 31124 29794 31136
rect 30190 31124 30196 31136
rect 29788 31096 30196 31124
rect 29788 31084 29794 31096
rect 30190 31084 30196 31096
rect 30248 31124 30254 31136
rect 30285 31127 30343 31133
rect 30285 31124 30297 31127
rect 30248 31096 30297 31124
rect 30248 31084 30254 31096
rect 30285 31093 30297 31096
rect 30331 31093 30343 31127
rect 30285 31087 30343 31093
rect 30466 31084 30472 31136
rect 30524 31084 30530 31136
rect 31202 31084 31208 31136
rect 31260 31124 31266 31136
rect 34146 31124 34152 31136
rect 31260 31096 34152 31124
rect 31260 31084 31266 31096
rect 34146 31084 34152 31096
rect 34204 31124 34210 31136
rect 34422 31124 34428 31136
rect 34204 31096 34428 31124
rect 34204 31084 34210 31096
rect 34422 31084 34428 31096
rect 34480 31084 34486 31136
rect 34609 31127 34667 31133
rect 34609 31093 34621 31127
rect 34655 31124 34667 31127
rect 34974 31124 34980 31136
rect 34655 31096 34980 31124
rect 34655 31093 34667 31096
rect 34609 31087 34667 31093
rect 34974 31084 34980 31096
rect 35032 31084 35038 31136
rect 35621 31127 35679 31133
rect 35621 31093 35633 31127
rect 35667 31124 35679 31127
rect 35710 31124 35716 31136
rect 35667 31096 35716 31124
rect 35667 31093 35679 31096
rect 35621 31087 35679 31093
rect 35710 31084 35716 31096
rect 35768 31084 35774 31136
rect 35820 31124 35848 31164
rect 36170 31152 36176 31204
rect 36228 31152 36234 31204
rect 36630 31152 36636 31204
rect 36688 31152 36694 31204
rect 36262 31124 36268 31136
rect 35820 31096 36268 31124
rect 36262 31084 36268 31096
rect 36320 31084 36326 31136
rect 36814 31084 36820 31136
rect 36872 31124 36878 31136
rect 37246 31124 37274 31300
rect 37921 31297 37933 31300
rect 37967 31297 37979 31331
rect 37921 31291 37979 31297
rect 38102 31220 38108 31272
rect 38160 31220 38166 31272
rect 36872 31096 37274 31124
rect 36872 31084 36878 31096
rect 37366 31084 37372 31136
rect 37424 31124 37430 31136
rect 37918 31124 37924 31136
rect 37424 31096 37924 31124
rect 37424 31084 37430 31096
rect 37918 31084 37924 31096
rect 37976 31084 37982 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 5905 30923 5963 30929
rect 5905 30889 5917 30923
rect 5951 30920 5963 30923
rect 5994 30920 6000 30932
rect 5951 30892 6000 30920
rect 5951 30889 5963 30892
rect 5905 30883 5963 30889
rect 5994 30880 6000 30892
rect 6052 30880 6058 30932
rect 6457 30923 6515 30929
rect 6457 30889 6469 30923
rect 6503 30920 6515 30923
rect 8202 30920 8208 30932
rect 6503 30892 8208 30920
rect 6503 30889 6515 30892
rect 6457 30883 6515 30889
rect 8202 30880 8208 30892
rect 8260 30880 8266 30932
rect 8573 30923 8631 30929
rect 8573 30889 8585 30923
rect 8619 30920 8631 30923
rect 11054 30920 11060 30932
rect 8619 30892 11060 30920
rect 8619 30889 8631 30892
rect 8573 30883 8631 30889
rect 11054 30880 11060 30892
rect 11112 30880 11118 30932
rect 11517 30923 11575 30929
rect 11517 30889 11529 30923
rect 11563 30920 11575 30923
rect 12158 30920 12164 30932
rect 11563 30892 12164 30920
rect 11563 30889 11575 30892
rect 11517 30883 11575 30889
rect 12158 30880 12164 30892
rect 12216 30880 12222 30932
rect 14458 30920 14464 30932
rect 12360 30892 14464 30920
rect 9030 30812 9036 30864
rect 9088 30852 9094 30864
rect 11701 30855 11759 30861
rect 11701 30852 11713 30855
rect 9088 30824 11713 30852
rect 9088 30812 9094 30824
rect 11701 30821 11713 30824
rect 11747 30852 11759 30855
rect 12250 30852 12256 30864
rect 11747 30824 12256 30852
rect 11747 30821 11759 30824
rect 11701 30815 11759 30821
rect 12250 30812 12256 30824
rect 12308 30812 12314 30864
rect 4893 30787 4951 30793
rect 4893 30753 4905 30787
rect 4939 30784 4951 30787
rect 7098 30784 7104 30796
rect 4939 30756 5396 30784
rect 4939 30753 4951 30756
rect 4893 30747 4951 30753
rect 5368 30728 5396 30756
rect 5828 30756 7104 30784
rect 5169 30719 5227 30725
rect 5169 30685 5181 30719
rect 5215 30685 5227 30719
rect 5169 30679 5227 30685
rect 5184 30648 5212 30679
rect 5350 30676 5356 30728
rect 5408 30676 5414 30728
rect 5828 30725 5856 30756
rect 7098 30744 7104 30756
rect 7156 30744 7162 30796
rect 8478 30744 8484 30796
rect 8536 30784 8542 30796
rect 8938 30784 8944 30796
rect 8536 30756 8944 30784
rect 8536 30744 8542 30756
rect 8938 30744 8944 30756
rect 8996 30784 9002 30796
rect 9585 30787 9643 30793
rect 8996 30756 9444 30784
rect 8996 30744 9002 30756
rect 5813 30719 5871 30725
rect 5813 30685 5825 30719
rect 5859 30685 5871 30719
rect 5813 30679 5871 30685
rect 6457 30719 6515 30725
rect 6457 30685 6469 30719
rect 6503 30716 6515 30719
rect 6638 30716 6644 30728
rect 6503 30688 6644 30716
rect 6503 30685 6515 30688
rect 6457 30679 6515 30685
rect 6638 30676 6644 30688
rect 6696 30676 6702 30728
rect 6733 30719 6791 30725
rect 6733 30685 6745 30719
rect 6779 30716 6791 30719
rect 6914 30716 6920 30728
rect 6779 30688 6920 30716
rect 6779 30685 6791 30688
rect 6733 30679 6791 30685
rect 6914 30676 6920 30688
rect 6972 30676 6978 30728
rect 7193 30719 7251 30725
rect 7193 30685 7205 30719
rect 7239 30716 7251 30719
rect 7282 30716 7288 30728
rect 7239 30688 7288 30716
rect 7239 30685 7251 30688
rect 7193 30679 7251 30685
rect 7282 30676 7288 30688
rect 7340 30676 7346 30728
rect 9416 30725 9444 30756
rect 9585 30753 9597 30787
rect 9631 30784 9643 30787
rect 9674 30784 9680 30796
rect 9631 30756 9680 30784
rect 9631 30753 9643 30756
rect 9585 30747 9643 30753
rect 9674 30744 9680 30756
rect 9732 30744 9738 30796
rect 10134 30744 10140 30796
rect 10192 30784 10198 30796
rect 10413 30787 10471 30793
rect 10413 30784 10425 30787
rect 10192 30756 10425 30784
rect 10192 30744 10198 30756
rect 10413 30753 10425 30756
rect 10459 30753 10471 30787
rect 10413 30747 10471 30753
rect 11422 30744 11428 30796
rect 11480 30784 11486 30796
rect 12360 30784 12388 30892
rect 14458 30880 14464 30892
rect 14516 30880 14522 30932
rect 14645 30923 14703 30929
rect 14645 30889 14657 30923
rect 14691 30920 14703 30923
rect 14826 30920 14832 30932
rect 14691 30892 14832 30920
rect 14691 30889 14703 30892
rect 14645 30883 14703 30889
rect 14826 30880 14832 30892
rect 14884 30880 14890 30932
rect 16132 30892 17172 30920
rect 12989 30855 13047 30861
rect 12989 30821 13001 30855
rect 13035 30852 13047 30855
rect 16132 30852 16160 30892
rect 13035 30824 16160 30852
rect 13035 30821 13047 30824
rect 12989 30815 13047 30821
rect 11480 30756 12388 30784
rect 11480 30744 11486 30756
rect 7460 30719 7518 30725
rect 7460 30685 7472 30719
rect 7506 30716 7518 30719
rect 9217 30719 9275 30725
rect 7506 30688 8524 30716
rect 7506 30685 7518 30688
rect 7460 30679 7518 30685
rect 8496 30660 8524 30688
rect 9217 30685 9229 30719
rect 9263 30685 9275 30719
rect 9217 30682 9275 30685
rect 9140 30679 9275 30682
rect 9401 30719 9459 30725
rect 9401 30685 9413 30719
rect 9447 30685 9459 30719
rect 9401 30679 9459 30685
rect 5721 30651 5779 30657
rect 5721 30648 5733 30651
rect 5184 30620 5733 30648
rect 5721 30617 5733 30620
rect 5767 30648 5779 30651
rect 5767 30620 7604 30648
rect 5767 30617 5779 30620
rect 5721 30611 5779 30617
rect 5074 30540 5080 30592
rect 5132 30580 5138 30592
rect 5261 30583 5319 30589
rect 5261 30580 5273 30583
rect 5132 30552 5273 30580
rect 5132 30540 5138 30552
rect 5261 30549 5273 30552
rect 5307 30549 5319 30583
rect 5261 30543 5319 30549
rect 6641 30583 6699 30589
rect 6641 30549 6653 30583
rect 6687 30580 6699 30583
rect 7466 30580 7472 30592
rect 6687 30552 7472 30580
rect 6687 30549 6699 30552
rect 6641 30543 6699 30549
rect 7466 30540 7472 30552
rect 7524 30540 7530 30592
rect 7576 30580 7604 30620
rect 8478 30608 8484 30660
rect 8536 30608 8542 30660
rect 8754 30608 8760 30660
rect 8812 30648 8818 30660
rect 9140 30654 9260 30679
rect 9490 30676 9496 30728
rect 9548 30716 9554 30728
rect 10045 30719 10103 30725
rect 10045 30716 10057 30719
rect 9548 30688 10057 30716
rect 9548 30676 9554 30688
rect 10045 30685 10057 30688
rect 10091 30685 10103 30719
rect 10045 30679 10103 30685
rect 10226 30676 10232 30728
rect 10284 30676 10290 30728
rect 12360 30725 12388 30756
rect 12618 30744 12624 30796
rect 12676 30784 12682 30796
rect 13633 30787 13691 30793
rect 13633 30784 13645 30787
rect 12676 30756 13645 30784
rect 12676 30744 12682 30756
rect 13633 30753 13645 30756
rect 13679 30753 13691 30787
rect 13633 30747 13691 30753
rect 14458 30744 14464 30796
rect 14516 30784 14522 30796
rect 15657 30787 15715 30793
rect 15657 30784 15669 30787
rect 14516 30756 15669 30784
rect 14516 30744 14522 30756
rect 15657 30753 15669 30756
rect 15703 30784 15715 30787
rect 15746 30784 15752 30796
rect 15703 30756 15752 30784
rect 15703 30753 15715 30756
rect 15657 30747 15715 30753
rect 15746 30744 15752 30756
rect 15804 30744 15810 30796
rect 17144 30784 17172 30892
rect 17586 30880 17592 30932
rect 17644 30920 17650 30932
rect 19613 30923 19671 30929
rect 19613 30920 19625 30923
rect 17644 30892 19625 30920
rect 17644 30880 17650 30892
rect 19613 30889 19625 30892
rect 19659 30889 19671 30923
rect 19613 30883 19671 30889
rect 20165 30923 20223 30929
rect 20165 30889 20177 30923
rect 20211 30920 20223 30923
rect 20254 30920 20260 30932
rect 20211 30892 20260 30920
rect 20211 30889 20223 30892
rect 20165 30883 20223 30889
rect 20254 30880 20260 30892
rect 20312 30880 20318 30932
rect 21082 30880 21088 30932
rect 21140 30920 21146 30932
rect 21726 30920 21732 30932
rect 21140 30892 21732 30920
rect 21140 30880 21146 30892
rect 21726 30880 21732 30892
rect 21784 30880 21790 30932
rect 23750 30920 23756 30932
rect 22112 30892 23756 30920
rect 18046 30812 18052 30864
rect 18104 30852 18110 30864
rect 22112 30852 22140 30892
rect 23750 30880 23756 30892
rect 23808 30880 23814 30932
rect 23934 30880 23940 30932
rect 23992 30920 23998 30932
rect 23992 30892 27476 30920
rect 23992 30880 23998 30892
rect 22278 30852 22284 30864
rect 18104 30824 22140 30852
rect 22204 30824 22284 30852
rect 18104 30812 18110 30824
rect 20625 30787 20683 30793
rect 20625 30784 20637 30787
rect 17144 30756 20637 30784
rect 20625 30753 20637 30756
rect 20671 30753 20683 30787
rect 20625 30747 20683 30753
rect 20717 30787 20775 30793
rect 20717 30753 20729 30787
rect 20763 30753 20775 30787
rect 22204 30784 22232 30824
rect 22278 30812 22284 30824
rect 22336 30852 22342 30864
rect 22646 30852 22652 30864
rect 22336 30824 22652 30852
rect 22336 30812 22342 30824
rect 22646 30812 22652 30824
rect 22704 30852 22710 30864
rect 23017 30855 23075 30861
rect 23017 30852 23029 30855
rect 22704 30824 23029 30852
rect 22704 30812 22710 30824
rect 23017 30821 23029 30824
rect 23063 30821 23075 30855
rect 23017 30815 23075 30821
rect 20717 30747 20775 30753
rect 21836 30756 22232 30784
rect 10321 30719 10379 30725
rect 10321 30685 10333 30719
rect 10367 30685 10379 30719
rect 10321 30679 10379 30685
rect 10597 30719 10655 30725
rect 10597 30685 10609 30719
rect 10643 30716 10655 30719
rect 12345 30719 12403 30725
rect 10643 30688 12296 30716
rect 10643 30685 10655 30688
rect 10597 30679 10655 30685
rect 9140 30648 9168 30654
rect 8812 30620 9168 30648
rect 8812 30608 8818 30620
rect 8386 30580 8392 30592
rect 7576 30552 8392 30580
rect 8386 30540 8392 30552
rect 8444 30540 8450 30592
rect 9140 30580 9168 30620
rect 9582 30608 9588 30660
rect 9640 30648 9646 30660
rect 10336 30648 10364 30679
rect 9640 30620 10364 30648
rect 9640 30608 9646 30620
rect 11330 30608 11336 30660
rect 11388 30608 11394 30660
rect 11514 30608 11520 30660
rect 11572 30657 11578 30660
rect 11572 30651 11591 30657
rect 11579 30617 11591 30651
rect 11572 30611 11591 30617
rect 11572 30608 11578 30611
rect 12066 30608 12072 30660
rect 12124 30648 12130 30660
rect 12161 30651 12219 30657
rect 12161 30648 12173 30651
rect 12124 30620 12173 30648
rect 12124 30608 12130 30620
rect 12161 30617 12173 30620
rect 12207 30617 12219 30651
rect 12268 30648 12296 30688
rect 12345 30685 12357 30719
rect 12391 30685 12403 30719
rect 12345 30679 12403 30685
rect 12529 30719 12587 30725
rect 12529 30685 12541 30719
rect 12575 30716 12587 30719
rect 12986 30716 12992 30728
rect 12575 30688 12992 30716
rect 12575 30685 12587 30688
rect 12529 30679 12587 30685
rect 12986 30676 12992 30688
rect 13044 30676 13050 30728
rect 13170 30676 13176 30728
rect 13228 30676 13234 30728
rect 13354 30676 13360 30728
rect 13412 30676 13418 30728
rect 13446 30676 13452 30728
rect 13504 30725 13510 30728
rect 13504 30719 13533 30725
rect 13521 30685 13533 30719
rect 13814 30716 13820 30728
rect 13504 30679 13533 30685
rect 13648 30688 13820 30716
rect 13504 30676 13510 30679
rect 12894 30648 12900 30660
rect 12268 30620 12900 30648
rect 12161 30611 12219 30617
rect 12894 30608 12900 30620
rect 12952 30608 12958 30660
rect 13265 30651 13323 30657
rect 13265 30617 13277 30651
rect 13311 30648 13323 30651
rect 13648 30648 13676 30688
rect 13814 30676 13820 30688
rect 13872 30676 13878 30728
rect 15286 30676 15292 30728
rect 15344 30676 15350 30728
rect 15378 30676 15384 30728
rect 15436 30716 15442 30728
rect 15473 30719 15531 30725
rect 15473 30716 15485 30719
rect 15436 30688 15485 30716
rect 15436 30676 15442 30688
rect 15473 30685 15485 30688
rect 15519 30685 15531 30719
rect 15473 30679 15531 30685
rect 16117 30719 16175 30725
rect 16117 30685 16129 30719
rect 16163 30716 16175 30719
rect 18138 30716 18144 30728
rect 16163 30688 18144 30716
rect 16163 30685 16175 30688
rect 16117 30679 16175 30685
rect 18138 30676 18144 30688
rect 18196 30716 18202 30728
rect 18693 30719 18751 30725
rect 18693 30716 18705 30719
rect 18196 30688 18705 30716
rect 18196 30676 18202 30688
rect 18693 30685 18705 30688
rect 18739 30685 18751 30719
rect 18693 30679 18751 30685
rect 20530 30676 20536 30728
rect 20588 30676 20594 30728
rect 20732 30716 20760 30747
rect 21836 30725 21864 30756
rect 22830 30744 22836 30796
rect 22888 30784 22894 30796
rect 22888 30756 23428 30784
rect 22888 30744 22894 30756
rect 20640 30688 20760 30716
rect 21821 30719 21879 30725
rect 20640 30660 20668 30688
rect 21821 30685 21833 30719
rect 21867 30685 21879 30719
rect 21821 30679 21879 30685
rect 21913 30719 21971 30725
rect 21913 30685 21925 30719
rect 21959 30685 21971 30719
rect 21913 30679 21971 30685
rect 13311 30620 13676 30648
rect 13311 30617 13323 30620
rect 13265 30611 13323 30617
rect 9490 30580 9496 30592
rect 9140 30552 9496 30580
rect 9490 30540 9496 30552
rect 9548 30540 9554 30592
rect 10226 30540 10232 30592
rect 10284 30580 10290 30592
rect 10781 30583 10839 30589
rect 10781 30580 10793 30583
rect 10284 30552 10793 30580
rect 10284 30540 10290 30552
rect 10781 30549 10793 30552
rect 10827 30549 10839 30583
rect 10781 30543 10839 30549
rect 11790 30540 11796 30592
rect 11848 30580 11854 30592
rect 13280 30580 13308 30611
rect 13722 30608 13728 30660
rect 13780 30648 13786 30660
rect 14461 30651 14519 30657
rect 14461 30648 14473 30651
rect 13780 30620 14473 30648
rect 13780 30608 13786 30620
rect 14461 30617 14473 30620
rect 14507 30617 14519 30651
rect 15010 30648 15016 30660
rect 14461 30611 14519 30617
rect 14752 30620 15016 30648
rect 11848 30552 13308 30580
rect 11848 30540 11854 30552
rect 13446 30540 13452 30592
rect 13504 30580 13510 30592
rect 14661 30583 14719 30589
rect 14661 30580 14673 30583
rect 13504 30552 14673 30580
rect 13504 30540 13510 30552
rect 14661 30549 14673 30552
rect 14707 30580 14719 30583
rect 14752 30580 14780 30620
rect 15010 30608 15016 30620
rect 15068 30608 15074 30660
rect 16384 30651 16442 30657
rect 16384 30617 16396 30651
rect 16430 30648 16442 30651
rect 16482 30648 16488 30660
rect 16430 30620 16488 30648
rect 16430 30617 16442 30620
rect 16384 30611 16442 30617
rect 16482 30608 16488 30620
rect 16540 30608 16546 30660
rect 16942 30608 16948 30660
rect 17000 30648 17006 30660
rect 17000 30620 17724 30648
rect 17000 30608 17006 30620
rect 14707 30552 14780 30580
rect 14707 30549 14719 30552
rect 14661 30543 14719 30549
rect 14826 30540 14832 30592
rect 14884 30540 14890 30592
rect 17497 30583 17555 30589
rect 17497 30549 17509 30583
rect 17543 30580 17555 30583
rect 17586 30580 17592 30592
rect 17543 30552 17592 30580
rect 17543 30549 17555 30552
rect 17497 30543 17555 30549
rect 17586 30540 17592 30552
rect 17644 30540 17650 30592
rect 17696 30580 17724 30620
rect 17954 30608 17960 30660
rect 18012 30608 18018 30660
rect 18322 30608 18328 30660
rect 18380 30648 18386 30660
rect 18506 30648 18512 30660
rect 18380 30620 18512 30648
rect 18380 30608 18386 30620
rect 18506 30608 18512 30620
rect 18564 30608 18570 30660
rect 19521 30651 19579 30657
rect 19521 30617 19533 30651
rect 19567 30617 19579 30651
rect 19521 30611 19579 30617
rect 19536 30580 19564 30611
rect 20622 30608 20628 30660
rect 20680 30608 20686 30660
rect 21928 30648 21956 30679
rect 22002 30676 22008 30728
rect 22060 30676 22066 30728
rect 22094 30676 22100 30728
rect 22152 30676 22158 30728
rect 22370 30676 22376 30728
rect 22428 30716 22434 30728
rect 22646 30716 22652 30728
rect 22428 30688 22652 30716
rect 22428 30676 22434 30688
rect 22646 30676 22652 30688
rect 22704 30676 22710 30728
rect 23201 30719 23259 30725
rect 23201 30685 23213 30719
rect 23247 30685 23259 30719
rect 23400 30716 23428 30756
rect 23474 30744 23480 30796
rect 23532 30784 23538 30796
rect 23569 30787 23627 30793
rect 23569 30784 23581 30787
rect 23532 30756 23581 30784
rect 23532 30744 23538 30756
rect 23569 30753 23581 30756
rect 23615 30753 23627 30787
rect 23569 30747 23627 30753
rect 24302 30744 24308 30796
rect 24360 30784 24366 30796
rect 24581 30787 24639 30793
rect 24581 30784 24593 30787
rect 24360 30756 24593 30784
rect 24360 30744 24366 30756
rect 24581 30753 24593 30756
rect 24627 30753 24639 30787
rect 24581 30747 24639 30753
rect 24762 30744 24768 30796
rect 24820 30744 24826 30796
rect 25056 30793 25084 30892
rect 26050 30812 26056 30864
rect 26108 30852 26114 30864
rect 26237 30855 26295 30861
rect 26237 30852 26249 30855
rect 26108 30824 26249 30852
rect 26108 30812 26114 30824
rect 26237 30821 26249 30824
rect 26283 30821 26295 30855
rect 27338 30852 27344 30864
rect 26237 30815 26295 30821
rect 26988 30824 27344 30852
rect 25041 30787 25099 30793
rect 25041 30753 25053 30787
rect 25087 30753 25099 30787
rect 25041 30747 25099 30753
rect 25774 30744 25780 30796
rect 25832 30784 25838 30796
rect 25832 30756 26372 30784
rect 25832 30744 25838 30756
rect 23661 30719 23719 30725
rect 23661 30716 23673 30719
rect 23400 30688 23673 30716
rect 23201 30679 23259 30685
rect 23661 30685 23673 30688
rect 23707 30685 23719 30719
rect 23661 30679 23719 30685
rect 25133 30719 25191 30725
rect 25133 30685 25145 30719
rect 25179 30685 25191 30719
rect 25133 30679 25191 30685
rect 22462 30648 22468 30660
rect 20732 30620 21772 30648
rect 21928 30620 22468 30648
rect 20732 30580 20760 30620
rect 17696 30552 20760 30580
rect 20898 30540 20904 30592
rect 20956 30580 20962 30592
rect 21637 30583 21695 30589
rect 21637 30580 21649 30583
rect 20956 30552 21649 30580
rect 20956 30540 20962 30552
rect 21637 30549 21649 30552
rect 21683 30549 21695 30583
rect 21744 30580 21772 30620
rect 22462 30608 22468 30620
rect 22520 30608 22526 30660
rect 22554 30608 22560 30660
rect 22612 30648 22618 30660
rect 23216 30648 23244 30679
rect 22612 30620 23244 30648
rect 22612 30608 22618 30620
rect 22186 30580 22192 30592
rect 21744 30552 22192 30580
rect 21637 30543 21695 30549
rect 22186 30540 22192 30552
rect 22244 30540 22250 30592
rect 23216 30580 23244 30620
rect 24762 30608 24768 30660
rect 24820 30648 24826 30660
rect 25148 30648 25176 30679
rect 25498 30676 25504 30728
rect 25556 30716 25562 30728
rect 26344 30725 26372 30756
rect 26053 30719 26111 30725
rect 26053 30716 26065 30719
rect 25556 30688 26065 30716
rect 25556 30676 25562 30688
rect 26053 30685 26065 30688
rect 26099 30685 26111 30719
rect 26053 30679 26111 30685
rect 26329 30719 26387 30725
rect 26329 30685 26341 30719
rect 26375 30685 26387 30719
rect 26329 30679 26387 30685
rect 26602 30676 26608 30728
rect 26660 30716 26666 30728
rect 26988 30716 27016 30824
rect 27338 30812 27344 30824
rect 27396 30812 27402 30864
rect 27062 30744 27068 30796
rect 27120 30784 27126 30796
rect 27249 30787 27307 30793
rect 27249 30784 27261 30787
rect 27120 30756 27261 30784
rect 27120 30744 27126 30756
rect 27249 30753 27261 30756
rect 27295 30753 27307 30787
rect 27448 30784 27476 30892
rect 27522 30880 27528 30932
rect 27580 30920 27586 30932
rect 28626 30920 28632 30932
rect 27580 30892 28632 30920
rect 27580 30880 27586 30892
rect 28626 30880 28632 30892
rect 28684 30880 28690 30932
rect 29270 30880 29276 30932
rect 29328 30920 29334 30932
rect 30834 30920 30840 30932
rect 29328 30892 30840 30920
rect 29328 30880 29334 30892
rect 30834 30880 30840 30892
rect 30892 30880 30898 30932
rect 31202 30880 31208 30932
rect 31260 30880 31266 30932
rect 31754 30880 31760 30932
rect 31812 30920 31818 30932
rect 32122 30920 32128 30932
rect 31812 30892 32128 30920
rect 31812 30880 31818 30892
rect 32122 30880 32128 30892
rect 32180 30880 32186 30932
rect 32490 30880 32496 30932
rect 32548 30920 32554 30932
rect 36078 30920 36084 30932
rect 32548 30892 36084 30920
rect 32548 30880 32554 30892
rect 36078 30880 36084 30892
rect 36136 30880 36142 30932
rect 36541 30923 36599 30929
rect 36541 30889 36553 30923
rect 36587 30920 36599 30923
rect 37550 30920 37556 30932
rect 36587 30892 37556 30920
rect 36587 30889 36599 30892
rect 36541 30883 36599 30889
rect 37550 30880 37556 30892
rect 37608 30880 37614 30932
rect 38105 30923 38163 30929
rect 38105 30889 38117 30923
rect 38151 30920 38163 30923
rect 38194 30920 38200 30932
rect 38151 30892 38200 30920
rect 38151 30889 38163 30892
rect 38105 30883 38163 30889
rect 38194 30880 38200 30892
rect 38252 30880 38258 30932
rect 28166 30812 28172 30864
rect 28224 30852 28230 30864
rect 28350 30852 28356 30864
rect 28224 30824 28356 30852
rect 28224 30812 28230 30824
rect 28350 30812 28356 30824
rect 28408 30812 28414 30864
rect 28537 30855 28595 30861
rect 28537 30821 28549 30855
rect 28583 30852 28595 30855
rect 28810 30852 28816 30864
rect 28583 30824 28816 30852
rect 28583 30821 28595 30824
rect 28537 30815 28595 30821
rect 28552 30784 28580 30815
rect 28810 30812 28816 30824
rect 28868 30812 28874 30864
rect 28994 30812 29000 30864
rect 29052 30852 29058 30864
rect 29052 30824 31432 30852
rect 29052 30812 29058 30824
rect 29546 30784 29552 30796
rect 27249 30747 27307 30753
rect 27356 30756 28580 30784
rect 28736 30756 29552 30784
rect 27356 30725 27384 30756
rect 27157 30719 27215 30725
rect 27157 30716 27169 30719
rect 26660 30688 27169 30716
rect 26660 30676 26666 30688
rect 27157 30685 27169 30688
rect 27203 30685 27215 30719
rect 27157 30679 27215 30685
rect 27341 30719 27399 30725
rect 27341 30685 27353 30719
rect 27387 30685 27399 30719
rect 27341 30679 27399 30685
rect 27430 30676 27436 30728
rect 27488 30676 27494 30728
rect 27525 30719 27583 30725
rect 27525 30685 27537 30719
rect 27571 30685 27583 30719
rect 27525 30679 27583 30685
rect 28445 30719 28503 30725
rect 28445 30685 28457 30719
rect 28491 30685 28503 30719
rect 28445 30679 28503 30685
rect 24820 30620 25176 30648
rect 24820 30608 24826 30620
rect 26418 30608 26424 30660
rect 26476 30648 26482 30660
rect 27540 30648 27568 30679
rect 28166 30648 28172 30660
rect 26476 30620 28172 30648
rect 26476 30608 26482 30620
rect 28166 30608 28172 30620
rect 28224 30608 28230 30660
rect 28460 30648 28488 30679
rect 28626 30676 28632 30728
rect 28684 30716 28690 30728
rect 28736 30725 28764 30756
rect 29546 30744 29552 30756
rect 29604 30784 29610 30796
rect 29733 30787 29791 30793
rect 29733 30784 29745 30787
rect 29604 30756 29745 30784
rect 29604 30744 29610 30756
rect 29733 30753 29745 30756
rect 29779 30784 29791 30787
rect 30006 30784 30012 30796
rect 29779 30756 30012 30784
rect 29779 30753 29791 30756
rect 29733 30747 29791 30753
rect 30006 30744 30012 30756
rect 30064 30744 30070 30796
rect 30098 30744 30104 30796
rect 30156 30784 30162 30796
rect 30193 30787 30251 30793
rect 30193 30784 30205 30787
rect 30156 30756 30205 30784
rect 30156 30744 30162 30756
rect 30193 30753 30205 30756
rect 30239 30753 30251 30787
rect 30193 30747 30251 30753
rect 30285 30787 30343 30793
rect 30285 30753 30297 30787
rect 30331 30784 30343 30787
rect 30374 30784 30380 30796
rect 30331 30756 30380 30784
rect 30331 30753 30343 30756
rect 30285 30747 30343 30753
rect 30374 30744 30380 30756
rect 30432 30744 30438 30796
rect 31404 30784 31432 30824
rect 31478 30812 31484 30864
rect 31536 30852 31542 30864
rect 32306 30852 32312 30864
rect 31536 30824 32168 30852
rect 31536 30812 31542 30824
rect 31662 30784 31668 30796
rect 31404 30756 31668 30784
rect 31662 30744 31668 30756
rect 31720 30744 31726 30796
rect 28721 30719 28779 30725
rect 28721 30716 28733 30719
rect 28684 30688 28733 30716
rect 28684 30676 28690 30688
rect 28721 30685 28733 30688
rect 28767 30685 28779 30719
rect 28721 30679 28779 30685
rect 28810 30676 28816 30728
rect 28868 30716 28874 30728
rect 29822 30716 29828 30728
rect 28868 30688 29828 30716
rect 28868 30676 28874 30688
rect 29822 30676 29828 30688
rect 29880 30676 29886 30728
rect 31754 30676 31760 30728
rect 31812 30676 31818 30728
rect 31846 30676 31852 30728
rect 31904 30676 31910 30728
rect 32140 30725 32168 30824
rect 32232 30824 32312 30852
rect 32232 30793 32260 30824
rect 32306 30812 32312 30824
rect 32364 30812 32370 30864
rect 32858 30852 32864 30864
rect 32784 30824 32864 30852
rect 32217 30787 32275 30793
rect 32217 30753 32229 30787
rect 32263 30753 32275 30787
rect 32217 30747 32275 30753
rect 32125 30719 32183 30725
rect 32125 30685 32137 30719
rect 32171 30685 32183 30719
rect 32125 30679 32183 30685
rect 32306 30676 32312 30728
rect 32364 30716 32370 30728
rect 32784 30725 32812 30824
rect 32858 30812 32864 30824
rect 32916 30812 32922 30864
rect 33134 30812 33140 30864
rect 33192 30852 33198 30864
rect 36814 30852 36820 30864
rect 33192 30824 36820 30852
rect 33192 30812 33198 30824
rect 36814 30812 36820 30824
rect 36872 30812 36878 30864
rect 32950 30744 32956 30796
rect 33008 30784 33014 30796
rect 33008 30756 33410 30784
rect 33008 30744 33014 30756
rect 32769 30719 32827 30725
rect 32769 30716 32781 30719
rect 32364 30688 32781 30716
rect 32364 30676 32370 30688
rect 32769 30685 32781 30688
rect 32815 30685 32827 30719
rect 32769 30679 32827 30685
rect 32862 30719 32920 30725
rect 32862 30685 32874 30719
rect 32908 30716 32920 30719
rect 32908 30688 32996 30716
rect 32908 30685 32920 30688
rect 32862 30679 32920 30685
rect 30374 30648 30380 30660
rect 28460 30620 30380 30648
rect 28736 30592 28764 30620
rect 30374 30608 30380 30620
rect 30432 30608 30438 30660
rect 24026 30580 24032 30592
rect 23216 30552 24032 30580
rect 24026 30540 24032 30552
rect 24084 30540 24090 30592
rect 25774 30540 25780 30592
rect 25832 30580 25838 30592
rect 25869 30583 25927 30589
rect 25869 30580 25881 30583
rect 25832 30552 25881 30580
rect 25832 30540 25838 30552
rect 25869 30549 25881 30552
rect 25915 30580 25927 30583
rect 26326 30580 26332 30592
rect 25915 30552 26332 30580
rect 25915 30549 25927 30552
rect 25869 30543 25927 30549
rect 26326 30540 26332 30552
rect 26384 30540 26390 30592
rect 26878 30540 26884 30592
rect 26936 30580 26942 30592
rect 27614 30580 27620 30592
rect 26936 30552 27620 30580
rect 26936 30540 26942 30552
rect 27614 30540 27620 30552
rect 27672 30540 27678 30592
rect 27706 30540 27712 30592
rect 27764 30580 27770 30592
rect 28534 30580 28540 30592
rect 27764 30552 28540 30580
rect 27764 30540 27770 30552
rect 28534 30540 28540 30552
rect 28592 30540 28598 30592
rect 28718 30540 28724 30592
rect 28776 30540 28782 30592
rect 28902 30540 28908 30592
rect 28960 30540 28966 30592
rect 29822 30540 29828 30592
rect 29880 30580 29886 30592
rect 29917 30583 29975 30589
rect 29917 30580 29929 30583
rect 29880 30552 29929 30580
rect 29880 30540 29886 30552
rect 29917 30549 29929 30552
rect 29963 30580 29975 30583
rect 31386 30580 31392 30592
rect 29963 30552 31392 30580
rect 29963 30549 29975 30552
rect 29917 30543 29975 30549
rect 31386 30540 31392 30552
rect 31444 30540 31450 30592
rect 32582 30540 32588 30592
rect 32640 30580 32646 30592
rect 32968 30580 32996 30688
rect 33226 30676 33232 30728
rect 33284 30725 33290 30728
rect 33284 30716 33292 30725
rect 33382 30716 33410 30756
rect 33962 30744 33968 30796
rect 34020 30784 34026 30796
rect 34241 30787 34299 30793
rect 34241 30784 34253 30787
rect 34020 30756 34253 30784
rect 34020 30744 34026 30756
rect 34241 30753 34253 30756
rect 34287 30753 34299 30787
rect 34241 30747 34299 30753
rect 37090 30744 37096 30796
rect 37148 30744 37154 30796
rect 37366 30744 37372 30796
rect 37424 30784 37430 30796
rect 37553 30787 37611 30793
rect 37553 30784 37565 30787
rect 37424 30756 37565 30784
rect 37424 30744 37430 30756
rect 37553 30753 37565 30756
rect 37599 30753 37611 30787
rect 37553 30747 37611 30753
rect 38286 30744 38292 30796
rect 38344 30744 38350 30796
rect 34057 30719 34115 30725
rect 34057 30716 34069 30719
rect 33284 30688 33325 30716
rect 33382 30688 34069 30716
rect 33284 30679 33292 30688
rect 34057 30685 34069 30688
rect 34103 30685 34115 30719
rect 34057 30679 34115 30685
rect 34333 30719 34391 30725
rect 34333 30685 34345 30719
rect 34379 30685 34391 30719
rect 34333 30679 34391 30685
rect 33284 30676 33290 30679
rect 33045 30651 33103 30657
rect 33045 30617 33057 30651
rect 33091 30617 33103 30651
rect 33045 30611 33103 30617
rect 32640 30552 32996 30580
rect 33060 30580 33088 30611
rect 33134 30608 33140 30660
rect 33192 30608 33198 30660
rect 33778 30608 33784 30660
rect 33836 30648 33842 30660
rect 34348 30648 34376 30679
rect 34882 30676 34888 30728
rect 34940 30676 34946 30728
rect 35161 30719 35219 30725
rect 35161 30716 35173 30719
rect 34992 30688 35173 30716
rect 34992 30648 35020 30688
rect 35161 30685 35173 30688
rect 35207 30685 35219 30719
rect 35161 30679 35219 30685
rect 35253 30719 35311 30725
rect 35253 30685 35265 30719
rect 35299 30716 35311 30719
rect 35434 30716 35440 30728
rect 35299 30688 35440 30716
rect 35299 30685 35311 30688
rect 35253 30679 35311 30685
rect 35434 30676 35440 30688
rect 35492 30676 35498 30728
rect 35894 30676 35900 30728
rect 35952 30676 35958 30728
rect 36078 30725 36084 30728
rect 36045 30719 36084 30725
rect 36045 30685 36057 30719
rect 36045 30679 36084 30685
rect 36078 30676 36084 30679
rect 36136 30676 36142 30728
rect 36403 30719 36461 30725
rect 36403 30685 36415 30719
rect 36449 30716 36461 30719
rect 36538 30716 36544 30728
rect 36449 30688 36544 30716
rect 36449 30685 36461 30688
rect 36403 30679 36461 30685
rect 36538 30676 36544 30688
rect 36596 30676 36602 30728
rect 36630 30676 36636 30728
rect 36688 30716 36694 30728
rect 36814 30716 36820 30728
rect 36688 30688 36820 30716
rect 36688 30676 36694 30688
rect 36814 30676 36820 30688
rect 36872 30676 36878 30728
rect 37182 30676 37188 30728
rect 37240 30676 37246 30728
rect 38013 30719 38071 30725
rect 38013 30685 38025 30719
rect 38059 30716 38071 30719
rect 38378 30716 38384 30728
rect 38059 30688 38384 30716
rect 38059 30685 38071 30688
rect 38013 30679 38071 30685
rect 38378 30676 38384 30688
rect 38436 30676 38442 30728
rect 33836 30620 34376 30648
rect 34420 30620 35020 30648
rect 35069 30651 35127 30657
rect 33836 30608 33842 30620
rect 33318 30580 33324 30592
rect 33060 30552 33324 30580
rect 32640 30540 32646 30552
rect 33318 30540 33324 30552
rect 33376 30540 33382 30592
rect 33413 30583 33471 30589
rect 33413 30549 33425 30583
rect 33459 30580 33471 30583
rect 33502 30580 33508 30592
rect 33459 30552 33508 30580
rect 33459 30549 33471 30552
rect 33413 30543 33471 30549
rect 33502 30540 33508 30552
rect 33560 30540 33566 30592
rect 33594 30540 33600 30592
rect 33652 30580 33658 30592
rect 33873 30583 33931 30589
rect 33873 30580 33885 30583
rect 33652 30552 33885 30580
rect 33652 30540 33658 30552
rect 33873 30549 33885 30552
rect 33919 30549 33931 30583
rect 33873 30543 33931 30549
rect 34054 30540 34060 30592
rect 34112 30580 34118 30592
rect 34420 30580 34448 30620
rect 35069 30617 35081 30651
rect 35115 30648 35127 30651
rect 36170 30648 36176 30660
rect 35115 30620 36176 30648
rect 35115 30617 35127 30620
rect 35069 30611 35127 30617
rect 36170 30608 36176 30620
rect 36228 30608 36234 30660
rect 36262 30608 36268 30660
rect 36320 30648 36326 30660
rect 36320 30620 38056 30648
rect 36320 30608 36326 30620
rect 38028 30592 38056 30620
rect 34112 30552 34448 30580
rect 35437 30583 35495 30589
rect 34112 30540 34118 30552
rect 35437 30549 35449 30583
rect 35483 30580 35495 30583
rect 37642 30580 37648 30592
rect 35483 30552 37648 30580
rect 35483 30549 35495 30552
rect 35437 30543 35495 30549
rect 37642 30540 37648 30552
rect 37700 30540 37706 30592
rect 38010 30540 38016 30592
rect 38068 30540 38074 30592
rect 38286 30540 38292 30592
rect 38344 30540 38350 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 5994 30336 6000 30388
rect 6052 30376 6058 30388
rect 11330 30376 11336 30388
rect 6052 30348 11336 30376
rect 6052 30336 6058 30348
rect 11330 30336 11336 30348
rect 11388 30336 11394 30388
rect 13170 30376 13176 30388
rect 12544 30348 13176 30376
rect 8018 30308 8024 30320
rect 6748 30280 8024 30308
rect 6748 30249 6776 30280
rect 8018 30268 8024 30280
rect 8076 30268 8082 30320
rect 8478 30268 8484 30320
rect 8536 30308 8542 30320
rect 9122 30308 9128 30320
rect 8536 30280 9128 30308
rect 8536 30268 8542 30280
rect 9122 30268 9128 30280
rect 9180 30268 9186 30320
rect 9214 30268 9220 30320
rect 9272 30308 9278 30320
rect 10965 30311 11023 30317
rect 9272 30280 10916 30308
rect 9272 30268 9278 30280
rect 6733 30243 6791 30249
rect 6733 30209 6745 30243
rect 6779 30209 6791 30243
rect 6733 30203 6791 30209
rect 6917 30243 6975 30249
rect 6917 30209 6929 30243
rect 6963 30240 6975 30243
rect 7644 30243 7702 30249
rect 6963 30212 7328 30240
rect 6963 30209 6975 30212
rect 6917 30203 6975 30209
rect 6638 29996 6644 30048
rect 6696 30036 6702 30048
rect 6733 30039 6791 30045
rect 6733 30036 6745 30039
rect 6696 30008 6745 30036
rect 6696 29996 6702 30008
rect 6733 30005 6745 30008
rect 6779 30005 6791 30039
rect 7300 30036 7328 30212
rect 7644 30209 7656 30243
rect 7690 30240 7702 30243
rect 8110 30240 8116 30252
rect 7690 30212 8116 30240
rect 7690 30209 7702 30212
rect 7644 30203 7702 30209
rect 8110 30200 8116 30212
rect 8168 30200 8174 30252
rect 8938 30200 8944 30252
rect 8996 30240 9002 30252
rect 9677 30243 9735 30249
rect 9677 30240 9689 30243
rect 8996 30212 9689 30240
rect 8996 30200 9002 30212
rect 9677 30209 9689 30212
rect 9723 30209 9735 30243
rect 9677 30203 9735 30209
rect 9766 30200 9772 30252
rect 9824 30200 9830 30252
rect 9968 30249 9996 30280
rect 9953 30243 10011 30249
rect 9953 30209 9965 30243
rect 9999 30209 10011 30243
rect 9953 30203 10011 30209
rect 10137 30243 10195 30249
rect 10137 30209 10149 30243
rect 10183 30240 10195 30243
rect 10888 30240 10916 30280
rect 10965 30277 10977 30311
rect 11011 30308 11023 30311
rect 11146 30308 11152 30320
rect 11011 30280 11152 30308
rect 11011 30277 11023 30280
rect 10965 30271 11023 30277
rect 11146 30268 11152 30280
rect 11204 30268 11210 30320
rect 11238 30268 11244 30320
rect 11296 30308 11302 30320
rect 11793 30311 11851 30317
rect 11296 30280 11744 30308
rect 11296 30268 11302 30280
rect 11716 30252 11744 30280
rect 11793 30277 11805 30311
rect 11839 30308 11851 30311
rect 12544 30308 12572 30348
rect 13170 30336 13176 30348
rect 13228 30336 13234 30388
rect 15102 30376 15108 30388
rect 13572 30348 15108 30376
rect 11839 30280 12572 30308
rect 11839 30277 11851 30280
rect 11793 30271 11851 30277
rect 12894 30268 12900 30320
rect 12952 30308 12958 30320
rect 13357 30311 13415 30317
rect 13357 30308 13369 30311
rect 12952 30280 13369 30308
rect 12952 30268 12958 30280
rect 13357 30277 13369 30280
rect 13403 30277 13415 30311
rect 13357 30271 13415 30277
rect 11514 30240 11520 30252
rect 10183 30212 10824 30240
rect 10888 30212 11520 30240
rect 10183 30209 10195 30212
rect 10137 30203 10195 30209
rect 7374 30132 7380 30184
rect 7432 30132 7438 30184
rect 8570 30132 8576 30184
rect 8628 30172 8634 30184
rect 9784 30172 9812 30200
rect 8628 30144 9812 30172
rect 8628 30132 8634 30144
rect 10152 30104 10180 30203
rect 10597 30175 10655 30181
rect 10597 30172 10609 30175
rect 8303 30076 10180 30104
rect 10428 30144 10609 30172
rect 7742 30036 7748 30048
rect 7300 30008 7748 30036
rect 6733 29999 6791 30005
rect 7742 29996 7748 30008
rect 7800 29996 7806 30048
rect 8018 29996 8024 30048
rect 8076 30036 8082 30048
rect 8303 30036 8331 30076
rect 8076 30008 8331 30036
rect 8076 29996 8082 30008
rect 8754 29996 8760 30048
rect 8812 29996 8818 30048
rect 9122 29996 9128 30048
rect 9180 30036 9186 30048
rect 9401 30039 9459 30045
rect 9401 30036 9413 30039
rect 9180 30008 9413 30036
rect 9180 29996 9186 30008
rect 9401 30005 9413 30008
rect 9447 30005 9459 30039
rect 9401 29999 9459 30005
rect 9490 29996 9496 30048
rect 9548 30036 9554 30048
rect 9674 30036 9680 30048
rect 9548 30008 9680 30036
rect 9548 29996 9554 30008
rect 9674 29996 9680 30008
rect 9732 29996 9738 30048
rect 9861 30039 9919 30045
rect 9861 30005 9873 30039
rect 9907 30036 9919 30039
rect 10428 30036 10456 30144
rect 10597 30141 10609 30144
rect 10643 30141 10655 30175
rect 10796 30172 10824 30212
rect 11514 30200 11520 30212
rect 11572 30200 11578 30252
rect 11698 30200 11704 30252
rect 11756 30200 11762 30252
rect 11885 30243 11943 30249
rect 11885 30209 11897 30243
rect 11931 30240 11943 30243
rect 12434 30240 12440 30252
rect 11931 30212 12440 30240
rect 11931 30209 11943 30212
rect 11885 30203 11943 30209
rect 12434 30200 12440 30212
rect 12492 30200 12498 30252
rect 13572 30240 13600 30348
rect 15102 30336 15108 30348
rect 15160 30336 15166 30388
rect 20162 30336 20168 30388
rect 20220 30376 20226 30388
rect 21174 30376 21180 30388
rect 20220 30348 21180 30376
rect 20220 30336 20226 30348
rect 21174 30336 21180 30348
rect 21232 30336 21238 30388
rect 22097 30379 22155 30385
rect 22097 30345 22109 30379
rect 22143 30345 22155 30379
rect 22097 30339 22155 30345
rect 14369 30311 14427 30317
rect 14369 30277 14381 30311
rect 14415 30308 14427 30311
rect 17129 30311 17187 30317
rect 14415 30280 16988 30308
rect 14415 30277 14427 30280
rect 14369 30271 14427 30277
rect 12728 30212 13600 30240
rect 12728 30184 12756 30212
rect 13630 30200 13636 30252
rect 13688 30200 13694 30252
rect 14277 30243 14335 30249
rect 14277 30209 14289 30243
rect 14323 30240 14335 30243
rect 14826 30240 14832 30252
rect 14323 30212 14832 30240
rect 14323 30209 14335 30212
rect 14277 30203 14335 30209
rect 14826 30200 14832 30212
rect 14884 30200 14890 30252
rect 14921 30243 14979 30249
rect 14921 30209 14933 30243
rect 14967 30240 14979 30243
rect 15010 30240 15016 30252
rect 14967 30212 15016 30240
rect 14967 30209 14979 30212
rect 14921 30203 14979 30209
rect 15010 30200 15016 30212
rect 15068 30200 15074 30252
rect 15188 30243 15246 30249
rect 15188 30209 15200 30243
rect 15234 30240 15246 30243
rect 16206 30240 16212 30252
rect 15234 30212 16212 30240
rect 15234 30209 15246 30212
rect 15188 30203 15246 30209
rect 16206 30200 16212 30212
rect 16264 30200 16270 30252
rect 16390 30200 16396 30252
rect 16448 30240 16454 30252
rect 16853 30243 16911 30249
rect 16853 30240 16865 30243
rect 16448 30212 16865 30240
rect 16448 30200 16454 30212
rect 16853 30209 16865 30212
rect 16899 30209 16911 30243
rect 16853 30203 16911 30209
rect 11790 30172 11796 30184
rect 10796 30144 11796 30172
rect 10597 30135 10655 30141
rect 11790 30132 11796 30144
rect 11848 30132 11854 30184
rect 12529 30175 12587 30181
rect 12529 30141 12541 30175
rect 12575 30141 12587 30175
rect 12529 30135 12587 30141
rect 10502 30064 10508 30116
rect 10560 30104 10566 30116
rect 12544 30104 12572 30135
rect 12618 30132 12624 30184
rect 12676 30132 12682 30184
rect 12710 30132 12716 30184
rect 12768 30132 12774 30184
rect 12802 30132 12808 30184
rect 12860 30132 12866 30184
rect 13541 30175 13599 30181
rect 13541 30141 13553 30175
rect 13587 30172 13599 30175
rect 13722 30172 13728 30184
rect 13587 30144 13728 30172
rect 13587 30141 13599 30144
rect 13541 30135 13599 30141
rect 13722 30132 13728 30144
rect 13780 30132 13786 30184
rect 16960 30172 16988 30280
rect 17129 30277 17141 30311
rect 17175 30308 17187 30311
rect 17586 30308 17592 30320
rect 17175 30280 17592 30308
rect 17175 30277 17187 30280
rect 17129 30271 17187 30277
rect 17586 30268 17592 30280
rect 17644 30268 17650 30320
rect 20622 30268 20628 30320
rect 20680 30308 20686 30320
rect 20680 30280 21404 30308
rect 20680 30268 20686 30280
rect 17034 30200 17040 30252
rect 17092 30200 17098 30252
rect 17218 30200 17224 30252
rect 17276 30200 17282 30252
rect 17310 30200 17316 30252
rect 17368 30240 17374 30252
rect 18141 30243 18199 30249
rect 18141 30240 18153 30243
rect 17368 30212 18153 30240
rect 17368 30200 17374 30212
rect 18141 30209 18153 30212
rect 18187 30240 18199 30243
rect 19334 30240 19340 30252
rect 18187 30212 19340 30240
rect 18187 30209 18199 30212
rect 18141 30203 18199 30209
rect 19334 30200 19340 30212
rect 19392 30200 19398 30252
rect 20257 30243 20315 30249
rect 20257 30209 20269 30243
rect 20303 30240 20315 30243
rect 20303 30212 20852 30240
rect 20303 30209 20315 30212
rect 20257 30203 20315 30209
rect 18322 30172 18328 30184
rect 16960 30144 18328 30172
rect 18322 30132 18328 30144
rect 18380 30132 18386 30184
rect 18414 30132 18420 30184
rect 18472 30132 18478 30184
rect 20824 30172 20852 30212
rect 20898 30200 20904 30252
rect 20956 30200 20962 30252
rect 20993 30243 21051 30249
rect 20993 30209 21005 30243
rect 21039 30240 21051 30243
rect 21082 30240 21088 30252
rect 21039 30212 21088 30240
rect 21039 30209 21051 30212
rect 20993 30203 21051 30209
rect 21082 30200 21088 30212
rect 21140 30200 21146 30252
rect 21266 30200 21272 30252
rect 21324 30200 21330 30252
rect 21376 30249 21404 30280
rect 21450 30268 21456 30320
rect 21508 30308 21514 30320
rect 22112 30308 22140 30339
rect 23750 30336 23756 30388
rect 23808 30376 23814 30388
rect 26234 30376 26240 30388
rect 23808 30348 26240 30376
rect 23808 30336 23814 30348
rect 26234 30336 26240 30348
rect 26292 30376 26298 30388
rect 26292 30348 26924 30376
rect 26292 30336 26298 30348
rect 22186 30308 22192 30320
rect 21508 30280 22192 30308
rect 21508 30268 21514 30280
rect 22186 30268 22192 30280
rect 22244 30268 22250 30320
rect 22554 30268 22560 30320
rect 22612 30308 22618 30320
rect 23106 30308 23112 30320
rect 22612 30280 23112 30308
rect 22612 30268 22618 30280
rect 23106 30268 23112 30280
rect 23164 30308 23170 30320
rect 23164 30280 23244 30308
rect 23164 30268 23170 30280
rect 21361 30243 21419 30249
rect 21361 30209 21373 30243
rect 21407 30209 21419 30243
rect 21361 30203 21419 30209
rect 21174 30172 21180 30184
rect 20824 30144 21180 30172
rect 21174 30132 21180 30144
rect 21232 30132 21238 30184
rect 21376 30172 21404 30203
rect 22002 30200 22008 30252
rect 22060 30240 22066 30252
rect 22060 30212 22232 30240
rect 22060 30200 22066 30212
rect 22204 30172 22232 30212
rect 22278 30200 22284 30252
rect 22336 30200 22342 30252
rect 22462 30200 22468 30252
rect 22520 30200 22526 30252
rect 23216 30249 23244 30280
rect 24578 30268 24584 30320
rect 24636 30268 24642 30320
rect 25038 30268 25044 30320
rect 25096 30308 25102 30320
rect 25133 30311 25191 30317
rect 25133 30308 25145 30311
rect 25096 30280 25145 30308
rect 25096 30268 25102 30280
rect 25133 30277 25145 30280
rect 25179 30308 25191 30311
rect 25590 30308 25596 30320
rect 25179 30280 25596 30308
rect 25179 30277 25191 30280
rect 25133 30271 25191 30277
rect 25590 30268 25596 30280
rect 25648 30268 25654 30320
rect 26050 30268 26056 30320
rect 26108 30308 26114 30320
rect 26786 30308 26792 30320
rect 26108 30280 26792 30308
rect 26108 30268 26114 30280
rect 26786 30268 26792 30280
rect 26844 30268 26850 30320
rect 23017 30243 23075 30249
rect 23017 30209 23029 30243
rect 23063 30209 23075 30243
rect 23017 30203 23075 30209
rect 23201 30243 23259 30249
rect 23201 30209 23213 30243
rect 23247 30209 23259 30243
rect 23201 30203 23259 30209
rect 23032 30172 23060 30203
rect 23474 30200 23480 30252
rect 23532 30240 23538 30252
rect 23937 30243 23995 30249
rect 23937 30240 23949 30243
rect 23532 30212 23949 30240
rect 23532 30200 23538 30212
rect 23937 30209 23949 30212
rect 23983 30209 23995 30243
rect 23937 30203 23995 30209
rect 24486 30200 24492 30252
rect 24544 30240 24550 30252
rect 24765 30243 24823 30249
rect 24765 30240 24777 30243
rect 24544 30212 24777 30240
rect 24544 30200 24550 30212
rect 24765 30209 24777 30212
rect 24811 30209 24823 30243
rect 24765 30203 24823 30209
rect 24854 30200 24860 30252
rect 24912 30240 24918 30252
rect 26896 30240 26924 30348
rect 27338 30336 27344 30388
rect 27396 30376 27402 30388
rect 29822 30376 29828 30388
rect 27396 30348 29828 30376
rect 27396 30336 27402 30348
rect 29822 30336 29828 30348
rect 29880 30336 29886 30388
rect 30098 30336 30104 30388
rect 30156 30336 30162 30388
rect 30190 30336 30196 30388
rect 30248 30376 30254 30388
rect 34149 30379 34207 30385
rect 34149 30376 34161 30379
rect 30248 30348 34161 30376
rect 30248 30336 30254 30348
rect 34149 30345 34161 30348
rect 34195 30376 34207 30379
rect 34606 30376 34612 30388
rect 34195 30348 34612 30376
rect 34195 30345 34207 30348
rect 34149 30339 34207 30345
rect 34606 30336 34612 30348
rect 34664 30336 34670 30388
rect 36078 30336 36084 30388
rect 36136 30376 36142 30388
rect 37829 30379 37887 30385
rect 37829 30376 37841 30379
rect 36136 30348 37841 30376
rect 36136 30336 36142 30348
rect 37829 30345 37841 30348
rect 37875 30376 37887 30379
rect 38194 30376 38200 30388
rect 37875 30348 38200 30376
rect 37875 30345 37887 30348
rect 37829 30339 37887 30345
rect 38194 30336 38200 30348
rect 38252 30336 38258 30388
rect 27062 30268 27068 30320
rect 27120 30308 27126 30320
rect 27706 30308 27712 30320
rect 27120 30280 27712 30308
rect 27120 30268 27126 30280
rect 27706 30268 27712 30280
rect 27764 30268 27770 30320
rect 30116 30308 30144 30336
rect 28552 30280 30144 30308
rect 31205 30311 31263 30317
rect 27433 30243 27491 30249
rect 27433 30240 27445 30243
rect 24912 30212 26096 30240
rect 26896 30212 27445 30240
rect 24912 30200 24918 30212
rect 23566 30172 23572 30184
rect 21376 30144 22140 30172
rect 22204 30144 23572 30172
rect 10560 30076 12572 30104
rect 10560 30064 10566 30076
rect 16482 30064 16488 30116
rect 16540 30104 16546 30116
rect 17405 30107 17463 30113
rect 17405 30104 17417 30107
rect 16540 30076 17417 30104
rect 16540 30064 16546 30076
rect 17405 30073 17417 30076
rect 17451 30073 17463 30107
rect 22002 30104 22008 30116
rect 17405 30067 17463 30073
rect 19076 30076 22008 30104
rect 10870 30036 10876 30048
rect 9907 30008 10876 30036
rect 9907 30005 9919 30008
rect 9861 29999 9919 30005
rect 10870 29996 10876 30008
rect 10928 29996 10934 30048
rect 10962 29996 10968 30048
rect 11020 29996 11026 30048
rect 11149 30039 11207 30045
rect 11149 30005 11161 30039
rect 11195 30036 11207 30039
rect 11238 30036 11244 30048
rect 11195 30008 11244 30036
rect 11195 30005 11207 30008
rect 11149 29999 11207 30005
rect 11238 29996 11244 30008
rect 11296 29996 11302 30048
rect 12342 29996 12348 30048
rect 12400 29996 12406 30048
rect 13078 29996 13084 30048
rect 13136 30036 13142 30048
rect 13357 30039 13415 30045
rect 13357 30036 13369 30039
rect 13136 30008 13369 30036
rect 13136 29996 13142 30008
rect 13357 30005 13369 30008
rect 13403 30005 13415 30039
rect 13357 29999 13415 30005
rect 13814 29996 13820 30048
rect 13872 29996 13878 30048
rect 15930 29996 15936 30048
rect 15988 30036 15994 30048
rect 16301 30039 16359 30045
rect 16301 30036 16313 30039
rect 15988 30008 16313 30036
rect 15988 29996 15994 30008
rect 16301 30005 16313 30008
rect 16347 30036 16359 30039
rect 19076 30036 19104 30076
rect 22002 30064 22008 30076
rect 22060 30064 22066 30116
rect 22112 30104 22140 30144
rect 23566 30132 23572 30144
rect 23624 30132 23630 30184
rect 25590 30132 25596 30184
rect 25648 30132 25654 30184
rect 26068 30181 26096 30212
rect 27433 30209 27445 30212
rect 27479 30209 27491 30243
rect 27433 30203 27491 30209
rect 27525 30243 27583 30249
rect 27525 30209 27537 30243
rect 27571 30240 27583 30243
rect 28442 30240 28448 30252
rect 27571 30212 28448 30240
rect 27571 30209 27583 30212
rect 27525 30203 27583 30209
rect 28442 30200 28448 30212
rect 28500 30200 28506 30252
rect 26053 30175 26111 30181
rect 26053 30141 26065 30175
rect 26099 30141 26111 30175
rect 27338 30172 27344 30184
rect 26053 30135 26111 30141
rect 26140 30144 27344 30172
rect 22554 30104 22560 30116
rect 22112 30076 22560 30104
rect 22554 30064 22560 30076
rect 22612 30064 22618 30116
rect 23106 30064 23112 30116
rect 23164 30104 23170 30116
rect 25222 30104 25228 30116
rect 23164 30076 25228 30104
rect 23164 30064 23170 30076
rect 25222 30064 25228 30076
rect 25280 30064 25286 30116
rect 25314 30064 25320 30116
rect 25372 30104 25378 30116
rect 25866 30104 25872 30116
rect 25372 30076 25872 30104
rect 25372 30064 25378 30076
rect 25866 30064 25872 30076
rect 25924 30064 25930 30116
rect 16347 30008 19104 30036
rect 16347 30005 16359 30008
rect 16301 29999 16359 30005
rect 19702 29996 19708 30048
rect 19760 29996 19766 30048
rect 21082 29996 21088 30048
rect 21140 30036 21146 30048
rect 21450 30036 21456 30048
rect 21140 30008 21456 30036
rect 21140 29996 21146 30008
rect 21450 29996 21456 30008
rect 21508 29996 21514 30048
rect 22462 29996 22468 30048
rect 22520 30036 22526 30048
rect 24029 30039 24087 30045
rect 24029 30036 24041 30039
rect 22520 30008 24041 30036
rect 22520 29996 22526 30008
rect 24029 30005 24041 30008
rect 24075 30005 24087 30039
rect 24029 29999 24087 30005
rect 24578 29996 24584 30048
rect 24636 30036 24642 30048
rect 25406 30036 25412 30048
rect 24636 30008 25412 30036
rect 24636 29996 24642 30008
rect 25406 29996 25412 30008
rect 25464 30036 25470 30048
rect 26140 30036 26168 30144
rect 27338 30132 27344 30144
rect 27396 30132 27402 30184
rect 27617 30175 27675 30181
rect 27617 30141 27629 30175
rect 27663 30172 27675 30175
rect 27706 30172 27712 30184
rect 27663 30144 27712 30172
rect 27663 30141 27675 30144
rect 27617 30135 27675 30141
rect 27706 30132 27712 30144
rect 27764 30172 27770 30184
rect 28074 30172 28080 30184
rect 27764 30144 28080 30172
rect 27764 30132 27770 30144
rect 28074 30132 28080 30144
rect 28132 30132 28138 30184
rect 28166 30132 28172 30184
rect 28224 30132 28230 30184
rect 26326 30064 26332 30116
rect 26384 30104 26390 30116
rect 27798 30104 27804 30116
rect 26384 30076 27804 30104
rect 26384 30064 26390 30076
rect 27356 30048 27384 30076
rect 27798 30064 27804 30076
rect 27856 30064 27862 30116
rect 28552 30113 28580 30280
rect 31205 30277 31217 30311
rect 31251 30308 31263 30311
rect 31251 30280 31616 30308
rect 31251 30277 31263 30280
rect 31205 30271 31263 30277
rect 29733 30243 29791 30249
rect 29733 30240 29745 30243
rect 28736 30212 29745 30240
rect 28736 30181 28764 30212
rect 29733 30209 29745 30212
rect 29779 30240 29791 30243
rect 30282 30240 30288 30252
rect 29779 30238 30052 30240
rect 30208 30238 30288 30240
rect 29779 30212 30288 30238
rect 29779 30209 29791 30212
rect 30024 30210 30236 30212
rect 29733 30203 29791 30209
rect 30282 30200 30288 30212
rect 30340 30200 30346 30252
rect 31481 30243 31539 30249
rect 31481 30240 31493 30243
rect 31312 30212 31493 30240
rect 28721 30175 28779 30181
rect 28721 30141 28733 30175
rect 28767 30141 28779 30175
rect 28721 30135 28779 30141
rect 28537 30107 28595 30113
rect 28537 30073 28549 30107
rect 28583 30073 28595 30107
rect 28537 30067 28595 30073
rect 28626 30064 28632 30116
rect 28684 30064 28690 30116
rect 25464 30008 26168 30036
rect 25464 29996 25470 30008
rect 27154 29996 27160 30048
rect 27212 29996 27218 30048
rect 27338 29996 27344 30048
rect 27396 29996 27402 30048
rect 27430 29996 27436 30048
rect 27488 30036 27494 30048
rect 28736 30036 28764 30135
rect 29086 30132 29092 30184
rect 29144 30132 29150 30184
rect 29546 30132 29552 30184
rect 29604 30172 29610 30184
rect 29641 30175 29699 30181
rect 29641 30172 29653 30175
rect 29604 30144 29653 30172
rect 29604 30132 29610 30144
rect 29641 30141 29653 30144
rect 29687 30141 29699 30175
rect 29641 30135 29699 30141
rect 29822 30132 29828 30184
rect 29880 30172 29886 30184
rect 30193 30175 30251 30181
rect 30193 30172 30205 30175
rect 29880 30144 30205 30172
rect 29880 30132 29886 30144
rect 30193 30141 30205 30144
rect 30239 30141 30251 30175
rect 30193 30135 30251 30141
rect 30098 30064 30104 30116
rect 30156 30064 30162 30116
rect 31312 30104 31340 30212
rect 31481 30209 31493 30212
rect 31527 30209 31539 30243
rect 31588 30240 31616 30280
rect 31662 30268 31668 30320
rect 31720 30308 31726 30320
rect 32309 30311 32367 30317
rect 32309 30308 32321 30311
rect 31720 30280 32321 30308
rect 31720 30268 31726 30280
rect 32309 30277 32321 30280
rect 32355 30277 32367 30311
rect 32309 30271 32367 30277
rect 33781 30311 33839 30317
rect 33781 30277 33793 30311
rect 33827 30308 33839 30311
rect 34238 30308 34244 30320
rect 33827 30280 34244 30308
rect 33827 30277 33839 30280
rect 33781 30271 33839 30277
rect 34238 30268 34244 30280
rect 34296 30268 34302 30320
rect 36722 30308 36728 30320
rect 35084 30280 36728 30308
rect 33226 30240 33232 30252
rect 31588 30212 33232 30240
rect 31481 30203 31539 30209
rect 33226 30200 33232 30212
rect 33284 30200 33290 30252
rect 33502 30200 33508 30252
rect 33560 30200 33566 30252
rect 33653 30243 33711 30249
rect 33653 30209 33665 30243
rect 33699 30209 33711 30243
rect 33653 30203 33711 30209
rect 31389 30175 31447 30181
rect 31389 30141 31401 30175
rect 31435 30172 31447 30175
rect 31754 30172 31760 30184
rect 31435 30144 31760 30172
rect 31435 30141 31447 30144
rect 31389 30135 31447 30141
rect 31754 30132 31760 30144
rect 31812 30132 31818 30184
rect 31938 30132 31944 30184
rect 31996 30172 32002 30184
rect 32677 30175 32735 30181
rect 32677 30172 32689 30175
rect 31996 30144 32689 30172
rect 31996 30132 32002 30144
rect 32677 30141 32689 30144
rect 32723 30141 32735 30175
rect 32677 30135 32735 30141
rect 32950 30132 32956 30184
rect 33008 30172 33014 30184
rect 33668 30172 33696 30203
rect 33870 30200 33876 30252
rect 33928 30200 33934 30252
rect 34011 30243 34069 30249
rect 34011 30209 34023 30243
rect 34057 30240 34069 30243
rect 34146 30240 34152 30252
rect 34057 30212 34152 30240
rect 34057 30209 34069 30212
rect 34011 30203 34069 30209
rect 34146 30200 34152 30212
rect 34204 30240 34210 30252
rect 34422 30240 34428 30252
rect 34204 30212 34428 30240
rect 34204 30200 34210 30212
rect 34422 30200 34428 30212
rect 34480 30200 34486 30252
rect 35084 30249 35112 30280
rect 36722 30268 36728 30280
rect 36780 30268 36786 30320
rect 37550 30268 37556 30320
rect 37608 30308 37614 30320
rect 37921 30311 37979 30317
rect 37921 30308 37933 30311
rect 37608 30280 37933 30308
rect 37608 30268 37614 30280
rect 37921 30277 37933 30280
rect 37967 30277 37979 30311
rect 37921 30271 37979 30277
rect 35342 30249 35348 30252
rect 35069 30243 35127 30249
rect 35069 30209 35081 30243
rect 35115 30209 35127 30243
rect 35336 30240 35348 30249
rect 35303 30212 35348 30240
rect 35069 30203 35127 30209
rect 35336 30203 35348 30212
rect 35342 30200 35348 30203
rect 35400 30200 35406 30252
rect 33008 30144 33640 30172
rect 33668 30144 34013 30172
rect 33008 30132 33014 30144
rect 32306 30104 32312 30116
rect 30208 30076 32312 30104
rect 30208 30048 30236 30076
rect 32306 30064 32312 30076
rect 32364 30064 32370 30116
rect 32585 30107 32643 30113
rect 32585 30073 32597 30107
rect 32631 30104 32643 30107
rect 33502 30104 33508 30116
rect 32631 30076 33508 30104
rect 32631 30073 32643 30076
rect 32585 30067 32643 30073
rect 33502 30064 33508 30076
rect 33560 30064 33566 30116
rect 33612 30104 33640 30144
rect 33686 30104 33692 30116
rect 33612 30076 33692 30104
rect 33686 30064 33692 30076
rect 33744 30064 33750 30116
rect 33985 30104 34013 30144
rect 38102 30132 38108 30184
rect 38160 30132 38166 30184
rect 33985 30076 35112 30104
rect 27488 30008 28764 30036
rect 27488 29996 27494 30008
rect 30190 29996 30196 30048
rect 30248 29996 30254 30048
rect 30469 30039 30527 30045
rect 30469 30005 30481 30039
rect 30515 30036 30527 30039
rect 30650 30036 30656 30048
rect 30515 30008 30656 30036
rect 30515 30005 30527 30008
rect 30469 29999 30527 30005
rect 30650 29996 30656 30008
rect 30708 29996 30714 30048
rect 31202 29996 31208 30048
rect 31260 29996 31266 30048
rect 31662 29996 31668 30048
rect 31720 29996 31726 30048
rect 32122 29996 32128 30048
rect 32180 30036 32186 30048
rect 32447 30039 32505 30045
rect 32447 30036 32459 30039
rect 32180 30008 32459 30036
rect 32180 29996 32186 30008
rect 32447 30005 32459 30008
rect 32493 30005 32505 30039
rect 32447 29999 32505 30005
rect 32769 30039 32827 30045
rect 32769 30005 32781 30039
rect 32815 30036 32827 30039
rect 32858 30036 32864 30048
rect 32815 30008 32864 30036
rect 32815 30005 32827 30008
rect 32769 29999 32827 30005
rect 32858 29996 32864 30008
rect 32916 29996 32922 30048
rect 33134 29996 33140 30048
rect 33192 30036 33198 30048
rect 34882 30036 34888 30048
rect 33192 30008 34888 30036
rect 33192 29996 33198 30008
rect 34882 29996 34888 30008
rect 34940 29996 34946 30048
rect 35084 30036 35112 30076
rect 35802 30036 35808 30048
rect 35084 30008 35808 30036
rect 35802 29996 35808 30008
rect 35860 30036 35866 30048
rect 36354 30036 36360 30048
rect 35860 30008 36360 30036
rect 35860 29996 35866 30008
rect 36354 29996 36360 30008
rect 36412 30036 36418 30048
rect 36449 30039 36507 30045
rect 36449 30036 36461 30039
rect 36412 30008 36461 30036
rect 36412 29996 36418 30008
rect 36449 30005 36461 30008
rect 36495 30005 36507 30039
rect 36449 29999 36507 30005
rect 37458 29996 37464 30048
rect 37516 29996 37522 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 3970 29792 3976 29844
rect 4028 29832 4034 29844
rect 4522 29832 4528 29844
rect 4028 29804 4528 29832
rect 4028 29792 4034 29804
rect 4522 29792 4528 29804
rect 4580 29792 4586 29844
rect 8110 29792 8116 29844
rect 8168 29792 8174 29844
rect 8202 29792 8208 29844
rect 8260 29832 8266 29844
rect 10321 29835 10379 29841
rect 10321 29832 10333 29835
rect 8260 29804 10333 29832
rect 8260 29792 8266 29804
rect 10321 29801 10333 29804
rect 10367 29801 10379 29835
rect 10321 29795 10379 29801
rect 10410 29792 10416 29844
rect 10468 29832 10474 29844
rect 11425 29835 11483 29841
rect 11425 29832 11437 29835
rect 10468 29804 11437 29832
rect 10468 29792 10474 29804
rect 11425 29801 11437 29804
rect 11471 29801 11483 29835
rect 12710 29832 12716 29844
rect 11425 29795 11483 29801
rect 11548 29804 12716 29832
rect 6825 29767 6883 29773
rect 6825 29733 6837 29767
rect 6871 29764 6883 29767
rect 9398 29764 9404 29776
rect 6871 29736 9404 29764
rect 6871 29733 6883 29736
rect 6825 29727 6883 29733
rect 9398 29724 9404 29736
rect 9456 29724 9462 29776
rect 9490 29724 9496 29776
rect 9548 29764 9554 29776
rect 10873 29767 10931 29773
rect 10873 29764 10885 29767
rect 9548 29736 10885 29764
rect 9548 29724 9554 29736
rect 10873 29733 10885 29736
rect 10919 29733 10931 29767
rect 10873 29727 10931 29733
rect 11146 29724 11152 29776
rect 11204 29764 11210 29776
rect 11548 29764 11576 29804
rect 12710 29792 12716 29804
rect 12768 29792 12774 29844
rect 13262 29792 13268 29844
rect 13320 29832 13326 29844
rect 13541 29835 13599 29841
rect 13541 29832 13553 29835
rect 13320 29804 13553 29832
rect 13320 29792 13326 29804
rect 13541 29801 13553 29804
rect 13587 29801 13599 29835
rect 16022 29832 16028 29844
rect 13541 29795 13599 29801
rect 13648 29804 16028 29832
rect 11974 29764 11980 29776
rect 11204 29736 11576 29764
rect 11624 29736 11980 29764
rect 11204 29724 11210 29736
rect 7190 29696 7196 29708
rect 6840 29668 7196 29696
rect 6840 29637 6868 29668
rect 7190 29656 7196 29668
rect 7248 29656 7254 29708
rect 7558 29696 7564 29708
rect 7392 29668 7564 29696
rect 6825 29631 6883 29637
rect 6825 29597 6837 29631
rect 6871 29597 6883 29631
rect 6825 29591 6883 29597
rect 7006 29588 7012 29640
rect 7064 29588 7070 29640
rect 7098 29588 7104 29640
rect 7156 29628 7162 29640
rect 7392 29628 7420 29668
rect 7558 29656 7564 29668
rect 7616 29696 7622 29708
rect 8573 29699 8631 29705
rect 7616 29668 7696 29696
rect 7616 29656 7622 29668
rect 7668 29637 7696 29668
rect 8573 29665 8585 29699
rect 8619 29696 8631 29699
rect 8754 29696 8760 29708
rect 8619 29668 8760 29696
rect 8619 29665 8631 29668
rect 8573 29659 8631 29665
rect 8754 29656 8760 29668
rect 8812 29656 8818 29708
rect 9122 29656 9128 29708
rect 9180 29656 9186 29708
rect 9582 29656 9588 29708
rect 9640 29696 9646 29708
rect 10502 29696 10508 29708
rect 9640 29668 10508 29696
rect 9640 29656 9646 29668
rect 10502 29656 10508 29668
rect 10560 29656 10566 29708
rect 11624 29705 11652 29736
rect 11974 29724 11980 29736
rect 12032 29724 12038 29776
rect 12434 29724 12440 29776
rect 12492 29764 12498 29776
rect 13648 29764 13676 29804
rect 16022 29792 16028 29804
rect 16080 29792 16086 29844
rect 16206 29792 16212 29844
rect 16264 29792 16270 29844
rect 16482 29792 16488 29844
rect 16540 29832 16546 29844
rect 16540 29804 21220 29832
rect 16540 29792 16546 29804
rect 12492 29736 13676 29764
rect 13725 29767 13783 29773
rect 12492 29724 12498 29736
rect 13725 29733 13737 29767
rect 13771 29764 13783 29767
rect 15378 29764 15384 29776
rect 13771 29736 15384 29764
rect 13771 29733 13783 29736
rect 13725 29727 13783 29733
rect 15378 29724 15384 29736
rect 15436 29764 15442 29776
rect 17034 29764 17040 29776
rect 15436 29736 17040 29764
rect 15436 29724 15442 29736
rect 17034 29724 17040 29736
rect 17092 29724 17098 29776
rect 18598 29724 18604 29776
rect 18656 29764 18662 29776
rect 19702 29764 19708 29776
rect 18656 29736 19708 29764
rect 18656 29724 18662 29736
rect 19702 29724 19708 29736
rect 19760 29764 19766 29776
rect 20898 29764 20904 29776
rect 19760 29736 20904 29764
rect 19760 29724 19766 29736
rect 20898 29724 20904 29736
rect 20956 29724 20962 29776
rect 11609 29699 11667 29705
rect 11609 29665 11621 29699
rect 11655 29665 11667 29699
rect 11609 29659 11667 29665
rect 11701 29699 11759 29705
rect 11701 29665 11713 29699
rect 11747 29696 11759 29699
rect 12805 29699 12863 29705
rect 12805 29696 12817 29699
rect 11747 29668 12817 29696
rect 11747 29665 11759 29668
rect 11701 29659 11759 29665
rect 12805 29665 12817 29668
rect 12851 29665 12863 29699
rect 12805 29659 12863 29665
rect 13630 29656 13636 29708
rect 13688 29696 13694 29708
rect 13688 29668 16528 29696
rect 13688 29656 13694 29668
rect 7156 29600 7420 29628
rect 7469 29631 7527 29637
rect 7156 29588 7162 29600
rect 7469 29597 7481 29631
rect 7515 29597 7527 29631
rect 7469 29591 7527 29597
rect 7653 29631 7711 29637
rect 7653 29597 7665 29631
rect 7699 29597 7711 29631
rect 7653 29591 7711 29597
rect 7484 29492 7512 29591
rect 8294 29588 8300 29640
rect 8352 29588 8358 29640
rect 8478 29588 8484 29640
rect 8536 29628 8542 29640
rect 9306 29628 9312 29640
rect 8536 29600 9312 29628
rect 8536 29588 8542 29600
rect 9306 29588 9312 29600
rect 9364 29588 9370 29640
rect 9493 29631 9551 29637
rect 9493 29597 9505 29631
rect 9539 29628 9551 29631
rect 10134 29628 10140 29640
rect 9539 29600 10140 29628
rect 9539 29597 9551 29600
rect 9493 29591 9551 29597
rect 7561 29563 7619 29569
rect 7561 29529 7573 29563
rect 7607 29560 7619 29563
rect 9508 29560 9536 29591
rect 10134 29588 10140 29600
rect 10192 29588 10198 29640
rect 10226 29588 10232 29640
rect 10284 29588 10290 29640
rect 10686 29588 10692 29640
rect 10744 29588 10750 29640
rect 11793 29631 11851 29637
rect 11793 29628 11805 29631
rect 10796 29600 11805 29628
rect 7607 29532 9536 29560
rect 10152 29560 10180 29588
rect 10796 29560 10824 29600
rect 11793 29597 11805 29600
rect 11839 29597 11851 29631
rect 11793 29591 11851 29597
rect 11885 29631 11943 29637
rect 11885 29597 11897 29631
rect 11931 29628 11943 29631
rect 12986 29628 12992 29640
rect 11931 29600 12992 29628
rect 11931 29597 11943 29600
rect 11885 29591 11943 29597
rect 12986 29588 12992 29600
rect 13044 29628 13050 29640
rect 13722 29628 13728 29640
rect 13044 29600 13728 29628
rect 13044 29588 13050 29600
rect 13722 29588 13728 29600
rect 13780 29588 13786 29640
rect 14734 29588 14740 29640
rect 14792 29628 14798 29640
rect 15657 29631 15715 29637
rect 15657 29628 15669 29631
rect 14792 29600 15669 29628
rect 14792 29588 14798 29600
rect 15657 29597 15669 29600
rect 15703 29597 15715 29631
rect 15657 29591 15715 29597
rect 15930 29588 15936 29640
rect 15988 29588 15994 29640
rect 16022 29588 16028 29640
rect 16080 29588 16086 29640
rect 10152 29532 10824 29560
rect 7607 29529 7619 29532
rect 7561 29523 7619 29529
rect 10870 29520 10876 29572
rect 10928 29560 10934 29572
rect 11238 29560 11244 29572
rect 10928 29532 11244 29560
rect 10928 29520 10934 29532
rect 11238 29520 11244 29532
rect 11296 29520 11302 29572
rect 12250 29520 12256 29572
rect 12308 29560 12314 29572
rect 12434 29560 12440 29572
rect 12308 29532 12440 29560
rect 12308 29520 12314 29532
rect 12434 29520 12440 29532
rect 12492 29520 12498 29572
rect 12618 29520 12624 29572
rect 12676 29520 12682 29572
rect 13078 29520 13084 29572
rect 13136 29560 13142 29572
rect 13357 29563 13415 29569
rect 13357 29560 13369 29563
rect 13136 29532 13369 29560
rect 13136 29520 13142 29532
rect 13357 29529 13369 29532
rect 13403 29529 13415 29563
rect 13357 29523 13415 29529
rect 14274 29520 14280 29572
rect 14332 29520 14338 29572
rect 15010 29520 15016 29572
rect 15068 29520 15074 29572
rect 15470 29520 15476 29572
rect 15528 29560 15534 29572
rect 15841 29563 15899 29569
rect 15841 29560 15853 29563
rect 15528 29532 15853 29560
rect 15528 29520 15534 29532
rect 15841 29529 15853 29532
rect 15887 29560 15899 29563
rect 16390 29560 16396 29572
rect 15887 29532 16396 29560
rect 15887 29529 15899 29532
rect 15841 29523 15899 29529
rect 16390 29520 16396 29532
rect 16448 29520 16454 29572
rect 16500 29560 16528 29668
rect 16942 29588 16948 29640
rect 17000 29628 17006 29640
rect 17221 29631 17279 29637
rect 17221 29628 17233 29631
rect 17000 29600 17233 29628
rect 17000 29588 17006 29600
rect 17221 29597 17233 29600
rect 17267 29628 17279 29631
rect 17310 29628 17316 29640
rect 17267 29600 17316 29628
rect 17267 29597 17279 29600
rect 17221 29591 17279 29597
rect 17310 29588 17316 29600
rect 17368 29588 17374 29640
rect 17954 29588 17960 29640
rect 18012 29628 18018 29640
rect 19150 29628 19156 29640
rect 18012 29600 19156 29628
rect 18012 29588 18018 29600
rect 19150 29588 19156 29600
rect 19208 29628 19214 29640
rect 21192 29637 21220 29804
rect 21284 29804 23612 29832
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 19208 29600 19441 29628
rect 19208 29588 19214 29600
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 21177 29631 21235 29637
rect 21177 29597 21189 29631
rect 21223 29597 21235 29631
rect 21177 29591 21235 29597
rect 17466 29563 17524 29569
rect 17466 29560 17478 29563
rect 16500 29532 17478 29560
rect 17466 29529 17478 29532
rect 17512 29529 17524 29563
rect 17466 29523 17524 29529
rect 17586 29520 17592 29572
rect 17644 29560 17650 29572
rect 17644 29532 19104 29560
rect 17644 29520 17650 29532
rect 8202 29492 8208 29504
rect 7484 29464 8208 29492
rect 8202 29452 8208 29464
rect 8260 29492 8266 29504
rect 8662 29492 8668 29504
rect 8260 29464 8668 29492
rect 8260 29452 8266 29464
rect 8662 29452 8668 29464
rect 8720 29452 8726 29504
rect 9766 29452 9772 29504
rect 9824 29452 9830 29504
rect 12710 29452 12716 29504
rect 12768 29492 12774 29504
rect 13446 29492 13452 29504
rect 12768 29464 13452 29492
rect 12768 29452 12774 29464
rect 13446 29452 13452 29464
rect 13504 29492 13510 29504
rect 13557 29495 13615 29501
rect 13557 29492 13569 29495
rect 13504 29464 13569 29492
rect 13504 29452 13510 29464
rect 13557 29461 13569 29464
rect 13603 29461 13615 29495
rect 13557 29455 13615 29461
rect 13722 29452 13728 29504
rect 13780 29492 13786 29504
rect 16850 29492 16856 29504
rect 13780 29464 16856 29492
rect 13780 29452 13786 29464
rect 16850 29452 16856 29464
rect 16908 29452 16914 29504
rect 18601 29495 18659 29501
rect 18601 29461 18613 29495
rect 18647 29492 18659 29495
rect 18966 29492 18972 29504
rect 18647 29464 18972 29492
rect 18647 29461 18659 29464
rect 18601 29455 18659 29461
rect 18966 29452 18972 29464
rect 19024 29452 19030 29504
rect 19076 29492 19104 29532
rect 19334 29520 19340 29572
rect 19392 29560 19398 29572
rect 20254 29560 20260 29572
rect 19392 29532 20260 29560
rect 19392 29520 19398 29532
rect 20254 29520 20260 29532
rect 20312 29520 20318 29572
rect 21284 29492 21312 29804
rect 21542 29724 21548 29776
rect 21600 29764 21606 29776
rect 22646 29764 22652 29776
rect 21600 29736 22652 29764
rect 21600 29724 21606 29736
rect 22646 29724 22652 29736
rect 22704 29764 22710 29776
rect 23584 29773 23612 29804
rect 24486 29792 24492 29844
rect 24544 29832 24550 29844
rect 27062 29832 27068 29844
rect 24544 29804 27068 29832
rect 24544 29792 24550 29804
rect 27062 29792 27068 29804
rect 27120 29792 27126 29844
rect 27338 29792 27344 29844
rect 27396 29792 27402 29844
rect 28166 29792 28172 29844
rect 28224 29832 28230 29844
rect 29822 29832 29828 29844
rect 28224 29804 29828 29832
rect 28224 29792 28230 29804
rect 29822 29792 29828 29804
rect 29880 29792 29886 29844
rect 30282 29792 30288 29844
rect 30340 29792 30346 29844
rect 30466 29792 30472 29844
rect 30524 29832 30530 29844
rect 34514 29832 34520 29844
rect 30524 29804 34520 29832
rect 30524 29792 30530 29804
rect 34514 29792 34520 29804
rect 34572 29792 34578 29844
rect 34974 29792 34980 29844
rect 35032 29792 35038 29844
rect 36078 29792 36084 29844
rect 36136 29832 36142 29844
rect 36446 29832 36452 29844
rect 36136 29804 36452 29832
rect 36136 29792 36142 29804
rect 36446 29792 36452 29804
rect 36504 29792 36510 29844
rect 36832 29804 38148 29832
rect 23569 29767 23627 29773
rect 22704 29736 23520 29764
rect 22704 29724 22710 29736
rect 21910 29656 21916 29708
rect 21968 29656 21974 29708
rect 22002 29656 22008 29708
rect 22060 29696 22066 29708
rect 23492 29696 23520 29736
rect 23569 29733 23581 29767
rect 23615 29733 23627 29767
rect 23569 29727 23627 29733
rect 25774 29724 25780 29776
rect 25832 29764 25838 29776
rect 30558 29764 30564 29776
rect 25832 29736 30564 29764
rect 25832 29724 25838 29736
rect 30558 29724 30564 29736
rect 30616 29724 30622 29776
rect 30745 29767 30803 29773
rect 30745 29733 30757 29767
rect 30791 29733 30803 29767
rect 30745 29727 30803 29733
rect 22060 29668 23244 29696
rect 23492 29668 24624 29696
rect 22060 29656 22066 29668
rect 21450 29588 21456 29640
rect 21508 29628 21514 29640
rect 21729 29631 21787 29637
rect 21729 29628 21741 29631
rect 21508 29600 21741 29628
rect 21508 29588 21514 29600
rect 21729 29597 21741 29600
rect 21775 29597 21787 29631
rect 21729 29591 21787 29597
rect 22186 29588 22192 29640
rect 22244 29588 22250 29640
rect 22741 29631 22799 29637
rect 22741 29597 22753 29631
rect 22787 29597 22799 29631
rect 23216 29628 23244 29668
rect 23474 29628 23480 29640
rect 23216 29600 23480 29628
rect 22741 29591 22799 29597
rect 21634 29520 21640 29572
rect 21692 29560 21698 29572
rect 22756 29560 22784 29591
rect 23474 29588 23480 29600
rect 23532 29588 23538 29640
rect 23658 29588 23664 29640
rect 23716 29588 23722 29640
rect 23750 29588 23756 29640
rect 23808 29588 23814 29640
rect 23934 29588 23940 29640
rect 23992 29588 23998 29640
rect 24596 29637 24624 29668
rect 24762 29656 24768 29708
rect 24820 29696 24826 29708
rect 25130 29696 25136 29708
rect 24820 29668 25136 29696
rect 24820 29656 24826 29668
rect 25130 29656 25136 29668
rect 25188 29656 25194 29708
rect 25222 29656 25228 29708
rect 25280 29696 25286 29708
rect 25958 29696 25964 29708
rect 25280 29668 25964 29696
rect 25280 29656 25286 29668
rect 25958 29656 25964 29668
rect 26016 29696 26022 29708
rect 30190 29696 30196 29708
rect 26016 29668 27108 29696
rect 26016 29656 26022 29668
rect 24581 29631 24639 29637
rect 24581 29597 24593 29631
rect 24627 29628 24639 29631
rect 24854 29628 24860 29640
rect 24627 29600 24860 29628
rect 24627 29597 24639 29600
rect 24581 29591 24639 29597
rect 24854 29588 24860 29600
rect 24912 29588 24918 29640
rect 25041 29631 25099 29637
rect 25041 29597 25053 29631
rect 25087 29628 25099 29631
rect 25590 29628 25596 29640
rect 25087 29600 25596 29628
rect 25087 29597 25099 29600
rect 25041 29591 25099 29597
rect 25590 29588 25596 29600
rect 25648 29588 25654 29640
rect 26053 29631 26111 29637
rect 26053 29597 26065 29631
rect 26099 29628 26111 29631
rect 26970 29628 26976 29640
rect 26099 29600 26976 29628
rect 26099 29597 26111 29600
rect 26053 29591 26111 29597
rect 26970 29588 26976 29600
rect 27028 29588 27034 29640
rect 26237 29563 26295 29569
rect 26237 29560 26249 29563
rect 21692 29532 26249 29560
rect 21692 29520 21698 29532
rect 26237 29529 26249 29532
rect 26283 29529 26295 29563
rect 26237 29523 26295 29529
rect 26602 29520 26608 29572
rect 26660 29520 26666 29572
rect 26789 29563 26847 29569
rect 26789 29529 26801 29563
rect 26835 29560 26847 29563
rect 27080 29560 27108 29668
rect 27632 29668 30196 29696
rect 27246 29588 27252 29640
rect 27304 29628 27310 29640
rect 27632 29637 27660 29668
rect 30190 29656 30196 29668
rect 30248 29656 30254 29708
rect 30374 29656 30380 29708
rect 30432 29656 30438 29708
rect 30760 29696 30788 29727
rect 33134 29724 33140 29776
rect 33192 29724 33198 29776
rect 33318 29724 33324 29776
rect 33376 29764 33382 29776
rect 33376 29736 34376 29764
rect 33376 29724 33382 29736
rect 32582 29696 32588 29708
rect 30760 29668 32588 29696
rect 32582 29656 32588 29668
rect 32640 29656 32646 29708
rect 27525 29631 27583 29637
rect 27525 29628 27537 29631
rect 27304 29600 27537 29628
rect 27304 29588 27310 29600
rect 27525 29597 27537 29600
rect 27571 29597 27583 29631
rect 27525 29591 27583 29597
rect 27617 29631 27675 29637
rect 27617 29597 27629 29631
rect 27663 29597 27675 29631
rect 27617 29591 27675 29597
rect 28166 29588 28172 29640
rect 28224 29628 28230 29640
rect 28442 29628 28448 29640
rect 28224 29600 28448 29628
rect 28224 29588 28230 29600
rect 28442 29588 28448 29600
rect 28500 29628 28506 29640
rect 28718 29628 28724 29640
rect 28500 29600 28724 29628
rect 28500 29588 28506 29600
rect 28718 29588 28724 29600
rect 28776 29628 28782 29640
rect 28902 29628 28908 29640
rect 28776 29600 28908 29628
rect 28776 29588 28782 29600
rect 28902 29588 28908 29600
rect 28960 29588 28966 29640
rect 28997 29631 29055 29637
rect 28997 29597 29009 29631
rect 29043 29628 29055 29631
rect 29362 29628 29368 29640
rect 29043 29600 29368 29628
rect 29043 29597 29055 29600
rect 28997 29591 29055 29597
rect 26835 29532 27108 29560
rect 26835 29529 26847 29532
rect 26789 29523 26847 29529
rect 27154 29520 27160 29572
rect 27212 29560 27218 29572
rect 27341 29563 27399 29569
rect 27341 29560 27353 29563
rect 27212 29532 27353 29560
rect 27212 29520 27218 29532
rect 27341 29529 27353 29532
rect 27387 29529 27399 29563
rect 27341 29523 27399 29529
rect 27430 29520 27436 29572
rect 27488 29560 27494 29572
rect 27488 29532 28580 29560
rect 27488 29520 27494 29532
rect 19076 29464 21312 29492
rect 23290 29452 23296 29504
rect 23348 29452 23354 29504
rect 23566 29452 23572 29504
rect 23624 29492 23630 29504
rect 24673 29495 24731 29501
rect 24673 29492 24685 29495
rect 23624 29464 24685 29492
rect 23624 29452 23630 29464
rect 24673 29461 24685 29464
rect 24719 29461 24731 29495
rect 24673 29455 24731 29461
rect 26697 29495 26755 29501
rect 26697 29461 26709 29495
rect 26743 29492 26755 29495
rect 27706 29492 27712 29504
rect 26743 29464 27712 29492
rect 26743 29461 26755 29464
rect 26697 29455 26755 29461
rect 27706 29452 27712 29464
rect 27764 29452 27770 29504
rect 27798 29452 27804 29504
rect 27856 29452 27862 29504
rect 28552 29501 28580 29532
rect 28626 29520 28632 29572
rect 28684 29560 28690 29572
rect 29012 29560 29040 29591
rect 29362 29588 29368 29600
rect 29420 29588 29426 29640
rect 30558 29588 30564 29640
rect 30616 29588 30622 29640
rect 31294 29588 31300 29640
rect 31352 29588 31358 29640
rect 31386 29588 31392 29640
rect 31444 29628 31450 29640
rect 31941 29631 31999 29637
rect 31941 29628 31953 29631
rect 31444 29600 31953 29628
rect 31444 29588 31450 29600
rect 31941 29597 31953 29600
rect 31987 29597 31999 29631
rect 31941 29591 31999 29597
rect 32306 29588 32312 29640
rect 32364 29628 32370 29640
rect 33153 29637 33181 29724
rect 33045 29631 33103 29637
rect 33045 29628 33057 29631
rect 32364 29600 33057 29628
rect 32364 29588 32370 29600
rect 33045 29597 33057 29600
rect 33091 29597 33103 29631
rect 33045 29591 33103 29597
rect 33138 29631 33196 29637
rect 33138 29597 33150 29631
rect 33184 29597 33196 29631
rect 33138 29591 33196 29597
rect 33321 29631 33379 29637
rect 33321 29597 33333 29631
rect 33367 29628 33379 29631
rect 33436 29628 33464 29736
rect 33686 29656 33692 29708
rect 33744 29696 33750 29708
rect 34241 29699 34299 29705
rect 34241 29696 34253 29699
rect 33744 29668 34253 29696
rect 33744 29656 33750 29668
rect 34241 29665 34253 29668
rect 34287 29665 34299 29699
rect 34348 29696 34376 29736
rect 34606 29724 34612 29776
rect 34664 29764 34670 29776
rect 36832 29764 36860 29804
rect 34664 29736 36860 29764
rect 38120 29764 38148 29804
rect 38194 29792 38200 29844
rect 38252 29792 38258 29844
rect 38286 29764 38292 29776
rect 38120 29736 38292 29764
rect 34664 29724 34670 29736
rect 34790 29696 34796 29708
rect 34348 29668 34796 29696
rect 34241 29659 34299 29665
rect 34790 29656 34796 29668
rect 34848 29656 34854 29708
rect 34992 29705 35020 29736
rect 38286 29724 38292 29736
rect 38344 29724 38350 29776
rect 34977 29699 35035 29705
rect 34977 29665 34989 29699
rect 35023 29665 35035 29699
rect 34977 29659 35035 29665
rect 35526 29656 35532 29708
rect 35584 29696 35590 29708
rect 36354 29696 36360 29708
rect 35584 29668 35848 29696
rect 35584 29656 35590 29668
rect 33367 29600 33464 29628
rect 33510 29631 33568 29637
rect 33367 29597 33379 29600
rect 33321 29591 33379 29597
rect 33510 29597 33522 29631
rect 33556 29597 33568 29631
rect 33510 29591 33568 29597
rect 28684 29532 29040 29560
rect 28684 29520 28690 29532
rect 29178 29520 29184 29572
rect 29236 29560 29242 29572
rect 29822 29560 29828 29572
rect 29236 29532 29828 29560
rect 29236 29520 29242 29532
rect 29822 29520 29828 29532
rect 29880 29520 29886 29572
rect 30098 29520 30104 29572
rect 30156 29560 30162 29572
rect 30650 29560 30656 29572
rect 30156 29532 30656 29560
rect 30156 29520 30162 29532
rect 30650 29520 30656 29532
rect 30708 29520 30714 29572
rect 30742 29520 30748 29572
rect 30800 29560 30806 29572
rect 33413 29563 33471 29569
rect 33413 29560 33425 29563
rect 30800 29532 33425 29560
rect 30800 29520 30806 29532
rect 33413 29529 33425 29532
rect 33459 29529 33471 29563
rect 33413 29523 33471 29529
rect 33525 29560 33553 29591
rect 33870 29588 33876 29640
rect 33928 29628 33934 29640
rect 34149 29631 34207 29637
rect 34149 29628 34161 29631
rect 33928 29600 34161 29628
rect 33928 29588 33934 29600
rect 34149 29597 34161 29600
rect 34195 29597 34207 29631
rect 34149 29591 34207 29597
rect 34422 29588 34428 29640
rect 34480 29628 34486 29640
rect 34885 29631 34943 29637
rect 34885 29628 34897 29631
rect 34480 29600 34897 29628
rect 34480 29588 34486 29600
rect 34885 29597 34897 29600
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 35710 29588 35716 29640
rect 35768 29588 35774 29640
rect 35820 29637 35848 29668
rect 36096 29668 36360 29696
rect 36096 29637 36124 29668
rect 36354 29656 36360 29668
rect 36412 29656 36418 29708
rect 35806 29631 35864 29637
rect 35806 29597 35818 29631
rect 35852 29597 35864 29631
rect 35806 29591 35864 29597
rect 36081 29631 36139 29637
rect 36081 29597 36093 29631
rect 36127 29597 36139 29631
rect 36081 29591 36139 29597
rect 36219 29631 36277 29637
rect 36219 29597 36231 29631
rect 36265 29628 36277 29631
rect 36538 29628 36544 29640
rect 36265 29600 36544 29628
rect 36265 29597 36277 29600
rect 36219 29591 36277 29597
rect 36538 29588 36544 29600
rect 36596 29588 36602 29640
rect 36630 29588 36636 29640
rect 36688 29628 36694 29640
rect 36817 29631 36875 29637
rect 36817 29628 36829 29631
rect 36688 29600 36829 29628
rect 36688 29588 36694 29600
rect 36817 29597 36829 29600
rect 36863 29628 36875 29631
rect 36906 29628 36912 29640
rect 36863 29600 36912 29628
rect 36863 29597 36875 29600
rect 36817 29591 36875 29597
rect 36906 29588 36912 29600
rect 36964 29588 36970 29640
rect 37084 29631 37142 29637
rect 37084 29597 37096 29631
rect 37130 29628 37142 29631
rect 37458 29628 37464 29640
rect 37130 29600 37464 29628
rect 37130 29597 37142 29600
rect 37084 29591 37142 29597
rect 37458 29588 37464 29600
rect 37516 29588 37522 29640
rect 34698 29560 34704 29572
rect 33525 29532 34704 29560
rect 28537 29495 28595 29501
rect 28537 29461 28549 29495
rect 28583 29461 28595 29495
rect 28537 29455 28595 29461
rect 29730 29452 29736 29504
rect 29788 29452 29794 29504
rect 30466 29452 30472 29504
rect 30524 29492 30530 29504
rect 31478 29492 31484 29504
rect 30524 29464 31484 29492
rect 30524 29452 30530 29464
rect 31478 29452 31484 29464
rect 31536 29452 31542 29504
rect 32309 29495 32367 29501
rect 32309 29461 32321 29495
rect 32355 29492 32367 29495
rect 33226 29492 33232 29504
rect 32355 29464 33232 29492
rect 32355 29461 32367 29464
rect 32309 29455 32367 29461
rect 33226 29452 33232 29464
rect 33284 29492 33290 29504
rect 33525 29492 33553 29532
rect 34698 29520 34704 29532
rect 34756 29520 34762 29572
rect 35989 29563 36047 29569
rect 35989 29529 36001 29563
rect 36035 29560 36047 29563
rect 36556 29560 36584 29588
rect 37550 29560 37556 29572
rect 36035 29532 36492 29560
rect 36556 29532 37556 29560
rect 36035 29529 36047 29532
rect 35989 29523 36047 29529
rect 36188 29504 36216 29532
rect 33284 29464 33553 29492
rect 33284 29452 33290 29464
rect 33686 29452 33692 29504
rect 33744 29452 33750 29504
rect 34606 29452 34612 29504
rect 34664 29492 34670 29504
rect 35253 29495 35311 29501
rect 35253 29492 35265 29495
rect 34664 29464 35265 29492
rect 34664 29452 34670 29464
rect 35253 29461 35265 29464
rect 35299 29461 35311 29495
rect 35253 29455 35311 29461
rect 36170 29452 36176 29504
rect 36228 29452 36234 29504
rect 36354 29452 36360 29504
rect 36412 29452 36418 29504
rect 36464 29492 36492 29532
rect 37550 29520 37556 29532
rect 37608 29520 37614 29572
rect 36538 29492 36544 29504
rect 36464 29464 36544 29492
rect 36538 29452 36544 29464
rect 36596 29452 36602 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 7466 29248 7472 29300
rect 7524 29248 7530 29300
rect 8110 29248 8116 29300
rect 8168 29248 8174 29300
rect 8386 29248 8392 29300
rect 8444 29288 8450 29300
rect 9582 29288 9588 29300
rect 8444 29260 9588 29288
rect 8444 29248 8450 29260
rect 9582 29248 9588 29260
rect 9640 29248 9646 29300
rect 9674 29248 9680 29300
rect 9732 29288 9738 29300
rect 12710 29288 12716 29300
rect 9732 29260 12716 29288
rect 9732 29248 9738 29260
rect 12710 29248 12716 29260
rect 12768 29248 12774 29300
rect 13906 29288 13912 29300
rect 12912 29260 13912 29288
rect 7374 29180 7380 29232
rect 7432 29220 7438 29232
rect 12912 29229 12940 29260
rect 13906 29248 13912 29260
rect 13964 29248 13970 29300
rect 14826 29248 14832 29300
rect 14884 29288 14890 29300
rect 14884 29260 15792 29288
rect 14884 29248 14890 29260
rect 12897 29223 12955 29229
rect 7432 29192 10916 29220
rect 7432 29180 7438 29192
rect 7285 29155 7343 29161
rect 7285 29121 7297 29155
rect 7331 29121 7343 29155
rect 7285 29115 7343 29121
rect 7469 29155 7527 29161
rect 7469 29121 7481 29155
rect 7515 29152 7527 29155
rect 7558 29152 7564 29164
rect 7515 29124 7564 29152
rect 7515 29121 7527 29124
rect 7469 29115 7527 29121
rect 7300 29084 7328 29115
rect 7558 29112 7564 29124
rect 7616 29112 7622 29164
rect 7926 29112 7932 29164
rect 7984 29112 7990 29164
rect 8113 29155 8171 29161
rect 8113 29121 8125 29155
rect 8159 29152 8171 29155
rect 8202 29152 8208 29164
rect 8159 29124 8208 29152
rect 8159 29121 8171 29124
rect 8113 29115 8171 29121
rect 8202 29112 8208 29124
rect 8260 29112 8266 29164
rect 8573 29155 8631 29161
rect 8573 29121 8585 29155
rect 8619 29121 8631 29155
rect 8573 29115 8631 29121
rect 8386 29084 8392 29096
rect 7300 29056 8392 29084
rect 8386 29044 8392 29056
rect 8444 29044 8450 29096
rect 4614 28976 4620 29028
rect 4672 29016 4678 29028
rect 7006 29016 7012 29028
rect 4672 28988 7012 29016
rect 4672 28976 4678 28988
rect 7006 28976 7012 28988
rect 7064 28976 7070 29028
rect 4522 28908 4528 28960
rect 4580 28948 4586 28960
rect 7190 28948 7196 28960
rect 4580 28920 7196 28948
rect 4580 28908 4586 28920
rect 7190 28908 7196 28920
rect 7248 28908 7254 28960
rect 7834 28908 7840 28960
rect 7892 28948 7898 28960
rect 8588 28948 8616 29115
rect 8754 29112 8760 29164
rect 8812 29112 8818 29164
rect 8846 29112 8852 29164
rect 8904 29152 8910 29164
rect 9493 29155 9551 29161
rect 9493 29152 9505 29155
rect 8904 29124 9505 29152
rect 8904 29112 8910 29124
rect 9493 29121 9505 29124
rect 9539 29121 9551 29155
rect 9493 29115 9551 29121
rect 9677 29155 9735 29161
rect 9677 29121 9689 29155
rect 9723 29152 9735 29155
rect 9766 29152 9772 29164
rect 9723 29124 9772 29152
rect 9723 29121 9735 29124
rect 9677 29115 9735 29121
rect 9766 29112 9772 29124
rect 9824 29112 9830 29164
rect 10410 29112 10416 29164
rect 10468 29152 10474 29164
rect 10594 29152 10600 29164
rect 10468 29124 10600 29152
rect 10468 29112 10474 29124
rect 10594 29112 10600 29124
rect 10652 29112 10658 29164
rect 10689 29155 10747 29161
rect 10689 29121 10701 29155
rect 10735 29152 10747 29155
rect 10778 29152 10784 29164
rect 10735 29124 10784 29152
rect 10735 29121 10747 29124
rect 10689 29115 10747 29121
rect 10778 29112 10784 29124
rect 10836 29112 10842 29164
rect 10888 29152 10916 29192
rect 11348 29192 12434 29220
rect 11348 29152 11376 29192
rect 10888 29124 11376 29152
rect 11698 29112 11704 29164
rect 11756 29152 11762 29164
rect 11977 29155 12035 29161
rect 11977 29152 11989 29155
rect 11756 29124 11989 29152
rect 11756 29112 11762 29124
rect 11977 29121 11989 29124
rect 12023 29121 12035 29155
rect 12406 29152 12434 29192
rect 12897 29189 12909 29223
rect 12943 29189 12955 29223
rect 15010 29220 15016 29232
rect 12897 29183 12955 29189
rect 13004 29192 15016 29220
rect 13004 29152 13032 29192
rect 12406 29124 13032 29152
rect 13081 29155 13139 29161
rect 11977 29115 12035 29121
rect 13081 29121 13093 29155
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 13173 29155 13231 29161
rect 13173 29121 13185 29155
rect 13219 29152 13231 29155
rect 13262 29152 13268 29164
rect 13219 29124 13268 29152
rect 13219 29121 13231 29124
rect 13173 29115 13231 29121
rect 9214 29044 9220 29096
rect 9272 29044 9278 29096
rect 9398 29044 9404 29096
rect 9456 29044 9462 29096
rect 9582 29084 9588 29096
rect 9508 29056 9588 29084
rect 8662 28976 8668 29028
rect 8720 28976 8726 29028
rect 8846 29016 8852 29028
rect 8772 28988 8852 29016
rect 8772 28948 8800 28988
rect 8846 28976 8852 28988
rect 8904 28976 8910 29028
rect 8938 28976 8944 29028
rect 8996 29016 9002 29028
rect 9508 29016 9536 29056
rect 9582 29044 9588 29056
rect 9640 29044 9646 29096
rect 11514 29044 11520 29096
rect 11572 29084 11578 29096
rect 12161 29087 12219 29093
rect 12161 29084 12173 29087
rect 11572 29056 12173 29084
rect 11572 29044 11578 29056
rect 12161 29053 12173 29056
rect 12207 29053 12219 29087
rect 12161 29047 12219 29053
rect 12618 29044 12624 29096
rect 12676 29084 12682 29096
rect 13096 29084 13124 29115
rect 13262 29112 13268 29124
rect 13320 29112 13326 29164
rect 13648 29161 13676 29192
rect 15010 29180 15016 29192
rect 15068 29180 15074 29232
rect 15764 29229 15792 29260
rect 17770 29248 17776 29300
rect 17828 29288 17834 29300
rect 20533 29291 20591 29297
rect 17828 29260 20392 29288
rect 17828 29248 17834 29260
rect 15749 29223 15807 29229
rect 15749 29189 15761 29223
rect 15795 29220 15807 29223
rect 17034 29220 17040 29232
rect 15795 29192 17040 29220
rect 15795 29189 15807 29192
rect 15749 29183 15807 29189
rect 17034 29180 17040 29192
rect 17092 29220 17098 29232
rect 20254 29220 20260 29232
rect 17092 29192 18368 29220
rect 17092 29180 17098 29192
rect 13633 29155 13691 29161
rect 13633 29121 13645 29155
rect 13679 29121 13691 29155
rect 13889 29155 13947 29161
rect 13889 29152 13901 29155
rect 13633 29115 13691 29121
rect 13740 29124 13901 29152
rect 13740 29084 13768 29124
rect 13889 29121 13901 29124
rect 13935 29121 13947 29155
rect 13889 29115 13947 29121
rect 14734 29112 14740 29164
rect 14792 29152 14798 29164
rect 15473 29155 15531 29161
rect 15473 29152 15485 29155
rect 14792 29124 15485 29152
rect 14792 29112 14798 29124
rect 15473 29121 15485 29124
rect 15519 29121 15531 29155
rect 15473 29115 15531 29121
rect 15562 29112 15568 29164
rect 15620 29152 15626 29164
rect 15657 29155 15715 29161
rect 15657 29152 15669 29155
rect 15620 29124 15669 29152
rect 15620 29112 15626 29124
rect 15657 29121 15669 29124
rect 15703 29121 15715 29155
rect 15657 29115 15715 29121
rect 15841 29155 15899 29161
rect 15841 29121 15853 29155
rect 15887 29152 15899 29155
rect 16022 29152 16028 29164
rect 15887 29124 16028 29152
rect 15887 29121 15899 29124
rect 15841 29115 15899 29121
rect 16022 29112 16028 29124
rect 16080 29112 16086 29164
rect 16850 29112 16856 29164
rect 16908 29112 16914 29164
rect 17126 29112 17132 29164
rect 17184 29152 17190 29164
rect 18340 29161 18368 29192
rect 19168 29192 20260 29220
rect 18141 29155 18199 29161
rect 18141 29152 18153 29155
rect 17184 29124 18153 29152
rect 17184 29112 17190 29124
rect 18141 29121 18153 29124
rect 18187 29121 18199 29155
rect 18141 29115 18199 29121
rect 18325 29155 18383 29161
rect 18325 29121 18337 29155
rect 18371 29121 18383 29155
rect 18325 29115 18383 29121
rect 18417 29155 18475 29161
rect 18417 29121 18429 29155
rect 18463 29152 18475 29155
rect 18506 29152 18512 29164
rect 18463 29124 18512 29152
rect 18463 29121 18475 29124
rect 18417 29115 18475 29121
rect 18506 29112 18512 29124
rect 18564 29112 18570 29164
rect 19168 29161 19196 29192
rect 20254 29180 20260 29192
rect 20312 29180 20318 29232
rect 19153 29155 19211 29161
rect 19153 29121 19165 29155
rect 19199 29121 19211 29155
rect 19153 29115 19211 29121
rect 19242 29112 19248 29164
rect 19300 29152 19306 29164
rect 19409 29155 19467 29161
rect 19409 29152 19421 29155
rect 19300 29124 19421 29152
rect 19300 29112 19306 29124
rect 19409 29121 19421 29124
rect 19455 29121 19467 29155
rect 20364 29152 20392 29260
rect 20533 29257 20545 29291
rect 20579 29257 20591 29291
rect 20533 29251 20591 29257
rect 20548 29220 20576 29251
rect 20714 29248 20720 29300
rect 20772 29288 20778 29300
rect 20993 29291 21051 29297
rect 20993 29288 21005 29291
rect 20772 29260 21005 29288
rect 20772 29248 20778 29260
rect 20993 29257 21005 29260
rect 21039 29257 21051 29291
rect 20993 29251 21051 29257
rect 21266 29248 21272 29300
rect 21324 29288 21330 29300
rect 21361 29291 21419 29297
rect 21361 29288 21373 29291
rect 21324 29260 21373 29288
rect 21324 29248 21330 29260
rect 21361 29257 21373 29260
rect 21407 29257 21419 29291
rect 21361 29251 21419 29257
rect 22462 29248 22468 29300
rect 22520 29248 22526 29300
rect 22922 29248 22928 29300
rect 22980 29288 22986 29300
rect 23753 29291 23811 29297
rect 23753 29288 23765 29291
rect 22980 29260 23765 29288
rect 22980 29248 22986 29260
rect 23753 29257 23765 29260
rect 23799 29257 23811 29291
rect 23753 29251 23811 29257
rect 24121 29291 24179 29297
rect 24121 29257 24133 29291
rect 24167 29288 24179 29291
rect 24578 29288 24584 29300
rect 24167 29260 24584 29288
rect 24167 29257 24179 29260
rect 24121 29251 24179 29257
rect 24578 29248 24584 29260
rect 24636 29248 24642 29300
rect 24673 29291 24731 29297
rect 24673 29257 24685 29291
rect 24719 29288 24731 29291
rect 24762 29288 24768 29300
rect 24719 29260 24768 29288
rect 24719 29257 24731 29260
rect 24673 29251 24731 29257
rect 24762 29248 24768 29260
rect 24820 29248 24826 29300
rect 24946 29248 24952 29300
rect 25004 29288 25010 29300
rect 26418 29288 26424 29300
rect 25004 29260 26424 29288
rect 25004 29248 25010 29260
rect 26418 29248 26424 29260
rect 26476 29248 26482 29300
rect 26513 29291 26571 29297
rect 26513 29257 26525 29291
rect 26559 29288 26571 29291
rect 26602 29288 26608 29300
rect 26559 29260 26608 29288
rect 26559 29257 26571 29260
rect 26513 29251 26571 29257
rect 26602 29248 26608 29260
rect 26660 29248 26666 29300
rect 29270 29288 29276 29300
rect 27724 29260 29276 29288
rect 21284 29220 21312 29248
rect 20548 29192 21312 29220
rect 21177 29155 21235 29161
rect 21177 29152 21189 29155
rect 20364 29124 21189 29152
rect 19409 29115 19467 29121
rect 21177 29121 21189 29124
rect 21223 29121 21235 29155
rect 21177 29115 21235 29121
rect 21266 29112 21272 29164
rect 21324 29152 21330 29164
rect 21453 29155 21511 29161
rect 21453 29152 21465 29155
rect 21324 29124 21465 29152
rect 21324 29112 21330 29124
rect 21453 29121 21465 29124
rect 21499 29152 21511 29155
rect 22094 29152 22100 29164
rect 21499 29124 22100 29152
rect 21499 29121 21511 29124
rect 21453 29115 21511 29121
rect 22094 29112 22100 29124
rect 22152 29112 22158 29164
rect 22370 29112 22376 29164
rect 22428 29112 22434 29164
rect 23937 29155 23995 29161
rect 23937 29152 23949 29155
rect 22572 29124 23949 29152
rect 12676 29056 13124 29084
rect 13648 29056 13768 29084
rect 16040 29084 16068 29112
rect 17037 29087 17095 29093
rect 17037 29084 17049 29087
rect 16040 29056 17049 29084
rect 12676 29044 12682 29056
rect 8996 28988 9536 29016
rect 8996 28976 9002 28988
rect 9674 28976 9680 29028
rect 9732 28976 9738 29028
rect 10502 28976 10508 29028
rect 10560 29016 10566 29028
rect 10597 29019 10655 29025
rect 10597 29016 10609 29019
rect 10560 28988 10609 29016
rect 10560 28976 10566 28988
rect 10597 28985 10609 28988
rect 10643 28985 10655 29019
rect 10597 28979 10655 28985
rect 11974 28976 11980 29028
rect 12032 29016 12038 29028
rect 12897 29019 12955 29025
rect 12897 29016 12909 29019
rect 12032 28988 12909 29016
rect 12032 28976 12038 28988
rect 12897 28985 12909 28988
rect 12943 28985 12955 29019
rect 12897 28979 12955 28985
rect 13078 28976 13084 29028
rect 13136 29016 13142 29028
rect 13648 29016 13676 29056
rect 17037 29053 17049 29056
rect 17083 29084 17095 29087
rect 17218 29084 17224 29096
rect 17083 29056 17224 29084
rect 17083 29053 17095 29056
rect 17037 29047 17095 29053
rect 17218 29044 17224 29056
rect 17276 29044 17282 29096
rect 20990 29044 20996 29096
rect 21048 29084 21054 29096
rect 22572 29084 22600 29124
rect 23937 29121 23949 29124
rect 23983 29121 23995 29155
rect 23937 29115 23995 29121
rect 21048 29056 22600 29084
rect 22649 29087 22707 29093
rect 21048 29044 21054 29056
rect 22649 29053 22661 29087
rect 22695 29084 22707 29087
rect 23474 29084 23480 29096
rect 22695 29056 23480 29084
rect 22695 29053 22707 29056
rect 22649 29047 22707 29053
rect 23474 29044 23480 29056
rect 23532 29044 23538 29096
rect 13136 28988 13676 29016
rect 15856 28988 16160 29016
rect 13136 28976 13142 28988
rect 9692 28948 9720 28976
rect 7892 28920 9720 28948
rect 7892 28908 7898 28920
rect 9858 28908 9864 28960
rect 9916 28948 9922 28960
rect 10229 28951 10287 28957
rect 10229 28948 10241 28951
rect 9916 28920 10241 28948
rect 9916 28908 9922 28920
rect 10229 28917 10241 28920
rect 10275 28917 10287 28951
rect 10229 28911 10287 28917
rect 10410 28908 10416 28960
rect 10468 28948 10474 28960
rect 10962 28948 10968 28960
rect 10468 28920 10968 28948
rect 10468 28908 10474 28920
rect 10962 28908 10968 28920
rect 11020 28908 11026 28960
rect 15010 28908 15016 28960
rect 15068 28908 15074 28960
rect 15194 28908 15200 28960
rect 15252 28948 15258 28960
rect 15856 28948 15884 28988
rect 15252 28920 15884 28948
rect 15252 28908 15258 28920
rect 15930 28908 15936 28960
rect 15988 28948 15994 28960
rect 16025 28951 16083 28957
rect 16025 28948 16037 28951
rect 15988 28920 16037 28948
rect 15988 28908 15994 28920
rect 16025 28917 16037 28920
rect 16071 28917 16083 28951
rect 16132 28948 16160 28988
rect 18598 28976 18604 29028
rect 18656 28976 18662 29028
rect 23750 29016 23756 29028
rect 20088 28988 23756 29016
rect 20088 28960 20116 28988
rect 23750 28976 23756 28988
rect 23808 28976 23814 29028
rect 23952 29016 23980 29115
rect 24210 29112 24216 29164
rect 24268 29112 24274 29164
rect 24854 29112 24860 29164
rect 24912 29112 24918 29164
rect 24964 29161 24992 29248
rect 25682 29180 25688 29232
rect 25740 29220 25746 29232
rect 26053 29223 26111 29229
rect 26053 29220 26065 29223
rect 25740 29192 26065 29220
rect 25740 29180 25746 29192
rect 26053 29189 26065 29192
rect 26099 29189 26111 29223
rect 27724 29220 27752 29260
rect 26053 29183 26111 29189
rect 26160 29192 27752 29220
rect 24949 29155 25007 29161
rect 24949 29121 24961 29155
rect 24995 29121 25007 29155
rect 24949 29115 25007 29121
rect 25038 29112 25044 29164
rect 25096 29112 25102 29164
rect 25133 29155 25191 29161
rect 25133 29121 25145 29155
rect 25179 29121 25191 29155
rect 25133 29115 25191 29121
rect 25317 29155 25375 29161
rect 25317 29121 25329 29155
rect 25363 29152 25375 29155
rect 25498 29152 25504 29164
rect 25363 29124 25504 29152
rect 25363 29121 25375 29124
rect 25317 29115 25375 29121
rect 25148 29084 25176 29115
rect 25498 29112 25504 29124
rect 25556 29112 25562 29164
rect 26160 29084 26188 29192
rect 27890 29180 27896 29232
rect 27948 29220 27954 29232
rect 28537 29223 28595 29229
rect 28537 29220 28549 29223
rect 27948 29192 28549 29220
rect 27948 29180 27954 29192
rect 28537 29189 28549 29192
rect 28583 29189 28595 29223
rect 28537 29183 28595 29189
rect 26329 29155 26387 29161
rect 26329 29121 26341 29155
rect 26375 29152 26387 29155
rect 26878 29152 26884 29164
rect 26375 29124 26884 29152
rect 26375 29121 26387 29124
rect 26329 29115 26387 29121
rect 26878 29112 26884 29124
rect 26936 29112 26942 29164
rect 27062 29112 27068 29164
rect 27120 29152 27126 29164
rect 27157 29155 27215 29161
rect 27157 29152 27169 29155
rect 27120 29124 27169 29152
rect 27120 29112 27126 29124
rect 27157 29121 27169 29124
rect 27203 29121 27215 29155
rect 27157 29115 27215 29121
rect 27338 29112 27344 29164
rect 27396 29112 27402 29164
rect 28166 29112 28172 29164
rect 28224 29112 28230 29164
rect 28258 29112 28264 29164
rect 28316 29152 28322 29164
rect 28353 29155 28411 29161
rect 28353 29152 28365 29155
rect 28316 29124 28365 29152
rect 28316 29112 28322 29124
rect 28353 29121 28365 29124
rect 28399 29121 28411 29155
rect 28353 29115 28411 29121
rect 25148 29056 26188 29084
rect 26234 29044 26240 29096
rect 26292 29084 26298 29096
rect 28828 29084 28856 29260
rect 29270 29248 29276 29260
rect 29328 29248 29334 29300
rect 31938 29288 31944 29300
rect 29472 29260 31944 29288
rect 29089 29223 29147 29229
rect 29089 29189 29101 29223
rect 29135 29220 29147 29223
rect 29178 29220 29184 29232
rect 29135 29192 29184 29220
rect 29135 29189 29147 29192
rect 29089 29183 29147 29189
rect 29178 29180 29184 29192
rect 29236 29180 29242 29232
rect 29362 29112 29368 29164
rect 29420 29112 29426 29164
rect 29472 29161 29500 29260
rect 31938 29248 31944 29260
rect 31996 29248 32002 29300
rect 32674 29248 32680 29300
rect 32732 29288 32738 29300
rect 33226 29288 33232 29300
rect 32732 29260 33232 29288
rect 32732 29248 32738 29260
rect 33226 29248 33232 29260
rect 33284 29248 33290 29300
rect 33870 29288 33876 29300
rect 33336 29260 33876 29288
rect 29822 29180 29828 29232
rect 29880 29220 29886 29232
rect 29880 29192 30880 29220
rect 29880 29180 29886 29192
rect 29457 29155 29515 29161
rect 29457 29121 29469 29155
rect 29503 29121 29515 29155
rect 29457 29115 29515 29121
rect 29549 29155 29607 29161
rect 29549 29121 29561 29155
rect 29595 29121 29607 29155
rect 29549 29115 29607 29121
rect 29733 29155 29791 29161
rect 29733 29121 29745 29155
rect 29779 29121 29791 29155
rect 29733 29115 29791 29121
rect 29564 29084 29592 29115
rect 26292 29056 28764 29084
rect 28828 29056 29592 29084
rect 29748 29084 29776 29115
rect 30466 29112 30472 29164
rect 30524 29112 30530 29164
rect 30558 29112 30564 29164
rect 30616 29112 30622 29164
rect 30650 29112 30656 29164
rect 30708 29112 30714 29164
rect 30852 29161 30880 29192
rect 30926 29180 30932 29232
rect 30984 29220 30990 29232
rect 31573 29223 31631 29229
rect 31573 29220 31585 29223
rect 30984 29192 31585 29220
rect 30984 29180 30990 29192
rect 31573 29189 31585 29192
rect 31619 29189 31631 29223
rect 31573 29183 31631 29189
rect 33042 29180 33048 29232
rect 33100 29180 33106 29232
rect 30837 29155 30895 29161
rect 30837 29121 30849 29155
rect 30883 29121 30895 29155
rect 30837 29115 30895 29121
rect 31294 29112 31300 29164
rect 31352 29112 31358 29164
rect 32585 29155 32643 29161
rect 32585 29121 32597 29155
rect 32631 29152 32643 29155
rect 32766 29152 32772 29164
rect 32631 29124 32772 29152
rect 32631 29121 32643 29124
rect 32585 29115 32643 29121
rect 32766 29112 32772 29124
rect 32824 29112 32830 29164
rect 31018 29084 31024 29096
rect 29748 29056 31024 29084
rect 26292 29044 26298 29056
rect 23952 28988 25268 29016
rect 16390 28948 16396 28960
rect 16132 28920 16396 28948
rect 16025 28911 16083 28917
rect 16390 28908 16396 28920
rect 16448 28948 16454 28960
rect 16666 28948 16672 28960
rect 16448 28920 16672 28948
rect 16448 28908 16454 28920
rect 16666 28908 16672 28920
rect 16724 28908 16730 28960
rect 17678 28908 17684 28960
rect 17736 28948 17742 28960
rect 18141 28951 18199 28957
rect 18141 28948 18153 28951
rect 17736 28920 18153 28948
rect 17736 28908 17742 28920
rect 18141 28917 18153 28920
rect 18187 28917 18199 28951
rect 18141 28911 18199 28917
rect 20070 28908 20076 28960
rect 20128 28908 20134 28960
rect 22002 28908 22008 28960
rect 22060 28908 22066 28960
rect 22278 28908 22284 28960
rect 22336 28948 22342 28960
rect 23658 28948 23664 28960
rect 22336 28920 23664 28948
rect 22336 28908 22342 28920
rect 23658 28908 23664 28920
rect 23716 28908 23722 28960
rect 25240 28948 25268 28988
rect 25682 28976 25688 29028
rect 25740 29016 25746 29028
rect 27433 29019 27491 29025
rect 27433 29016 27445 29019
rect 25740 28988 27445 29016
rect 25740 28976 25746 28988
rect 27433 28985 27445 28988
rect 27479 28985 27491 29019
rect 28736 29016 28764 29056
rect 31018 29044 31024 29056
rect 31076 29044 31082 29096
rect 31478 29044 31484 29096
rect 31536 29084 31542 29096
rect 33336 29084 33364 29260
rect 33870 29248 33876 29260
rect 33928 29248 33934 29300
rect 34238 29288 34244 29300
rect 33980 29260 34244 29288
rect 33502 29180 33508 29232
rect 33560 29220 33566 29232
rect 33980 29229 34008 29260
rect 34238 29248 34244 29260
rect 34296 29248 34302 29300
rect 34333 29291 34391 29297
rect 34333 29257 34345 29291
rect 34379 29257 34391 29291
rect 35526 29288 35532 29300
rect 34333 29251 34391 29257
rect 34992 29260 35532 29288
rect 33965 29223 34023 29229
rect 33965 29220 33977 29223
rect 33560 29192 33977 29220
rect 33560 29180 33566 29192
rect 33965 29189 33977 29192
rect 34011 29189 34023 29223
rect 33965 29183 34023 29189
rect 34054 29180 34060 29232
rect 34112 29180 34118 29232
rect 33686 29112 33692 29164
rect 33744 29112 33750 29164
rect 33782 29155 33840 29161
rect 33782 29121 33794 29155
rect 33828 29121 33840 29155
rect 33782 29115 33840 29121
rect 33797 29084 33825 29115
rect 34146 29112 34152 29164
rect 34204 29161 34210 29164
rect 34204 29152 34212 29161
rect 34204 29124 34249 29152
rect 34204 29115 34212 29124
rect 34204 29112 34210 29115
rect 31536 29056 33364 29084
rect 33704 29056 33825 29084
rect 31536 29044 31542 29056
rect 33704 29028 33732 29056
rect 34238 29044 34244 29096
rect 34296 29084 34302 29096
rect 34348 29084 34376 29251
rect 34992 29161 35020 29260
rect 35526 29248 35532 29260
rect 35584 29248 35590 29300
rect 36354 29248 36360 29300
rect 36412 29288 36418 29300
rect 37921 29291 37979 29297
rect 37921 29288 37933 29291
rect 36412 29260 37933 29288
rect 36412 29248 36418 29260
rect 37921 29257 37933 29260
rect 37967 29257 37979 29291
rect 37921 29251 37979 29257
rect 36446 29220 36452 29232
rect 35360 29192 36452 29220
rect 34977 29155 35035 29161
rect 34977 29121 34989 29155
rect 35023 29121 35035 29155
rect 34977 29115 35035 29121
rect 35066 29112 35072 29164
rect 35124 29112 35130 29164
rect 35360 29161 35388 29192
rect 36446 29180 36452 29192
rect 36504 29180 36510 29232
rect 37182 29180 37188 29232
rect 37240 29220 37246 29232
rect 37829 29223 37887 29229
rect 37829 29220 37841 29223
rect 37240 29192 37841 29220
rect 37240 29180 37246 29192
rect 37829 29189 37841 29192
rect 37875 29220 37887 29223
rect 38194 29220 38200 29232
rect 37875 29192 38200 29220
rect 37875 29189 37887 29192
rect 37829 29183 37887 29189
rect 38194 29180 38200 29192
rect 38252 29180 38258 29232
rect 35253 29155 35311 29161
rect 35253 29121 35265 29155
rect 35299 29121 35311 29155
rect 35253 29115 35311 29121
rect 35345 29155 35403 29161
rect 35345 29121 35357 29155
rect 35391 29121 35403 29155
rect 35345 29115 35403 29121
rect 34296 29056 34376 29084
rect 34296 29044 34302 29056
rect 34514 29044 34520 29096
rect 34572 29084 34578 29096
rect 34793 29087 34851 29093
rect 34793 29084 34805 29087
rect 34572 29056 34805 29084
rect 34572 29044 34578 29056
rect 34793 29053 34805 29056
rect 34839 29053 34851 29087
rect 34793 29047 34851 29053
rect 34882 29044 34888 29096
rect 34940 29044 34946 29096
rect 35268 29084 35296 29115
rect 35710 29112 35716 29164
rect 35768 29152 35774 29164
rect 35805 29155 35863 29161
rect 35805 29152 35817 29155
rect 35768 29124 35817 29152
rect 35768 29112 35774 29124
rect 35805 29121 35817 29124
rect 35851 29121 35863 29155
rect 35805 29115 35863 29121
rect 35986 29112 35992 29164
rect 36044 29112 36050 29164
rect 35894 29084 35900 29096
rect 35268 29056 35900 29084
rect 35894 29044 35900 29056
rect 35952 29044 35958 29096
rect 36004 29084 36032 29112
rect 37918 29084 37924 29096
rect 36004 29056 37924 29084
rect 37918 29044 37924 29056
rect 37976 29044 37982 29096
rect 38102 29044 38108 29096
rect 38160 29044 38166 29096
rect 30558 29016 30564 29028
rect 28736 28988 30564 29016
rect 27433 28979 27491 28985
rect 30558 28976 30564 28988
rect 30616 28976 30622 29028
rect 33686 28976 33692 29028
rect 33744 28976 33750 29028
rect 34900 29016 34928 29044
rect 35434 29016 35440 29028
rect 34900 28988 35440 29016
rect 35434 28976 35440 28988
rect 35492 29016 35498 29028
rect 35492 28988 36124 29016
rect 35492 28976 35498 28988
rect 26053 28951 26111 28957
rect 26053 28948 26065 28951
rect 25240 28920 26065 28948
rect 26053 28917 26065 28920
rect 26099 28917 26111 28951
rect 26053 28911 26111 28917
rect 26510 28908 26516 28960
rect 26568 28948 26574 28960
rect 27062 28948 27068 28960
rect 26568 28920 27068 28948
rect 26568 28908 26574 28920
rect 27062 28908 27068 28920
rect 27120 28908 27126 28960
rect 27338 28908 27344 28960
rect 27396 28948 27402 28960
rect 27890 28948 27896 28960
rect 27396 28920 27896 28948
rect 27396 28908 27402 28920
rect 27890 28908 27896 28920
rect 27948 28908 27954 28960
rect 28445 28951 28503 28957
rect 28445 28917 28457 28951
rect 28491 28948 28503 28951
rect 29270 28948 29276 28960
rect 28491 28920 29276 28948
rect 28491 28917 28503 28920
rect 28445 28911 28503 28917
rect 29270 28908 29276 28920
rect 29328 28908 29334 28960
rect 29362 28908 29368 28960
rect 29420 28948 29426 28960
rect 30193 28951 30251 28957
rect 30193 28948 30205 28951
rect 29420 28920 30205 28948
rect 29420 28908 29426 28920
rect 30193 28917 30205 28920
rect 30239 28917 30251 28951
rect 30193 28911 30251 28917
rect 30466 28908 30472 28960
rect 30524 28948 30530 28960
rect 31202 28948 31208 28960
rect 30524 28920 31208 28948
rect 30524 28908 30530 28920
rect 31202 28908 31208 28920
rect 31260 28908 31266 28960
rect 32766 28908 32772 28960
rect 32824 28948 32830 28960
rect 35710 28948 35716 28960
rect 32824 28920 35716 28948
rect 32824 28908 32830 28920
rect 35710 28908 35716 28920
rect 35768 28948 35774 28960
rect 35986 28948 35992 28960
rect 35768 28920 35992 28948
rect 35768 28908 35774 28920
rect 35986 28908 35992 28920
rect 36044 28908 36050 28960
rect 36096 28957 36124 28988
rect 36081 28951 36139 28957
rect 36081 28917 36093 28951
rect 36127 28917 36139 28951
rect 36081 28911 36139 28917
rect 37458 28908 37464 28960
rect 37516 28908 37522 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 5810 28704 5816 28756
rect 5868 28744 5874 28756
rect 10413 28747 10471 28753
rect 5868 28716 9444 28744
rect 5868 28704 5874 28716
rect 9416 28676 9444 28716
rect 10413 28713 10425 28747
rect 10459 28744 10471 28747
rect 12437 28747 12495 28753
rect 12437 28744 12449 28747
rect 10459 28716 12449 28744
rect 10459 28713 10471 28716
rect 10413 28707 10471 28713
rect 12437 28713 12449 28716
rect 12483 28713 12495 28747
rect 14366 28744 14372 28756
rect 12437 28707 12495 28713
rect 13372 28716 14372 28744
rect 10594 28676 10600 28688
rect 9416 28648 10600 28676
rect 7098 28500 7104 28552
rect 7156 28540 7162 28552
rect 7193 28543 7251 28549
rect 7193 28540 7205 28543
rect 7156 28512 7205 28540
rect 7156 28500 7162 28512
rect 7193 28509 7205 28512
rect 7239 28509 7251 28543
rect 7193 28503 7251 28509
rect 9306 28500 9312 28552
rect 9364 28500 9370 28552
rect 9416 28549 9444 28648
rect 10594 28636 10600 28648
rect 10652 28636 10658 28688
rect 10686 28636 10692 28688
rect 10744 28636 10750 28688
rect 9766 28608 9772 28620
rect 9600 28580 9772 28608
rect 9600 28549 9628 28580
rect 9766 28568 9772 28580
rect 9824 28568 9830 28620
rect 11425 28611 11483 28617
rect 11425 28608 11437 28611
rect 9968 28580 11437 28608
rect 9401 28543 9459 28549
rect 9401 28509 9413 28543
rect 9447 28509 9459 28543
rect 9401 28503 9459 28509
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28509 9643 28543
rect 9585 28503 9643 28509
rect 9677 28543 9735 28549
rect 9677 28509 9689 28543
rect 9723 28540 9735 28543
rect 9858 28540 9864 28552
rect 9723 28512 9864 28540
rect 9723 28509 9735 28512
rect 9677 28503 9735 28509
rect 9858 28500 9864 28512
rect 9916 28500 9922 28552
rect 7460 28475 7518 28481
rect 7460 28441 7472 28475
rect 7506 28472 7518 28475
rect 8018 28472 8024 28484
rect 7506 28444 8024 28472
rect 7506 28441 7518 28444
rect 7460 28435 7518 28441
rect 8018 28432 8024 28444
rect 8076 28432 8082 28484
rect 9766 28432 9772 28484
rect 9824 28472 9830 28484
rect 9968 28472 9996 28580
rect 11425 28577 11437 28580
rect 11471 28608 11483 28611
rect 12526 28608 12532 28620
rect 11471 28580 12532 28608
rect 11471 28577 11483 28580
rect 11425 28571 11483 28577
rect 12526 28568 12532 28580
rect 12584 28568 12590 28620
rect 12621 28611 12679 28617
rect 12621 28577 12633 28611
rect 12667 28608 12679 28611
rect 13372 28608 13400 28716
rect 14366 28704 14372 28716
rect 14424 28704 14430 28756
rect 15010 28704 15016 28756
rect 15068 28744 15074 28756
rect 18874 28744 18880 28756
rect 15068 28716 18880 28744
rect 15068 28704 15074 28716
rect 18874 28704 18880 28716
rect 18932 28704 18938 28756
rect 20073 28747 20131 28753
rect 20073 28713 20085 28747
rect 20119 28744 20131 28747
rect 24210 28744 24216 28756
rect 20119 28716 24216 28744
rect 20119 28713 20131 28716
rect 20073 28707 20131 28713
rect 24210 28704 24216 28716
rect 24268 28704 24274 28756
rect 24302 28704 24308 28756
rect 24360 28744 24366 28756
rect 26050 28744 26056 28756
rect 24360 28716 26056 28744
rect 24360 28704 24366 28716
rect 26050 28704 26056 28716
rect 26108 28704 26114 28756
rect 26145 28747 26203 28753
rect 26145 28713 26157 28747
rect 26191 28713 26203 28747
rect 26145 28707 26203 28713
rect 15194 28676 15200 28688
rect 12667 28580 13400 28608
rect 13464 28648 15200 28676
rect 12667 28577 12679 28580
rect 12621 28571 12679 28577
rect 10042 28500 10048 28552
rect 10100 28540 10106 28552
rect 10597 28543 10655 28549
rect 10597 28540 10609 28543
rect 10100 28512 10609 28540
rect 10100 28500 10106 28512
rect 10597 28509 10609 28512
rect 10643 28509 10655 28543
rect 10597 28503 10655 28509
rect 9824 28444 9996 28472
rect 9824 28432 9830 28444
rect 8386 28364 8392 28416
rect 8444 28404 8450 28416
rect 8573 28407 8631 28413
rect 8573 28404 8585 28407
rect 8444 28376 8585 28404
rect 8444 28364 8450 28376
rect 8573 28373 8585 28376
rect 8619 28373 8631 28407
rect 8573 28367 8631 28373
rect 9122 28364 9128 28416
rect 9180 28364 9186 28416
rect 10612 28404 10640 28503
rect 10778 28500 10784 28552
rect 10836 28500 10842 28552
rect 10873 28543 10931 28549
rect 10873 28509 10885 28543
rect 10919 28540 10931 28543
rect 10962 28540 10968 28552
rect 10919 28512 10968 28540
rect 10919 28509 10931 28512
rect 10873 28503 10931 28509
rect 10962 28500 10968 28512
rect 11020 28500 11026 28552
rect 11514 28540 11520 28552
rect 11072 28512 11520 28540
rect 10686 28432 10692 28484
rect 10744 28472 10750 28484
rect 11072 28472 11100 28512
rect 11514 28500 11520 28512
rect 11572 28540 11578 28552
rect 11609 28543 11667 28549
rect 11609 28540 11621 28543
rect 11572 28512 11621 28540
rect 11572 28500 11578 28512
rect 11609 28509 11621 28512
rect 11655 28509 11667 28543
rect 11609 28503 11667 28509
rect 11701 28543 11759 28549
rect 11701 28509 11713 28543
rect 11747 28540 11759 28543
rect 12250 28540 12256 28552
rect 11747 28512 12256 28540
rect 11747 28509 11759 28512
rect 11701 28503 11759 28509
rect 12250 28500 12256 28512
rect 12308 28500 12314 28552
rect 12342 28500 12348 28552
rect 12400 28540 12406 28552
rect 12437 28543 12495 28549
rect 12437 28540 12449 28543
rect 12400 28512 12449 28540
rect 12400 28500 12406 28512
rect 12437 28509 12449 28512
rect 12483 28509 12495 28543
rect 12437 28503 12495 28509
rect 12710 28500 12716 28552
rect 12768 28500 12774 28552
rect 13464 28549 13492 28648
rect 15194 28636 15200 28648
rect 15252 28636 15258 28688
rect 17034 28636 17040 28688
rect 17092 28636 17098 28688
rect 17678 28636 17684 28688
rect 17736 28676 17742 28688
rect 21726 28676 21732 28688
rect 17736 28648 21732 28676
rect 17736 28636 17742 28648
rect 21726 28636 21732 28648
rect 21784 28676 21790 28688
rect 24578 28676 24584 28688
rect 21784 28648 24584 28676
rect 21784 28636 21790 28648
rect 24578 28636 24584 28648
rect 24636 28636 24642 28688
rect 26160 28676 26188 28707
rect 26970 28704 26976 28756
rect 27028 28704 27034 28756
rect 27062 28704 27068 28756
rect 27120 28704 27126 28756
rect 30374 28744 30380 28756
rect 28368 28716 30380 28744
rect 27798 28676 27804 28688
rect 26160 28648 27804 28676
rect 27798 28636 27804 28648
rect 27856 28636 27862 28688
rect 15646 28611 15704 28617
rect 15646 28608 15658 28611
rect 15304 28580 15658 28608
rect 13449 28543 13507 28549
rect 13449 28509 13461 28543
rect 13495 28509 13507 28543
rect 13449 28503 13507 28509
rect 13541 28543 13599 28549
rect 13541 28509 13553 28543
rect 13587 28540 13599 28543
rect 14182 28540 14188 28552
rect 13587 28512 14188 28540
rect 13587 28509 13599 28512
rect 13541 28503 13599 28509
rect 14182 28500 14188 28512
rect 14240 28500 14246 28552
rect 14274 28500 14280 28552
rect 14332 28500 14338 28552
rect 15304 28484 15332 28580
rect 15646 28577 15658 28580
rect 15692 28577 15704 28611
rect 15646 28571 15704 28577
rect 18138 28568 18144 28620
rect 18196 28568 18202 28620
rect 19889 28611 19947 28617
rect 19889 28577 19901 28611
rect 19935 28608 19947 28611
rect 19978 28608 19984 28620
rect 19935 28580 19984 28608
rect 19935 28577 19947 28580
rect 19889 28571 19947 28577
rect 19978 28568 19984 28580
rect 20036 28568 20042 28620
rect 21818 28568 21824 28620
rect 21876 28608 21882 28620
rect 21913 28611 21971 28617
rect 21913 28608 21925 28611
rect 21876 28580 21925 28608
rect 21876 28568 21882 28580
rect 21913 28577 21925 28580
rect 21959 28577 21971 28611
rect 23937 28611 23995 28617
rect 23937 28608 23949 28611
rect 21913 28571 21971 28577
rect 22020 28580 23949 28608
rect 15930 28549 15936 28552
rect 15924 28540 15936 28549
rect 15891 28512 15936 28540
rect 15924 28503 15936 28512
rect 15930 28500 15936 28503
rect 15988 28500 15994 28552
rect 17862 28500 17868 28552
rect 17920 28540 17926 28552
rect 17957 28543 18015 28549
rect 17957 28540 17969 28543
rect 17920 28512 17969 28540
rect 17920 28500 17926 28512
rect 17957 28509 17969 28512
rect 18003 28509 18015 28543
rect 17957 28503 18015 28509
rect 18230 28500 18236 28552
rect 18288 28540 18294 28552
rect 18693 28543 18751 28549
rect 18693 28540 18705 28543
rect 18288 28512 18705 28540
rect 18288 28500 18294 28512
rect 18693 28509 18705 28512
rect 18739 28509 18751 28543
rect 18693 28503 18751 28509
rect 18874 28500 18880 28552
rect 18932 28540 18938 28552
rect 19797 28543 19855 28549
rect 19797 28540 19809 28543
rect 18932 28512 19809 28540
rect 18932 28500 18938 28512
rect 19797 28509 19809 28512
rect 19843 28509 19855 28543
rect 19797 28503 19855 28509
rect 20901 28543 20959 28549
rect 20901 28509 20913 28543
rect 20947 28540 20959 28543
rect 21082 28540 21088 28552
rect 20947 28512 21088 28540
rect 20947 28509 20959 28512
rect 20901 28503 20959 28509
rect 21082 28500 21088 28512
rect 21140 28500 21146 28552
rect 21177 28543 21235 28549
rect 21177 28509 21189 28543
rect 21223 28540 21235 28543
rect 21223 28512 21680 28540
rect 21223 28509 21235 28512
rect 21177 28503 21235 28509
rect 10744 28444 11100 28472
rect 10744 28432 10750 28444
rect 11422 28432 11428 28484
rect 11480 28472 11486 28484
rect 11793 28475 11851 28481
rect 11793 28472 11805 28475
rect 11480 28444 11805 28472
rect 11480 28432 11486 28444
rect 11716 28416 11744 28444
rect 11793 28441 11805 28444
rect 11839 28441 11851 28475
rect 11793 28435 11851 28441
rect 11977 28475 12035 28481
rect 11977 28441 11989 28475
rect 12023 28472 12035 28475
rect 12802 28472 12808 28484
rect 12023 28444 12808 28472
rect 12023 28441 12035 28444
rect 11977 28435 12035 28441
rect 12802 28432 12808 28444
rect 12860 28432 12866 28484
rect 13722 28432 13728 28484
rect 13780 28432 13786 28484
rect 15105 28475 15163 28481
rect 15105 28441 15117 28475
rect 15151 28472 15163 28475
rect 15286 28472 15292 28484
rect 15151 28444 15292 28472
rect 15151 28441 15163 28444
rect 15105 28435 15163 28441
rect 15286 28432 15292 28444
rect 15344 28432 15350 28484
rect 16114 28432 16120 28484
rect 16172 28472 16178 28484
rect 20625 28475 20683 28481
rect 20625 28472 20637 28475
rect 16172 28444 20637 28472
rect 16172 28432 16178 28444
rect 20625 28441 20637 28444
rect 20671 28441 20683 28475
rect 20625 28435 20683 28441
rect 20993 28475 21051 28481
rect 20993 28441 21005 28475
rect 21039 28472 21051 28475
rect 21652 28472 21680 28512
rect 21726 28500 21732 28552
rect 21784 28540 21790 28552
rect 22020 28540 22048 28580
rect 23937 28577 23949 28580
rect 23983 28577 23995 28611
rect 23937 28571 23995 28577
rect 24026 28568 24032 28620
rect 24084 28608 24090 28620
rect 26053 28611 26111 28617
rect 24084 28580 25544 28608
rect 24084 28568 24090 28580
rect 21784 28512 22048 28540
rect 21784 28500 21790 28512
rect 22186 28500 22192 28552
rect 22244 28500 22250 28552
rect 22465 28543 22523 28549
rect 22465 28509 22477 28543
rect 22511 28509 22523 28543
rect 22465 28503 22523 28509
rect 22480 28472 22508 28503
rect 22646 28500 22652 28552
rect 22704 28500 22710 28552
rect 22922 28500 22928 28552
rect 22980 28500 22986 28552
rect 23842 28500 23848 28552
rect 23900 28500 23906 28552
rect 24578 28500 24584 28552
rect 24636 28500 24642 28552
rect 25133 28543 25191 28549
rect 25133 28509 25145 28543
rect 25179 28540 25191 28543
rect 25406 28540 25412 28552
rect 25179 28512 25412 28540
rect 25179 28509 25191 28512
rect 25133 28503 25191 28509
rect 25406 28500 25412 28512
rect 25464 28500 25470 28552
rect 25516 28540 25544 28580
rect 26053 28577 26065 28611
rect 26099 28608 26111 28611
rect 26234 28608 26240 28620
rect 26099 28580 26240 28608
rect 26099 28577 26111 28580
rect 26053 28571 26111 28577
rect 26234 28568 26240 28580
rect 26292 28568 26298 28620
rect 26418 28568 26424 28620
rect 26476 28608 26482 28620
rect 26973 28611 27031 28617
rect 26973 28608 26985 28611
rect 26476 28580 26985 28608
rect 26476 28568 26482 28580
rect 26973 28577 26985 28580
rect 27019 28608 27031 28611
rect 28258 28608 28264 28620
rect 27019 28580 28264 28608
rect 27019 28577 27031 28580
rect 26973 28571 27031 28577
rect 28258 28568 28264 28580
rect 28316 28568 28322 28620
rect 25516 28512 26004 28540
rect 21039 28444 21588 28472
rect 21652 28444 22508 28472
rect 21039 28441 21051 28444
rect 20993 28435 21051 28441
rect 11054 28404 11060 28416
rect 10612 28376 11060 28404
rect 11054 28364 11060 28376
rect 11112 28364 11118 28416
rect 11698 28364 11704 28416
rect 11756 28364 11762 28416
rect 12342 28364 12348 28416
rect 12400 28404 12406 28416
rect 12897 28407 12955 28413
rect 12897 28404 12909 28407
rect 12400 28376 12909 28404
rect 12400 28364 12406 28376
rect 12897 28373 12909 28376
rect 12943 28373 12955 28407
rect 12897 28367 12955 28373
rect 13446 28364 13452 28416
rect 13504 28364 13510 28416
rect 13538 28364 13544 28416
rect 13596 28404 13602 28416
rect 16574 28404 16580 28416
rect 13596 28376 16580 28404
rect 13596 28364 13602 28376
rect 16574 28364 16580 28376
rect 16632 28364 16638 28416
rect 17494 28364 17500 28416
rect 17552 28364 17558 28416
rect 17586 28364 17592 28416
rect 17644 28404 17650 28416
rect 17865 28407 17923 28413
rect 17865 28404 17877 28407
rect 17644 28376 17877 28404
rect 17644 28364 17650 28376
rect 17865 28373 17877 28376
rect 17911 28373 17923 28407
rect 17865 28367 17923 28373
rect 18785 28407 18843 28413
rect 18785 28373 18797 28407
rect 18831 28404 18843 28407
rect 20530 28404 20536 28416
rect 18831 28376 20536 28404
rect 18831 28373 18843 28376
rect 18785 28367 18843 28373
rect 20530 28364 20536 28376
rect 20588 28364 20594 28416
rect 20806 28364 20812 28416
rect 20864 28404 20870 28416
rect 21450 28404 21456 28416
rect 20864 28376 21456 28404
rect 20864 28364 20870 28376
rect 21450 28364 21456 28376
rect 21508 28364 21514 28416
rect 21560 28404 21588 28444
rect 22554 28432 22560 28484
rect 22612 28472 22618 28484
rect 22940 28472 22968 28500
rect 22612 28444 22968 28472
rect 22612 28432 22618 28444
rect 23382 28432 23388 28484
rect 23440 28432 23446 28484
rect 23474 28432 23480 28484
rect 23532 28472 23538 28484
rect 24762 28472 24768 28484
rect 23532 28444 24768 28472
rect 23532 28432 23538 28444
rect 24762 28432 24768 28444
rect 24820 28472 24826 28484
rect 25682 28472 25688 28484
rect 24820 28444 25688 28472
rect 24820 28432 24826 28444
rect 25682 28432 25688 28444
rect 25740 28432 25746 28484
rect 25866 28432 25872 28484
rect 25924 28432 25930 28484
rect 25976 28472 26004 28512
rect 26142 28500 26148 28552
rect 26200 28500 26206 28552
rect 27154 28500 27160 28552
rect 27212 28540 27218 28552
rect 27522 28540 27528 28552
rect 27212 28512 27528 28540
rect 27212 28500 27218 28512
rect 27522 28500 27528 28512
rect 27580 28500 27586 28552
rect 28368 28540 28396 28716
rect 30374 28704 30380 28716
rect 30432 28704 30438 28756
rect 30837 28747 30895 28753
rect 30837 28713 30849 28747
rect 30883 28744 30895 28747
rect 31018 28744 31024 28756
rect 30883 28716 31024 28744
rect 30883 28713 30895 28716
rect 30837 28707 30895 28713
rect 31018 28704 31024 28716
rect 31076 28704 31082 28756
rect 31478 28704 31484 28756
rect 31536 28744 31542 28756
rect 33042 28744 33048 28756
rect 31536 28716 33048 28744
rect 31536 28704 31542 28716
rect 33042 28704 33048 28716
rect 33100 28704 33106 28756
rect 33502 28704 33508 28756
rect 33560 28744 33566 28756
rect 33870 28744 33876 28756
rect 33560 28716 33876 28744
rect 33560 28704 33566 28716
rect 33870 28704 33876 28716
rect 33928 28704 33934 28756
rect 36078 28744 36084 28756
rect 33980 28716 36084 28744
rect 32950 28676 32956 28688
rect 28828 28648 32956 28676
rect 28828 28549 28856 28648
rect 32950 28636 32956 28648
rect 33008 28636 33014 28688
rect 33686 28636 33692 28688
rect 33744 28676 33750 28688
rect 33980 28676 34008 28716
rect 36078 28704 36084 28716
rect 36136 28744 36142 28756
rect 36265 28747 36323 28753
rect 36265 28744 36277 28747
rect 36136 28716 36277 28744
rect 36136 28704 36142 28716
rect 36265 28713 36277 28716
rect 36311 28713 36323 28747
rect 36265 28707 36323 28713
rect 38194 28704 38200 28756
rect 38252 28704 38258 28756
rect 33744 28648 34008 28676
rect 33744 28636 33750 28648
rect 29178 28568 29184 28620
rect 29236 28568 29242 28620
rect 29270 28568 29276 28620
rect 29328 28608 29334 28620
rect 31294 28608 31300 28620
rect 29328 28580 31300 28608
rect 29328 28568 29334 28580
rect 31294 28568 31300 28580
rect 31352 28568 31358 28620
rect 32033 28611 32091 28617
rect 32033 28608 32045 28611
rect 31404 28580 32045 28608
rect 27908 28512 28396 28540
rect 28629 28543 28687 28549
rect 26789 28475 26847 28481
rect 26789 28472 26801 28475
rect 25976 28444 26801 28472
rect 26789 28441 26801 28444
rect 26835 28441 26847 28475
rect 26789 28435 26847 28441
rect 27709 28475 27767 28481
rect 27709 28441 27721 28475
rect 27755 28472 27767 28475
rect 27798 28472 27804 28484
rect 27755 28444 27804 28472
rect 27755 28441 27767 28444
rect 27709 28435 27767 28441
rect 27798 28432 27804 28444
rect 27856 28432 27862 28484
rect 21634 28404 21640 28416
rect 21560 28376 21640 28404
rect 21634 28364 21640 28376
rect 21692 28364 21698 28416
rect 23566 28364 23572 28416
rect 23624 28404 23630 28416
rect 24673 28407 24731 28413
rect 24673 28404 24685 28407
rect 23624 28376 24685 28404
rect 23624 28364 23630 28376
rect 24673 28373 24685 28376
rect 24719 28373 24731 28407
rect 24673 28367 24731 28373
rect 25406 28364 25412 28416
rect 25464 28404 25470 28416
rect 25958 28404 25964 28416
rect 25464 28376 25964 28404
rect 25464 28364 25470 28376
rect 25958 28364 25964 28376
rect 26016 28364 26022 28416
rect 26329 28407 26387 28413
rect 26329 28373 26341 28407
rect 26375 28404 26387 28407
rect 27908 28404 27936 28512
rect 28629 28509 28641 28543
rect 28675 28509 28687 28543
rect 28629 28503 28687 28509
rect 28813 28543 28871 28549
rect 28813 28509 28825 28543
rect 28859 28509 28871 28543
rect 28813 28503 28871 28509
rect 30285 28543 30343 28549
rect 30285 28509 30297 28543
rect 30331 28540 30343 28543
rect 30374 28540 30380 28552
rect 30331 28512 30380 28540
rect 30331 28509 30343 28512
rect 30285 28503 30343 28509
rect 28644 28472 28672 28503
rect 30374 28500 30380 28512
rect 30432 28500 30438 28552
rect 30650 28500 30656 28552
rect 30708 28540 30714 28552
rect 31404 28540 31432 28580
rect 32033 28577 32045 28580
rect 32079 28577 32091 28611
rect 32033 28571 32091 28577
rect 34882 28568 34888 28620
rect 34940 28568 34946 28620
rect 30708 28512 31432 28540
rect 31573 28543 31631 28549
rect 30708 28500 30714 28512
rect 31573 28509 31585 28543
rect 31619 28509 31631 28543
rect 31573 28503 31631 28509
rect 28902 28472 28908 28484
rect 28644 28444 28908 28472
rect 28902 28432 28908 28444
rect 28960 28432 28966 28484
rect 29089 28475 29147 28481
rect 29089 28441 29101 28475
rect 29135 28472 29147 28475
rect 31588 28472 31616 28503
rect 31662 28500 31668 28552
rect 31720 28540 31726 28552
rect 33413 28543 33471 28549
rect 33413 28540 33425 28543
rect 31720 28512 33425 28540
rect 31720 28500 31726 28512
rect 33413 28509 33425 28512
rect 33459 28509 33471 28543
rect 33413 28503 33471 28509
rect 33686 28500 33692 28552
rect 33744 28540 33750 28552
rect 33965 28543 34023 28549
rect 33965 28540 33977 28543
rect 33744 28512 33977 28540
rect 33744 28500 33750 28512
rect 33965 28509 33977 28512
rect 34011 28509 34023 28543
rect 34900 28540 34928 28568
rect 36817 28543 36875 28549
rect 36817 28540 36829 28543
rect 34900 28512 36829 28540
rect 33965 28503 34023 28509
rect 36817 28509 36829 28512
rect 36863 28509 36875 28543
rect 36817 28503 36875 28509
rect 37084 28543 37142 28549
rect 37084 28509 37096 28543
rect 37130 28540 37142 28543
rect 37458 28540 37464 28552
rect 37130 28512 37464 28540
rect 37130 28509 37142 28512
rect 37084 28503 37142 28509
rect 37458 28500 37464 28512
rect 37516 28500 37522 28552
rect 29135 28444 31616 28472
rect 29135 28441 29147 28444
rect 29089 28435 29147 28441
rect 32674 28432 32680 28484
rect 32732 28472 32738 28484
rect 35152 28475 35210 28481
rect 32732 28444 34376 28472
rect 32732 28432 32738 28444
rect 26375 28376 27936 28404
rect 27985 28407 28043 28413
rect 26375 28373 26387 28376
rect 26329 28367 26387 28373
rect 27985 28373 27997 28407
rect 28031 28404 28043 28407
rect 28810 28404 28816 28416
rect 28031 28376 28816 28404
rect 28031 28373 28043 28376
rect 27985 28367 28043 28373
rect 28810 28364 28816 28376
rect 28868 28364 28874 28416
rect 31018 28364 31024 28416
rect 31076 28404 31082 28416
rect 33686 28404 33692 28416
rect 31076 28376 33692 28404
rect 31076 28364 31082 28376
rect 33686 28364 33692 28376
rect 33744 28404 33750 28416
rect 34238 28404 34244 28416
rect 33744 28376 34244 28404
rect 33744 28364 33750 28376
rect 34238 28364 34244 28376
rect 34296 28364 34302 28416
rect 34348 28404 34376 28444
rect 35152 28441 35164 28475
rect 35198 28472 35210 28475
rect 38378 28472 38384 28484
rect 35198 28444 38384 28472
rect 35198 28441 35210 28444
rect 35152 28435 35210 28441
rect 38378 28432 38384 28444
rect 38436 28432 38442 28484
rect 35710 28404 35716 28416
rect 34348 28376 35716 28404
rect 35710 28364 35716 28376
rect 35768 28364 35774 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 8018 28160 8024 28212
rect 8076 28160 8082 28212
rect 8481 28203 8539 28209
rect 8481 28169 8493 28203
rect 8527 28200 8539 28203
rect 9122 28200 9128 28212
rect 8527 28172 9128 28200
rect 8527 28169 8539 28172
rect 8481 28163 8539 28169
rect 9122 28160 9128 28172
rect 9180 28160 9186 28212
rect 9953 28203 10011 28209
rect 9953 28169 9965 28203
rect 9999 28200 10011 28203
rect 10134 28200 10140 28212
rect 9999 28172 10140 28200
rect 9999 28169 10011 28172
rect 9953 28163 10011 28169
rect 10134 28160 10140 28172
rect 10192 28160 10198 28212
rect 10689 28203 10747 28209
rect 10689 28169 10701 28203
rect 10735 28200 10747 28203
rect 10778 28200 10784 28212
rect 10735 28172 10784 28200
rect 10735 28169 10747 28172
rect 10689 28163 10747 28169
rect 10778 28160 10784 28172
rect 10836 28160 10842 28212
rect 11793 28203 11851 28209
rect 11793 28169 11805 28203
rect 11839 28200 11851 28203
rect 12710 28200 12716 28212
rect 11839 28172 12716 28200
rect 11839 28169 11851 28172
rect 11793 28163 11851 28169
rect 12710 28160 12716 28172
rect 12768 28160 12774 28212
rect 17865 28203 17923 28209
rect 14752 28172 17816 28200
rect 8294 28092 8300 28144
rect 8352 28132 8358 28144
rect 10502 28132 10508 28144
rect 8352 28104 8708 28132
rect 8352 28092 8358 28104
rect 8386 28024 8392 28076
rect 8444 28024 8450 28076
rect 8478 27956 8484 28008
rect 8536 27996 8542 28008
rect 8573 27999 8631 28005
rect 8573 27996 8585 27999
rect 8536 27968 8585 27996
rect 8536 27956 8542 27968
rect 8573 27965 8585 27968
rect 8619 27965 8631 27999
rect 8680 27996 8708 28104
rect 9784 28104 10508 28132
rect 9784 28073 9812 28104
rect 10502 28092 10508 28104
rect 10560 28092 10566 28144
rect 14182 28132 14188 28144
rect 10796 28104 11192 28132
rect 9769 28067 9827 28073
rect 9769 28033 9781 28067
rect 9815 28033 9827 28067
rect 9769 28027 9827 28033
rect 10042 28024 10048 28076
rect 10100 28064 10106 28076
rect 10796 28064 10824 28104
rect 10100 28036 10824 28064
rect 10100 28024 10106 28036
rect 10870 28024 10876 28076
rect 10928 28024 10934 28076
rect 11164 28073 11192 28104
rect 12176 28104 14188 28132
rect 12176 28076 12204 28104
rect 14182 28092 14188 28104
rect 14240 28092 14246 28144
rect 12066 28073 12072 28076
rect 11057 28067 11115 28073
rect 11057 28033 11069 28067
rect 11103 28033 11115 28067
rect 11057 28027 11115 28033
rect 11149 28067 11207 28073
rect 11149 28033 11161 28067
rect 11195 28033 11207 28067
rect 11149 28027 11207 28033
rect 12049 28067 12072 28073
rect 12049 28033 12061 28067
rect 12049 28027 12072 28033
rect 10134 27996 10140 28008
rect 8680 27968 10140 27996
rect 8573 27959 8631 27965
rect 10134 27956 10140 27968
rect 10192 27956 10198 28008
rect 10686 27956 10692 28008
rect 10744 27996 10750 28008
rect 11072 27996 11100 28027
rect 12066 28024 12072 28027
rect 12124 28024 12130 28076
rect 12158 28024 12164 28076
rect 12216 28024 12222 28076
rect 12250 28024 12256 28076
rect 12308 28024 12314 28076
rect 12434 28024 12440 28076
rect 12492 28024 12498 28076
rect 13170 28073 13176 28076
rect 13164 28027 13176 28073
rect 13170 28024 13176 28027
rect 13228 28024 13234 28076
rect 13630 28024 13636 28076
rect 13688 28064 13694 28076
rect 14752 28073 14780 28172
rect 15562 28132 15568 28144
rect 14844 28104 15568 28132
rect 14737 28067 14795 28073
rect 13688 28036 14688 28064
rect 13688 28024 13694 28036
rect 10744 27968 11100 27996
rect 10744 27956 10750 27968
rect 12894 27956 12900 28008
rect 12952 27956 12958 28008
rect 14660 27996 14688 28036
rect 14737 28033 14749 28067
rect 14783 28033 14795 28067
rect 14737 28027 14795 28033
rect 14844 27996 14872 28104
rect 15562 28092 15568 28104
rect 15620 28092 15626 28144
rect 15657 28135 15715 28141
rect 15657 28101 15669 28135
rect 15703 28132 15715 28135
rect 17126 28132 17132 28144
rect 15703 28104 17132 28132
rect 15703 28101 15715 28104
rect 15657 28095 15715 28101
rect 17126 28092 17132 28104
rect 17184 28092 17190 28144
rect 17788 28132 17816 28172
rect 17865 28169 17877 28203
rect 17911 28200 17923 28203
rect 18693 28203 18751 28209
rect 18693 28200 18705 28203
rect 17911 28172 18705 28200
rect 17911 28169 17923 28172
rect 17865 28163 17923 28169
rect 18693 28169 18705 28172
rect 18739 28169 18751 28203
rect 20714 28200 20720 28212
rect 18693 28163 18751 28169
rect 19306 28172 20720 28200
rect 19306 28132 19334 28172
rect 20714 28160 20720 28172
rect 20772 28160 20778 28212
rect 21082 28160 21088 28212
rect 21140 28200 21146 28212
rect 21542 28200 21548 28212
rect 21140 28172 21548 28200
rect 21140 28160 21146 28172
rect 21542 28160 21548 28172
rect 21600 28160 21606 28212
rect 22002 28160 22008 28212
rect 22060 28200 22066 28212
rect 22465 28203 22523 28209
rect 22465 28200 22477 28203
rect 22060 28172 22477 28200
rect 22060 28160 22066 28172
rect 22465 28169 22477 28172
rect 22511 28169 22523 28203
rect 22465 28163 22523 28169
rect 23198 28160 23204 28212
rect 23256 28200 23262 28212
rect 23256 28172 23796 28200
rect 23256 28160 23262 28172
rect 17788 28104 19334 28132
rect 20625 28135 20683 28141
rect 20625 28101 20637 28135
rect 20671 28132 20683 28135
rect 20671 28104 23244 28132
rect 20671 28101 20683 28104
rect 20625 28095 20683 28101
rect 14921 28067 14979 28073
rect 14921 28033 14933 28067
rect 14967 28033 14979 28067
rect 14921 28027 14979 28033
rect 14660 27968 14872 27996
rect 14936 27996 14964 28027
rect 15010 28024 15016 28076
rect 15068 28064 15074 28076
rect 15378 28064 15384 28076
rect 15068 28036 15384 28064
rect 15068 28024 15074 28036
rect 15378 28024 15384 28036
rect 15436 28024 15442 28076
rect 15749 28067 15807 28073
rect 15749 28033 15761 28067
rect 15795 28064 15807 28067
rect 16022 28064 16028 28076
rect 15795 28036 16028 28064
rect 15795 28033 15807 28036
rect 15749 28027 15807 28033
rect 16022 28024 16028 28036
rect 16080 28024 16086 28076
rect 16850 28024 16856 28076
rect 16908 28024 16914 28076
rect 17310 28024 17316 28076
rect 17368 28064 17374 28076
rect 17957 28067 18015 28073
rect 17957 28064 17969 28067
rect 17368 28036 17969 28064
rect 17368 28024 17374 28036
rect 17957 28033 17969 28036
rect 18003 28033 18015 28067
rect 17957 28027 18015 28033
rect 18322 28024 18328 28076
rect 18380 28064 18386 28076
rect 19061 28067 19119 28073
rect 19061 28064 19073 28067
rect 18380 28036 19073 28064
rect 18380 28024 18386 28036
rect 19061 28033 19073 28036
rect 19107 28033 19119 28067
rect 20070 28064 20076 28076
rect 19061 28027 19119 28033
rect 19260 28036 20076 28064
rect 17678 27996 17684 28008
rect 14936 27968 17684 27996
rect 17678 27956 17684 27968
rect 17736 27956 17742 28008
rect 18141 27999 18199 28005
rect 18141 27965 18153 27999
rect 18187 27996 18199 27999
rect 18874 27996 18880 28008
rect 18187 27968 18880 27996
rect 18187 27965 18199 27968
rect 18141 27959 18199 27965
rect 18874 27956 18880 27968
rect 18932 27956 18938 28008
rect 19150 27956 19156 28008
rect 19208 27956 19214 28008
rect 19260 28005 19288 28036
rect 20070 28024 20076 28036
rect 20128 28024 20134 28076
rect 20257 28067 20315 28073
rect 20257 28033 20269 28067
rect 20303 28033 20315 28067
rect 20257 28027 20315 28033
rect 20441 28067 20499 28073
rect 20441 28033 20453 28067
rect 20487 28064 20499 28067
rect 21082 28064 21088 28076
rect 20487 28036 21088 28064
rect 20487 28033 20499 28036
rect 20441 28027 20499 28033
rect 19245 27999 19303 28005
rect 19245 27965 19257 27999
rect 19291 27965 19303 27999
rect 19245 27959 19303 27965
rect 19518 27956 19524 28008
rect 19576 27996 19582 28008
rect 20272 27996 20300 28027
rect 21082 28024 21088 28036
rect 21140 28024 21146 28076
rect 21269 28067 21327 28073
rect 21269 28033 21281 28067
rect 21315 28033 21327 28067
rect 21269 28027 21327 28033
rect 21284 27996 21312 28027
rect 21358 28024 21364 28076
rect 21416 28064 21422 28076
rect 22373 28067 22431 28073
rect 22373 28064 22385 28067
rect 21416 28036 22385 28064
rect 21416 28024 21422 28036
rect 22373 28033 22385 28036
rect 22419 28064 22431 28067
rect 22922 28064 22928 28076
rect 22419 28036 22928 28064
rect 22419 28033 22431 28036
rect 22373 28027 22431 28033
rect 22922 28024 22928 28036
rect 22980 28024 22986 28076
rect 22094 27996 22100 28008
rect 19576 27968 22100 27996
rect 19576 27956 19582 27968
rect 22094 27956 22100 27968
rect 22152 27956 22158 28008
rect 22649 27999 22707 28005
rect 22649 27965 22661 27999
rect 22695 27996 22707 27999
rect 22738 27996 22744 28008
rect 22695 27968 22744 27996
rect 22695 27965 22707 27968
rect 22649 27959 22707 27965
rect 7558 27888 7564 27940
rect 7616 27928 7622 27940
rect 9766 27928 9772 27940
rect 7616 27900 9772 27928
rect 7616 27888 7622 27900
rect 9766 27888 9772 27900
rect 9824 27888 9830 27940
rect 10042 27888 10048 27940
rect 10100 27928 10106 27940
rect 12526 27928 12532 27940
rect 10100 27900 12532 27928
rect 10100 27888 10106 27900
rect 12526 27888 12532 27900
rect 12584 27888 12590 27940
rect 14090 27888 14096 27940
rect 14148 27928 14154 27940
rect 14277 27931 14335 27937
rect 14277 27928 14289 27931
rect 14148 27900 14289 27928
rect 14148 27888 14154 27900
rect 14277 27897 14289 27900
rect 14323 27928 14335 27931
rect 16850 27928 16856 27940
rect 14323 27900 16856 27928
rect 14323 27897 14335 27900
rect 14277 27891 14335 27897
rect 16850 27888 16856 27900
rect 16908 27888 16914 27940
rect 16945 27931 17003 27937
rect 16945 27897 16957 27931
rect 16991 27928 17003 27931
rect 19886 27928 19892 27940
rect 16991 27900 19892 27928
rect 16991 27897 17003 27900
rect 16945 27891 17003 27897
rect 19886 27888 19892 27900
rect 19944 27888 19950 27940
rect 21358 27888 21364 27940
rect 21416 27888 21422 27940
rect 22664 27928 22692 27959
rect 22738 27956 22744 27968
rect 22796 27956 22802 28008
rect 23216 27996 23244 28104
rect 23290 28092 23296 28144
rect 23348 28132 23354 28144
rect 23348 28104 23704 28132
rect 23348 28092 23354 28104
rect 23385 28067 23443 28073
rect 23385 28033 23397 28067
rect 23431 28064 23443 28067
rect 23474 28064 23480 28076
rect 23431 28036 23480 28064
rect 23431 28033 23443 28036
rect 23385 28027 23443 28033
rect 23474 28024 23480 28036
rect 23532 28024 23538 28076
rect 23566 28024 23572 28076
rect 23624 28024 23630 28076
rect 23676 28073 23704 28104
rect 23661 28067 23719 28073
rect 23661 28033 23673 28067
rect 23707 28033 23719 28067
rect 23768 28064 23796 28172
rect 24118 28160 24124 28212
rect 24176 28200 24182 28212
rect 25590 28200 25596 28212
rect 24176 28172 25596 28200
rect 24176 28160 24182 28172
rect 25590 28160 25596 28172
rect 25648 28160 25654 28212
rect 27522 28200 27528 28212
rect 27264 28172 27528 28200
rect 23842 28092 23848 28144
rect 23900 28132 23906 28144
rect 23900 28104 25728 28132
rect 23900 28092 23906 28104
rect 24673 28067 24731 28073
rect 24673 28064 24685 28067
rect 23768 28036 24685 28064
rect 23661 28027 23719 28033
rect 24673 28033 24685 28036
rect 24719 28064 24731 28067
rect 24854 28064 24860 28076
rect 24719 28036 24860 28064
rect 24719 28033 24731 28036
rect 24673 28027 24731 28033
rect 24854 28024 24860 28036
rect 24912 28024 24918 28076
rect 24949 28067 25007 28073
rect 24949 28033 24961 28067
rect 24995 28064 25007 28067
rect 25314 28064 25320 28076
rect 24995 28036 25320 28064
rect 24995 28033 25007 28036
rect 24949 28027 25007 28033
rect 25314 28024 25320 28036
rect 25372 28024 25378 28076
rect 25406 28024 25412 28076
rect 25464 28024 25470 28076
rect 25700 28073 25728 28104
rect 26050 28092 26056 28144
rect 26108 28132 26114 28144
rect 27264 28132 27292 28172
rect 27522 28160 27528 28172
rect 27580 28200 27586 28212
rect 28626 28200 28632 28212
rect 27580 28172 28632 28200
rect 27580 28160 27586 28172
rect 28626 28160 28632 28172
rect 28684 28160 28690 28212
rect 30558 28160 30564 28212
rect 30616 28200 30622 28212
rect 30616 28172 34928 28200
rect 30616 28160 30622 28172
rect 26108 28104 27292 28132
rect 26108 28092 26114 28104
rect 25593 28067 25651 28073
rect 25593 28033 25605 28067
rect 25639 28033 25651 28067
rect 25593 28027 25651 28033
rect 25685 28067 25743 28073
rect 25685 28033 25697 28067
rect 25731 28033 25743 28067
rect 25685 28027 25743 28033
rect 25961 28067 26019 28073
rect 25961 28033 25973 28067
rect 26007 28064 26019 28067
rect 27154 28064 27160 28076
rect 26007 28036 27160 28064
rect 26007 28033 26019 28036
rect 25961 28027 26019 28033
rect 25498 27996 25504 28008
rect 23216 27968 25504 27996
rect 25498 27956 25504 27968
rect 25556 27996 25562 28008
rect 25608 27996 25636 28027
rect 27154 28024 27160 28036
rect 27212 28024 27218 28076
rect 27264 28073 27292 28104
rect 28718 28092 28724 28144
rect 28776 28132 28782 28144
rect 31662 28132 31668 28144
rect 28776 28104 31668 28132
rect 28776 28092 28782 28104
rect 31662 28092 31668 28104
rect 31720 28092 31726 28144
rect 31846 28092 31852 28144
rect 31904 28132 31910 28144
rect 33045 28135 33103 28141
rect 33045 28132 33057 28135
rect 31904 28104 33057 28132
rect 31904 28092 31910 28104
rect 33045 28101 33057 28104
rect 33091 28101 33103 28135
rect 34790 28132 34796 28144
rect 33045 28095 33103 28101
rect 33704 28104 34796 28132
rect 27249 28067 27307 28073
rect 27249 28033 27261 28067
rect 27295 28033 27307 28067
rect 27249 28027 27307 28033
rect 28166 28024 28172 28076
rect 28224 28064 28230 28076
rect 28353 28067 28411 28073
rect 28353 28064 28365 28067
rect 28224 28036 28365 28064
rect 28224 28024 28230 28036
rect 28353 28033 28365 28036
rect 28399 28064 28411 28067
rect 28534 28064 28540 28076
rect 28399 28036 28540 28064
rect 28399 28033 28411 28036
rect 28353 28027 28411 28033
rect 28534 28024 28540 28036
rect 28592 28024 28598 28076
rect 28994 28024 29000 28076
rect 29052 28024 29058 28076
rect 29086 28024 29092 28076
rect 29144 28064 29150 28076
rect 29365 28067 29423 28073
rect 29365 28064 29377 28067
rect 29144 28036 29377 28064
rect 29144 28024 29150 28036
rect 29365 28033 29377 28036
rect 29411 28033 29423 28067
rect 29365 28027 29423 28033
rect 29641 28067 29699 28073
rect 29641 28033 29653 28067
rect 29687 28033 29699 28067
rect 29641 28027 29699 28033
rect 25556 27968 25636 27996
rect 25777 27999 25835 28005
rect 25556 27956 25562 27968
rect 25777 27965 25789 27999
rect 25823 27996 25835 27999
rect 26050 27996 26056 28008
rect 25823 27968 26056 27996
rect 25823 27965 25835 27968
rect 25777 27959 25835 27965
rect 21468 27900 22692 27928
rect 9582 27820 9588 27872
rect 9640 27820 9646 27872
rect 10134 27820 10140 27872
rect 10192 27860 10198 27872
rect 12710 27860 12716 27872
rect 10192 27832 12716 27860
rect 10192 27820 10198 27832
rect 12710 27820 12716 27832
rect 12768 27820 12774 27872
rect 14737 27863 14795 27869
rect 14737 27829 14749 27863
rect 14783 27860 14795 27863
rect 15102 27860 15108 27872
rect 14783 27832 15108 27860
rect 14783 27829 14795 27832
rect 14737 27823 14795 27829
rect 15102 27820 15108 27832
rect 15160 27820 15166 27872
rect 15930 27820 15936 27872
rect 15988 27820 15994 27872
rect 17497 27863 17555 27869
rect 17497 27829 17509 27863
rect 17543 27860 17555 27863
rect 18322 27860 18328 27872
rect 17543 27832 18328 27860
rect 17543 27829 17555 27832
rect 17497 27823 17555 27829
rect 18322 27820 18328 27832
rect 18380 27820 18386 27872
rect 18414 27820 18420 27872
rect 18472 27860 18478 27872
rect 18690 27860 18696 27872
rect 18472 27832 18696 27860
rect 18472 27820 18478 27832
rect 18690 27820 18696 27832
rect 18748 27860 18754 27872
rect 21468 27860 21496 27900
rect 23014 27888 23020 27940
rect 23072 27928 23078 27940
rect 23072 27900 23428 27928
rect 23072 27888 23078 27900
rect 18748 27832 21496 27860
rect 18748 27820 18754 27832
rect 22002 27820 22008 27872
rect 22060 27820 22066 27872
rect 23198 27820 23204 27872
rect 23256 27820 23262 27872
rect 23400 27860 23428 27900
rect 23474 27888 23480 27940
rect 23532 27888 23538 27940
rect 24857 27931 24915 27937
rect 24857 27928 24869 27931
rect 23676 27900 24869 27928
rect 23676 27860 23704 27900
rect 24857 27897 24869 27900
rect 24903 27897 24915 27931
rect 24857 27891 24915 27897
rect 25590 27888 25596 27940
rect 25648 27928 25654 27940
rect 25792 27928 25820 27959
rect 26050 27956 26056 27968
rect 26108 27956 26114 28008
rect 26142 27956 26148 28008
rect 26200 27996 26206 28008
rect 27706 27996 27712 28008
rect 26200 27968 27712 27996
rect 26200 27956 26206 27968
rect 27706 27956 27712 27968
rect 27764 27956 27770 28008
rect 27985 27999 28043 28005
rect 27985 27965 27997 27999
rect 28031 27965 28043 27999
rect 27985 27959 28043 27965
rect 28000 27928 28028 27959
rect 28258 27956 28264 28008
rect 28316 27996 28322 28008
rect 29656 27996 29684 28027
rect 30650 28024 30656 28076
rect 30708 28024 30714 28076
rect 31570 28024 31576 28076
rect 31628 28024 31634 28076
rect 32306 28024 32312 28076
rect 32364 28024 32370 28076
rect 33704 28073 33732 28104
rect 34790 28092 34796 28104
rect 34848 28092 34854 28144
rect 33689 28067 33747 28073
rect 33689 28033 33701 28067
rect 33735 28033 33747 28067
rect 33689 28027 33747 28033
rect 33782 28067 33840 28073
rect 33782 28033 33794 28067
rect 33828 28033 33840 28067
rect 33782 28027 33840 28033
rect 28316 27968 29684 27996
rect 28316 27956 28322 27968
rect 30466 27956 30472 28008
rect 30524 27996 30530 28008
rect 30834 27996 30840 28008
rect 30524 27968 30840 27996
rect 30524 27956 30530 27968
rect 30834 27956 30840 27968
rect 30892 27956 30898 28008
rect 31757 27999 31815 28005
rect 31757 27965 31769 27999
rect 31803 27996 31815 27999
rect 32766 27996 32772 28008
rect 31803 27968 32772 27996
rect 31803 27965 31815 27968
rect 31757 27959 31815 27965
rect 32766 27956 32772 27968
rect 32824 27956 32830 28008
rect 33797 27996 33825 28027
rect 33870 28024 33876 28076
rect 33928 28064 33934 28076
rect 33965 28067 34023 28073
rect 33965 28064 33977 28067
rect 33928 28036 33977 28064
rect 33928 28024 33934 28036
rect 33965 28033 33977 28036
rect 34011 28033 34023 28067
rect 33965 28027 34023 28033
rect 34054 28024 34060 28076
rect 34112 28024 34118 28076
rect 34146 28024 34152 28076
rect 34204 28073 34210 28076
rect 34204 28067 34253 28073
rect 34204 28033 34207 28067
rect 34241 28064 34253 28067
rect 34422 28064 34428 28076
rect 34241 28036 34428 28064
rect 34241 28033 34253 28036
rect 34204 28027 34253 28033
rect 34204 28024 34210 28027
rect 34422 28024 34428 28036
rect 34480 28024 34486 28076
rect 34900 28073 34928 28172
rect 35342 28160 35348 28212
rect 35400 28200 35406 28212
rect 36909 28203 36967 28209
rect 36909 28200 36921 28203
rect 35400 28172 36921 28200
rect 35400 28160 35406 28172
rect 36909 28169 36921 28172
rect 36955 28169 36967 28203
rect 36909 28163 36967 28169
rect 35360 28132 35388 28160
rect 34999 28104 35388 28132
rect 35796 28135 35854 28141
rect 34885 28067 34943 28073
rect 34885 28033 34897 28067
rect 34931 28033 34943 28067
rect 34885 28027 34943 28033
rect 34999 27996 35027 28104
rect 35796 28101 35808 28135
rect 35842 28132 35854 28135
rect 37366 28132 37372 28144
rect 35842 28104 37372 28132
rect 35842 28101 35854 28104
rect 35796 28095 35854 28101
rect 37366 28092 37372 28104
rect 37424 28092 37430 28144
rect 35069 28067 35127 28073
rect 35069 28033 35081 28067
rect 35115 28033 35127 28067
rect 35069 28027 35127 28033
rect 33797 27968 35027 27996
rect 25648 27900 25820 27928
rect 26068 27900 28028 27928
rect 29457 27931 29515 27937
rect 25648 27888 25654 27900
rect 23400 27832 23704 27860
rect 24486 27820 24492 27872
rect 24544 27820 24550 27872
rect 24670 27820 24676 27872
rect 24728 27860 24734 27872
rect 26068 27860 26096 27900
rect 29457 27897 29469 27931
rect 29503 27928 29515 27931
rect 33318 27928 33324 27940
rect 29503 27900 33324 27928
rect 29503 27897 29515 27900
rect 29457 27891 29515 27897
rect 33318 27888 33324 27900
rect 33376 27888 33382 27940
rect 35084 27928 35112 28027
rect 35158 28024 35164 28076
rect 35216 28064 35222 28076
rect 35529 28067 35587 28073
rect 35529 28064 35541 28067
rect 35216 28036 35541 28064
rect 35216 28024 35222 28036
rect 35529 28033 35541 28036
rect 35575 28033 35587 28067
rect 35529 28027 35587 28033
rect 37458 28024 37464 28076
rect 37516 28064 37522 28076
rect 37553 28067 37611 28073
rect 37553 28064 37565 28067
rect 37516 28036 37565 28064
rect 37516 28024 37522 28036
rect 37553 28033 37565 28036
rect 37599 28033 37611 28067
rect 37553 28027 37611 28033
rect 38010 27956 38016 28008
rect 38068 27956 38074 28008
rect 33428 27900 35112 27928
rect 24728 27832 26096 27860
rect 24728 27820 24734 27832
rect 26142 27820 26148 27872
rect 26200 27820 26206 27872
rect 26326 27820 26332 27872
rect 26384 27860 26390 27872
rect 29638 27860 29644 27872
rect 26384 27832 29644 27860
rect 26384 27820 26390 27832
rect 29638 27820 29644 27832
rect 29696 27820 29702 27872
rect 29730 27820 29736 27872
rect 29788 27860 29794 27872
rect 33428 27860 33456 27900
rect 29788 27832 33456 27860
rect 29788 27820 29794 27832
rect 33502 27820 33508 27872
rect 33560 27860 33566 27872
rect 34054 27860 34060 27872
rect 33560 27832 34060 27860
rect 33560 27820 33566 27832
rect 34054 27820 34060 27832
rect 34112 27820 34118 27872
rect 34333 27863 34391 27869
rect 34333 27829 34345 27863
rect 34379 27860 34391 27863
rect 34422 27860 34428 27872
rect 34379 27832 34428 27860
rect 34379 27829 34391 27832
rect 34333 27823 34391 27829
rect 34422 27820 34428 27832
rect 34480 27820 34486 27872
rect 34606 27820 34612 27872
rect 34664 27860 34670 27872
rect 34885 27863 34943 27869
rect 34885 27860 34897 27863
rect 34664 27832 34897 27860
rect 34664 27820 34670 27832
rect 34885 27829 34897 27832
rect 34931 27829 34943 27863
rect 34885 27823 34943 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 4706 27616 4712 27668
rect 4764 27656 4770 27668
rect 6914 27656 6920 27668
rect 4764 27628 6920 27656
rect 4764 27616 4770 27628
rect 6914 27616 6920 27628
rect 6972 27616 6978 27668
rect 9125 27659 9183 27665
rect 9125 27625 9137 27659
rect 9171 27656 9183 27659
rect 9306 27656 9312 27668
rect 9171 27628 9312 27656
rect 9171 27625 9183 27628
rect 9125 27619 9183 27625
rect 9306 27616 9312 27628
rect 9364 27616 9370 27668
rect 10042 27616 10048 27668
rect 10100 27616 10106 27668
rect 12250 27656 12256 27668
rect 11624 27628 12256 27656
rect 3510 27548 3516 27600
rect 3568 27588 3574 27600
rect 5350 27588 5356 27600
rect 3568 27560 5356 27588
rect 3568 27548 3574 27560
rect 5350 27548 5356 27560
rect 5408 27548 5414 27600
rect 7098 27480 7104 27532
rect 7156 27480 7162 27532
rect 10686 27520 10692 27532
rect 9692 27492 10692 27520
rect 7116 27452 7144 27480
rect 9692 27464 9720 27492
rect 10686 27480 10692 27492
rect 10744 27520 10750 27532
rect 10744 27492 11008 27520
rect 10744 27480 10750 27492
rect 8202 27452 8208 27464
rect 7116 27424 8208 27452
rect 8202 27412 8208 27424
rect 8260 27412 8266 27464
rect 8570 27412 8576 27464
rect 8628 27452 8634 27464
rect 9125 27455 9183 27461
rect 9125 27452 9137 27455
rect 8628 27424 9137 27452
rect 8628 27412 8634 27424
rect 9125 27421 9137 27424
rect 9171 27421 9183 27455
rect 9125 27415 9183 27421
rect 9309 27455 9367 27461
rect 9309 27421 9321 27455
rect 9355 27452 9367 27455
rect 9674 27452 9680 27464
rect 9355 27424 9680 27452
rect 9355 27421 9367 27424
rect 9309 27415 9367 27421
rect 9674 27412 9680 27424
rect 9732 27412 9738 27464
rect 9953 27455 10011 27461
rect 9953 27421 9965 27455
rect 9999 27421 10011 27455
rect 9953 27415 10011 27421
rect 10781 27455 10839 27461
rect 10781 27421 10793 27455
rect 10827 27452 10839 27455
rect 10870 27452 10876 27464
rect 10827 27424 10876 27452
rect 10827 27421 10839 27424
rect 10781 27415 10839 27421
rect 7368 27387 7426 27393
rect 7368 27353 7380 27387
rect 7414 27384 7426 27387
rect 8018 27384 8024 27396
rect 7414 27356 8024 27384
rect 7414 27353 7426 27356
rect 7368 27347 7426 27353
rect 8018 27344 8024 27356
rect 8076 27344 8082 27396
rect 9968 27384 9996 27415
rect 10870 27412 10876 27424
rect 10928 27412 10934 27464
rect 10980 27461 11008 27492
rect 10965 27455 11023 27461
rect 10965 27421 10977 27455
rect 11011 27421 11023 27455
rect 10965 27415 11023 27421
rect 11054 27412 11060 27464
rect 11112 27452 11118 27464
rect 11624 27452 11652 27628
rect 12250 27616 12256 27628
rect 12308 27656 12314 27668
rect 12308 27628 12572 27656
rect 12308 27616 12314 27628
rect 12066 27548 12072 27600
rect 12124 27548 12130 27600
rect 11698 27480 11704 27532
rect 11756 27520 11762 27532
rect 11885 27523 11943 27529
rect 11885 27520 11897 27523
rect 11756 27492 11897 27520
rect 11756 27480 11762 27492
rect 11885 27489 11897 27492
rect 11931 27489 11943 27523
rect 11885 27483 11943 27489
rect 11977 27523 12035 27529
rect 11977 27489 11989 27523
rect 12023 27520 12035 27523
rect 12084 27520 12112 27548
rect 12023 27492 12112 27520
rect 12161 27523 12219 27529
rect 12023 27489 12035 27492
rect 11977 27483 12035 27489
rect 12161 27489 12173 27523
rect 12207 27520 12219 27523
rect 12342 27520 12348 27532
rect 12207 27492 12348 27520
rect 12207 27489 12219 27492
rect 12161 27483 12219 27489
rect 11112 27424 11652 27452
rect 11112 27412 11118 27424
rect 11992 27384 12020 27483
rect 12342 27480 12348 27492
rect 12400 27480 12406 27532
rect 12544 27520 12572 27628
rect 12710 27616 12716 27668
rect 12768 27656 12774 27668
rect 13078 27656 13084 27668
rect 12768 27628 13084 27656
rect 12768 27616 12774 27628
rect 13078 27616 13084 27628
rect 13136 27616 13142 27668
rect 13170 27616 13176 27668
rect 13228 27656 13234 27668
rect 13265 27659 13323 27665
rect 13265 27656 13277 27659
rect 13228 27628 13277 27656
rect 13228 27616 13234 27628
rect 13265 27625 13277 27628
rect 13311 27625 13323 27659
rect 13265 27619 13323 27625
rect 17862 27616 17868 27668
rect 17920 27616 17926 27668
rect 19886 27616 19892 27668
rect 19944 27656 19950 27668
rect 22186 27656 22192 27668
rect 19944 27628 22192 27656
rect 19944 27616 19950 27628
rect 22186 27616 22192 27628
rect 22244 27616 22250 27668
rect 23106 27616 23112 27668
rect 23164 27616 23170 27668
rect 23290 27616 23296 27668
rect 23348 27656 23354 27668
rect 23474 27656 23480 27668
rect 23348 27628 23480 27656
rect 23348 27616 23354 27628
rect 23474 27616 23480 27628
rect 23532 27616 23538 27668
rect 24486 27616 24492 27668
rect 24544 27656 24550 27668
rect 24673 27659 24731 27665
rect 24673 27656 24685 27659
rect 24544 27628 24685 27656
rect 24544 27616 24550 27628
rect 24673 27625 24685 27628
rect 24719 27625 24731 27659
rect 24673 27619 24731 27625
rect 26050 27616 26056 27668
rect 26108 27656 26114 27668
rect 26108 27628 26188 27656
rect 26108 27616 26114 27628
rect 13354 27548 13360 27600
rect 13412 27588 13418 27600
rect 14550 27588 14556 27600
rect 13412 27560 14556 27588
rect 13412 27548 13418 27560
rect 14550 27548 14556 27560
rect 14608 27548 14614 27600
rect 17037 27591 17095 27597
rect 17037 27557 17049 27591
rect 17083 27588 17095 27591
rect 17126 27588 17132 27600
rect 17083 27560 17132 27588
rect 17083 27557 17095 27560
rect 17037 27551 17095 27557
rect 17126 27548 17132 27560
rect 17184 27548 17190 27600
rect 21266 27588 21272 27600
rect 20732 27560 21272 27588
rect 15562 27520 15568 27532
rect 12544 27492 15568 27520
rect 12069 27455 12127 27461
rect 12069 27421 12081 27455
rect 12115 27452 12127 27455
rect 12434 27452 12440 27464
rect 12115 27424 12440 27452
rect 12115 27421 12127 27424
rect 12069 27415 12127 27421
rect 12434 27412 12440 27424
rect 12492 27412 12498 27464
rect 12710 27412 12716 27464
rect 12768 27412 12774 27464
rect 12802 27412 12808 27464
rect 12860 27452 12866 27464
rect 12897 27455 12955 27461
rect 12897 27452 12909 27455
rect 12860 27424 12909 27452
rect 12860 27412 12866 27424
rect 12897 27421 12909 27424
rect 12943 27421 12955 27455
rect 12897 27415 12955 27421
rect 13078 27412 13084 27464
rect 13136 27412 13142 27464
rect 13446 27412 13452 27464
rect 13504 27452 13510 27464
rect 14476 27461 14504 27492
rect 15562 27480 15568 27492
rect 15620 27480 15626 27532
rect 18322 27480 18328 27532
rect 18380 27480 18386 27532
rect 18414 27480 18420 27532
rect 18472 27480 18478 27532
rect 19797 27523 19855 27529
rect 19797 27489 19809 27523
rect 19843 27520 19855 27523
rect 20162 27520 20168 27532
rect 19843 27492 20168 27520
rect 19843 27489 19855 27492
rect 19797 27483 19855 27489
rect 20162 27480 20168 27492
rect 20220 27480 20226 27532
rect 14277 27455 14335 27461
rect 14277 27452 14289 27455
rect 13504 27424 14289 27452
rect 13504 27412 13510 27424
rect 14277 27421 14289 27424
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 14461 27455 14519 27461
rect 14461 27421 14473 27455
rect 14507 27421 14519 27455
rect 14461 27415 14519 27421
rect 14550 27412 14556 27464
rect 14608 27412 14614 27464
rect 14645 27455 14703 27461
rect 14645 27421 14657 27455
rect 14691 27446 14703 27455
rect 15194 27452 15200 27464
rect 14752 27446 15200 27452
rect 14691 27424 15200 27446
rect 14691 27421 14780 27424
rect 14645 27418 14780 27421
rect 14645 27415 14703 27418
rect 15194 27412 15200 27424
rect 15252 27412 15258 27464
rect 15286 27412 15292 27464
rect 15344 27452 15350 27464
rect 15654 27452 15660 27464
rect 15344 27424 15660 27452
rect 15344 27412 15350 27424
rect 15654 27412 15660 27424
rect 15712 27412 15718 27464
rect 15930 27461 15936 27464
rect 15924 27452 15936 27461
rect 15891 27424 15936 27452
rect 15924 27415 15936 27424
rect 15930 27412 15936 27415
rect 15988 27412 15994 27464
rect 16482 27412 16488 27464
rect 16540 27452 16546 27464
rect 17954 27452 17960 27464
rect 16540 27424 17960 27452
rect 16540 27412 16546 27424
rect 17954 27412 17960 27424
rect 18012 27412 18018 27464
rect 18230 27412 18236 27464
rect 18288 27452 18294 27464
rect 19889 27455 19947 27461
rect 18288 27424 19840 27452
rect 18288 27412 18294 27424
rect 9968 27356 12020 27384
rect 12989 27387 13047 27393
rect 12989 27353 13001 27387
rect 13035 27384 13047 27387
rect 14090 27384 14096 27396
rect 13035 27356 14096 27384
rect 13035 27353 13047 27356
rect 12989 27347 13047 27353
rect 14090 27344 14096 27356
rect 14148 27344 14154 27396
rect 19242 27384 19248 27396
rect 14191 27356 19248 27384
rect 8481 27319 8539 27325
rect 8481 27285 8493 27319
rect 8527 27316 8539 27319
rect 8570 27316 8576 27328
rect 8527 27288 8576 27316
rect 8527 27285 8539 27288
rect 8481 27279 8539 27285
rect 8570 27276 8576 27288
rect 8628 27276 8634 27328
rect 10410 27276 10416 27328
rect 10468 27316 10474 27328
rect 10597 27319 10655 27325
rect 10597 27316 10609 27319
rect 10468 27288 10609 27316
rect 10468 27276 10474 27288
rect 10597 27285 10609 27288
rect 10643 27285 10655 27319
rect 10597 27279 10655 27285
rect 11701 27319 11759 27325
rect 11701 27285 11713 27319
rect 11747 27316 11759 27319
rect 11882 27316 11888 27328
rect 11747 27288 11888 27316
rect 11747 27285 11759 27288
rect 11701 27279 11759 27285
rect 11882 27276 11888 27288
rect 11940 27276 11946 27328
rect 11974 27276 11980 27328
rect 12032 27316 12038 27328
rect 14191 27316 14219 27356
rect 19242 27344 19248 27356
rect 19300 27344 19306 27396
rect 12032 27288 14219 27316
rect 12032 27276 12038 27288
rect 14826 27276 14832 27328
rect 14884 27276 14890 27328
rect 18046 27276 18052 27328
rect 18104 27316 18110 27328
rect 18233 27319 18291 27325
rect 18233 27316 18245 27319
rect 18104 27288 18245 27316
rect 18104 27276 18110 27288
rect 18233 27285 18245 27288
rect 18279 27316 18291 27319
rect 18690 27316 18696 27328
rect 18279 27288 18696 27316
rect 18279 27285 18291 27288
rect 18233 27279 18291 27285
rect 18690 27276 18696 27288
rect 18748 27276 18754 27328
rect 19058 27276 19064 27328
rect 19116 27316 19122 27328
rect 19613 27319 19671 27325
rect 19613 27316 19625 27319
rect 19116 27288 19625 27316
rect 19116 27276 19122 27288
rect 19613 27285 19625 27288
rect 19659 27285 19671 27319
rect 19812 27316 19840 27424
rect 19889 27421 19901 27455
rect 19935 27452 19947 27455
rect 20732 27452 20760 27560
rect 21266 27548 21272 27560
rect 21324 27548 21330 27600
rect 22370 27548 22376 27600
rect 22428 27588 22434 27600
rect 23385 27591 23443 27597
rect 22428 27560 23336 27588
rect 22428 27548 22434 27560
rect 20824 27492 21036 27520
rect 20824 27461 20852 27492
rect 19935 27424 20760 27452
rect 20809 27455 20867 27461
rect 19935 27421 19947 27424
rect 19889 27415 19947 27421
rect 20809 27421 20821 27455
rect 20855 27421 20867 27455
rect 20809 27415 20867 27421
rect 20901 27455 20959 27461
rect 20901 27421 20913 27455
rect 20947 27421 20959 27455
rect 21008 27452 21036 27492
rect 22002 27480 22008 27532
rect 22060 27520 22066 27532
rect 22281 27523 22339 27529
rect 22281 27520 22293 27523
rect 22060 27492 22293 27520
rect 22060 27480 22066 27492
rect 22281 27489 22293 27492
rect 22327 27489 22339 27523
rect 22281 27483 22339 27489
rect 22465 27523 22523 27529
rect 22465 27489 22477 27523
rect 22511 27520 22523 27523
rect 23198 27520 23204 27532
rect 22511 27492 23204 27520
rect 22511 27489 22523 27492
rect 22465 27483 22523 27489
rect 23198 27480 23204 27492
rect 23256 27480 23262 27532
rect 23308 27520 23336 27560
rect 23385 27557 23397 27591
rect 23431 27588 23443 27591
rect 25866 27588 25872 27600
rect 23431 27560 25872 27588
rect 23431 27557 23443 27560
rect 23385 27551 23443 27557
rect 25866 27548 25872 27560
rect 25924 27548 25930 27600
rect 26160 27588 26188 27628
rect 26786 27616 26792 27668
rect 26844 27656 26850 27668
rect 28350 27656 28356 27668
rect 26844 27628 28356 27656
rect 26844 27616 26850 27628
rect 28350 27616 28356 27628
rect 28408 27616 28414 27668
rect 28534 27616 28540 27668
rect 28592 27656 28598 27668
rect 30558 27656 30564 27668
rect 28592 27628 30564 27656
rect 28592 27616 28598 27628
rect 30558 27616 30564 27628
rect 30616 27616 30622 27668
rect 34790 27616 34796 27668
rect 34848 27656 34854 27668
rect 35529 27659 35587 27665
rect 35529 27656 35541 27659
rect 34848 27628 35541 27656
rect 34848 27616 34854 27628
rect 35529 27625 35541 27628
rect 35575 27625 35587 27659
rect 35529 27619 35587 27625
rect 35636 27628 36308 27656
rect 27890 27588 27896 27600
rect 26160 27560 27896 27588
rect 23308 27492 24440 27520
rect 22094 27452 22100 27464
rect 21008 27424 22100 27452
rect 20901 27415 20959 27421
rect 20165 27387 20223 27393
rect 20165 27353 20177 27387
rect 20211 27353 20223 27387
rect 20165 27347 20223 27353
rect 20257 27387 20315 27393
rect 20257 27353 20269 27387
rect 20303 27353 20315 27387
rect 20257 27347 20315 27353
rect 20180 27316 20208 27347
rect 19812 27288 20208 27316
rect 20272 27316 20300 27347
rect 20438 27344 20444 27396
rect 20496 27384 20502 27396
rect 20916 27384 20944 27415
rect 22094 27412 22100 27424
rect 22152 27412 22158 27464
rect 23014 27412 23020 27464
rect 23072 27412 23078 27464
rect 23106 27412 23112 27464
rect 23164 27412 23170 27464
rect 23845 27455 23903 27461
rect 23845 27421 23857 27455
rect 23891 27421 23903 27455
rect 23845 27415 23903 27421
rect 20496 27356 20944 27384
rect 21085 27387 21143 27393
rect 20496 27344 20502 27356
rect 21085 27353 21097 27387
rect 21131 27384 21143 27387
rect 21542 27384 21548 27396
rect 21131 27356 21548 27384
rect 21131 27353 21143 27356
rect 21085 27347 21143 27353
rect 21542 27344 21548 27356
rect 21600 27344 21606 27396
rect 22189 27387 22247 27393
rect 22189 27353 22201 27387
rect 22235 27384 22247 27387
rect 23566 27384 23572 27396
rect 22235 27356 23572 27384
rect 22235 27353 22247 27356
rect 22189 27347 22247 27353
rect 23566 27344 23572 27356
rect 23624 27344 23630 27396
rect 23860 27384 23888 27415
rect 24026 27412 24032 27464
rect 24084 27412 24090 27464
rect 24412 27452 24440 27492
rect 24486 27480 24492 27532
rect 24544 27520 24550 27532
rect 24857 27523 24915 27529
rect 24857 27520 24869 27523
rect 24544 27492 24869 27520
rect 24544 27480 24550 27492
rect 24857 27489 24869 27492
rect 24903 27489 24915 27523
rect 24857 27483 24915 27489
rect 25056 27492 26004 27520
rect 25056 27461 25084 27492
rect 25041 27455 25099 27461
rect 24412 27424 24992 27452
rect 24394 27384 24400 27396
rect 23860 27356 24400 27384
rect 24394 27344 24400 27356
rect 24452 27344 24458 27396
rect 24578 27344 24584 27396
rect 24636 27344 24642 27396
rect 24964 27384 24992 27424
rect 25041 27421 25053 27455
rect 25087 27421 25099 27455
rect 25041 27415 25099 27421
rect 25314 27412 25320 27464
rect 25372 27452 25378 27464
rect 25869 27455 25927 27461
rect 25869 27452 25881 27455
rect 25372 27424 25881 27452
rect 25372 27412 25378 27424
rect 25869 27421 25881 27424
rect 25915 27421 25927 27455
rect 25976 27452 26004 27492
rect 26050 27480 26056 27532
rect 26108 27520 26114 27532
rect 26145 27523 26203 27529
rect 26145 27520 26157 27523
rect 26108 27492 26157 27520
rect 26108 27480 26114 27492
rect 26145 27489 26157 27492
rect 26191 27489 26203 27523
rect 26145 27483 26203 27489
rect 26237 27523 26295 27529
rect 26237 27489 26249 27523
rect 26283 27520 26295 27523
rect 27338 27520 27344 27532
rect 26283 27492 27344 27520
rect 26283 27489 26295 27492
rect 26237 27483 26295 27489
rect 27338 27480 27344 27492
rect 27396 27480 27402 27532
rect 26602 27452 26608 27464
rect 25976 27424 26608 27452
rect 25869 27415 25927 27421
rect 26602 27412 26608 27424
rect 26660 27452 26666 27464
rect 27525 27455 27583 27461
rect 26660 27424 27476 27452
rect 26660 27412 26666 27424
rect 26234 27384 26240 27396
rect 24964 27356 26240 27384
rect 26234 27344 26240 27356
rect 26292 27344 26298 27396
rect 26326 27344 26332 27396
rect 26384 27393 26390 27396
rect 26384 27387 26412 27393
rect 26400 27353 26412 27387
rect 27448 27384 27476 27424
rect 27525 27421 27537 27455
rect 27571 27452 27583 27455
rect 27632 27452 27660 27560
rect 27890 27548 27896 27560
rect 27948 27548 27954 27600
rect 28074 27548 28080 27600
rect 28132 27588 28138 27600
rect 30006 27588 30012 27600
rect 28132 27560 30012 27588
rect 28132 27548 28138 27560
rect 30006 27548 30012 27560
rect 30064 27548 30070 27600
rect 30650 27548 30656 27600
rect 30708 27588 30714 27600
rect 35636 27588 35664 27628
rect 30708 27560 35664 27588
rect 30708 27548 30714 27560
rect 35986 27548 35992 27600
rect 36044 27548 36050 27600
rect 27798 27480 27804 27532
rect 27856 27520 27862 27532
rect 27985 27523 28043 27529
rect 27985 27520 27997 27523
rect 27856 27492 27997 27520
rect 27856 27480 27862 27492
rect 27985 27489 27997 27492
rect 28031 27520 28043 27523
rect 28718 27520 28724 27532
rect 28031 27492 28724 27520
rect 28031 27489 28043 27492
rect 27985 27483 28043 27489
rect 28718 27480 28724 27492
rect 28776 27480 28782 27532
rect 29178 27520 29184 27532
rect 28828 27492 29184 27520
rect 27571 27424 27660 27452
rect 27709 27455 27767 27461
rect 27571 27421 27583 27424
rect 27525 27415 27583 27421
rect 27709 27421 27721 27455
rect 27755 27452 27767 27455
rect 28074 27452 28080 27464
rect 27755 27424 28080 27452
rect 27755 27421 27767 27424
rect 27709 27415 27767 27421
rect 28074 27412 28080 27424
rect 28132 27412 28138 27464
rect 28828 27461 28856 27492
rect 29178 27480 29184 27492
rect 29236 27480 29242 27532
rect 32214 27480 32220 27532
rect 32272 27480 32278 27532
rect 33336 27492 36032 27520
rect 28813 27455 28871 27461
rect 28813 27421 28825 27455
rect 28859 27421 28871 27455
rect 28813 27415 28871 27421
rect 28902 27412 28908 27464
rect 28960 27412 28966 27464
rect 28997 27455 29055 27461
rect 28997 27421 29009 27455
rect 29043 27421 29055 27455
rect 28997 27415 29055 27421
rect 29089 27455 29147 27461
rect 29089 27421 29101 27455
rect 29135 27452 29147 27455
rect 29270 27452 29276 27464
rect 29135 27424 29276 27452
rect 29135 27421 29147 27424
rect 29089 27415 29147 27421
rect 29012 27384 29040 27415
rect 29270 27412 29276 27424
rect 29328 27412 29334 27464
rect 29917 27455 29975 27461
rect 29917 27421 29929 27455
rect 29963 27452 29975 27455
rect 30006 27452 30012 27464
rect 29963 27424 30012 27452
rect 29963 27421 29975 27424
rect 29917 27415 29975 27421
rect 30006 27412 30012 27424
rect 30064 27412 30070 27464
rect 30374 27412 30380 27464
rect 30432 27412 30438 27464
rect 30558 27412 30564 27464
rect 30616 27412 30622 27464
rect 32769 27455 32827 27461
rect 32769 27452 32781 27455
rect 31404 27424 32781 27452
rect 31018 27384 31024 27396
rect 27448 27356 28764 27384
rect 29012 27356 31024 27384
rect 26384 27347 26412 27353
rect 26384 27344 26390 27347
rect 20714 27316 20720 27328
rect 20272 27288 20720 27316
rect 19613 27279 19671 27285
rect 20714 27276 20720 27288
rect 20772 27276 20778 27328
rect 21818 27276 21824 27328
rect 21876 27276 21882 27328
rect 23474 27276 23480 27328
rect 23532 27316 23538 27328
rect 23937 27319 23995 27325
rect 23937 27316 23949 27319
rect 23532 27288 23949 27316
rect 23532 27276 23538 27288
rect 23937 27285 23949 27288
rect 23983 27285 23995 27319
rect 23937 27279 23995 27285
rect 25222 27276 25228 27328
rect 25280 27276 25286 27328
rect 26513 27319 26571 27325
rect 26513 27285 26525 27319
rect 26559 27316 26571 27319
rect 27246 27316 27252 27328
rect 26559 27288 27252 27316
rect 26559 27285 26571 27288
rect 26513 27279 26571 27285
rect 27246 27276 27252 27288
rect 27304 27276 27310 27328
rect 28626 27276 28632 27328
rect 28684 27276 28690 27328
rect 28736 27316 28764 27356
rect 31018 27344 31024 27356
rect 31076 27344 31082 27396
rect 31294 27344 31300 27396
rect 31352 27384 31358 27396
rect 31404 27393 31432 27424
rect 32769 27421 32781 27424
rect 32815 27421 32827 27455
rect 32769 27415 32827 27421
rect 31389 27387 31447 27393
rect 31389 27384 31401 27387
rect 31352 27356 31401 27384
rect 31352 27344 31358 27356
rect 31389 27353 31401 27356
rect 31435 27353 31447 27387
rect 31389 27347 31447 27353
rect 33134 27344 33140 27396
rect 33192 27384 33198 27396
rect 33336 27384 33364 27492
rect 33410 27412 33416 27464
rect 33468 27452 33474 27464
rect 33468 27424 33640 27452
rect 33468 27412 33474 27424
rect 33505 27387 33563 27393
rect 33505 27384 33517 27387
rect 33192 27356 33517 27384
rect 33192 27344 33198 27356
rect 33505 27353 33517 27356
rect 33551 27353 33563 27387
rect 33612 27384 33640 27424
rect 33686 27412 33692 27464
rect 33744 27452 33750 27464
rect 34149 27455 34207 27461
rect 34149 27452 34161 27455
rect 33744 27424 34161 27452
rect 33744 27412 33750 27424
rect 34149 27421 34161 27424
rect 34195 27421 34207 27455
rect 34149 27415 34207 27421
rect 34333 27455 34391 27461
rect 34333 27421 34345 27455
rect 34379 27421 34391 27455
rect 34333 27415 34391 27421
rect 34348 27384 34376 27415
rect 34882 27412 34888 27464
rect 34940 27412 34946 27464
rect 34978 27455 35036 27461
rect 34978 27421 34990 27455
rect 35024 27421 35036 27455
rect 34978 27415 35036 27421
rect 34422 27384 34428 27396
rect 33612 27356 34428 27384
rect 33505 27347 33563 27353
rect 34422 27344 34428 27356
rect 34480 27344 34486 27396
rect 34790 27344 34796 27396
rect 34848 27384 34854 27396
rect 34992 27384 35020 27415
rect 35066 27412 35072 27464
rect 35124 27452 35130 27464
rect 35350 27455 35408 27461
rect 35350 27454 35362 27455
rect 35222 27452 35362 27454
rect 35124 27426 35362 27452
rect 35124 27424 35250 27426
rect 35124 27412 35130 27424
rect 35350 27421 35362 27426
rect 35396 27421 35408 27455
rect 36004 27452 36032 27492
rect 36280 27461 36308 27628
rect 36265 27455 36323 27461
rect 36004 27424 36216 27452
rect 35350 27415 35408 27421
rect 34848 27356 35020 27384
rect 34848 27344 34854 27356
rect 35158 27344 35164 27396
rect 35216 27344 35222 27396
rect 35253 27387 35311 27393
rect 35253 27353 35265 27387
rect 35299 27353 35311 27387
rect 35253 27347 35311 27353
rect 35989 27387 36047 27393
rect 35989 27353 36001 27387
rect 36035 27384 36047 27387
rect 36078 27384 36084 27396
rect 36035 27356 36084 27384
rect 36035 27353 36047 27356
rect 35989 27347 36047 27353
rect 29825 27319 29883 27325
rect 29825 27316 29837 27319
rect 28736 27288 29837 27316
rect 29825 27285 29837 27288
rect 29871 27316 29883 27319
rect 32766 27316 32772 27328
rect 29871 27288 32772 27316
rect 29871 27285 29883 27288
rect 29825 27279 29883 27285
rect 32766 27276 32772 27288
rect 32824 27276 32830 27328
rect 33318 27276 33324 27328
rect 33376 27316 33382 27328
rect 34241 27319 34299 27325
rect 34241 27316 34253 27319
rect 33376 27288 34253 27316
rect 33376 27276 33382 27288
rect 34241 27285 34253 27288
rect 34287 27285 34299 27319
rect 34241 27279 34299 27285
rect 34514 27276 34520 27328
rect 34572 27316 34578 27328
rect 35268 27316 35296 27347
rect 36078 27344 36084 27356
rect 36136 27344 36142 27396
rect 36188 27384 36216 27424
rect 36265 27421 36277 27455
rect 36311 27421 36323 27455
rect 36265 27415 36323 27421
rect 36630 27412 36636 27464
rect 36688 27412 36694 27464
rect 36722 27412 36728 27464
rect 36780 27412 36786 27464
rect 36648 27384 36676 27412
rect 36188 27356 36676 27384
rect 36992 27387 37050 27393
rect 36992 27353 37004 27387
rect 37038 27384 37050 27387
rect 37458 27384 37464 27396
rect 37038 27356 37464 27384
rect 37038 27353 37050 27356
rect 36992 27347 37050 27353
rect 37458 27344 37464 27356
rect 37516 27344 37522 27396
rect 35802 27316 35808 27328
rect 34572 27288 35808 27316
rect 34572 27276 34578 27288
rect 35802 27276 35808 27288
rect 35860 27276 35866 27328
rect 36173 27319 36231 27325
rect 36173 27285 36185 27319
rect 36219 27316 36231 27319
rect 36630 27316 36636 27328
rect 36219 27288 36636 27316
rect 36219 27285 36231 27288
rect 36173 27279 36231 27285
rect 36630 27276 36636 27288
rect 36688 27276 36694 27328
rect 38102 27276 38108 27328
rect 38160 27276 38166 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 8018 27072 8024 27124
rect 8076 27072 8082 27124
rect 8481 27115 8539 27121
rect 8481 27081 8493 27115
rect 8527 27112 8539 27115
rect 9306 27112 9312 27124
rect 8527 27084 9312 27112
rect 8527 27081 8539 27084
rect 8481 27075 8539 27081
rect 9306 27072 9312 27084
rect 9364 27072 9370 27124
rect 12986 27112 12992 27124
rect 11247 27084 12992 27112
rect 8389 27047 8447 27053
rect 8389 27013 8401 27047
rect 8435 27044 8447 27047
rect 8570 27044 8576 27056
rect 8435 27016 8576 27044
rect 8435 27013 8447 27016
rect 8389 27007 8447 27013
rect 8570 27004 8576 27016
rect 8628 27044 8634 27056
rect 11054 27044 11060 27056
rect 8628 27016 11060 27044
rect 8628 27004 8634 27016
rect 11054 27004 11060 27016
rect 11112 27004 11118 27056
rect 9582 26936 9588 26988
rect 9640 26936 9646 26988
rect 9769 26979 9827 26985
rect 9769 26945 9781 26979
rect 9815 26945 9827 26979
rect 9769 26939 9827 26945
rect 8665 26911 8723 26917
rect 8665 26877 8677 26911
rect 8711 26877 8723 26911
rect 9784 26908 9812 26939
rect 9858 26936 9864 26988
rect 9916 26936 9922 26988
rect 9953 26979 10011 26985
rect 9953 26945 9965 26979
rect 9999 26976 10011 26979
rect 10781 26979 10839 26985
rect 9999 26948 10732 26976
rect 9999 26945 10011 26948
rect 9953 26939 10011 26945
rect 9784 26880 10088 26908
rect 8665 26871 8723 26877
rect 8680 26840 8708 26871
rect 9950 26840 9956 26852
rect 8680 26812 9956 26840
rect 9950 26800 9956 26812
rect 10008 26800 10014 26852
rect 10060 26840 10088 26880
rect 10134 26868 10140 26920
rect 10192 26908 10198 26920
rect 10502 26908 10508 26920
rect 10192 26880 10508 26908
rect 10192 26868 10198 26880
rect 10502 26868 10508 26880
rect 10560 26908 10566 26920
rect 10597 26911 10655 26917
rect 10597 26908 10609 26911
rect 10560 26880 10609 26908
rect 10560 26868 10566 26880
rect 10597 26877 10609 26880
rect 10643 26877 10655 26911
rect 10704 26908 10732 26948
rect 10781 26945 10793 26979
rect 10827 26976 10839 26979
rect 10962 26976 10968 26988
rect 10827 26948 10968 26976
rect 10827 26945 10839 26948
rect 10781 26939 10839 26945
rect 10962 26936 10968 26948
rect 11020 26936 11026 26988
rect 10870 26908 10876 26920
rect 10704 26880 10876 26908
rect 10597 26871 10655 26877
rect 10870 26868 10876 26880
rect 10928 26908 10934 26920
rect 11247 26908 11275 27084
rect 12802 27044 12808 27056
rect 12452 27016 12808 27044
rect 12452 26985 12480 27016
rect 12802 27004 12808 27016
rect 12860 27004 12866 27056
rect 12437 26979 12495 26985
rect 12437 26945 12449 26979
rect 12483 26945 12495 26979
rect 12437 26939 12495 26945
rect 12621 26979 12679 26985
rect 12621 26945 12633 26979
rect 12667 26945 12679 26979
rect 12621 26939 12679 26945
rect 12713 26979 12771 26985
rect 12713 26945 12725 26979
rect 12759 26976 12771 26979
rect 12912 26976 12940 27084
rect 12986 27072 12992 27084
rect 13044 27072 13050 27124
rect 13446 27072 13452 27124
rect 13504 27112 13510 27124
rect 15949 27115 16007 27121
rect 15949 27112 15961 27115
rect 13504 27084 15961 27112
rect 13504 27072 13510 27084
rect 15949 27081 15961 27084
rect 15995 27081 16007 27115
rect 15949 27075 16007 27081
rect 18138 27072 18144 27124
rect 18196 27112 18202 27124
rect 18877 27115 18935 27121
rect 18877 27112 18889 27115
rect 18196 27084 18889 27112
rect 18196 27072 18202 27084
rect 18877 27081 18889 27084
rect 18923 27081 18935 27115
rect 18877 27075 18935 27081
rect 19242 27072 19248 27124
rect 19300 27112 19306 27124
rect 19300 27084 20034 27112
rect 19300 27072 19306 27084
rect 14176 27047 14234 27053
rect 14176 27013 14188 27047
rect 14222 27044 14234 27047
rect 14826 27044 14832 27056
rect 14222 27016 14832 27044
rect 14222 27013 14234 27016
rect 14176 27007 14234 27013
rect 14826 27004 14832 27016
rect 14884 27004 14890 27056
rect 15749 27047 15807 27053
rect 15749 27013 15761 27047
rect 15795 27013 15807 27047
rect 19334 27044 19340 27056
rect 15749 27007 15807 27013
rect 18892 27016 19340 27044
rect 12759 26948 12940 26976
rect 13265 26979 13323 26985
rect 12759 26945 12771 26948
rect 12713 26939 12771 26945
rect 13265 26945 13277 26979
rect 13311 26976 13323 26979
rect 13354 26976 13360 26988
rect 13311 26948 13360 26976
rect 13311 26945 13323 26948
rect 13265 26939 13323 26945
rect 10928 26880 11275 26908
rect 12636 26908 12664 26939
rect 13354 26936 13360 26948
rect 13412 26936 13418 26988
rect 13446 26936 13452 26988
rect 13504 26936 13510 26988
rect 14458 26936 14464 26988
rect 14516 26976 14522 26988
rect 15764 26976 15792 27007
rect 18892 26988 18920 27016
rect 19334 27004 19340 27016
rect 19392 27044 19398 27056
rect 19392 27016 19472 27044
rect 19392 27004 19398 27016
rect 14516 26948 15792 26976
rect 14516 26936 14522 26948
rect 16942 26936 16948 26988
rect 17000 26936 17006 26988
rect 17212 26979 17270 26985
rect 17212 26945 17224 26979
rect 17258 26976 17270 26979
rect 17494 26976 17500 26988
rect 17258 26948 17500 26976
rect 17258 26945 17270 26948
rect 17212 26939 17270 26945
rect 17494 26936 17500 26948
rect 17552 26936 17558 26988
rect 17586 26936 17592 26988
rect 17644 26976 17650 26988
rect 17644 26948 18368 26976
rect 17644 26936 17650 26948
rect 13170 26908 13176 26920
rect 12636 26880 13176 26908
rect 10928 26868 10934 26880
rect 13170 26868 13176 26880
rect 13228 26868 13234 26920
rect 13906 26868 13912 26920
rect 13964 26868 13970 26920
rect 15378 26868 15384 26920
rect 15436 26908 15442 26920
rect 16022 26908 16028 26920
rect 15436 26880 16028 26908
rect 15436 26868 15442 26880
rect 16022 26868 16028 26880
rect 16080 26868 16086 26920
rect 10965 26843 11023 26849
rect 10060 26812 10640 26840
rect 10612 26784 10640 26812
rect 10965 26809 10977 26843
rect 11011 26840 11023 26843
rect 11011 26812 13952 26840
rect 11011 26809 11023 26812
rect 10965 26803 11023 26809
rect 10134 26732 10140 26784
rect 10192 26732 10198 26784
rect 10594 26732 10600 26784
rect 10652 26772 10658 26784
rect 10980 26772 11008 26803
rect 10652 26744 11008 26772
rect 10652 26732 10658 26744
rect 12250 26732 12256 26784
rect 12308 26732 12314 26784
rect 13262 26732 13268 26784
rect 13320 26732 13326 26784
rect 13924 26772 13952 26812
rect 15194 26800 15200 26852
rect 15252 26840 15258 26852
rect 15252 26812 16988 26840
rect 15252 26800 15258 26812
rect 14918 26772 14924 26784
rect 13924 26744 14924 26772
rect 14918 26732 14924 26744
rect 14976 26732 14982 26784
rect 15286 26732 15292 26784
rect 15344 26732 15350 26784
rect 15562 26732 15568 26784
rect 15620 26772 15626 26784
rect 15933 26775 15991 26781
rect 15933 26772 15945 26775
rect 15620 26744 15945 26772
rect 15620 26732 15626 26744
rect 15933 26741 15945 26744
rect 15979 26741 15991 26775
rect 15933 26735 15991 26741
rect 16114 26732 16120 26784
rect 16172 26732 16178 26784
rect 16960 26772 16988 26812
rect 18230 26772 18236 26784
rect 16960 26744 18236 26772
rect 18230 26732 18236 26744
rect 18288 26732 18294 26784
rect 18340 26781 18368 26948
rect 18598 26936 18604 26988
rect 18656 26936 18662 26988
rect 18874 26936 18880 26988
rect 18932 26936 18938 26988
rect 19058 26936 19064 26988
rect 19116 26936 19122 26988
rect 19153 26979 19211 26985
rect 19153 26945 19165 26979
rect 19199 26976 19211 26979
rect 19242 26976 19248 26988
rect 19199 26948 19248 26976
rect 19199 26945 19211 26948
rect 19153 26939 19211 26945
rect 19242 26936 19248 26948
rect 19300 26936 19306 26988
rect 19444 26985 19472 27016
rect 19429 26979 19487 26985
rect 19429 26945 19441 26979
rect 19475 26945 19487 26979
rect 19429 26939 19487 26945
rect 20006 26966 20034 27084
rect 20070 27072 20076 27124
rect 20128 27112 20134 27124
rect 21358 27112 21364 27124
rect 20128 27084 21364 27112
rect 20128 27072 20134 27084
rect 20533 27047 20591 27053
rect 20533 27044 20545 27047
rect 20364 27016 20545 27044
rect 20364 26966 20392 27016
rect 20533 27013 20545 27016
rect 20579 27013 20591 27047
rect 20533 27007 20591 27013
rect 20622 27004 20628 27056
rect 20680 27004 20686 27056
rect 20732 27053 20760 27084
rect 21358 27072 21364 27084
rect 21416 27072 21422 27124
rect 22002 27072 22008 27124
rect 22060 27112 22066 27124
rect 25222 27112 25228 27124
rect 22060 27084 25228 27112
rect 22060 27072 22066 27084
rect 25222 27072 25228 27084
rect 25280 27072 25286 27124
rect 26418 27112 26424 27124
rect 25992 27084 26424 27112
rect 20732 27047 20801 27053
rect 20732 27016 20755 27047
rect 20743 27013 20755 27016
rect 20789 27013 20801 27047
rect 20743 27007 20801 27013
rect 21818 27004 21824 27056
rect 21876 27044 21882 27056
rect 23385 27047 23443 27053
rect 23385 27044 23397 27047
rect 21876 27016 23397 27044
rect 21876 27004 21882 27016
rect 23385 27013 23397 27016
rect 23431 27013 23443 27047
rect 23842 27044 23848 27056
rect 23385 27007 23443 27013
rect 23492 27016 23848 27044
rect 20006 26938 20392 26966
rect 20441 26979 20499 26985
rect 20441 26945 20453 26979
rect 20487 26976 20499 26979
rect 22373 26979 22431 26985
rect 22373 26976 22385 26979
rect 20487 26948 22385 26976
rect 20487 26945 20499 26948
rect 20441 26939 20499 26945
rect 22373 26945 22385 26948
rect 22419 26976 22431 26979
rect 22462 26976 22468 26988
rect 22419 26948 22468 26976
rect 22419 26945 22431 26948
rect 22373 26939 22431 26945
rect 22462 26936 22468 26948
rect 22520 26936 22526 26988
rect 22557 26979 22615 26985
rect 22557 26945 22569 26979
rect 22603 26945 22615 26979
rect 22557 26939 22615 26945
rect 22925 26979 22983 26985
rect 22925 26945 22937 26979
rect 22971 26976 22983 26979
rect 23290 26976 23296 26988
rect 22971 26948 23296 26976
rect 22971 26945 22983 26948
rect 22925 26939 22983 26945
rect 18616 26908 18644 26936
rect 19337 26911 19395 26917
rect 19337 26908 19349 26911
rect 18616 26880 19349 26908
rect 19337 26877 19349 26880
rect 19383 26877 19395 26911
rect 19337 26871 19395 26877
rect 19886 26868 19892 26920
rect 19944 26908 19950 26920
rect 20530 26908 20536 26920
rect 19944 26880 20536 26908
rect 19944 26868 19950 26880
rect 20530 26868 20536 26880
rect 20588 26868 20594 26920
rect 20898 26908 20904 26920
rect 20640 26880 20904 26908
rect 18506 26800 18512 26852
rect 18564 26840 18570 26852
rect 20640 26840 20668 26880
rect 20898 26868 20904 26880
rect 20956 26868 20962 26920
rect 21358 26868 21364 26920
rect 21416 26908 21422 26920
rect 22572 26908 22600 26939
rect 23290 26936 23296 26948
rect 23348 26976 23354 26988
rect 23492 26976 23520 27016
rect 23842 27004 23848 27016
rect 23900 27004 23906 27056
rect 24118 27004 24124 27056
rect 24176 27044 24182 27056
rect 24176 27016 24440 27044
rect 24176 27004 24182 27016
rect 24412 26985 24440 27016
rect 24486 27004 24492 27056
rect 24544 27044 24550 27056
rect 24673 27047 24731 27053
rect 24673 27044 24685 27047
rect 24544 27016 24685 27044
rect 24544 27004 24550 27016
rect 24673 27013 24685 27016
rect 24719 27013 24731 27047
rect 25992 27044 26020 27084
rect 26418 27072 26424 27084
rect 26476 27072 26482 27124
rect 26605 27115 26663 27121
rect 26605 27081 26617 27115
rect 26651 27112 26663 27115
rect 27982 27112 27988 27124
rect 26651 27084 27988 27112
rect 26651 27081 26663 27084
rect 26605 27075 26663 27081
rect 27982 27072 27988 27084
rect 28040 27072 28046 27124
rect 28074 27072 28080 27124
rect 28132 27112 28138 27124
rect 28132 27084 31754 27112
rect 28132 27072 28138 27084
rect 24673 27007 24731 27013
rect 25240 27016 26020 27044
rect 25240 26988 25268 27016
rect 26050 27004 26056 27056
rect 26108 27044 26114 27056
rect 27617 27047 27675 27053
rect 27617 27044 27629 27047
rect 26108 27016 27629 27044
rect 26108 27004 26114 27016
rect 27617 27013 27629 27016
rect 27663 27013 27675 27047
rect 27617 27007 27675 27013
rect 27706 27004 27712 27056
rect 27764 27004 27770 27056
rect 27890 27004 27896 27056
rect 27948 27044 27954 27056
rect 27948 27016 28672 27044
rect 27948 27004 27954 27016
rect 23348 26948 23520 26976
rect 23569 26979 23627 26985
rect 23348 26936 23354 26948
rect 23569 26945 23581 26979
rect 23615 26976 23627 26979
rect 24397 26979 24455 26985
rect 23615 26948 24348 26976
rect 23615 26945 23627 26948
rect 23569 26939 23627 26945
rect 21416 26880 22600 26908
rect 21416 26868 21422 26880
rect 23750 26868 23756 26920
rect 23808 26908 23814 26920
rect 24213 26911 24271 26917
rect 24213 26908 24225 26911
rect 23808 26880 24225 26908
rect 23808 26868 23814 26880
rect 24213 26877 24225 26880
rect 24259 26877 24271 26911
rect 24320 26908 24348 26948
rect 24397 26945 24409 26979
rect 24443 26945 24455 26979
rect 24397 26939 24455 26945
rect 24765 26979 24823 26985
rect 24765 26945 24777 26979
rect 24811 26976 24823 26979
rect 25222 26976 25228 26988
rect 24811 26948 25228 26976
rect 24811 26945 24823 26948
rect 24765 26939 24823 26945
rect 25222 26936 25228 26948
rect 25280 26936 25286 26988
rect 25590 26936 25596 26988
rect 25648 26936 25654 26988
rect 26329 26979 26387 26985
rect 26329 26945 26341 26979
rect 26375 26945 26387 26979
rect 26329 26939 26387 26945
rect 26513 26979 26571 26985
rect 26513 26945 26525 26979
rect 26559 26976 26571 26979
rect 26694 26976 26700 26988
rect 26559 26948 26700 26976
rect 26559 26945 26571 26948
rect 26513 26939 26571 26945
rect 26344 26908 26372 26939
rect 26694 26936 26700 26948
rect 26752 26936 26758 26988
rect 27246 26936 27252 26988
rect 27304 26936 27310 26988
rect 28166 26936 28172 26988
rect 28224 26976 28230 26988
rect 28537 26979 28595 26985
rect 28537 26976 28549 26979
rect 28224 26948 28549 26976
rect 28224 26936 28230 26948
rect 28537 26945 28549 26948
rect 28583 26945 28595 26979
rect 28644 26976 28672 27016
rect 28994 27004 29000 27056
rect 29052 27044 29058 27056
rect 31389 27047 31447 27053
rect 29052 27016 31340 27044
rect 29052 27004 29058 27016
rect 29086 26976 29092 26988
rect 28644 26948 29092 26976
rect 28537 26939 28595 26945
rect 29086 26936 29092 26948
rect 29144 26976 29150 26988
rect 29181 26979 29239 26985
rect 29181 26976 29193 26979
rect 29144 26948 29193 26976
rect 29144 26936 29150 26948
rect 29181 26945 29193 26948
rect 29227 26945 29239 26979
rect 29181 26939 29239 26945
rect 31018 26936 31024 26988
rect 31076 26936 31082 26988
rect 31312 26976 31340 27016
rect 31389 27013 31401 27047
rect 31435 27044 31447 27047
rect 31726 27044 31754 27084
rect 34882 27072 34888 27124
rect 34940 27112 34946 27124
rect 37090 27112 37096 27124
rect 34940 27084 37096 27112
rect 34940 27072 34946 27084
rect 37090 27072 37096 27084
rect 37148 27072 37154 27124
rect 37458 27072 37464 27124
rect 37516 27072 37522 27124
rect 37734 27072 37740 27124
rect 37792 27112 37798 27124
rect 37921 27115 37979 27121
rect 37921 27112 37933 27115
rect 37792 27084 37933 27112
rect 37792 27072 37798 27084
rect 37921 27081 37933 27084
rect 37967 27081 37979 27115
rect 37921 27075 37979 27081
rect 31435 27016 31616 27044
rect 31726 27016 33916 27044
rect 31435 27013 31447 27016
rect 31389 27007 31447 27013
rect 31588 26976 31616 27016
rect 31846 26976 31852 26988
rect 31312 26948 31432 26976
rect 31588 26948 31852 26976
rect 27430 26908 27436 26920
rect 24320 26880 27436 26908
rect 24213 26871 24271 26877
rect 27430 26868 27436 26880
rect 27488 26868 27494 26920
rect 28994 26868 29000 26920
rect 29052 26908 29058 26920
rect 29273 26911 29331 26917
rect 29273 26908 29285 26911
rect 29052 26880 29285 26908
rect 29052 26868 29058 26880
rect 29273 26877 29285 26880
rect 29319 26877 29331 26911
rect 29273 26871 29331 26877
rect 30742 26868 30748 26920
rect 30800 26868 30806 26920
rect 30929 26911 30987 26917
rect 30929 26877 30941 26911
rect 30975 26908 30987 26911
rect 31110 26908 31116 26920
rect 30975 26880 31116 26908
rect 30975 26877 30987 26880
rect 30929 26871 30987 26877
rect 31110 26868 31116 26880
rect 31168 26868 31174 26920
rect 31297 26911 31355 26917
rect 31297 26877 31309 26911
rect 31343 26877 31355 26911
rect 31404 26908 31432 26948
rect 31846 26936 31852 26948
rect 31904 26976 31910 26988
rect 32398 26976 32404 26988
rect 31904 26948 32404 26976
rect 31904 26936 31910 26948
rect 32398 26936 32404 26948
rect 32456 26936 32462 26988
rect 32490 26936 32496 26988
rect 32548 26976 32554 26988
rect 32692 26985 32720 27016
rect 32585 26979 32643 26985
rect 32585 26976 32597 26979
rect 32548 26948 32597 26976
rect 32548 26936 32554 26948
rect 32585 26945 32597 26948
rect 32631 26945 32643 26979
rect 32585 26939 32643 26945
rect 32677 26979 32735 26985
rect 32677 26945 32689 26979
rect 32723 26945 32735 26979
rect 32677 26939 32735 26945
rect 32861 26979 32919 26985
rect 32861 26945 32873 26979
rect 32907 26945 32919 26979
rect 32861 26939 32919 26945
rect 33321 26979 33379 26985
rect 33321 26945 33333 26979
rect 33367 26976 33379 26979
rect 33410 26976 33416 26988
rect 33367 26948 33416 26976
rect 33367 26945 33379 26948
rect 33321 26939 33379 26945
rect 31404 26880 31754 26908
rect 31297 26871 31355 26877
rect 25866 26840 25872 26852
rect 18564 26812 20668 26840
rect 22066 26812 25872 26840
rect 18564 26800 18570 26812
rect 18325 26775 18383 26781
rect 18325 26741 18337 26775
rect 18371 26772 18383 26775
rect 18874 26772 18880 26784
rect 18371 26744 18880 26772
rect 18371 26741 18383 26744
rect 18325 26735 18383 26741
rect 18874 26732 18880 26744
rect 18932 26732 18938 26784
rect 20257 26775 20315 26781
rect 20257 26741 20269 26775
rect 20303 26772 20315 26775
rect 20622 26772 20628 26784
rect 20303 26744 20628 26772
rect 20303 26741 20315 26744
rect 20257 26735 20315 26741
rect 20622 26732 20628 26744
rect 20680 26732 20686 26784
rect 20806 26732 20812 26784
rect 20864 26772 20870 26784
rect 22066 26772 22094 26812
rect 25866 26800 25872 26812
rect 25924 26800 25930 26852
rect 26878 26800 26884 26852
rect 26936 26840 26942 26852
rect 29730 26840 29736 26852
rect 26936 26812 29736 26840
rect 26936 26800 26942 26812
rect 29730 26800 29736 26812
rect 29788 26800 29794 26852
rect 30006 26800 30012 26852
rect 30064 26840 30070 26852
rect 30760 26840 30788 26868
rect 31312 26840 31340 26871
rect 30064 26812 31340 26840
rect 31726 26840 31754 26880
rect 32214 26868 32220 26920
rect 32272 26908 32278 26920
rect 32876 26908 32904 26939
rect 33410 26936 33416 26948
rect 33468 26936 33474 26988
rect 33778 26936 33784 26988
rect 33836 26936 33842 26988
rect 33888 26985 33916 27016
rect 34606 27004 34612 27056
rect 34664 27044 34670 27056
rect 35161 27047 35219 27053
rect 35161 27044 35173 27047
rect 34664 27016 35173 27044
rect 34664 27004 34670 27016
rect 35161 27013 35173 27016
rect 35207 27013 35219 27047
rect 35161 27007 35219 27013
rect 35253 27047 35311 27053
rect 35253 27013 35265 27047
rect 35299 27044 35311 27047
rect 35710 27044 35716 27056
rect 35299 27016 35716 27044
rect 35299 27013 35311 27016
rect 35253 27007 35311 27013
rect 35710 27004 35716 27016
rect 35768 27004 35774 27056
rect 35802 27004 35808 27056
rect 35860 27044 35866 27056
rect 35860 27016 36308 27044
rect 35860 27004 35866 27016
rect 33873 26979 33931 26985
rect 33873 26945 33885 26979
rect 33919 26945 33931 26979
rect 33873 26939 33931 26945
rect 34054 26936 34060 26988
rect 34112 26936 34118 26988
rect 34974 26936 34980 26988
rect 35032 26936 35038 26988
rect 35345 26979 35403 26985
rect 35345 26945 35357 26979
rect 35391 26976 35403 26979
rect 35434 26976 35440 26988
rect 35391 26948 35440 26976
rect 35391 26945 35403 26948
rect 35345 26939 35403 26945
rect 35434 26936 35440 26948
rect 35492 26936 35498 26988
rect 35894 26936 35900 26988
rect 35952 26976 35958 26988
rect 36280 26985 36308 27016
rect 36354 27004 36360 27056
rect 36412 27004 36418 27056
rect 35989 26979 36047 26985
rect 35989 26976 36001 26979
rect 35952 26948 36001 26976
rect 35952 26936 35958 26948
rect 35989 26945 36001 26948
rect 36035 26945 36047 26979
rect 35989 26939 36047 26945
rect 36173 26979 36231 26985
rect 36173 26945 36185 26979
rect 36219 26945 36231 26979
rect 36173 26939 36231 26945
rect 36265 26979 36323 26985
rect 36265 26945 36277 26979
rect 36311 26945 36323 26979
rect 36372 26976 36400 27004
rect 36449 26979 36507 26985
rect 36449 26976 36461 26979
rect 36372 26948 36461 26976
rect 36265 26939 36323 26945
rect 36449 26945 36461 26948
rect 36495 26945 36507 26979
rect 36449 26939 36507 26945
rect 36541 26979 36599 26985
rect 36541 26945 36553 26979
rect 36587 26945 36599 26979
rect 36541 26939 36599 26945
rect 37829 26979 37887 26985
rect 37829 26945 37841 26979
rect 37875 26976 37887 26979
rect 38102 26976 38108 26988
rect 37875 26948 38108 26976
rect 37875 26945 37887 26948
rect 37829 26939 37887 26945
rect 34072 26908 34100 26936
rect 32272 26880 34100 26908
rect 34517 26911 34575 26917
rect 32272 26868 32278 26880
rect 34517 26877 34529 26911
rect 34563 26908 34575 26911
rect 35802 26908 35808 26920
rect 34563 26880 35808 26908
rect 34563 26877 34575 26880
rect 34517 26871 34575 26877
rect 35802 26868 35808 26880
rect 35860 26868 35866 26920
rect 36188 26908 36216 26939
rect 36188 26880 36308 26908
rect 33870 26840 33876 26852
rect 31726 26812 33876 26840
rect 30064 26800 30070 26812
rect 33870 26800 33876 26812
rect 33928 26800 33934 26852
rect 36280 26840 36308 26880
rect 36354 26868 36360 26920
rect 36412 26908 36418 26920
rect 36556 26908 36584 26939
rect 36412 26880 36584 26908
rect 36412 26868 36418 26880
rect 36630 26840 36636 26852
rect 33980 26812 36636 26840
rect 20864 26744 22094 26772
rect 20864 26732 20870 26744
rect 23750 26732 23756 26784
rect 23808 26732 23814 26784
rect 24486 26732 24492 26784
rect 24544 26772 24550 26784
rect 24854 26772 24860 26784
rect 24544 26744 24860 26772
rect 24544 26732 24550 26744
rect 24854 26732 24860 26744
rect 24912 26732 24918 26784
rect 27430 26732 27436 26784
rect 27488 26772 27494 26784
rect 30374 26772 30380 26784
rect 27488 26744 30380 26772
rect 27488 26732 27494 26744
rect 30374 26732 30380 26744
rect 30432 26732 30438 26784
rect 30745 26775 30803 26781
rect 30745 26741 30757 26775
rect 30791 26772 30803 26775
rect 31846 26772 31852 26784
rect 30791 26744 31852 26772
rect 30791 26741 30803 26744
rect 30745 26735 30803 26741
rect 31846 26732 31852 26744
rect 31904 26732 31910 26784
rect 32490 26732 32496 26784
rect 32548 26772 32554 26784
rect 33980 26772 34008 26812
rect 36630 26800 36636 26812
rect 36688 26800 36694 26852
rect 32548 26744 34008 26772
rect 32548 26732 32554 26744
rect 34146 26732 34152 26784
rect 34204 26772 34210 26784
rect 34422 26772 34428 26784
rect 34204 26744 34428 26772
rect 34204 26732 34210 26744
rect 34422 26732 34428 26744
rect 34480 26732 34486 26784
rect 34698 26732 34704 26784
rect 34756 26772 34762 26784
rect 35529 26775 35587 26781
rect 35529 26772 35541 26775
rect 34756 26744 35541 26772
rect 34756 26732 34762 26744
rect 35529 26741 35541 26744
rect 35575 26741 35587 26775
rect 35529 26735 35587 26741
rect 35802 26732 35808 26784
rect 35860 26772 35866 26784
rect 37844 26772 37872 26939
rect 38102 26936 38108 26948
rect 38160 26936 38166 26988
rect 38010 26868 38016 26920
rect 38068 26868 38074 26920
rect 38470 26868 38476 26920
rect 38528 26908 38534 26920
rect 39114 26908 39120 26920
rect 38528 26880 39120 26908
rect 38528 26868 38534 26880
rect 39114 26868 39120 26880
rect 39172 26868 39178 26920
rect 35860 26744 37872 26772
rect 35860 26732 35866 26744
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 11330 26528 11336 26580
rect 11388 26568 11394 26580
rect 18506 26568 18512 26580
rect 11388 26540 18512 26568
rect 11388 26528 11394 26540
rect 18506 26528 18512 26540
rect 18564 26528 18570 26580
rect 20254 26528 20260 26580
rect 20312 26568 20318 26580
rect 20312 26540 22508 26568
rect 20312 26528 20318 26540
rect 13170 26460 13176 26512
rect 13228 26500 13234 26512
rect 15194 26500 15200 26512
rect 13228 26472 15200 26500
rect 13228 26460 13234 26472
rect 15194 26460 15200 26472
rect 15252 26460 15258 26512
rect 15289 26503 15347 26509
rect 15289 26469 15301 26503
rect 15335 26500 15347 26503
rect 15562 26500 15568 26512
rect 15335 26472 15568 26500
rect 15335 26469 15347 26472
rect 15289 26463 15347 26469
rect 15562 26460 15568 26472
rect 15620 26460 15626 26512
rect 16850 26460 16856 26512
rect 16908 26500 16914 26512
rect 18877 26503 18935 26509
rect 16908 26472 18828 26500
rect 16908 26460 16914 26472
rect 8202 26392 8208 26444
rect 8260 26432 8266 26444
rect 9953 26435 10011 26441
rect 9953 26432 9965 26435
rect 8260 26404 9965 26432
rect 8260 26392 8266 26404
rect 9953 26401 9965 26404
rect 9999 26401 10011 26435
rect 15654 26432 15660 26444
rect 9953 26395 10011 26401
rect 13924 26404 15660 26432
rect 9968 26364 9996 26395
rect 13924 26376 13952 26404
rect 15654 26392 15660 26404
rect 15712 26432 15718 26444
rect 15749 26435 15807 26441
rect 15749 26432 15761 26435
rect 15712 26404 15761 26432
rect 15712 26392 15718 26404
rect 15749 26401 15761 26404
rect 15795 26401 15807 26435
rect 15749 26395 15807 26401
rect 17402 26392 17408 26444
rect 17460 26432 17466 26444
rect 17460 26404 18000 26432
rect 17460 26392 17466 26404
rect 11698 26364 11704 26376
rect 9968 26336 11704 26364
rect 11698 26324 11704 26336
rect 11756 26364 11762 26376
rect 11793 26367 11851 26373
rect 11793 26364 11805 26367
rect 11756 26336 11805 26364
rect 11756 26324 11762 26336
rect 11793 26333 11805 26336
rect 11839 26364 11851 26367
rect 12894 26364 12900 26376
rect 11839 26336 12900 26364
rect 11839 26333 11851 26336
rect 11793 26327 11851 26333
rect 12894 26324 12900 26336
rect 12952 26364 12958 26376
rect 13906 26364 13912 26376
rect 12952 26336 13912 26364
rect 12952 26324 12958 26336
rect 13906 26324 13912 26336
rect 13964 26324 13970 26376
rect 14734 26324 14740 26376
rect 14792 26324 14798 26376
rect 14826 26324 14832 26376
rect 14884 26364 14890 26376
rect 15013 26367 15071 26373
rect 15013 26364 15025 26367
rect 14884 26336 15025 26364
rect 14884 26324 14890 26336
rect 15013 26333 15025 26336
rect 15059 26333 15071 26367
rect 15013 26327 15071 26333
rect 15105 26367 15163 26373
rect 15105 26333 15117 26367
rect 15151 26364 15163 26367
rect 15194 26364 15200 26376
rect 15151 26336 15200 26364
rect 15151 26333 15163 26336
rect 15105 26327 15163 26333
rect 10220 26299 10278 26305
rect 10220 26265 10232 26299
rect 10266 26296 10278 26299
rect 10962 26296 10968 26308
rect 10266 26268 10968 26296
rect 10266 26265 10278 26268
rect 10220 26259 10278 26265
rect 10962 26256 10968 26268
rect 11020 26256 11026 26308
rect 12060 26299 12118 26305
rect 12060 26265 12072 26299
rect 12106 26296 12118 26299
rect 12250 26296 12256 26308
rect 12106 26268 12256 26296
rect 12106 26265 12118 26268
rect 12060 26259 12118 26265
rect 12250 26256 12256 26268
rect 12308 26256 12314 26308
rect 12434 26256 12440 26308
rect 12492 26296 12498 26308
rect 14458 26296 14464 26308
rect 12492 26268 14464 26296
rect 12492 26256 12498 26268
rect 14458 26256 14464 26268
rect 14516 26256 14522 26308
rect 14918 26256 14924 26308
rect 14976 26256 14982 26308
rect 15028 26296 15056 26327
rect 15194 26324 15200 26336
rect 15252 26324 15258 26376
rect 15562 26324 15568 26376
rect 15620 26364 15626 26376
rect 16005 26367 16063 26373
rect 16005 26364 16017 26367
rect 15620 26336 16017 26364
rect 15620 26324 15626 26336
rect 16005 26333 16017 26336
rect 16051 26333 16063 26367
rect 16005 26327 16063 26333
rect 17770 26324 17776 26376
rect 17828 26324 17834 26376
rect 17862 26324 17868 26376
rect 17920 26324 17926 26376
rect 17972 26364 18000 26404
rect 18046 26392 18052 26444
rect 18104 26392 18110 26444
rect 18601 26435 18659 26441
rect 18601 26432 18613 26435
rect 18156 26404 18613 26432
rect 18156 26364 18184 26404
rect 18601 26401 18613 26404
rect 18647 26432 18659 26435
rect 18690 26432 18696 26444
rect 18647 26404 18696 26432
rect 18647 26401 18659 26404
rect 18601 26395 18659 26401
rect 18690 26392 18696 26404
rect 18748 26392 18754 26444
rect 18800 26432 18828 26472
rect 18877 26469 18889 26503
rect 18923 26500 18935 26503
rect 19334 26500 19340 26512
rect 18923 26472 19340 26500
rect 18923 26469 18935 26472
rect 18877 26463 18935 26469
rect 19334 26460 19340 26472
rect 19392 26460 19398 26512
rect 20364 26472 20760 26500
rect 20364 26432 20392 26472
rect 18800 26404 20392 26432
rect 17972 26336 18184 26364
rect 18230 26324 18236 26376
rect 18288 26364 18294 26376
rect 18509 26367 18567 26373
rect 18509 26364 18521 26367
rect 18288 26336 18521 26364
rect 18288 26324 18294 26336
rect 18509 26333 18521 26336
rect 18555 26333 18567 26367
rect 18509 26327 18567 26333
rect 19334 26324 19340 26376
rect 19392 26364 19398 26376
rect 19981 26367 20039 26373
rect 19981 26364 19993 26367
rect 19392 26336 19993 26364
rect 19392 26324 19398 26336
rect 19981 26333 19993 26336
rect 20027 26333 20039 26367
rect 19981 26327 20039 26333
rect 20070 26324 20076 26376
rect 20128 26364 20134 26376
rect 20530 26373 20536 26376
rect 20165 26367 20223 26373
rect 20165 26364 20177 26367
rect 20128 26336 20177 26364
rect 20128 26324 20134 26336
rect 20165 26333 20177 26336
rect 20211 26333 20223 26367
rect 20165 26327 20223 26333
rect 20487 26367 20536 26373
rect 20487 26333 20499 26367
rect 20533 26333 20536 26367
rect 20487 26327 20536 26333
rect 20530 26324 20536 26327
rect 20588 26324 20594 26376
rect 20625 26367 20683 26373
rect 20625 26333 20637 26367
rect 20671 26364 20683 26367
rect 20732 26364 20760 26472
rect 21726 26432 21732 26444
rect 20671 26336 20760 26364
rect 21560 26404 21732 26432
rect 20671 26333 20683 26336
rect 20625 26327 20683 26333
rect 16574 26296 16580 26308
rect 15028 26268 16580 26296
rect 16574 26256 16580 26268
rect 16632 26256 16638 26308
rect 19886 26256 19892 26308
rect 19944 26296 19950 26308
rect 20257 26299 20315 26305
rect 20257 26296 20269 26299
rect 19944 26268 20269 26296
rect 19944 26256 19950 26268
rect 20257 26265 20269 26268
rect 20303 26265 20315 26299
rect 20257 26259 20315 26265
rect 20349 26299 20407 26305
rect 20349 26265 20361 26299
rect 20395 26296 20407 26299
rect 21560 26296 21588 26404
rect 21726 26392 21732 26404
rect 21784 26392 21790 26444
rect 22480 26441 22508 26540
rect 22646 26528 22652 26580
rect 22704 26568 22710 26580
rect 25958 26568 25964 26580
rect 22704 26540 25964 26568
rect 22704 26528 22710 26540
rect 25958 26528 25964 26540
rect 26016 26568 26022 26580
rect 28074 26568 28080 26580
rect 26016 26540 28080 26568
rect 26016 26528 26022 26540
rect 28074 26528 28080 26540
rect 28132 26528 28138 26580
rect 28258 26528 28264 26580
rect 28316 26568 28322 26580
rect 30466 26568 30472 26580
rect 28316 26540 30472 26568
rect 28316 26528 28322 26540
rect 30466 26528 30472 26540
rect 30524 26528 30530 26580
rect 30742 26528 30748 26580
rect 30800 26568 30806 26580
rect 30800 26540 32904 26568
rect 30800 26528 30806 26540
rect 23566 26460 23572 26512
rect 23624 26500 23630 26512
rect 23842 26500 23848 26512
rect 23624 26472 23848 26500
rect 23624 26460 23630 26472
rect 23842 26460 23848 26472
rect 23900 26460 23906 26512
rect 24578 26460 24584 26512
rect 24636 26500 24642 26512
rect 30650 26500 30656 26512
rect 24636 26472 27844 26500
rect 24636 26460 24642 26472
rect 22465 26435 22523 26441
rect 22465 26401 22477 26435
rect 22511 26401 22523 26435
rect 22465 26395 22523 26401
rect 26142 26392 26148 26444
rect 26200 26432 26206 26444
rect 27816 26441 27844 26472
rect 28184 26472 30656 26500
rect 27801 26435 27859 26441
rect 26200 26404 26280 26432
rect 26200 26392 26206 26404
rect 21634 26324 21640 26376
rect 21692 26324 21698 26376
rect 21821 26367 21879 26373
rect 21821 26364 21833 26367
rect 21744 26336 21833 26364
rect 20395 26268 21588 26296
rect 20395 26265 20407 26268
rect 20349 26259 20407 26265
rect 5258 26188 5264 26240
rect 5316 26228 5322 26240
rect 11054 26228 11060 26240
rect 5316 26200 11060 26228
rect 5316 26188 5322 26200
rect 11054 26188 11060 26200
rect 11112 26188 11118 26240
rect 11974 26188 11980 26240
rect 12032 26228 12038 26240
rect 12526 26228 12532 26240
rect 12032 26200 12532 26228
rect 12032 26188 12038 26200
rect 12526 26188 12532 26200
rect 12584 26188 12590 26240
rect 12986 26188 12992 26240
rect 13044 26228 13050 26240
rect 16482 26228 16488 26240
rect 13044 26200 16488 26228
rect 13044 26188 13050 26200
rect 16482 26188 16488 26200
rect 16540 26188 16546 26240
rect 16592 26228 16620 26256
rect 17129 26231 17187 26237
rect 17129 26228 17141 26231
rect 16592 26200 17141 26228
rect 17129 26197 17141 26200
rect 17175 26197 17187 26231
rect 17129 26191 17187 26197
rect 17218 26188 17224 26240
rect 17276 26228 17282 26240
rect 17862 26228 17868 26240
rect 17276 26200 17868 26228
rect 17276 26188 17282 26200
rect 17862 26188 17868 26200
rect 17920 26188 17926 26240
rect 18506 26188 18512 26240
rect 18564 26228 18570 26240
rect 21450 26228 21456 26240
rect 18564 26200 21456 26228
rect 18564 26188 18570 26200
rect 21450 26188 21456 26200
rect 21508 26228 21514 26240
rect 21744 26228 21772 26336
rect 21821 26333 21833 26336
rect 21867 26333 21879 26367
rect 21821 26327 21879 26333
rect 22732 26367 22790 26373
rect 22732 26333 22744 26367
rect 22778 26364 22790 26367
rect 23750 26364 23756 26376
rect 22778 26336 23756 26364
rect 22778 26333 22790 26336
rect 22732 26327 22790 26333
rect 23750 26324 23756 26336
rect 23808 26324 23814 26376
rect 24670 26324 24676 26376
rect 24728 26324 24734 26376
rect 24854 26324 24860 26376
rect 24912 26324 24918 26376
rect 26252 26364 26280 26404
rect 27801 26401 27813 26435
rect 27847 26401 27859 26435
rect 27801 26395 27859 26401
rect 28074 26392 28080 26444
rect 28132 26432 28138 26444
rect 28184 26441 28212 26472
rect 30650 26460 30656 26472
rect 30708 26460 30714 26512
rect 31018 26460 31024 26512
rect 31076 26500 31082 26512
rect 32033 26503 32091 26509
rect 32033 26500 32045 26503
rect 31076 26472 32045 26500
rect 31076 26460 31082 26472
rect 32033 26469 32045 26472
rect 32079 26469 32091 26503
rect 32876 26500 32904 26540
rect 32950 26528 32956 26580
rect 33008 26568 33014 26580
rect 35802 26568 35808 26580
rect 33008 26540 35808 26568
rect 33008 26528 33014 26540
rect 35802 26528 35808 26540
rect 35860 26528 35866 26580
rect 36446 26528 36452 26580
rect 36504 26528 36510 26580
rect 35437 26503 35495 26509
rect 32876 26472 35393 26500
rect 32033 26463 32091 26469
rect 28169 26435 28227 26441
rect 28169 26432 28181 26435
rect 28132 26404 28181 26432
rect 28132 26392 28138 26404
rect 28169 26401 28181 26404
rect 28215 26401 28227 26435
rect 28169 26395 28227 26401
rect 28258 26392 28264 26444
rect 28316 26392 28322 26444
rect 28353 26435 28411 26441
rect 28353 26401 28365 26435
rect 28399 26432 28411 26435
rect 28534 26432 28540 26444
rect 28399 26404 28540 26432
rect 28399 26401 28411 26404
rect 28353 26395 28411 26401
rect 28534 26392 28540 26404
rect 28592 26392 28598 26444
rect 28810 26392 28816 26444
rect 28868 26432 28874 26444
rect 33594 26432 33600 26444
rect 28868 26404 30236 26432
rect 28868 26392 28874 26404
rect 26421 26367 26479 26373
rect 26421 26364 26433 26367
rect 26252 26336 26433 26364
rect 26421 26333 26433 26336
rect 26467 26333 26479 26367
rect 26421 26327 26479 26333
rect 28442 26324 28448 26376
rect 28500 26364 28506 26376
rect 28997 26367 29055 26373
rect 28997 26364 29009 26367
rect 28500 26336 29009 26364
rect 28500 26324 28506 26336
rect 28997 26333 29009 26336
rect 29043 26333 29055 26367
rect 28997 26327 29055 26333
rect 29178 26324 29184 26376
rect 29236 26324 29242 26376
rect 29270 26324 29276 26376
rect 29328 26364 29334 26376
rect 30101 26367 30159 26373
rect 30101 26364 30113 26367
rect 29328 26336 30113 26364
rect 29328 26324 29334 26336
rect 30101 26333 30113 26336
rect 30147 26333 30159 26367
rect 30101 26327 30159 26333
rect 22005 26299 22063 26305
rect 22005 26265 22017 26299
rect 22051 26296 22063 26299
rect 22462 26296 22468 26308
rect 22051 26268 22468 26296
rect 22051 26265 22063 26268
rect 22005 26259 22063 26265
rect 22462 26256 22468 26268
rect 22520 26256 22526 26308
rect 23566 26256 23572 26308
rect 23624 26296 23630 26308
rect 25130 26296 25136 26308
rect 23624 26268 25136 26296
rect 23624 26256 23630 26268
rect 25130 26256 25136 26268
rect 25188 26256 25194 26308
rect 25222 26256 25228 26308
rect 25280 26256 25286 26308
rect 25866 26256 25872 26308
rect 25924 26296 25930 26308
rect 26145 26299 26203 26305
rect 26145 26296 26157 26299
rect 25924 26268 26157 26296
rect 25924 26256 25930 26268
rect 26145 26265 26157 26268
rect 26191 26296 26203 26299
rect 26234 26296 26240 26308
rect 26191 26268 26240 26296
rect 26191 26265 26203 26268
rect 26145 26259 26203 26265
rect 26234 26256 26240 26268
rect 26292 26256 26298 26308
rect 26326 26256 26332 26308
rect 26384 26256 26390 26308
rect 26510 26256 26516 26308
rect 26568 26256 26574 26308
rect 26881 26299 26939 26305
rect 26881 26265 26893 26299
rect 26927 26296 26939 26299
rect 26970 26296 26976 26308
rect 26927 26268 26976 26296
rect 26927 26265 26939 26268
rect 26881 26259 26939 26265
rect 26970 26256 26976 26268
rect 27028 26256 27034 26308
rect 27062 26256 27068 26308
rect 27120 26296 27126 26308
rect 29089 26299 29147 26305
rect 29089 26296 29101 26299
rect 27120 26268 29101 26296
rect 27120 26256 27126 26268
rect 29089 26265 29101 26268
rect 29135 26265 29147 26299
rect 29089 26259 29147 26265
rect 29730 26256 29736 26308
rect 29788 26256 29794 26308
rect 29917 26299 29975 26305
rect 29917 26265 29929 26299
rect 29963 26296 29975 26299
rect 30208 26296 30236 26404
rect 30576 26404 33600 26432
rect 30576 26373 30604 26404
rect 33594 26392 33600 26404
rect 33652 26392 33658 26444
rect 33778 26392 33784 26444
rect 33836 26432 33842 26444
rect 34057 26435 34115 26441
rect 34057 26432 34069 26435
rect 33836 26404 34069 26432
rect 33836 26392 33842 26404
rect 34057 26401 34069 26404
rect 34103 26401 34115 26435
rect 34057 26395 34115 26401
rect 30742 26373 30748 26376
rect 30561 26367 30619 26373
rect 30561 26333 30573 26367
rect 30607 26333 30619 26367
rect 30561 26327 30619 26333
rect 30709 26367 30748 26373
rect 30709 26333 30721 26367
rect 30709 26327 30748 26333
rect 30742 26324 30748 26327
rect 30800 26324 30806 26376
rect 30926 26324 30932 26376
rect 30984 26324 30990 26376
rect 31067 26367 31125 26373
rect 31067 26333 31079 26367
rect 31113 26364 31125 26367
rect 31202 26364 31208 26376
rect 31113 26336 31208 26364
rect 31113 26333 31125 26336
rect 31067 26327 31125 26333
rect 31202 26324 31208 26336
rect 31260 26324 31266 26376
rect 31386 26324 31392 26376
rect 31444 26364 31450 26376
rect 31849 26367 31907 26373
rect 31849 26364 31861 26367
rect 31444 26336 31861 26364
rect 31444 26324 31450 26336
rect 31849 26333 31861 26336
rect 31895 26333 31907 26367
rect 31849 26327 31907 26333
rect 32858 26324 32864 26376
rect 32916 26364 32922 26376
rect 33502 26364 33508 26376
rect 32916 26336 33508 26364
rect 32916 26324 32922 26336
rect 33502 26324 33508 26336
rect 33560 26324 33566 26376
rect 33870 26324 33876 26376
rect 33928 26324 33934 26376
rect 34882 26324 34888 26376
rect 34940 26324 34946 26376
rect 35253 26367 35311 26373
rect 35253 26333 35265 26367
rect 35299 26333 35311 26367
rect 35365 26364 35393 26472
rect 35437 26469 35449 26503
rect 35483 26469 35495 26503
rect 35437 26463 35495 26469
rect 35452 26432 35480 26463
rect 35894 26460 35900 26512
rect 35952 26500 35958 26512
rect 35952 26472 36124 26500
rect 35952 26460 35958 26472
rect 35802 26432 35808 26444
rect 35452 26404 35808 26432
rect 35802 26392 35808 26404
rect 35860 26392 35866 26444
rect 36096 26432 36124 26472
rect 36538 26432 36544 26444
rect 36096 26404 36544 26432
rect 35365 26336 35849 26364
rect 35253 26327 35311 26333
rect 30837 26299 30895 26305
rect 30837 26296 30849 26299
rect 29963 26268 30236 26296
rect 30760 26268 30849 26296
rect 29963 26265 29975 26268
rect 29917 26259 29975 26265
rect 30760 26240 30788 26268
rect 30837 26265 30849 26268
rect 30883 26265 30895 26299
rect 30837 26259 30895 26265
rect 31570 26256 31576 26308
rect 31628 26296 31634 26308
rect 31665 26299 31723 26305
rect 31665 26296 31677 26299
rect 31628 26268 31677 26296
rect 31628 26256 31634 26268
rect 31665 26265 31677 26268
rect 31711 26265 31723 26299
rect 31665 26259 31723 26265
rect 32398 26256 32404 26308
rect 32456 26296 32462 26308
rect 32493 26299 32551 26305
rect 32493 26296 32505 26299
rect 32456 26268 32505 26296
rect 32456 26256 32462 26268
rect 32493 26265 32505 26268
rect 32539 26265 32551 26299
rect 32493 26259 32551 26265
rect 33042 26256 33048 26308
rect 33100 26296 33106 26308
rect 33229 26299 33287 26305
rect 33229 26296 33241 26299
rect 33100 26268 33241 26296
rect 33100 26256 33106 26268
rect 33229 26265 33241 26268
rect 33275 26265 33287 26299
rect 33229 26259 33287 26265
rect 35066 26256 35072 26308
rect 35124 26256 35130 26308
rect 35158 26256 35164 26308
rect 35216 26256 35222 26308
rect 35268 26296 35296 26327
rect 35342 26296 35348 26308
rect 35268 26268 35348 26296
rect 35342 26256 35348 26268
rect 35400 26256 35406 26308
rect 35821 26296 35849 26336
rect 35894 26324 35900 26376
rect 35952 26324 35958 26376
rect 36096 26373 36124 26404
rect 36538 26392 36544 26404
rect 36596 26392 36602 26444
rect 36081 26367 36139 26373
rect 36081 26333 36093 26367
rect 36127 26333 36139 26367
rect 36081 26327 36139 26333
rect 36170 26324 36176 26376
rect 36228 26324 36234 26376
rect 36262 26324 36268 26376
rect 36320 26324 36326 26376
rect 36906 26324 36912 26376
rect 36964 26324 36970 26376
rect 36814 26296 36820 26308
rect 35821 26268 36820 26296
rect 36814 26256 36820 26268
rect 36872 26256 36878 26308
rect 37176 26299 37234 26305
rect 37176 26265 37188 26299
rect 37222 26296 37234 26299
rect 37458 26296 37464 26308
rect 37222 26268 37464 26296
rect 37222 26265 37234 26268
rect 37176 26259 37234 26265
rect 37458 26256 37464 26268
rect 37516 26256 37522 26308
rect 21508 26200 21772 26228
rect 21508 26188 21514 26200
rect 25498 26188 25504 26240
rect 25556 26228 25562 26240
rect 27706 26228 27712 26240
rect 25556 26200 27712 26228
rect 25556 26188 25562 26200
rect 27706 26188 27712 26200
rect 27764 26188 27770 26240
rect 27890 26188 27896 26240
rect 27948 26228 27954 26240
rect 28902 26228 28908 26240
rect 27948 26200 28908 26228
rect 27948 26188 27954 26200
rect 28902 26188 28908 26200
rect 28960 26228 28966 26240
rect 30466 26228 30472 26240
rect 28960 26200 30472 26228
rect 28960 26188 28966 26200
rect 30466 26188 30472 26200
rect 30524 26188 30530 26240
rect 30742 26188 30748 26240
rect 30800 26188 30806 26240
rect 31202 26188 31208 26240
rect 31260 26188 31266 26240
rect 32858 26188 32864 26240
rect 32916 26228 32922 26240
rect 34790 26228 34796 26240
rect 32916 26200 34796 26228
rect 32916 26188 32922 26200
rect 34790 26188 34796 26200
rect 34848 26228 34854 26240
rect 35894 26228 35900 26240
rect 34848 26200 35900 26228
rect 34848 26188 34854 26200
rect 35894 26188 35900 26200
rect 35952 26228 35958 26240
rect 37734 26228 37740 26240
rect 35952 26200 37740 26228
rect 35952 26188 35958 26200
rect 37734 26188 37740 26200
rect 37792 26228 37798 26240
rect 38289 26231 38347 26237
rect 38289 26228 38301 26231
rect 37792 26200 38301 26228
rect 37792 26188 37798 26200
rect 38289 26197 38301 26200
rect 38335 26197 38347 26231
rect 38289 26191 38347 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 2406 25984 2412 26036
rect 2464 26024 2470 26036
rect 2464 25996 10272 26024
rect 2464 25984 2470 25996
rect 8656 25959 8714 25965
rect 8656 25925 8668 25959
rect 8702 25956 8714 25959
rect 10134 25956 10140 25968
rect 8702 25928 10140 25956
rect 8702 25925 8714 25928
rect 8656 25919 8714 25925
rect 10134 25916 10140 25928
rect 10192 25916 10198 25968
rect 10244 25956 10272 25996
rect 10962 25984 10968 26036
rect 11020 25984 11026 26036
rect 11054 25984 11060 26036
rect 11112 26024 11118 26036
rect 12986 26024 12992 26036
rect 11112 25996 12992 26024
rect 11112 25984 11118 25996
rect 12986 25984 12992 25996
rect 13044 25984 13050 26036
rect 13081 26027 13139 26033
rect 13081 25993 13093 26027
rect 13127 26024 13139 26027
rect 15838 26024 15844 26036
rect 13127 25996 15844 26024
rect 13127 25993 13139 25996
rect 13081 25987 13139 25993
rect 15838 25984 15844 25996
rect 15896 25984 15902 26036
rect 16482 25984 16488 26036
rect 16540 26024 16546 26036
rect 18506 26024 18512 26036
rect 16540 25996 18512 26024
rect 16540 25984 16546 25996
rect 18506 25984 18512 25996
rect 18564 25984 18570 26036
rect 18782 25984 18788 26036
rect 18840 25984 18846 26036
rect 19058 25984 19064 26036
rect 19116 26024 19122 26036
rect 19116 25996 20484 26024
rect 19116 25984 19122 25996
rect 10244 25928 12434 25956
rect 8294 25848 8300 25900
rect 8352 25888 8358 25900
rect 8389 25891 8447 25897
rect 8389 25888 8401 25891
rect 8352 25860 8401 25888
rect 8352 25848 8358 25860
rect 8389 25857 8401 25860
rect 8435 25857 8447 25891
rect 8389 25851 8447 25857
rect 10410 25848 10416 25900
rect 10468 25848 10474 25900
rect 10594 25848 10600 25900
rect 10652 25848 10658 25900
rect 10689 25891 10747 25897
rect 10689 25857 10701 25891
rect 10735 25857 10747 25891
rect 10689 25851 10747 25857
rect 10781 25891 10839 25897
rect 10781 25857 10793 25891
rect 10827 25888 10839 25891
rect 10870 25888 10876 25900
rect 10827 25860 10876 25888
rect 10827 25857 10839 25860
rect 10781 25851 10839 25857
rect 10704 25820 10732 25851
rect 10870 25848 10876 25860
rect 10928 25848 10934 25900
rect 11698 25848 11704 25900
rect 11756 25848 11762 25900
rect 11974 25897 11980 25900
rect 11968 25888 11980 25897
rect 11935 25860 11980 25888
rect 11968 25851 11980 25860
rect 11974 25848 11980 25851
rect 12032 25848 12038 25900
rect 12406 25888 12434 25928
rect 12710 25916 12716 25968
rect 12768 25956 12774 25968
rect 13633 25959 13691 25965
rect 13633 25956 13645 25959
rect 12768 25928 13645 25956
rect 12768 25916 12774 25928
rect 13633 25925 13645 25928
rect 13679 25925 13691 25959
rect 13633 25919 13691 25925
rect 14734 25916 14740 25968
rect 14792 25956 14798 25968
rect 14792 25928 17724 25956
rect 14792 25916 14798 25928
rect 13541 25891 13599 25897
rect 12406 25860 12756 25888
rect 11330 25820 11336 25832
rect 10704 25792 11336 25820
rect 11330 25780 11336 25792
rect 11388 25780 11394 25832
rect 12728 25820 12756 25860
rect 13541 25857 13553 25891
rect 13587 25888 13599 25891
rect 13722 25888 13728 25900
rect 13587 25860 13728 25888
rect 13587 25857 13599 25860
rect 13541 25851 13599 25857
rect 13722 25848 13728 25860
rect 13780 25848 13786 25900
rect 14090 25888 14096 25900
rect 13832 25860 14096 25888
rect 13832 25820 13860 25860
rect 14090 25848 14096 25860
rect 14148 25848 14154 25900
rect 14182 25848 14188 25900
rect 14240 25848 14246 25900
rect 14369 25891 14427 25897
rect 14369 25857 14381 25891
rect 14415 25888 14427 25891
rect 14458 25888 14464 25900
rect 14415 25860 14464 25888
rect 14415 25857 14427 25860
rect 14369 25851 14427 25857
rect 14458 25848 14464 25860
rect 14516 25848 14522 25900
rect 15096 25891 15154 25897
rect 15096 25857 15108 25891
rect 15142 25888 15154 25891
rect 15562 25888 15568 25900
rect 15142 25860 15568 25888
rect 15142 25857 15154 25860
rect 15096 25851 15154 25857
rect 15562 25848 15568 25860
rect 15620 25848 15626 25900
rect 17034 25848 17040 25900
rect 17092 25888 17098 25900
rect 17589 25891 17647 25897
rect 17589 25888 17601 25891
rect 17092 25860 17601 25888
rect 17092 25848 17098 25860
rect 17589 25857 17601 25860
rect 17635 25857 17647 25891
rect 17589 25851 17647 25857
rect 12728 25792 13860 25820
rect 13906 25780 13912 25832
rect 13964 25820 13970 25832
rect 14829 25823 14887 25829
rect 14829 25820 14841 25823
rect 13964 25792 14841 25820
rect 13964 25780 13970 25792
rect 14829 25789 14841 25792
rect 14875 25789 14887 25823
rect 14829 25783 14887 25789
rect 9769 25755 9827 25761
rect 9769 25721 9781 25755
rect 9815 25752 9827 25755
rect 9858 25752 9864 25764
rect 9815 25724 9864 25752
rect 9815 25721 9827 25724
rect 9769 25715 9827 25721
rect 9858 25712 9864 25724
rect 9916 25712 9922 25764
rect 14277 25755 14335 25761
rect 14277 25752 14289 25755
rect 13004 25724 14289 25752
rect 11698 25644 11704 25696
rect 11756 25684 11762 25696
rect 13004 25684 13032 25724
rect 14277 25721 14289 25724
rect 14323 25721 14335 25755
rect 17586 25752 17592 25764
rect 14277 25715 14335 25721
rect 15764 25724 17592 25752
rect 11756 25656 13032 25684
rect 11756 25644 11762 25656
rect 14090 25644 14096 25696
rect 14148 25684 14154 25696
rect 15764 25684 15792 25724
rect 17586 25712 17592 25724
rect 17644 25712 17650 25764
rect 14148 25656 15792 25684
rect 14148 25644 14154 25656
rect 16206 25644 16212 25696
rect 16264 25644 16270 25696
rect 17402 25644 17408 25696
rect 17460 25644 17466 25696
rect 17696 25684 17724 25928
rect 17954 25916 17960 25968
rect 18012 25956 18018 25968
rect 20456 25965 20484 25996
rect 21928 25996 22140 26024
rect 19245 25959 19303 25965
rect 19245 25956 19257 25959
rect 18012 25928 19257 25956
rect 18012 25916 18018 25928
rect 19245 25925 19257 25928
rect 19291 25925 19303 25959
rect 19245 25919 19303 25925
rect 20441 25959 20499 25965
rect 20441 25925 20453 25959
rect 20487 25956 20499 25959
rect 20530 25956 20536 25968
rect 20487 25928 20536 25956
rect 20487 25925 20499 25928
rect 20441 25919 20499 25925
rect 20530 25916 20536 25928
rect 20588 25916 20594 25968
rect 20901 25959 20959 25965
rect 20901 25925 20913 25959
rect 20947 25956 20959 25959
rect 21928 25956 21956 25996
rect 20947 25928 21956 25956
rect 20947 25925 20959 25928
rect 20901 25919 20959 25925
rect 22002 25916 22008 25968
rect 22060 25916 22066 25968
rect 22112 25956 22140 25996
rect 22186 25984 22192 26036
rect 22244 25984 22250 26036
rect 22925 26027 22983 26033
rect 22925 25993 22937 26027
rect 22971 26024 22983 26027
rect 32858 26024 32864 26036
rect 22971 25996 27200 26024
rect 22971 25993 22983 25996
rect 22925 25987 22983 25993
rect 23753 25959 23811 25965
rect 23753 25956 23765 25959
rect 22112 25928 23765 25956
rect 23753 25925 23765 25928
rect 23799 25925 23811 25959
rect 23753 25919 23811 25925
rect 24673 25959 24731 25965
rect 24673 25925 24685 25959
rect 24719 25956 24731 25959
rect 26694 25956 26700 25968
rect 24719 25928 26700 25956
rect 24719 25925 24731 25928
rect 24673 25919 24731 25925
rect 26694 25916 26700 25928
rect 26752 25916 26758 25968
rect 17773 25891 17831 25897
rect 17773 25857 17785 25891
rect 17819 25857 17831 25891
rect 17773 25851 17831 25857
rect 17788 25820 17816 25851
rect 17862 25848 17868 25900
rect 17920 25848 17926 25900
rect 18598 25848 18604 25900
rect 18656 25848 18662 25900
rect 19426 25848 19432 25900
rect 19484 25848 19490 25900
rect 19610 25848 19616 25900
rect 19668 25848 19674 25900
rect 20162 25848 20168 25900
rect 20220 25848 20226 25900
rect 20346 25848 20352 25900
rect 20404 25848 20410 25900
rect 20622 25848 20628 25900
rect 20680 25888 20686 25900
rect 21177 25891 21235 25897
rect 20680 25860 21128 25888
rect 20680 25848 20686 25860
rect 17788 25792 17954 25820
rect 17926 25752 17954 25792
rect 18414 25780 18420 25832
rect 18472 25780 18478 25832
rect 19058 25780 19064 25832
rect 19116 25820 19122 25832
rect 19334 25820 19340 25832
rect 19116 25792 19340 25820
rect 19116 25780 19122 25792
rect 19334 25780 19340 25792
rect 19392 25780 19398 25832
rect 19886 25820 19892 25832
rect 19444 25792 19892 25820
rect 19242 25752 19248 25764
rect 17926 25724 19248 25752
rect 19242 25712 19248 25724
rect 19300 25752 19306 25764
rect 19444 25752 19472 25792
rect 19886 25780 19892 25792
rect 19944 25780 19950 25832
rect 20990 25780 20996 25832
rect 21048 25780 21054 25832
rect 21100 25820 21128 25860
rect 21177 25857 21189 25891
rect 21223 25888 21235 25891
rect 21726 25888 21732 25900
rect 21223 25860 21732 25888
rect 21223 25857 21235 25860
rect 21177 25851 21235 25857
rect 21726 25848 21732 25860
rect 21784 25848 21790 25900
rect 22281 25891 22339 25897
rect 22281 25857 22293 25891
rect 22327 25857 22339 25891
rect 23937 25891 23995 25897
rect 23937 25888 23949 25891
rect 22281 25851 22339 25857
rect 22756 25860 23949 25888
rect 22296 25820 22324 25851
rect 22756 25829 22784 25860
rect 23937 25857 23949 25860
rect 23983 25857 23995 25891
rect 23937 25851 23995 25857
rect 25958 25848 25964 25900
rect 26016 25888 26022 25900
rect 27172 25897 27200 25996
rect 28828 25996 32864 26024
rect 26053 25891 26111 25897
rect 26053 25888 26065 25891
rect 26016 25860 26065 25888
rect 26016 25848 26022 25860
rect 26053 25857 26065 25860
rect 26099 25857 26111 25891
rect 27157 25891 27215 25897
rect 26053 25851 26111 25857
rect 26160 25860 27108 25888
rect 22741 25823 22799 25829
rect 22741 25820 22753 25823
rect 21100 25792 22324 25820
rect 22388 25792 22753 25820
rect 20346 25752 20352 25764
rect 19300 25724 19472 25752
rect 19536 25724 20352 25752
rect 19300 25712 19306 25724
rect 19536 25684 19564 25724
rect 20346 25712 20352 25724
rect 20404 25712 20410 25764
rect 20530 25712 20536 25764
rect 20588 25752 20594 25764
rect 21361 25755 21419 25761
rect 21361 25752 21373 25755
rect 20588 25724 21373 25752
rect 20588 25712 20594 25724
rect 21361 25721 21373 25724
rect 21407 25721 21419 25755
rect 21361 25715 21419 25721
rect 22005 25755 22063 25761
rect 22005 25721 22017 25755
rect 22051 25752 22063 25755
rect 22094 25752 22100 25764
rect 22051 25724 22100 25752
rect 22051 25721 22063 25724
rect 22005 25715 22063 25721
rect 22094 25712 22100 25724
rect 22152 25712 22158 25764
rect 22186 25712 22192 25764
rect 22244 25752 22250 25764
rect 22388 25752 22416 25792
rect 22741 25789 22753 25792
rect 22787 25789 22799 25823
rect 22741 25783 22799 25789
rect 23109 25823 23167 25829
rect 23109 25789 23121 25823
rect 23155 25789 23167 25823
rect 23109 25783 23167 25789
rect 23124 25752 23152 25783
rect 23198 25780 23204 25832
rect 23256 25820 23262 25832
rect 24213 25823 24271 25829
rect 24213 25820 24225 25823
rect 23256 25792 24225 25820
rect 23256 25780 23262 25792
rect 24213 25789 24225 25792
rect 24259 25789 24271 25823
rect 24213 25783 24271 25789
rect 24762 25780 24768 25832
rect 24820 25820 24826 25832
rect 24857 25823 24915 25829
rect 24857 25820 24869 25823
rect 24820 25792 24869 25820
rect 24820 25780 24826 25792
rect 24857 25789 24869 25792
rect 24903 25789 24915 25823
rect 24857 25783 24915 25789
rect 25041 25823 25099 25829
rect 25041 25789 25053 25823
rect 25087 25820 25099 25823
rect 26160 25820 26188 25860
rect 25087 25792 26188 25820
rect 26237 25823 26295 25829
rect 25087 25789 25099 25792
rect 25041 25783 25099 25789
rect 26237 25789 26249 25823
rect 26283 25820 26295 25823
rect 26694 25820 26700 25832
rect 26283 25792 26700 25820
rect 26283 25789 26295 25792
rect 26237 25783 26295 25789
rect 26694 25780 26700 25792
rect 26752 25780 26758 25832
rect 27080 25820 27108 25860
rect 27157 25857 27169 25891
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 27614 25848 27620 25900
rect 27672 25848 27678 25900
rect 27982 25848 27988 25900
rect 28040 25848 28046 25900
rect 28828 25897 28856 25996
rect 32858 25984 32864 25996
rect 32916 25984 32922 26036
rect 32950 25984 32956 26036
rect 33008 26024 33014 26036
rect 35066 26024 35072 26036
rect 33008 25996 35072 26024
rect 33008 25984 33014 25996
rect 35066 25984 35072 25996
rect 35124 25984 35130 26036
rect 35158 25984 35164 26036
rect 35216 26024 35222 26036
rect 36354 26024 36360 26036
rect 35216 25996 36360 26024
rect 35216 25984 35222 25996
rect 36354 25984 36360 25996
rect 36412 25984 36418 26036
rect 37458 25984 37464 26036
rect 37516 25984 37522 26036
rect 29089 25959 29147 25965
rect 29089 25925 29101 25959
rect 29135 25956 29147 25959
rect 29638 25956 29644 25968
rect 29135 25928 29644 25956
rect 29135 25925 29147 25928
rect 29089 25919 29147 25925
rect 29638 25916 29644 25928
rect 29696 25916 29702 25968
rect 30190 25956 30196 25968
rect 30024 25928 30196 25956
rect 28813 25891 28871 25897
rect 28813 25857 28825 25891
rect 28859 25857 28871 25891
rect 28813 25851 28871 25857
rect 28902 25848 28908 25900
rect 28960 25888 28966 25900
rect 28997 25891 29055 25897
rect 28997 25888 29009 25891
rect 28960 25860 29009 25888
rect 28960 25848 28966 25860
rect 28997 25857 29009 25860
rect 29043 25857 29055 25891
rect 28997 25851 29055 25857
rect 29178 25848 29184 25900
rect 29236 25848 29242 25900
rect 30024 25897 30052 25928
rect 30190 25916 30196 25928
rect 30248 25956 30254 25968
rect 31754 25956 31760 25968
rect 30248 25928 31760 25956
rect 30248 25916 30254 25928
rect 31754 25916 31760 25928
rect 31812 25956 31818 25968
rect 32214 25956 32220 25968
rect 31812 25928 32220 25956
rect 31812 25916 31818 25928
rect 32214 25916 32220 25928
rect 32272 25916 32278 25968
rect 32398 25916 32404 25968
rect 32456 25956 32462 25968
rect 32456 25928 32628 25956
rect 32456 25916 32462 25928
rect 30009 25891 30067 25897
rect 30009 25857 30021 25891
rect 30055 25857 30067 25891
rect 30837 25891 30895 25897
rect 30837 25888 30849 25891
rect 30009 25851 30067 25857
rect 30668 25860 30849 25888
rect 27706 25820 27712 25832
rect 27080 25792 27712 25820
rect 27706 25780 27712 25792
rect 27764 25820 27770 25832
rect 27890 25820 27896 25832
rect 27764 25792 27896 25820
rect 27764 25780 27770 25792
rect 27890 25780 27896 25792
rect 27948 25780 27954 25832
rect 28166 25780 28172 25832
rect 28224 25780 28230 25832
rect 28718 25780 28724 25832
rect 28776 25820 28782 25832
rect 30668 25820 30696 25860
rect 30837 25857 30849 25860
rect 30883 25888 30895 25891
rect 32490 25888 32496 25900
rect 30883 25860 32496 25888
rect 30883 25857 30895 25860
rect 30837 25851 30895 25857
rect 32490 25848 32496 25860
rect 32548 25848 32554 25900
rect 28776 25792 30696 25820
rect 28776 25780 28782 25792
rect 30742 25780 30748 25832
rect 30800 25780 30806 25832
rect 31297 25823 31355 25829
rect 31297 25789 31309 25823
rect 31343 25789 31355 25823
rect 31297 25783 31355 25789
rect 22244 25724 22416 25752
rect 22572 25724 23152 25752
rect 22244 25712 22250 25724
rect 17696 25656 19564 25684
rect 19978 25644 19984 25696
rect 20036 25684 20042 25696
rect 20162 25684 20168 25696
rect 20036 25656 20168 25684
rect 20036 25644 20042 25656
rect 20162 25644 20168 25656
rect 20220 25644 20226 25696
rect 20898 25644 20904 25696
rect 20956 25644 20962 25696
rect 20990 25644 20996 25696
rect 21048 25684 21054 25696
rect 21266 25684 21272 25696
rect 21048 25656 21272 25684
rect 21048 25644 21054 25656
rect 21266 25644 21272 25656
rect 21324 25684 21330 25696
rect 22572 25684 22600 25724
rect 23382 25712 23388 25764
rect 23440 25752 23446 25764
rect 24118 25752 24124 25764
rect 23440 25724 24124 25752
rect 23440 25712 23446 25724
rect 24118 25712 24124 25724
rect 24176 25712 24182 25764
rect 24673 25755 24731 25761
rect 24673 25721 24685 25755
rect 24719 25752 24731 25755
rect 26326 25752 26332 25764
rect 24719 25724 26332 25752
rect 24719 25721 24731 25724
rect 24673 25715 24731 25721
rect 26326 25712 26332 25724
rect 26384 25712 26390 25764
rect 26712 25752 26740 25780
rect 30190 25752 30196 25764
rect 26712 25724 30196 25752
rect 30190 25712 30196 25724
rect 30248 25712 30254 25764
rect 30558 25712 30564 25764
rect 30616 25752 30622 25764
rect 31312 25752 31340 25783
rect 31386 25780 31392 25832
rect 31444 25820 31450 25832
rect 32600 25820 32628 25928
rect 33042 25916 33048 25968
rect 33100 25956 33106 25968
rect 36906 25956 36912 25968
rect 33100 25928 35204 25956
rect 33100 25916 33106 25928
rect 32766 25848 32772 25900
rect 32824 25888 32830 25900
rect 33781 25891 33839 25897
rect 33781 25888 33793 25891
rect 32824 25860 33793 25888
rect 32824 25848 32830 25860
rect 33781 25857 33793 25860
rect 33827 25857 33839 25891
rect 33781 25851 33839 25857
rect 33962 25848 33968 25900
rect 34020 25888 34026 25900
rect 34057 25891 34115 25897
rect 34057 25888 34069 25891
rect 34020 25860 34069 25888
rect 34020 25848 34026 25860
rect 34057 25857 34069 25860
rect 34103 25857 34115 25891
rect 34057 25851 34115 25857
rect 31444 25792 32628 25820
rect 33229 25823 33287 25829
rect 31444 25780 31450 25792
rect 33229 25789 33241 25823
rect 33275 25820 33287 25823
rect 33275 25792 34376 25820
rect 33275 25789 33287 25792
rect 33229 25783 33287 25789
rect 30616 25724 31340 25752
rect 30616 25712 30622 25724
rect 32398 25712 32404 25764
rect 32456 25752 32462 25764
rect 33870 25752 33876 25764
rect 32456 25724 33876 25752
rect 32456 25712 32462 25724
rect 33870 25712 33876 25724
rect 33928 25712 33934 25764
rect 21324 25656 22600 25684
rect 21324 25644 21330 25656
rect 22738 25644 22744 25696
rect 22796 25684 22802 25696
rect 23109 25687 23167 25693
rect 23109 25684 23121 25687
rect 22796 25656 23121 25684
rect 22796 25644 22802 25656
rect 23109 25653 23121 25656
rect 23155 25653 23167 25687
rect 23109 25647 23167 25653
rect 24949 25687 25007 25693
rect 24949 25653 24961 25687
rect 24995 25684 25007 25687
rect 26878 25684 26884 25696
rect 24995 25656 26884 25684
rect 24995 25653 25007 25656
rect 24949 25647 25007 25653
rect 26878 25644 26884 25656
rect 26936 25644 26942 25696
rect 27982 25644 27988 25696
rect 28040 25684 28046 25696
rect 28350 25684 28356 25696
rect 28040 25656 28356 25684
rect 28040 25644 28046 25656
rect 28350 25644 28356 25656
rect 28408 25644 28414 25696
rect 29365 25687 29423 25693
rect 29365 25653 29377 25687
rect 29411 25684 29423 25687
rect 30374 25684 30380 25696
rect 29411 25656 30380 25684
rect 29411 25653 29423 25656
rect 29365 25647 29423 25653
rect 30374 25644 30380 25656
rect 30432 25644 30438 25696
rect 30466 25644 30472 25696
rect 30524 25684 30530 25696
rect 32214 25684 32220 25696
rect 30524 25656 32220 25684
rect 30524 25644 30530 25656
rect 32214 25644 32220 25656
rect 32272 25684 32278 25696
rect 33962 25684 33968 25696
rect 32272 25656 33968 25684
rect 32272 25644 32278 25656
rect 33962 25644 33968 25656
rect 34020 25644 34026 25696
rect 34348 25684 34376 25792
rect 34422 25780 34428 25832
rect 34480 25820 34486 25832
rect 35066 25820 35072 25832
rect 34480 25792 35072 25820
rect 34480 25780 34486 25792
rect 35066 25780 35072 25792
rect 35124 25780 35130 25832
rect 35176 25820 35204 25928
rect 35452 25928 36912 25956
rect 35452 25897 35480 25928
rect 36906 25916 36912 25928
rect 36964 25916 36970 25968
rect 37366 25916 37372 25968
rect 37424 25956 37430 25968
rect 37424 25928 37596 25956
rect 37424 25916 37430 25928
rect 35437 25891 35495 25897
rect 35437 25857 35449 25891
rect 35483 25857 35495 25891
rect 35437 25851 35495 25857
rect 35704 25891 35762 25897
rect 35704 25857 35716 25891
rect 35750 25888 35762 25891
rect 37568 25888 37596 25928
rect 37734 25916 37740 25968
rect 37792 25956 37798 25968
rect 37829 25959 37887 25965
rect 37829 25956 37841 25959
rect 37792 25928 37841 25956
rect 37792 25916 37798 25928
rect 37829 25925 37841 25928
rect 37875 25925 37887 25959
rect 37829 25919 37887 25925
rect 37921 25891 37979 25897
rect 37921 25888 37933 25891
rect 35750 25860 37504 25888
rect 37568 25860 37933 25888
rect 35750 25857 35762 25860
rect 35704 25851 35762 25857
rect 35452 25820 35480 25851
rect 35176 25792 35480 25820
rect 37476 25752 37504 25860
rect 37921 25857 37933 25860
rect 37967 25857 37979 25891
rect 37921 25851 37979 25857
rect 38010 25780 38016 25832
rect 38068 25780 38074 25832
rect 38562 25752 38568 25764
rect 37476 25724 38568 25752
rect 38562 25712 38568 25724
rect 38620 25712 38626 25764
rect 36722 25684 36728 25696
rect 34348 25656 36728 25684
rect 36722 25644 36728 25656
rect 36780 25644 36786 25696
rect 36814 25644 36820 25696
rect 36872 25644 36878 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 13265 25483 13323 25489
rect 13265 25449 13277 25483
rect 13311 25480 13323 25483
rect 15470 25480 15476 25492
rect 13311 25452 15476 25480
rect 13311 25449 13323 25452
rect 13265 25443 13323 25449
rect 15470 25440 15476 25452
rect 15528 25440 15534 25492
rect 15562 25440 15568 25492
rect 15620 25440 15626 25492
rect 16574 25440 16580 25492
rect 16632 25440 16638 25492
rect 17034 25440 17040 25492
rect 17092 25440 17098 25492
rect 18785 25483 18843 25489
rect 18785 25449 18797 25483
rect 18831 25480 18843 25483
rect 20438 25480 20444 25492
rect 18831 25452 20444 25480
rect 18831 25449 18843 25452
rect 18785 25443 18843 25449
rect 20438 25440 20444 25452
rect 20496 25440 20502 25492
rect 20622 25440 20628 25492
rect 20680 25480 20686 25492
rect 23566 25480 23572 25492
rect 20680 25452 23572 25480
rect 20680 25440 20686 25452
rect 23566 25440 23572 25452
rect 23624 25440 23630 25492
rect 23753 25483 23811 25489
rect 23753 25449 23765 25483
rect 23799 25480 23811 25483
rect 25682 25480 25688 25492
rect 23799 25452 25688 25480
rect 23799 25449 23811 25452
rect 23753 25443 23811 25449
rect 25682 25440 25688 25452
rect 25740 25440 25746 25492
rect 25866 25440 25872 25492
rect 25924 25440 25930 25492
rect 28092 25452 28488 25480
rect 10134 25372 10140 25424
rect 10192 25412 10198 25424
rect 10192 25384 12572 25412
rect 10192 25372 10198 25384
rect 9490 25304 9496 25356
rect 9548 25344 9554 25356
rect 9585 25347 9643 25353
rect 9585 25344 9597 25347
rect 9548 25316 9597 25344
rect 9548 25304 9554 25316
rect 9585 25313 9597 25316
rect 9631 25313 9643 25347
rect 9585 25307 9643 25313
rect 9769 25347 9827 25353
rect 9769 25313 9781 25347
rect 9815 25344 9827 25347
rect 10502 25344 10508 25356
rect 9815 25316 10508 25344
rect 9815 25313 9827 25316
rect 9769 25307 9827 25313
rect 10502 25304 10508 25316
rect 10560 25344 10566 25356
rect 10560 25316 10640 25344
rect 10560 25304 10566 25316
rect 8846 25236 8852 25288
rect 8904 25276 8910 25288
rect 10612 25285 10640 25316
rect 11422 25304 11428 25356
rect 11480 25344 11486 25356
rect 12544 25344 12572 25384
rect 13906 25372 13912 25424
rect 13964 25412 13970 25424
rect 14734 25412 14740 25424
rect 13964 25384 14740 25412
rect 13964 25372 13970 25384
rect 14734 25372 14740 25384
rect 14792 25372 14798 25424
rect 15102 25372 15108 25424
rect 15160 25412 15166 25424
rect 19794 25412 19800 25424
rect 15160 25384 19800 25412
rect 15160 25372 15166 25384
rect 19794 25372 19800 25384
rect 19852 25372 19858 25424
rect 19886 25372 19892 25424
rect 19944 25412 19950 25424
rect 23658 25412 23664 25424
rect 19944 25384 23664 25412
rect 19944 25372 19950 25384
rect 15194 25344 15200 25356
rect 11480 25316 12434 25344
rect 12544 25316 15200 25344
rect 11480 25304 11486 25316
rect 10413 25279 10471 25285
rect 10413 25276 10425 25279
rect 8904 25248 10425 25276
rect 8904 25236 8910 25248
rect 10413 25245 10425 25248
rect 10459 25245 10471 25279
rect 10413 25239 10471 25245
rect 10597 25279 10655 25285
rect 10597 25245 10609 25279
rect 10643 25245 10655 25279
rect 10597 25239 10655 25245
rect 10612 25208 10640 25239
rect 10870 25236 10876 25288
rect 10928 25276 10934 25288
rect 11517 25279 11575 25285
rect 11517 25276 11529 25279
rect 10928 25248 11529 25276
rect 10928 25236 10934 25248
rect 11517 25245 11529 25248
rect 11563 25245 11575 25279
rect 11517 25239 11575 25245
rect 11054 25208 11060 25220
rect 10612 25180 11060 25208
rect 11054 25168 11060 25180
rect 11112 25168 11118 25220
rect 11532 25208 11560 25239
rect 11606 25236 11612 25288
rect 11664 25276 11670 25288
rect 11701 25279 11759 25285
rect 11701 25276 11713 25279
rect 11664 25248 11713 25276
rect 11664 25236 11670 25248
rect 11701 25245 11713 25248
rect 11747 25245 11759 25279
rect 12406 25276 12434 25316
rect 13265 25279 13323 25285
rect 13265 25276 13277 25279
rect 12406 25248 13277 25276
rect 11701 25239 11759 25245
rect 13265 25245 13277 25248
rect 13311 25245 13323 25279
rect 13265 25239 13323 25245
rect 13446 25236 13452 25288
rect 13504 25236 13510 25288
rect 14384 25285 14412 25316
rect 15194 25304 15200 25316
rect 15252 25304 15258 25356
rect 16206 25344 16212 25356
rect 15304 25316 16212 25344
rect 14369 25279 14427 25285
rect 14369 25245 14381 25279
rect 14415 25245 14427 25279
rect 14369 25239 14427 25245
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25276 14611 25279
rect 14642 25276 14648 25288
rect 14599 25248 14648 25276
rect 14599 25245 14611 25248
rect 14553 25239 14611 25245
rect 14642 25236 14648 25248
rect 14700 25236 14706 25288
rect 15010 25236 15016 25288
rect 15068 25236 15074 25288
rect 15304 25285 15332 25316
rect 16206 25304 16212 25316
rect 16264 25344 16270 25356
rect 16669 25347 16727 25353
rect 16669 25344 16681 25347
rect 16264 25316 16681 25344
rect 16264 25304 16270 25316
rect 16669 25313 16681 25316
rect 16715 25313 16727 25347
rect 17586 25344 17592 25356
rect 16669 25307 16727 25313
rect 16868 25316 17592 25344
rect 16868 25288 16896 25316
rect 17586 25304 17592 25316
rect 17644 25344 17650 25356
rect 18141 25347 18199 25353
rect 18141 25344 18153 25347
rect 17644 25316 18153 25344
rect 17644 25304 17650 25316
rect 18141 25313 18153 25316
rect 18187 25344 18199 25347
rect 18598 25344 18604 25356
rect 18187 25316 18604 25344
rect 18187 25313 18199 25316
rect 18141 25307 18199 25313
rect 18598 25304 18604 25316
rect 18656 25304 18662 25356
rect 19058 25344 19064 25356
rect 18708 25316 19064 25344
rect 15289 25279 15347 25285
rect 15289 25245 15301 25279
rect 15335 25245 15347 25279
rect 15289 25239 15347 25245
rect 15378 25236 15384 25288
rect 15436 25276 15442 25288
rect 16574 25276 16580 25288
rect 15436 25248 16580 25276
rect 15436 25236 15442 25248
rect 16574 25236 16580 25248
rect 16632 25236 16638 25288
rect 16850 25236 16856 25288
rect 16908 25236 16914 25288
rect 16942 25236 16948 25288
rect 17000 25276 17006 25288
rect 18708 25285 18736 25316
rect 19058 25304 19064 25316
rect 19116 25304 19122 25356
rect 19429 25347 19487 25353
rect 19429 25313 19441 25347
rect 19475 25313 19487 25347
rect 19812 25344 19840 25372
rect 19429 25307 19487 25313
rect 19793 25316 19840 25344
rect 17957 25279 18015 25285
rect 17957 25276 17969 25279
rect 17000 25248 17969 25276
rect 17000 25236 17006 25248
rect 17957 25245 17969 25248
rect 18003 25245 18015 25279
rect 17957 25239 18015 25245
rect 18693 25279 18751 25285
rect 18693 25245 18705 25279
rect 18739 25245 18751 25279
rect 18693 25239 18751 25245
rect 18782 25236 18788 25288
rect 18840 25276 18846 25288
rect 18877 25279 18935 25285
rect 18877 25276 18889 25279
rect 18840 25248 18889 25276
rect 18840 25236 18846 25248
rect 18877 25245 18889 25248
rect 18923 25245 18935 25279
rect 19444 25276 19472 25307
rect 19793 25285 19821 25316
rect 18877 25239 18935 25245
rect 19260 25248 19472 25276
rect 19613 25279 19671 25285
rect 19613 25270 19625 25279
rect 12066 25208 12072 25220
rect 11532 25180 12072 25208
rect 12066 25168 12072 25180
rect 12124 25168 12130 25220
rect 14458 25168 14464 25220
rect 14516 25168 14522 25220
rect 14918 25168 14924 25220
rect 14976 25208 14982 25220
rect 15197 25211 15255 25217
rect 15197 25208 15209 25211
rect 14976 25180 15209 25208
rect 14976 25168 14982 25180
rect 15197 25177 15209 25180
rect 15243 25177 15255 25211
rect 17865 25211 17923 25217
rect 17865 25208 17877 25211
rect 15197 25171 15255 25177
rect 16684 25180 17877 25208
rect 9122 25100 9128 25152
rect 9180 25100 9186 25152
rect 9490 25100 9496 25152
rect 9548 25100 9554 25152
rect 10226 25100 10232 25152
rect 10284 25140 10290 25152
rect 10505 25143 10563 25149
rect 10505 25140 10517 25143
rect 10284 25112 10517 25140
rect 10284 25100 10290 25112
rect 10505 25109 10517 25112
rect 10551 25109 10563 25143
rect 10505 25103 10563 25109
rect 11609 25143 11667 25149
rect 11609 25109 11621 25143
rect 11655 25140 11667 25143
rect 11698 25140 11704 25152
rect 11655 25112 11704 25140
rect 11655 25109 11667 25112
rect 11609 25103 11667 25109
rect 11698 25100 11704 25112
rect 11756 25100 11762 25152
rect 15286 25100 15292 25152
rect 15344 25140 15350 25152
rect 16684 25140 16712 25180
rect 17865 25177 17877 25180
rect 17911 25177 17923 25211
rect 17865 25171 17923 25177
rect 18506 25168 18512 25220
rect 18564 25208 18570 25220
rect 19260 25208 19288 25248
rect 18564 25180 19288 25208
rect 19536 25245 19625 25270
rect 19659 25245 19671 25279
rect 19536 25242 19671 25245
rect 18564 25168 18570 25180
rect 15344 25112 16712 25140
rect 15344 25100 15350 25112
rect 17494 25100 17500 25152
rect 17552 25100 17558 25152
rect 19536 25140 19564 25242
rect 19613 25239 19671 25242
rect 19778 25279 19836 25285
rect 19778 25245 19790 25279
rect 19824 25245 19836 25279
rect 19778 25239 19836 25245
rect 19874 25279 19932 25285
rect 19874 25245 19886 25279
rect 19920 25245 19932 25279
rect 19874 25239 19932 25245
rect 19981 25279 20039 25285
rect 19981 25245 19993 25279
rect 20027 25270 20039 25279
rect 20088 25270 20116 25384
rect 20346 25304 20352 25356
rect 20404 25344 20410 25356
rect 21450 25344 21456 25356
rect 20404 25316 21456 25344
rect 20404 25304 20410 25316
rect 21450 25304 21456 25316
rect 21508 25304 21514 25356
rect 21637 25347 21695 25353
rect 21637 25313 21649 25347
rect 21683 25344 21695 25347
rect 22646 25344 22652 25356
rect 21683 25316 22652 25344
rect 21683 25313 21695 25316
rect 21637 25307 21695 25313
rect 22646 25304 22652 25316
rect 22704 25304 22710 25356
rect 22373 25279 22431 25285
rect 22373 25276 22385 25279
rect 20027 25245 20116 25270
rect 19981 25242 20116 25245
rect 22112 25248 22385 25276
rect 19981 25239 20039 25242
rect 19889 25208 19917 25239
rect 20346 25208 20352 25220
rect 19889 25180 20352 25208
rect 20346 25168 20352 25180
rect 20404 25168 20410 25220
rect 20622 25168 20628 25220
rect 20680 25208 20686 25220
rect 22112 25208 22140 25248
rect 22373 25245 22385 25248
rect 22419 25245 22431 25279
rect 22373 25239 22431 25245
rect 22462 25236 22468 25288
rect 22520 25236 22526 25288
rect 22741 25279 22799 25285
rect 22741 25245 22753 25279
rect 22787 25276 22799 25279
rect 22848 25276 22876 25384
rect 23658 25372 23664 25384
rect 23716 25372 23722 25424
rect 23937 25415 23995 25421
rect 23937 25381 23949 25415
rect 23983 25412 23995 25415
rect 24026 25412 24032 25424
rect 23983 25384 24032 25412
rect 23983 25381 23995 25384
rect 23937 25375 23995 25381
rect 24026 25372 24032 25384
rect 24084 25372 24090 25424
rect 24946 25412 24952 25424
rect 24136 25384 24952 25412
rect 23566 25304 23572 25356
rect 23624 25304 23630 25356
rect 23676 25344 23704 25372
rect 24136 25344 24164 25384
rect 24946 25372 24952 25384
rect 25004 25372 25010 25424
rect 25038 25372 25044 25424
rect 25096 25412 25102 25424
rect 25133 25415 25191 25421
rect 25133 25412 25145 25415
rect 25096 25384 25145 25412
rect 25096 25372 25102 25384
rect 25133 25381 25145 25384
rect 25179 25381 25191 25415
rect 25133 25375 25191 25381
rect 26234 25372 26240 25424
rect 26292 25412 26298 25424
rect 26697 25415 26755 25421
rect 26697 25412 26709 25415
rect 26292 25384 26709 25412
rect 26292 25372 26298 25384
rect 26697 25381 26709 25384
rect 26743 25381 26755 25415
rect 27982 25412 27988 25424
rect 26697 25375 26755 25381
rect 26804 25384 27988 25412
rect 23676 25316 24164 25344
rect 24578 25304 24584 25356
rect 24636 25344 24642 25356
rect 24673 25347 24731 25353
rect 24673 25344 24685 25347
rect 24636 25316 24685 25344
rect 24636 25304 24642 25316
rect 24673 25313 24685 25316
rect 24719 25313 24731 25347
rect 24673 25307 24731 25313
rect 24854 25304 24860 25356
rect 24912 25344 24918 25356
rect 24912 25316 25820 25344
rect 24912 25304 24918 25316
rect 22787 25248 22876 25276
rect 22787 25245 22799 25248
rect 22741 25239 22799 25245
rect 23106 25236 23112 25288
rect 23164 25276 23170 25288
rect 23753 25279 23811 25285
rect 23753 25276 23765 25279
rect 23164 25248 23765 25276
rect 23164 25236 23170 25248
rect 23753 25245 23765 25248
rect 23799 25245 23811 25279
rect 23753 25239 23811 25245
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25276 24823 25279
rect 25314 25276 25320 25288
rect 24811 25248 25320 25276
rect 24811 25245 24823 25248
rect 24765 25239 24823 25245
rect 25314 25236 25320 25248
rect 25372 25236 25378 25288
rect 25792 25285 25820 25316
rect 25866 25304 25872 25356
rect 25924 25344 25930 25356
rect 26804 25344 26832 25384
rect 27982 25372 27988 25384
rect 28040 25372 28046 25424
rect 28092 25344 28120 25452
rect 28460 25412 28488 25452
rect 28902 25440 28908 25492
rect 28960 25480 28966 25492
rect 29546 25480 29552 25492
rect 28960 25452 29552 25480
rect 28960 25440 28966 25452
rect 29546 25440 29552 25452
rect 29604 25440 29610 25492
rect 29841 25452 30052 25480
rect 28721 25415 28779 25421
rect 28721 25412 28733 25415
rect 28460 25384 28733 25412
rect 28721 25381 28733 25384
rect 28767 25381 28779 25415
rect 28721 25375 28779 25381
rect 28902 25344 28908 25356
rect 25924 25316 26832 25344
rect 27448 25316 28120 25344
rect 28184 25316 28908 25344
rect 25924 25304 25930 25316
rect 25777 25279 25835 25285
rect 25777 25245 25789 25279
rect 25823 25245 25835 25279
rect 25777 25239 25835 25245
rect 26510 25236 26516 25288
rect 26568 25236 26574 25288
rect 26602 25236 26608 25288
rect 26660 25236 26666 25288
rect 27448 25285 27476 25316
rect 27433 25279 27491 25285
rect 27433 25245 27445 25279
rect 27479 25245 27491 25279
rect 27433 25239 27491 25245
rect 27614 25236 27620 25288
rect 27672 25236 27678 25288
rect 27709 25279 27767 25285
rect 27709 25245 27721 25279
rect 27755 25276 27767 25279
rect 28074 25276 28080 25288
rect 27755 25248 28080 25276
rect 27755 25245 27767 25248
rect 27709 25239 27767 25245
rect 28074 25236 28080 25248
rect 28132 25236 28138 25288
rect 28184 25285 28212 25316
rect 28902 25304 28908 25316
rect 28960 25304 28966 25356
rect 28169 25279 28227 25285
rect 28169 25245 28181 25279
rect 28215 25245 28227 25279
rect 28445 25279 28503 25285
rect 28445 25276 28457 25279
rect 28169 25239 28227 25245
rect 28276 25248 28457 25276
rect 20680 25180 22140 25208
rect 22189 25211 22247 25217
rect 20680 25168 20686 25180
rect 22189 25177 22201 25211
rect 22235 25208 22247 25211
rect 22554 25208 22560 25220
rect 22235 25180 22560 25208
rect 22235 25177 22247 25180
rect 22189 25171 22247 25177
rect 22554 25168 22560 25180
rect 22612 25168 22618 25220
rect 23477 25211 23535 25217
rect 23477 25177 23489 25211
rect 23523 25177 23535 25211
rect 23477 25171 23535 25177
rect 20070 25140 20076 25152
rect 19536 25112 20076 25140
rect 20070 25100 20076 25112
rect 20128 25100 20134 25152
rect 20990 25100 20996 25152
rect 21048 25100 21054 25152
rect 21358 25100 21364 25152
rect 21416 25100 21422 25152
rect 21450 25100 21456 25152
rect 21508 25140 21514 25152
rect 23492 25140 23520 25171
rect 24854 25168 24860 25220
rect 24912 25208 24918 25220
rect 25593 25211 25651 25217
rect 25593 25208 25605 25211
rect 24912 25180 25605 25208
rect 24912 25168 24918 25180
rect 25593 25177 25605 25180
rect 25639 25177 25651 25211
rect 27632 25208 27660 25236
rect 25593 25171 25651 25177
rect 25700 25180 27660 25208
rect 25038 25140 25044 25152
rect 21508 25112 25044 25140
rect 21508 25100 21514 25112
rect 25038 25100 25044 25112
rect 25096 25100 25102 25152
rect 25130 25100 25136 25152
rect 25188 25140 25194 25152
rect 25700 25140 25728 25180
rect 27982 25168 27988 25220
rect 28040 25208 28046 25220
rect 28276 25208 28304 25248
rect 28445 25245 28457 25248
rect 28491 25245 28503 25279
rect 28445 25239 28503 25245
rect 28537 25279 28595 25285
rect 28537 25245 28549 25279
rect 28583 25245 28595 25279
rect 28537 25239 28595 25245
rect 29733 25279 29791 25285
rect 29733 25245 29745 25279
rect 29779 25276 29791 25279
rect 29841 25276 29869 25452
rect 30024 25412 30052 25452
rect 30282 25440 30288 25492
rect 30340 25440 30346 25492
rect 30466 25440 30472 25492
rect 30524 25480 30530 25492
rect 31386 25480 31392 25492
rect 30524 25452 31392 25480
rect 30524 25440 30530 25452
rect 31386 25440 31392 25452
rect 31444 25440 31450 25492
rect 33502 25440 33508 25492
rect 33560 25480 33566 25492
rect 33781 25483 33839 25489
rect 33781 25480 33793 25483
rect 33560 25452 33793 25480
rect 33560 25440 33566 25452
rect 33781 25449 33793 25452
rect 33827 25449 33839 25483
rect 33781 25443 33839 25449
rect 36078 25440 36084 25492
rect 36136 25480 36142 25492
rect 36630 25480 36636 25492
rect 36136 25452 36636 25480
rect 36136 25440 36142 25452
rect 36630 25440 36636 25452
rect 36688 25440 36694 25492
rect 36722 25440 36728 25492
rect 36780 25480 36786 25492
rect 39298 25480 39304 25492
rect 36780 25452 39304 25480
rect 36780 25440 36786 25452
rect 39298 25440 39304 25452
rect 39356 25440 39362 25492
rect 30926 25412 30932 25424
rect 30024 25384 30932 25412
rect 30926 25372 30932 25384
rect 30984 25372 30990 25424
rect 33410 25372 33416 25424
rect 33468 25412 33474 25424
rect 33670 25415 33728 25421
rect 33670 25412 33682 25415
rect 33468 25384 33682 25412
rect 33468 25372 33474 25384
rect 33670 25381 33682 25384
rect 33716 25381 33728 25415
rect 33670 25375 33728 25381
rect 29914 25304 29920 25356
rect 29972 25344 29978 25356
rect 30837 25347 30895 25353
rect 29972 25316 30052 25344
rect 29972 25304 29978 25316
rect 30024 25285 30052 25316
rect 30837 25313 30849 25347
rect 30883 25344 30895 25347
rect 31386 25344 31392 25356
rect 30883 25316 31392 25344
rect 30883 25313 30895 25316
rect 30837 25307 30895 25313
rect 31386 25304 31392 25316
rect 31444 25344 31450 25356
rect 32950 25344 32956 25356
rect 31444 25316 32956 25344
rect 31444 25304 31450 25316
rect 32950 25304 32956 25316
rect 33008 25304 33014 25356
rect 33685 25344 33713 25375
rect 35526 25372 35532 25424
rect 35584 25412 35590 25424
rect 35584 25384 36400 25412
rect 35584 25372 35590 25384
rect 33778 25344 33784 25356
rect 33685 25316 33784 25344
rect 33778 25304 33784 25316
rect 33836 25304 33842 25356
rect 33873 25347 33931 25353
rect 33873 25313 33885 25347
rect 33919 25344 33931 25347
rect 34422 25344 34428 25356
rect 33919 25316 34428 25344
rect 33919 25313 33931 25316
rect 33873 25307 33931 25313
rect 29779 25248 29869 25276
rect 30009 25279 30067 25285
rect 29779 25245 29791 25248
rect 29733 25239 29791 25245
rect 30009 25245 30021 25279
rect 30055 25245 30067 25279
rect 30009 25239 30067 25245
rect 30101 25279 30159 25285
rect 30101 25245 30113 25279
rect 30147 25276 30159 25279
rect 30190 25276 30196 25288
rect 30147 25248 30196 25276
rect 30147 25245 30159 25248
rect 30101 25239 30159 25245
rect 28040 25180 28304 25208
rect 28040 25168 28046 25180
rect 28350 25168 28356 25220
rect 28408 25168 28414 25220
rect 25188 25112 25728 25140
rect 25188 25100 25194 25112
rect 27246 25100 27252 25152
rect 27304 25100 27310 25152
rect 27890 25100 27896 25152
rect 27948 25140 27954 25152
rect 28552 25140 28580 25239
rect 30190 25236 30196 25248
rect 30248 25236 30254 25288
rect 30282 25236 30288 25288
rect 30340 25276 30346 25288
rect 31021 25279 31079 25285
rect 31021 25276 31033 25279
rect 30340 25248 31033 25276
rect 30340 25236 30346 25248
rect 31021 25245 31033 25248
rect 31067 25276 31079 25279
rect 31478 25276 31484 25288
rect 31067 25248 31484 25276
rect 31067 25245 31079 25248
rect 31021 25239 31079 25245
rect 31478 25236 31484 25248
rect 31536 25236 31542 25288
rect 32214 25236 32220 25288
rect 32272 25236 32278 25288
rect 32398 25276 32404 25288
rect 32324 25248 32404 25276
rect 29178 25208 29184 25220
rect 28828 25180 29184 25208
rect 28828 25140 28856 25180
rect 29178 25168 29184 25180
rect 29236 25208 29242 25220
rect 29236 25180 29500 25208
rect 29236 25168 29242 25180
rect 27948 25112 28856 25140
rect 27948 25100 27954 25112
rect 28902 25100 28908 25152
rect 28960 25140 28966 25152
rect 28994 25140 29000 25152
rect 28960 25112 29000 25140
rect 28960 25100 28966 25112
rect 28994 25100 29000 25112
rect 29052 25100 29058 25152
rect 29472 25140 29500 25180
rect 29546 25168 29552 25220
rect 29604 25208 29610 25220
rect 29917 25211 29975 25217
rect 29917 25208 29929 25211
rect 29604 25180 29929 25208
rect 29604 25168 29610 25180
rect 29917 25177 29929 25180
rect 29963 25208 29975 25211
rect 30466 25208 30472 25220
rect 29963 25180 30472 25208
rect 29963 25177 29975 25180
rect 29917 25171 29975 25177
rect 30466 25168 30472 25180
rect 30524 25168 30530 25220
rect 30558 25168 30564 25220
rect 30616 25208 30622 25220
rect 31205 25211 31263 25217
rect 31205 25208 31217 25211
rect 30616 25180 31217 25208
rect 30616 25168 30622 25180
rect 31205 25177 31217 25180
rect 31251 25177 31263 25211
rect 31205 25171 31263 25177
rect 31297 25211 31355 25217
rect 31297 25177 31309 25211
rect 31343 25208 31355 25211
rect 31570 25208 31576 25220
rect 31343 25180 31576 25208
rect 31343 25177 31355 25180
rect 31297 25171 31355 25177
rect 31570 25168 31576 25180
rect 31628 25208 31634 25220
rect 32232 25208 32260 25236
rect 31628 25180 32260 25208
rect 31628 25168 31634 25180
rect 30190 25140 30196 25152
rect 29472 25112 30196 25140
rect 30190 25100 30196 25112
rect 30248 25100 30254 25152
rect 31110 25100 31116 25152
rect 31168 25140 31174 25152
rect 32324 25140 32352 25248
rect 32398 25236 32404 25248
rect 32456 25236 32462 25288
rect 32769 25279 32827 25285
rect 32769 25245 32781 25279
rect 32815 25276 32827 25279
rect 32858 25276 32864 25288
rect 32815 25248 32864 25276
rect 32815 25245 32827 25248
rect 32769 25239 32827 25245
rect 32858 25236 32864 25248
rect 32916 25236 32922 25288
rect 33226 25236 33232 25288
rect 33284 25276 33290 25288
rect 33888 25276 33916 25307
rect 34422 25304 34428 25316
rect 34480 25304 34486 25356
rect 35618 25344 35624 25356
rect 34900 25316 35624 25344
rect 34900 25285 34928 25316
rect 35618 25304 35624 25316
rect 35676 25304 35682 25356
rect 33284 25248 33916 25276
rect 34885 25279 34943 25285
rect 33284 25236 33290 25248
rect 34885 25245 34897 25279
rect 34931 25245 34943 25279
rect 34885 25239 34943 25245
rect 35250 25236 35256 25288
rect 35308 25236 35314 25288
rect 36078 25236 36084 25288
rect 36136 25236 36142 25288
rect 36170 25236 36176 25288
rect 36228 25236 36234 25288
rect 36372 25285 36400 25384
rect 36906 25304 36912 25356
rect 36964 25304 36970 25356
rect 36357 25279 36415 25285
rect 36357 25245 36369 25279
rect 36403 25245 36415 25279
rect 36357 25239 36415 25245
rect 36449 25279 36507 25285
rect 36449 25245 36461 25279
rect 36495 25276 36507 25279
rect 37642 25276 37648 25288
rect 36495 25248 37648 25276
rect 36495 25245 36507 25248
rect 36449 25239 36507 25245
rect 37642 25236 37648 25248
rect 37700 25236 37706 25288
rect 33505 25211 33563 25217
rect 33505 25177 33517 25211
rect 33551 25208 33563 25211
rect 33594 25208 33600 25220
rect 33551 25180 33600 25208
rect 33551 25177 33563 25180
rect 33505 25171 33563 25177
rect 33594 25168 33600 25180
rect 33652 25168 33658 25220
rect 34241 25211 34299 25217
rect 34241 25177 34253 25211
rect 34287 25208 34299 25211
rect 34974 25208 34980 25220
rect 34287 25180 34980 25208
rect 34287 25177 34299 25180
rect 34241 25171 34299 25177
rect 34974 25168 34980 25180
rect 35032 25168 35038 25220
rect 35069 25211 35127 25217
rect 35069 25177 35081 25211
rect 35115 25177 35127 25211
rect 35069 25171 35127 25177
rect 35161 25211 35219 25217
rect 35161 25177 35173 25211
rect 35207 25208 35219 25211
rect 35802 25208 35808 25220
rect 35207 25180 35808 25208
rect 35207 25177 35219 25180
rect 35161 25171 35219 25177
rect 31168 25112 32352 25140
rect 33045 25143 33103 25149
rect 31168 25100 31174 25112
rect 33045 25109 33057 25143
rect 33091 25140 33103 25143
rect 33134 25140 33140 25152
rect 33091 25112 33140 25140
rect 33091 25109 33103 25112
rect 33045 25103 33103 25109
rect 33134 25100 33140 25112
rect 33192 25100 33198 25152
rect 33870 25100 33876 25152
rect 33928 25140 33934 25152
rect 34790 25140 34796 25152
rect 33928 25112 34796 25140
rect 33928 25100 33934 25112
rect 34790 25100 34796 25112
rect 34848 25140 34854 25152
rect 35084 25140 35112 25171
rect 35802 25168 35808 25180
rect 35860 25168 35866 25220
rect 35897 25211 35955 25217
rect 35897 25177 35909 25211
rect 35943 25208 35955 25211
rect 36998 25208 37004 25220
rect 35943 25180 37004 25208
rect 35943 25177 35955 25180
rect 35897 25171 35955 25177
rect 36998 25168 37004 25180
rect 37056 25168 37062 25220
rect 37182 25217 37188 25220
rect 37176 25171 37188 25217
rect 37182 25168 37188 25171
rect 37240 25168 37246 25220
rect 35342 25140 35348 25152
rect 34848 25112 35348 25140
rect 34848 25100 34854 25112
rect 35342 25100 35348 25112
rect 35400 25100 35406 25152
rect 35434 25100 35440 25152
rect 35492 25100 35498 25152
rect 35820 25140 35848 25168
rect 36814 25140 36820 25152
rect 35820 25112 36820 25140
rect 36814 25100 36820 25112
rect 36872 25100 36878 25152
rect 37826 25100 37832 25152
rect 37884 25140 37890 25152
rect 38289 25143 38347 25149
rect 38289 25140 38301 25143
rect 37884 25112 38301 25140
rect 37884 25100 37890 25112
rect 38289 25109 38301 25112
rect 38335 25109 38347 25143
rect 38289 25103 38347 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 9490 24896 9496 24948
rect 9548 24936 9554 24948
rect 9585 24939 9643 24945
rect 9585 24936 9597 24939
rect 9548 24908 9597 24936
rect 9548 24896 9554 24908
rect 9585 24905 9597 24908
rect 9631 24905 9643 24939
rect 9585 24899 9643 24905
rect 14277 24939 14335 24945
rect 14277 24905 14289 24939
rect 14323 24936 14335 24939
rect 15102 24936 15108 24948
rect 14323 24908 15108 24936
rect 14323 24905 14335 24908
rect 14277 24899 14335 24905
rect 8472 24871 8530 24877
rect 8472 24837 8484 24871
rect 8518 24868 8530 24871
rect 9122 24868 9128 24880
rect 8518 24840 9128 24868
rect 8518 24837 8530 24840
rect 8472 24831 8530 24837
rect 9122 24828 9128 24840
rect 9180 24828 9186 24880
rect 9600 24868 9628 24899
rect 15102 24896 15108 24908
rect 15160 24896 15166 24948
rect 16298 24896 16304 24948
rect 16356 24936 16362 24948
rect 16945 24939 17003 24945
rect 16945 24936 16957 24939
rect 16356 24908 16957 24936
rect 16356 24896 16362 24908
rect 16945 24905 16957 24908
rect 16991 24936 17003 24939
rect 17310 24936 17316 24948
rect 16991 24908 17316 24936
rect 16991 24905 17003 24908
rect 16945 24899 17003 24905
rect 17310 24896 17316 24908
rect 17368 24896 17374 24948
rect 17494 24896 17500 24948
rect 17552 24936 17558 24948
rect 17773 24939 17831 24945
rect 17773 24936 17785 24939
rect 17552 24908 17785 24936
rect 17552 24896 17558 24908
rect 17773 24905 17785 24908
rect 17819 24905 17831 24939
rect 19518 24936 19524 24948
rect 17773 24899 17831 24905
rect 17880 24908 19524 24936
rect 17880 24868 17908 24908
rect 19518 24896 19524 24908
rect 19576 24896 19582 24948
rect 19720 24908 20024 24936
rect 9600 24840 17908 24868
rect 18693 24871 18751 24877
rect 18693 24837 18705 24871
rect 18739 24868 18751 24871
rect 18782 24868 18788 24880
rect 18739 24840 18788 24868
rect 18739 24837 18751 24840
rect 18693 24831 18751 24837
rect 18782 24828 18788 24840
rect 18840 24828 18846 24880
rect 19720 24868 19748 24908
rect 18984 24840 19748 24868
rect 5350 24760 5356 24812
rect 5408 24800 5414 24812
rect 10134 24800 10140 24812
rect 5408 24772 10140 24800
rect 5408 24760 5414 24772
rect 10134 24760 10140 24772
rect 10192 24760 10198 24812
rect 10226 24760 10232 24812
rect 10284 24760 10290 24812
rect 10318 24760 10324 24812
rect 10376 24760 10382 24812
rect 10597 24803 10655 24809
rect 10597 24769 10609 24803
rect 10643 24800 10655 24803
rect 10870 24800 10876 24812
rect 10643 24772 10876 24800
rect 10643 24769 10655 24772
rect 10597 24763 10655 24769
rect 10870 24760 10876 24772
rect 10928 24760 10934 24812
rect 11698 24760 11704 24812
rect 11756 24760 11762 24812
rect 11882 24760 11888 24812
rect 11940 24760 11946 24812
rect 11974 24760 11980 24812
rect 12032 24760 12038 24812
rect 12066 24760 12072 24812
rect 12124 24760 12130 24812
rect 13164 24803 13222 24809
rect 13164 24769 13176 24803
rect 13210 24800 13222 24803
rect 16117 24803 16175 24809
rect 16117 24800 16129 24803
rect 13210 24772 13952 24800
rect 13210 24769 13222 24772
rect 13164 24763 13222 24769
rect 8202 24692 8208 24744
rect 8260 24692 8266 24744
rect 10689 24735 10747 24741
rect 10689 24701 10701 24735
rect 10735 24701 10747 24735
rect 10689 24695 10747 24701
rect 10704 24664 10732 24695
rect 11422 24692 11428 24744
rect 11480 24732 11486 24744
rect 12894 24732 12900 24744
rect 11480 24704 12900 24732
rect 11480 24692 11486 24704
rect 12894 24692 12900 24704
rect 12952 24692 12958 24744
rect 10870 24664 10876 24676
rect 10704 24636 10876 24664
rect 10870 24624 10876 24636
rect 10928 24664 10934 24676
rect 13924 24664 13952 24772
rect 15672 24772 16129 24800
rect 14366 24692 14372 24744
rect 14424 24732 14430 24744
rect 15197 24735 15255 24741
rect 15197 24732 15209 24735
rect 14424 24704 15209 24732
rect 14424 24692 14430 24704
rect 15197 24701 15209 24704
rect 15243 24701 15255 24735
rect 15197 24695 15255 24701
rect 15289 24735 15347 24741
rect 15289 24701 15301 24735
rect 15335 24701 15347 24735
rect 15289 24695 15347 24701
rect 14737 24667 14795 24673
rect 14737 24664 14749 24667
rect 10928 24636 12434 24664
rect 13924 24636 14749 24664
rect 10928 24624 10934 24636
rect 10042 24556 10048 24608
rect 10100 24556 10106 24608
rect 12250 24556 12256 24608
rect 12308 24556 12314 24608
rect 12406 24596 12434 24636
rect 14737 24633 14749 24636
rect 14783 24633 14795 24667
rect 14737 24627 14795 24633
rect 15010 24624 15016 24676
rect 15068 24664 15074 24676
rect 15304 24664 15332 24695
rect 15068 24636 15332 24664
rect 15068 24624 15074 24636
rect 15672 24596 15700 24772
rect 16117 24769 16129 24772
rect 16163 24800 16175 24803
rect 16206 24800 16212 24812
rect 16163 24772 16212 24800
rect 16163 24769 16175 24772
rect 16117 24763 16175 24769
rect 16206 24760 16212 24772
rect 16264 24760 16270 24812
rect 16301 24803 16359 24809
rect 16301 24769 16313 24803
rect 16347 24800 16359 24803
rect 16850 24800 16856 24812
rect 16347 24772 16856 24800
rect 16347 24769 16359 24772
rect 16301 24763 16359 24769
rect 16850 24760 16856 24772
rect 16908 24760 16914 24812
rect 17310 24760 17316 24812
rect 17368 24800 17374 24812
rect 17678 24800 17684 24812
rect 17368 24772 17684 24800
rect 17368 24760 17374 24772
rect 17678 24760 17684 24772
rect 17736 24760 17742 24812
rect 18984 24809 19012 24840
rect 19794 24828 19800 24880
rect 19852 24828 19858 24880
rect 18969 24803 19027 24809
rect 18969 24769 18981 24803
rect 19015 24769 19027 24803
rect 18969 24763 19027 24769
rect 19058 24760 19064 24812
rect 19116 24760 19122 24812
rect 19429 24803 19487 24809
rect 19429 24769 19441 24803
rect 19475 24800 19487 24803
rect 19610 24800 19616 24812
rect 19475 24772 19616 24800
rect 19475 24769 19487 24772
rect 19429 24763 19487 24769
rect 19610 24760 19616 24772
rect 19668 24760 19674 24812
rect 19996 24800 20024 24908
rect 20990 24896 20996 24948
rect 21048 24896 21054 24948
rect 22646 24896 22652 24948
rect 22704 24936 22710 24948
rect 26142 24936 26148 24948
rect 22704 24908 26148 24936
rect 22704 24896 22710 24908
rect 26142 24896 26148 24908
rect 26200 24896 26206 24948
rect 27614 24896 27620 24948
rect 27672 24936 27678 24948
rect 28350 24936 28356 24948
rect 27672 24908 28356 24936
rect 27672 24896 27678 24908
rect 28350 24896 28356 24908
rect 28408 24896 28414 24948
rect 29178 24936 29184 24948
rect 28966 24908 29184 24936
rect 21358 24828 21364 24880
rect 21416 24868 21422 24880
rect 24204 24871 24262 24877
rect 24204 24868 24216 24871
rect 21416 24840 24216 24868
rect 21416 24828 21422 24840
rect 24204 24837 24216 24840
rect 24250 24868 24262 24871
rect 24250 24840 25728 24868
rect 24250 24837 24262 24840
rect 24204 24831 24262 24837
rect 20254 24800 20260 24812
rect 19996 24772 20260 24800
rect 20254 24760 20260 24772
rect 20312 24760 20318 24812
rect 20898 24800 20904 24812
rect 20364 24772 20904 24800
rect 17957 24735 18015 24741
rect 17957 24701 17969 24735
rect 18003 24732 18015 24735
rect 18322 24732 18328 24744
rect 18003 24704 18328 24732
rect 18003 24701 18015 24704
rect 17957 24695 18015 24701
rect 18322 24692 18328 24704
rect 18380 24692 18386 24744
rect 15838 24624 15844 24676
rect 15896 24664 15902 24676
rect 18524 24664 18552 24718
rect 19794 24692 19800 24744
rect 19852 24732 19858 24744
rect 20364 24732 20392 24772
rect 20898 24760 20904 24772
rect 20956 24760 20962 24812
rect 21818 24760 21824 24812
rect 21876 24800 21882 24812
rect 22261 24803 22319 24809
rect 22261 24800 22273 24803
rect 21876 24772 22273 24800
rect 21876 24760 21882 24772
rect 22261 24769 22273 24772
rect 22307 24769 22319 24803
rect 22261 24763 22319 24769
rect 23934 24760 23940 24812
rect 23992 24760 23998 24812
rect 24670 24760 24676 24812
rect 24728 24800 24734 24812
rect 25700 24800 25728 24840
rect 25774 24828 25780 24880
rect 25832 24868 25838 24880
rect 25832 24840 27016 24868
rect 25832 24828 25838 24840
rect 25958 24800 25964 24812
rect 24728 24772 25636 24800
rect 25700 24772 25964 24800
rect 24728 24760 24734 24772
rect 19852 24704 20392 24732
rect 19852 24692 19858 24704
rect 20530 24692 20536 24744
rect 20588 24732 20594 24744
rect 21085 24735 21143 24741
rect 21085 24732 21097 24735
rect 20588 24704 21097 24732
rect 20588 24692 20594 24704
rect 21085 24701 21097 24704
rect 21131 24701 21143 24735
rect 21085 24695 21143 24701
rect 22002 24692 22008 24744
rect 22060 24692 22066 24744
rect 25608 24732 25636 24772
rect 25958 24760 25964 24772
rect 26016 24760 26022 24812
rect 26050 24760 26056 24812
rect 26108 24800 26114 24812
rect 26145 24803 26203 24809
rect 26145 24800 26157 24803
rect 26108 24772 26157 24800
rect 26108 24760 26114 24772
rect 26145 24769 26157 24772
rect 26191 24769 26203 24803
rect 26145 24763 26203 24769
rect 26234 24760 26240 24812
rect 26292 24760 26298 24812
rect 26334 24803 26392 24809
rect 26334 24769 26346 24803
rect 26380 24769 26392 24803
rect 26988 24800 27016 24840
rect 27338 24828 27344 24880
rect 27396 24868 27402 24880
rect 28966 24868 28994 24908
rect 29178 24896 29184 24908
rect 29236 24896 29242 24948
rect 30561 24939 30619 24945
rect 30561 24905 30573 24939
rect 30607 24936 30619 24939
rect 31202 24936 31208 24948
rect 30607 24908 31208 24936
rect 30607 24905 30619 24908
rect 30561 24899 30619 24905
rect 31202 24896 31208 24908
rect 31260 24896 31266 24948
rect 31478 24896 31484 24948
rect 31536 24936 31542 24948
rect 31536 24908 34652 24936
rect 31536 24896 31542 24908
rect 27396 24840 28994 24868
rect 27396 24828 27402 24840
rect 29086 24828 29092 24880
rect 29144 24868 29150 24880
rect 29144 24840 29316 24868
rect 29144 24828 29150 24840
rect 29288 24834 29316 24840
rect 27433 24803 27491 24809
rect 27433 24800 27445 24803
rect 26988 24772 27445 24800
rect 26334 24763 26392 24769
rect 27433 24769 27445 24772
rect 27479 24769 27491 24803
rect 27433 24763 27491 24769
rect 26349 24732 26377 24763
rect 27614 24760 27620 24812
rect 27672 24760 27678 24812
rect 27709 24803 27767 24809
rect 27709 24769 27721 24803
rect 27755 24769 27767 24803
rect 27709 24763 27767 24769
rect 27801 24803 27859 24809
rect 27801 24769 27813 24803
rect 27847 24800 27859 24803
rect 27890 24800 27896 24812
rect 27847 24772 27896 24800
rect 27847 24769 27859 24772
rect 27801 24763 27859 24769
rect 26878 24732 26884 24744
rect 25608 24704 26884 24732
rect 26878 24692 26884 24704
rect 26936 24692 26942 24744
rect 27724 24732 27752 24763
rect 27890 24760 27896 24772
rect 27948 24760 27954 24812
rect 28261 24803 28319 24809
rect 28261 24769 28273 24803
rect 28307 24800 28319 24803
rect 29178 24800 29184 24812
rect 28307 24772 29184 24800
rect 28307 24769 28319 24772
rect 28261 24763 28319 24769
rect 29178 24760 29184 24772
rect 29236 24760 29242 24812
rect 29288 24809 29408 24834
rect 29454 24828 29460 24880
rect 29512 24868 29518 24880
rect 30282 24868 30288 24880
rect 29512 24840 30288 24868
rect 29512 24828 29518 24840
rect 30282 24828 30288 24840
rect 30340 24828 30346 24880
rect 30466 24828 30472 24880
rect 30524 24868 30530 24880
rect 31294 24868 31300 24880
rect 30524 24840 31300 24868
rect 30524 24828 30530 24840
rect 31294 24828 31300 24840
rect 31352 24828 31358 24880
rect 32858 24828 32864 24880
rect 32916 24828 32922 24880
rect 33134 24828 33140 24880
rect 33192 24828 33198 24880
rect 33502 24828 33508 24880
rect 33560 24868 33566 24880
rect 34057 24871 34115 24877
rect 34057 24868 34069 24871
rect 33560 24840 34069 24868
rect 33560 24828 33566 24840
rect 34057 24837 34069 24840
rect 34103 24837 34115 24871
rect 34057 24831 34115 24837
rect 29288 24806 29423 24809
rect 29365 24803 29423 24806
rect 29365 24769 29377 24803
rect 29411 24769 29423 24803
rect 29365 24763 29423 24769
rect 29546 24760 29552 24812
rect 29604 24760 29610 24812
rect 29638 24760 29644 24812
rect 29696 24760 29702 24812
rect 29733 24803 29791 24809
rect 29733 24769 29745 24803
rect 29779 24800 29791 24803
rect 30190 24800 30196 24812
rect 29779 24772 30196 24800
rect 29779 24769 29791 24772
rect 29733 24763 29791 24769
rect 30190 24760 30196 24772
rect 30248 24760 30254 24812
rect 30374 24760 30380 24812
rect 30432 24760 30438 24812
rect 30650 24760 30656 24812
rect 30708 24760 30714 24812
rect 31386 24760 31392 24812
rect 31444 24760 31450 24812
rect 31481 24803 31539 24809
rect 31481 24769 31493 24803
rect 31527 24769 31539 24803
rect 31481 24763 31539 24769
rect 31665 24803 31723 24809
rect 31665 24769 31677 24803
rect 31711 24769 31723 24803
rect 31665 24763 31723 24769
rect 31757 24803 31815 24809
rect 31757 24769 31769 24803
rect 31803 24800 31815 24803
rect 32585 24803 32643 24809
rect 31803 24772 32352 24800
rect 31803 24769 31815 24772
rect 31757 24763 31815 24769
rect 27982 24732 27988 24744
rect 27724 24704 27988 24732
rect 27982 24692 27988 24704
rect 28040 24692 28046 24744
rect 28534 24692 28540 24744
rect 28592 24732 28598 24744
rect 31110 24732 31116 24744
rect 28592 24704 31116 24732
rect 28592 24692 28598 24704
rect 31110 24692 31116 24704
rect 31168 24692 31174 24744
rect 15896 24636 18552 24664
rect 19981 24667 20039 24673
rect 15896 24624 15902 24636
rect 19981 24633 19993 24667
rect 20027 24664 20039 24667
rect 20162 24664 20168 24676
rect 20027 24636 20168 24664
rect 20027 24633 20039 24636
rect 19981 24627 20039 24633
rect 20162 24624 20168 24636
rect 20220 24624 20226 24676
rect 25498 24624 25504 24676
rect 25556 24664 25562 24676
rect 31496 24664 31524 24763
rect 25556 24636 31524 24664
rect 25556 24624 25562 24636
rect 12406 24568 15700 24596
rect 16117 24599 16175 24605
rect 16117 24565 16129 24599
rect 16163 24596 16175 24599
rect 16758 24596 16764 24608
rect 16163 24568 16764 24596
rect 16163 24565 16175 24568
rect 16117 24559 16175 24565
rect 16758 24556 16764 24568
rect 16816 24556 16822 24608
rect 17310 24556 17316 24608
rect 17368 24556 17374 24608
rect 20530 24556 20536 24608
rect 20588 24556 20594 24608
rect 20714 24556 20720 24608
rect 20772 24596 20778 24608
rect 22646 24596 22652 24608
rect 20772 24568 22652 24596
rect 20772 24556 20778 24568
rect 22646 24556 22652 24568
rect 22704 24556 22710 24608
rect 23385 24599 23443 24605
rect 23385 24565 23397 24599
rect 23431 24596 23443 24599
rect 23842 24596 23848 24608
rect 23431 24568 23848 24596
rect 23431 24565 23443 24568
rect 23385 24559 23443 24565
rect 23842 24556 23848 24568
rect 23900 24556 23906 24608
rect 25314 24556 25320 24608
rect 25372 24596 25378 24608
rect 25958 24596 25964 24608
rect 25372 24568 25964 24596
rect 25372 24556 25378 24568
rect 25958 24556 25964 24568
rect 26016 24556 26022 24608
rect 26418 24556 26424 24608
rect 26476 24596 26482 24608
rect 26513 24599 26571 24605
rect 26513 24596 26525 24599
rect 26476 24568 26525 24596
rect 26476 24556 26482 24568
rect 26513 24565 26525 24568
rect 26559 24565 26571 24599
rect 26513 24559 26571 24565
rect 27890 24556 27896 24608
rect 27948 24596 27954 24608
rect 27985 24599 28043 24605
rect 27985 24596 27997 24599
rect 27948 24568 27997 24596
rect 27948 24556 27954 24568
rect 27985 24565 27997 24568
rect 28031 24565 28043 24599
rect 27985 24559 28043 24565
rect 28994 24556 29000 24608
rect 29052 24596 29058 24608
rect 29089 24599 29147 24605
rect 29089 24596 29101 24599
rect 29052 24568 29101 24596
rect 29052 24556 29058 24568
rect 29089 24565 29101 24568
rect 29135 24596 29147 24599
rect 29638 24596 29644 24608
rect 29135 24568 29644 24596
rect 29135 24565 29147 24568
rect 29089 24559 29147 24565
rect 29638 24556 29644 24568
rect 29696 24556 29702 24608
rect 29917 24599 29975 24605
rect 29917 24565 29929 24599
rect 29963 24596 29975 24599
rect 30282 24596 30288 24608
rect 29963 24568 30288 24596
rect 29963 24565 29975 24568
rect 29917 24559 29975 24565
rect 30282 24556 30288 24568
rect 30340 24556 30346 24608
rect 30374 24556 30380 24608
rect 30432 24556 30438 24608
rect 30466 24556 30472 24608
rect 30524 24596 30530 24608
rect 30834 24596 30840 24608
rect 30524 24568 30840 24596
rect 30524 24556 30530 24568
rect 30834 24556 30840 24568
rect 30892 24556 30898 24608
rect 31202 24556 31208 24608
rect 31260 24556 31266 24608
rect 31680 24596 31708 24763
rect 31754 24624 31760 24676
rect 31812 24664 31818 24676
rect 32214 24664 32220 24676
rect 31812 24636 32220 24664
rect 31812 24624 31818 24636
rect 32214 24624 32220 24636
rect 32272 24624 32278 24676
rect 32324 24673 32352 24772
rect 32585 24769 32597 24803
rect 32631 24769 32643 24803
rect 33152 24800 33180 24828
rect 34624 24812 34652 24908
rect 34974 24896 34980 24948
rect 35032 24936 35038 24948
rect 35618 24936 35624 24948
rect 35032 24908 35624 24936
rect 35032 24896 35038 24908
rect 35618 24896 35624 24908
rect 35676 24896 35682 24948
rect 35986 24896 35992 24948
rect 36044 24936 36050 24948
rect 37550 24936 37556 24948
rect 36044 24908 37556 24936
rect 36044 24896 36050 24908
rect 37550 24896 37556 24908
rect 37608 24896 37614 24948
rect 37826 24896 37832 24948
rect 37884 24896 37890 24948
rect 36081 24871 36139 24877
rect 36081 24868 36093 24871
rect 34772 24840 36093 24868
rect 33689 24803 33747 24809
rect 33689 24800 33701 24803
rect 33152 24772 33701 24800
rect 32585 24763 32643 24769
rect 33689 24769 33701 24772
rect 33735 24800 33747 24803
rect 33870 24800 33876 24812
rect 33735 24772 33876 24800
rect 33735 24769 33747 24772
rect 33689 24763 33747 24769
rect 32398 24692 32404 24744
rect 32456 24732 32462 24744
rect 32493 24735 32551 24741
rect 32493 24732 32505 24735
rect 32456 24704 32505 24732
rect 32456 24692 32462 24704
rect 32493 24701 32505 24704
rect 32539 24701 32551 24735
rect 32493 24695 32551 24701
rect 32309 24667 32367 24673
rect 32309 24633 32321 24667
rect 32355 24633 32367 24667
rect 32600 24664 32628 24763
rect 33870 24760 33876 24772
rect 33928 24760 33934 24812
rect 34606 24760 34612 24812
rect 34664 24760 34670 24812
rect 34772 24809 34800 24840
rect 36081 24837 36093 24840
rect 36127 24868 36139 24871
rect 37844 24868 37872 24896
rect 36127 24840 37872 24868
rect 36127 24837 36139 24840
rect 36081 24831 36139 24837
rect 34757 24803 34815 24809
rect 34757 24769 34769 24803
rect 34803 24769 34815 24803
rect 34757 24763 34815 24769
rect 34882 24760 34888 24812
rect 34940 24760 34946 24812
rect 34985 24803 35043 24809
rect 34985 24769 34997 24803
rect 35031 24769 35043 24803
rect 34985 24763 35043 24769
rect 35115 24803 35173 24809
rect 35115 24769 35127 24803
rect 35161 24800 35173 24803
rect 35342 24800 35348 24812
rect 35161 24772 35348 24800
rect 35161 24769 35173 24772
rect 35115 24763 35173 24769
rect 32950 24692 32956 24744
rect 33008 24692 33014 24744
rect 33134 24692 33140 24744
rect 33192 24732 33198 24744
rect 33597 24735 33655 24741
rect 33597 24732 33609 24735
rect 33192 24704 33609 24732
rect 33192 24692 33198 24704
rect 33597 24701 33609 24704
rect 33643 24701 33655 24735
rect 33597 24695 33655 24701
rect 33965 24735 34023 24741
rect 33965 24701 33977 24735
rect 34011 24732 34023 24735
rect 34054 24732 34060 24744
rect 34011 24704 34060 24732
rect 34011 24701 34023 24704
rect 33965 24695 34023 24701
rect 34054 24692 34060 24704
rect 34112 24732 34118 24744
rect 34999 24732 35027 24763
rect 35342 24760 35348 24772
rect 35400 24760 35406 24812
rect 35526 24760 35532 24812
rect 35584 24800 35590 24812
rect 35713 24803 35771 24809
rect 35713 24800 35725 24803
rect 35584 24772 35725 24800
rect 35584 24760 35590 24772
rect 35713 24769 35725 24772
rect 35759 24769 35771 24803
rect 35713 24763 35771 24769
rect 35802 24760 35808 24812
rect 35860 24760 35866 24812
rect 35986 24760 35992 24812
rect 36044 24760 36050 24812
rect 36262 24809 36268 24812
rect 36219 24803 36268 24809
rect 36219 24769 36231 24803
rect 36265 24769 36268 24803
rect 36219 24763 36268 24769
rect 36262 24760 36268 24763
rect 36320 24760 36326 24812
rect 39574 24800 39580 24812
rect 36372 24772 39580 24800
rect 36372 24732 36400 24772
rect 39574 24760 39580 24772
rect 39632 24760 39638 24812
rect 34112 24704 36400 24732
rect 34112 24692 34118 24704
rect 36446 24692 36452 24744
rect 36504 24732 36510 24744
rect 37921 24735 37979 24741
rect 37921 24732 37933 24735
rect 36504 24704 37933 24732
rect 36504 24692 36510 24704
rect 37921 24701 37933 24704
rect 37967 24701 37979 24735
rect 37921 24695 37979 24701
rect 38010 24692 38016 24744
rect 38068 24692 38074 24744
rect 33152 24664 33180 24692
rect 35434 24664 35440 24676
rect 32600 24636 33180 24664
rect 33336 24636 35440 24664
rect 32309 24627 32367 24633
rect 33336 24596 33364 24636
rect 35434 24624 35440 24636
rect 35492 24624 35498 24676
rect 35728 24636 37127 24664
rect 31680 24568 33364 24596
rect 33410 24556 33416 24608
rect 33468 24556 33474 24608
rect 33870 24556 33876 24608
rect 33928 24596 33934 24608
rect 34238 24596 34244 24608
rect 33928 24568 34244 24596
rect 33928 24556 33934 24568
rect 34238 24556 34244 24568
rect 34296 24556 34302 24608
rect 35253 24599 35311 24605
rect 35253 24565 35265 24599
rect 35299 24596 35311 24599
rect 35728 24596 35756 24636
rect 35299 24568 35756 24596
rect 35299 24565 35311 24568
rect 35253 24559 35311 24565
rect 35802 24556 35808 24608
rect 35860 24596 35866 24608
rect 36357 24599 36415 24605
rect 36357 24596 36369 24599
rect 35860 24568 36369 24596
rect 35860 24556 35866 24568
rect 36357 24565 36369 24568
rect 36403 24565 36415 24599
rect 37099 24596 37127 24636
rect 37182 24624 37188 24676
rect 37240 24664 37246 24676
rect 37461 24667 37519 24673
rect 37461 24664 37473 24667
rect 37240 24636 37473 24664
rect 37240 24624 37246 24636
rect 37461 24633 37473 24636
rect 37507 24633 37519 24667
rect 37461 24627 37519 24633
rect 37366 24596 37372 24608
rect 37099 24568 37372 24596
rect 36357 24559 36415 24565
rect 37366 24556 37372 24568
rect 37424 24556 37430 24608
rect 37642 24556 37648 24608
rect 37700 24596 37706 24608
rect 37918 24596 37924 24608
rect 37700 24568 37924 24596
rect 37700 24556 37706 24568
rect 37918 24556 37924 24568
rect 37976 24556 37982 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 2682 24352 2688 24404
rect 2740 24392 2746 24404
rect 14461 24395 14519 24401
rect 2740 24352 2774 24392
rect 14461 24361 14473 24395
rect 14507 24392 14519 24395
rect 15286 24392 15292 24404
rect 14507 24364 15292 24392
rect 14507 24361 14519 24364
rect 14461 24355 14519 24361
rect 15286 24352 15292 24364
rect 15344 24352 15350 24404
rect 16206 24352 16212 24404
rect 16264 24392 16270 24404
rect 18601 24395 18659 24401
rect 18601 24392 18613 24395
rect 16264 24364 18613 24392
rect 16264 24352 16270 24364
rect 18601 24361 18613 24364
rect 18647 24361 18659 24395
rect 18601 24355 18659 24361
rect 18690 24352 18696 24404
rect 18748 24352 18754 24404
rect 18874 24352 18880 24404
rect 18932 24392 18938 24404
rect 19610 24392 19616 24404
rect 18932 24364 19616 24392
rect 18932 24352 18938 24364
rect 19610 24352 19616 24364
rect 19668 24392 19674 24404
rect 19668 24364 20760 24392
rect 19668 24352 19674 24364
rect 2746 24052 2774 24352
rect 12161 24327 12219 24333
rect 12161 24293 12173 24327
rect 12207 24324 12219 24327
rect 14734 24324 14740 24336
rect 12207 24296 14740 24324
rect 12207 24293 12219 24296
rect 12161 24287 12219 24293
rect 11974 24216 11980 24268
rect 12032 24256 12038 24268
rect 12176 24256 12204 24287
rect 14734 24284 14740 24296
rect 14792 24284 14798 24336
rect 16393 24327 16451 24333
rect 16393 24293 16405 24327
rect 16439 24324 16451 24327
rect 19334 24324 19340 24336
rect 16439 24296 19340 24324
rect 16439 24293 16451 24296
rect 16393 24287 16451 24293
rect 12032 24228 12204 24256
rect 12032 24216 12038 24228
rect 12894 24216 12900 24268
rect 12952 24256 12958 24268
rect 13446 24256 13452 24268
rect 12952 24228 13452 24256
rect 12952 24216 12958 24228
rect 13446 24216 13452 24228
rect 13504 24256 13510 24268
rect 15013 24259 15071 24265
rect 15013 24256 15025 24259
rect 13504 24228 15025 24256
rect 13504 24216 13510 24228
rect 15013 24225 15025 24228
rect 15059 24225 15071 24259
rect 15013 24219 15071 24225
rect 8202 24148 8208 24200
rect 8260 24188 8266 24200
rect 10781 24191 10839 24197
rect 10781 24188 10793 24191
rect 8260 24160 10793 24188
rect 8260 24148 8266 24160
rect 10781 24157 10793 24160
rect 10827 24188 10839 24191
rect 11422 24188 11428 24200
rect 10827 24160 11428 24188
rect 10827 24157 10839 24160
rect 10781 24151 10839 24157
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 13206 24191 13264 24197
rect 13206 24188 13218 24191
rect 12400 24160 13218 24188
rect 12400 24148 12406 24160
rect 13206 24157 13218 24160
rect 13252 24157 13264 24191
rect 13206 24151 13264 24157
rect 13633 24191 13691 24197
rect 13633 24157 13645 24191
rect 13679 24157 13691 24191
rect 13633 24151 13691 24157
rect 11048 24123 11106 24129
rect 11048 24089 11060 24123
rect 11094 24120 11106 24123
rect 12250 24120 12256 24132
rect 11094 24092 12256 24120
rect 11094 24089 11106 24092
rect 11048 24083 11106 24089
rect 12250 24080 12256 24092
rect 12308 24080 12314 24132
rect 13648 24120 13676 24151
rect 13722 24148 13728 24200
rect 13780 24148 13786 24200
rect 14369 24191 14427 24197
rect 14369 24157 14381 24191
rect 14415 24188 14427 24191
rect 14826 24188 14832 24200
rect 14415 24160 14832 24188
rect 14415 24157 14427 24160
rect 14369 24151 14427 24157
rect 14826 24148 14832 24160
rect 14884 24148 14890 24200
rect 15654 24148 15660 24200
rect 15712 24188 15718 24200
rect 16408 24188 16436 24287
rect 19334 24284 19340 24296
rect 19392 24284 19398 24336
rect 17310 24216 17316 24268
rect 17368 24216 17374 24268
rect 17402 24216 17408 24268
rect 17460 24216 17466 24268
rect 18509 24259 18567 24265
rect 18509 24256 18521 24259
rect 17512 24228 18521 24256
rect 15712 24160 16436 24188
rect 15712 24148 15718 24160
rect 16574 24148 16580 24200
rect 16632 24188 16638 24200
rect 17512 24188 17540 24228
rect 18509 24225 18521 24228
rect 18555 24225 18567 24259
rect 20732 24256 20760 24364
rect 20898 24352 20904 24404
rect 20956 24392 20962 24404
rect 20993 24395 21051 24401
rect 20993 24392 21005 24395
rect 20956 24364 21005 24392
rect 20956 24352 20962 24364
rect 20993 24361 21005 24364
rect 21039 24361 21051 24395
rect 20993 24355 21051 24361
rect 21818 24352 21824 24404
rect 21876 24392 21882 24404
rect 21913 24395 21971 24401
rect 21913 24392 21925 24395
rect 21876 24364 21925 24392
rect 21876 24352 21882 24364
rect 21913 24361 21925 24364
rect 21959 24361 21971 24395
rect 21913 24355 21971 24361
rect 22462 24352 22468 24404
rect 22520 24392 22526 24404
rect 30374 24392 30380 24404
rect 22520 24364 30380 24392
rect 22520 24352 22526 24364
rect 30374 24352 30380 24364
rect 30432 24352 30438 24404
rect 31754 24352 31760 24404
rect 31812 24352 31818 24404
rect 32674 24352 32680 24404
rect 32732 24352 32738 24404
rect 33226 24352 33232 24404
rect 33284 24392 33290 24404
rect 33284 24364 33364 24392
rect 33284 24352 33290 24364
rect 20806 24284 20812 24336
rect 20864 24324 20870 24336
rect 26694 24324 26700 24336
rect 20864 24296 26700 24324
rect 20864 24284 20870 24296
rect 22462 24256 22468 24268
rect 20732 24228 22468 24256
rect 18509 24219 18567 24225
rect 22462 24216 22468 24228
rect 22520 24216 22526 24268
rect 22554 24216 22560 24268
rect 22612 24216 22618 24268
rect 23753 24259 23811 24265
rect 23753 24225 23765 24259
rect 23799 24256 23811 24259
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 23799 24228 24593 24256
rect 23799 24225 23811 24228
rect 23753 24219 23811 24225
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 16632 24160 17540 24188
rect 16632 24148 16638 24160
rect 18414 24148 18420 24200
rect 18472 24188 18478 24200
rect 18472 24160 18552 24188
rect 18472 24148 18478 24160
rect 13998 24120 14004 24132
rect 13648 24092 14004 24120
rect 13998 24080 14004 24092
rect 14056 24120 14062 24132
rect 15010 24120 15016 24132
rect 14056 24092 15016 24120
rect 14056 24080 14062 24092
rect 15010 24080 15016 24092
rect 15068 24080 15074 24132
rect 15280 24123 15338 24129
rect 15280 24089 15292 24123
rect 15326 24120 15338 24123
rect 15930 24120 15936 24132
rect 15326 24092 15936 24120
rect 15326 24089 15338 24092
rect 15280 24083 15338 24089
rect 15930 24080 15936 24092
rect 15988 24080 15994 24132
rect 12986 24052 12992 24064
rect 2746 24024 12992 24052
rect 12986 24012 12992 24024
rect 13044 24012 13050 24064
rect 13078 24012 13084 24064
rect 13136 24012 13142 24064
rect 13265 24055 13323 24061
rect 13265 24021 13277 24055
rect 13311 24052 13323 24055
rect 13354 24052 13360 24064
rect 13311 24024 13360 24052
rect 13311 24021 13323 24024
rect 13265 24015 13323 24021
rect 13354 24012 13360 24024
rect 13412 24012 13418 24064
rect 16850 24012 16856 24064
rect 16908 24012 16914 24064
rect 17126 24012 17132 24064
rect 17184 24052 17190 24064
rect 17221 24055 17279 24061
rect 17221 24052 17233 24055
rect 17184 24024 17233 24052
rect 17184 24012 17190 24024
rect 17221 24021 17233 24024
rect 17267 24021 17279 24055
rect 17221 24015 17279 24021
rect 18141 24055 18199 24061
rect 18141 24021 18153 24055
rect 18187 24052 18199 24055
rect 18414 24052 18420 24064
rect 18187 24024 18420 24052
rect 18187 24021 18199 24024
rect 18141 24015 18199 24021
rect 18414 24012 18420 24024
rect 18472 24012 18478 24064
rect 18524 24052 18552 24160
rect 18598 24148 18604 24200
rect 18656 24188 18662 24200
rect 18877 24191 18935 24197
rect 18877 24188 18889 24191
rect 18656 24160 18889 24188
rect 18656 24148 18662 24160
rect 18877 24157 18889 24160
rect 18923 24188 18935 24191
rect 19058 24188 19064 24200
rect 18923 24160 19064 24188
rect 18923 24157 18935 24160
rect 18877 24151 18935 24157
rect 19058 24148 19064 24160
rect 19116 24148 19122 24200
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24188 19671 24191
rect 22002 24188 22008 24200
rect 19659 24160 22008 24188
rect 19659 24157 19671 24160
rect 19613 24151 19671 24157
rect 22002 24148 22008 24160
rect 22060 24148 22066 24200
rect 23474 24148 23480 24200
rect 23532 24148 23538 24200
rect 24780 24197 24808 24296
rect 26694 24284 26700 24296
rect 26752 24324 26758 24336
rect 28350 24324 28356 24336
rect 26752 24296 28356 24324
rect 26752 24284 26758 24296
rect 28350 24284 28356 24296
rect 28408 24284 28414 24336
rect 28905 24327 28963 24333
rect 28905 24293 28917 24327
rect 28951 24324 28963 24327
rect 29638 24324 29644 24336
rect 28951 24296 29644 24324
rect 28951 24293 28963 24296
rect 28905 24287 28963 24293
rect 29638 24284 29644 24296
rect 29696 24284 29702 24336
rect 29841 24296 30144 24324
rect 24854 24216 24860 24268
rect 24912 24256 24918 24268
rect 24912 24228 25268 24256
rect 24912 24216 24918 24228
rect 24765 24191 24823 24197
rect 24765 24157 24777 24191
rect 24811 24157 24823 24191
rect 24765 24151 24823 24157
rect 24946 24148 24952 24200
rect 25004 24188 25010 24200
rect 25240 24197 25268 24228
rect 25682 24216 25688 24268
rect 25740 24256 25746 24268
rect 27154 24256 27160 24268
rect 25740 24228 27160 24256
rect 25740 24216 25746 24228
rect 27154 24216 27160 24228
rect 27212 24216 27218 24268
rect 27798 24216 27804 24268
rect 27856 24256 27862 24268
rect 27856 24228 28304 24256
rect 27856 24216 27862 24228
rect 25041 24191 25099 24197
rect 25041 24188 25053 24191
rect 25004 24160 25053 24188
rect 25004 24148 25010 24160
rect 25041 24157 25053 24160
rect 25087 24157 25099 24191
rect 25041 24151 25099 24157
rect 25225 24191 25283 24197
rect 25225 24157 25237 24191
rect 25271 24157 25283 24191
rect 25866 24188 25872 24200
rect 25225 24151 25283 24157
rect 25332 24160 25872 24188
rect 19880 24123 19938 24129
rect 19880 24089 19892 24123
rect 19926 24120 19938 24123
rect 20530 24120 20536 24132
rect 19926 24092 20536 24120
rect 19926 24089 19938 24092
rect 19880 24083 19938 24089
rect 20530 24080 20536 24092
rect 20588 24080 20594 24132
rect 22281 24123 22339 24129
rect 22281 24089 22293 24123
rect 22327 24120 22339 24123
rect 23842 24120 23848 24132
rect 22327 24092 23848 24120
rect 22327 24089 22339 24092
rect 22281 24083 22339 24089
rect 20070 24052 20076 24064
rect 18524 24024 20076 24052
rect 20070 24012 20076 24024
rect 20128 24012 20134 24064
rect 20254 24012 20260 24064
rect 20312 24052 20318 24064
rect 22296 24052 22324 24083
rect 23842 24080 23848 24092
rect 23900 24080 23906 24132
rect 23934 24080 23940 24132
rect 23992 24120 23998 24132
rect 25332 24120 25360 24160
rect 25866 24148 25872 24160
rect 25924 24148 25930 24200
rect 26234 24148 26240 24200
rect 26292 24188 26298 24200
rect 26329 24191 26387 24197
rect 26329 24188 26341 24191
rect 26292 24160 26341 24188
rect 26292 24148 26298 24160
rect 26329 24157 26341 24160
rect 26375 24157 26387 24191
rect 26329 24151 26387 24157
rect 26421 24191 26479 24197
rect 26421 24157 26433 24191
rect 26467 24157 26479 24191
rect 26421 24151 26479 24157
rect 26513 24191 26571 24197
rect 26513 24157 26525 24191
rect 26559 24157 26571 24191
rect 26513 24151 26571 24157
rect 23992 24092 25360 24120
rect 23992 24080 23998 24092
rect 25682 24080 25688 24132
rect 25740 24120 25746 24132
rect 26436 24120 26464 24151
rect 25740 24092 26464 24120
rect 25740 24080 25746 24092
rect 26527 24064 26555 24151
rect 26602 24148 26608 24200
rect 26660 24148 26666 24200
rect 26789 24191 26847 24197
rect 26789 24157 26801 24191
rect 26835 24188 26847 24191
rect 27062 24188 27068 24200
rect 26835 24160 27068 24188
rect 26835 24157 26847 24160
rect 26789 24151 26847 24157
rect 27062 24148 27068 24160
rect 27120 24148 27126 24200
rect 27890 24148 27896 24200
rect 27948 24148 27954 24200
rect 27982 24148 27988 24200
rect 28040 24148 28046 24200
rect 28276 24197 28304 24228
rect 28261 24191 28319 24197
rect 28261 24157 28273 24191
rect 28307 24157 28319 24191
rect 28261 24151 28319 24157
rect 28445 24191 28503 24197
rect 28445 24157 28457 24191
rect 28491 24188 28503 24191
rect 29181 24191 29239 24197
rect 29181 24188 29193 24191
rect 28491 24160 29193 24188
rect 28491 24157 28503 24160
rect 28445 24151 28503 24157
rect 29181 24157 29193 24160
rect 29227 24188 29239 24191
rect 29270 24188 29276 24200
rect 29227 24160 29276 24188
rect 29227 24157 29239 24160
rect 29181 24151 29239 24157
rect 29270 24148 29276 24160
rect 29328 24148 29334 24200
rect 29546 24148 29552 24200
rect 29604 24188 29610 24200
rect 29733 24191 29791 24197
rect 29604 24160 29684 24188
rect 29604 24148 29610 24160
rect 26694 24080 26700 24132
rect 26752 24120 26758 24132
rect 27249 24123 27307 24129
rect 27249 24120 27261 24123
rect 26752 24092 27261 24120
rect 26752 24080 26758 24092
rect 27249 24089 27261 24092
rect 27295 24089 27307 24123
rect 27249 24083 27307 24089
rect 28905 24123 28963 24129
rect 28905 24089 28917 24123
rect 28951 24120 28963 24123
rect 29656 24120 29684 24160
rect 29733 24157 29745 24191
rect 29779 24188 29791 24191
rect 29841 24188 29869 24296
rect 30116 24256 30144 24296
rect 30466 24284 30472 24336
rect 30524 24324 30530 24336
rect 30745 24327 30803 24333
rect 30745 24324 30757 24327
rect 30524 24296 30757 24324
rect 30524 24284 30530 24296
rect 30745 24293 30757 24296
rect 30791 24293 30803 24327
rect 30745 24287 30803 24293
rect 32122 24256 32128 24268
rect 30116 24228 32128 24256
rect 32122 24216 32128 24228
rect 32180 24216 32186 24268
rect 29779 24160 29869 24188
rect 30101 24191 30159 24197
rect 29779 24157 29791 24160
rect 29733 24151 29791 24157
rect 30101 24157 30113 24191
rect 30147 24188 30159 24191
rect 30190 24188 30196 24200
rect 30147 24160 30196 24188
rect 30147 24157 30159 24160
rect 30101 24151 30159 24157
rect 30190 24148 30196 24160
rect 30248 24148 30254 24200
rect 30282 24148 30288 24200
rect 30340 24188 30346 24200
rect 30745 24191 30803 24197
rect 30745 24188 30757 24191
rect 30340 24160 30757 24188
rect 30340 24148 30346 24160
rect 30745 24157 30757 24160
rect 30791 24157 30803 24191
rect 30745 24151 30803 24157
rect 31021 24191 31079 24197
rect 31021 24157 31033 24191
rect 31067 24157 31079 24191
rect 31021 24151 31079 24157
rect 31665 24191 31723 24197
rect 31665 24157 31677 24191
rect 31711 24188 31723 24191
rect 31846 24188 31852 24200
rect 31711 24160 31852 24188
rect 31711 24157 31723 24160
rect 31665 24151 31723 24157
rect 29917 24123 29975 24129
rect 29917 24120 29929 24123
rect 28951 24092 29592 24120
rect 29656 24092 29929 24120
rect 28951 24089 28963 24092
rect 28905 24083 28963 24089
rect 20312 24024 22324 24052
rect 22373 24055 22431 24061
rect 20312 24012 20318 24024
rect 22373 24021 22385 24055
rect 22419 24052 22431 24055
rect 23109 24055 23167 24061
rect 23109 24052 23121 24055
rect 22419 24024 23121 24052
rect 22419 24021 22431 24024
rect 22373 24015 22431 24021
rect 23109 24021 23121 24024
rect 23155 24021 23167 24055
rect 23109 24015 23167 24021
rect 23566 24012 23572 24064
rect 23624 24012 23630 24064
rect 25866 24012 25872 24064
rect 25924 24052 25930 24064
rect 26145 24055 26203 24061
rect 26145 24052 26157 24055
rect 25924 24024 26157 24052
rect 25924 24012 25930 24024
rect 26145 24021 26157 24024
rect 26191 24021 26203 24055
rect 26145 24015 26203 24021
rect 26510 24012 26516 24064
rect 26568 24012 26574 24064
rect 29086 24012 29092 24064
rect 29144 24012 29150 24064
rect 29564 24052 29592 24092
rect 29917 24089 29929 24092
rect 29963 24089 29975 24123
rect 29917 24083 29975 24089
rect 30009 24123 30067 24129
rect 30009 24089 30021 24123
rect 30055 24120 30067 24123
rect 30055 24092 30512 24120
rect 30055 24089 30067 24092
rect 30009 24083 30067 24089
rect 30285 24055 30343 24061
rect 30285 24052 30297 24055
rect 29564 24024 30297 24052
rect 30285 24021 30297 24024
rect 30331 24021 30343 24055
rect 30484 24052 30512 24092
rect 30650 24080 30656 24132
rect 30708 24120 30714 24132
rect 31036 24120 31064 24151
rect 31846 24148 31852 24160
rect 31904 24148 31910 24200
rect 33336 24197 33364 24364
rect 33778 24352 33784 24404
rect 33836 24392 33842 24404
rect 35342 24392 35348 24404
rect 33836 24364 35348 24392
rect 33836 24352 33842 24364
rect 35342 24352 35348 24364
rect 35400 24392 35406 24404
rect 36262 24392 36268 24404
rect 35400 24364 36268 24392
rect 35400 24352 35406 24364
rect 36262 24352 36268 24364
rect 36320 24352 36326 24404
rect 33594 24284 33600 24336
rect 33652 24284 33658 24336
rect 34422 24324 34428 24336
rect 33889 24296 34428 24324
rect 33612 24256 33640 24284
rect 33889 24256 33917 24296
rect 34422 24284 34428 24296
rect 34480 24284 34486 24336
rect 34885 24327 34943 24333
rect 34885 24293 34897 24327
rect 34931 24324 34943 24327
rect 35618 24324 35624 24336
rect 34931 24296 35624 24324
rect 34931 24293 34943 24296
rect 34885 24287 34943 24293
rect 35618 24284 35624 24296
rect 35676 24284 35682 24336
rect 35710 24284 35716 24336
rect 35768 24324 35774 24336
rect 36081 24327 36139 24333
rect 36081 24324 36093 24327
rect 35768 24296 36093 24324
rect 35768 24284 35774 24296
rect 36081 24293 36093 24296
rect 36127 24324 36139 24327
rect 36722 24324 36728 24336
rect 36127 24296 36728 24324
rect 36127 24293 36139 24296
rect 36081 24287 36139 24293
rect 36722 24284 36728 24296
rect 36780 24284 36786 24336
rect 33612 24228 33917 24256
rect 33321 24191 33379 24197
rect 33321 24157 33333 24191
rect 33367 24157 33379 24191
rect 33321 24151 33379 24157
rect 33502 24148 33508 24200
rect 33560 24188 33566 24200
rect 33597 24191 33655 24197
rect 33597 24188 33609 24191
rect 33560 24160 33609 24188
rect 33560 24148 33566 24160
rect 33597 24157 33609 24160
rect 33643 24157 33655 24191
rect 33597 24151 33655 24157
rect 33778 24148 33784 24200
rect 33836 24148 33842 24200
rect 33889 24188 33917 24228
rect 34072 24228 35940 24256
rect 33965 24191 34023 24197
rect 33965 24188 33977 24191
rect 33889 24160 33977 24188
rect 33965 24157 33977 24160
rect 34011 24157 34023 24191
rect 33965 24151 34023 24157
rect 30708 24092 31064 24120
rect 31481 24123 31539 24129
rect 30708 24080 30714 24092
rect 31481 24089 31493 24123
rect 31527 24120 31539 24123
rect 32214 24120 32220 24132
rect 31527 24092 32220 24120
rect 31527 24089 31539 24092
rect 31481 24083 31539 24089
rect 32214 24080 32220 24092
rect 32272 24080 32278 24132
rect 32490 24080 32496 24132
rect 32548 24080 32554 24132
rect 32582 24080 32588 24132
rect 32640 24120 32646 24132
rect 32693 24123 32751 24129
rect 32693 24120 32705 24123
rect 32640 24092 32705 24120
rect 32640 24080 32646 24092
rect 32693 24089 32705 24092
rect 32739 24089 32751 24123
rect 32693 24083 32751 24089
rect 32784 24092 33364 24120
rect 30834 24052 30840 24064
rect 30484 24024 30840 24052
rect 30285 24015 30343 24021
rect 30834 24012 30840 24024
rect 30892 24012 30898 24064
rect 30929 24055 30987 24061
rect 30929 24021 30941 24055
rect 30975 24052 30987 24055
rect 31110 24052 31116 24064
rect 30975 24024 31116 24052
rect 30975 24021 30987 24024
rect 30929 24015 30987 24021
rect 31110 24012 31116 24024
rect 31168 24052 31174 24064
rect 31662 24052 31668 24064
rect 31168 24024 31668 24052
rect 31168 24012 31174 24024
rect 31662 24012 31668 24024
rect 31720 24012 31726 24064
rect 32122 24012 32128 24064
rect 32180 24052 32186 24064
rect 32784 24052 32812 24092
rect 32180 24024 32812 24052
rect 32180 24012 32186 24024
rect 32858 24012 32864 24064
rect 32916 24012 32922 24064
rect 33336 24052 33364 24092
rect 33410 24080 33416 24132
rect 33468 24120 33474 24132
rect 34072 24120 34100 24228
rect 34882 24148 34888 24200
rect 34940 24148 34946 24200
rect 35066 24148 35072 24200
rect 35124 24188 35130 24200
rect 35161 24191 35219 24197
rect 35161 24188 35173 24191
rect 35124 24160 35173 24188
rect 35124 24148 35130 24160
rect 35161 24157 35173 24160
rect 35207 24157 35219 24191
rect 35161 24151 35219 24157
rect 35802 24148 35808 24200
rect 35860 24148 35866 24200
rect 35912 24197 35940 24228
rect 36906 24216 36912 24268
rect 36964 24216 36970 24268
rect 35897 24191 35955 24197
rect 35897 24157 35909 24191
rect 35943 24157 35955 24191
rect 35897 24151 35955 24157
rect 35986 24148 35992 24200
rect 36044 24188 36050 24200
rect 36173 24191 36231 24197
rect 36173 24188 36185 24191
rect 36044 24160 36185 24188
rect 36044 24148 36050 24160
rect 36173 24157 36185 24160
rect 36219 24188 36231 24191
rect 36262 24188 36268 24200
rect 36219 24160 36268 24188
rect 36219 24157 36231 24160
rect 36173 24151 36231 24157
rect 36262 24148 36268 24160
rect 36320 24148 36326 24200
rect 33468 24092 34100 24120
rect 34149 24123 34207 24129
rect 33468 24080 33474 24092
rect 34149 24089 34161 24123
rect 34195 24120 34207 24123
rect 35250 24120 35256 24132
rect 34195 24092 35256 24120
rect 34195 24089 34207 24092
rect 34149 24083 34207 24089
rect 35250 24080 35256 24092
rect 35308 24080 35314 24132
rect 35621 24123 35679 24129
rect 35621 24089 35633 24123
rect 35667 24120 35679 24123
rect 36446 24120 36452 24132
rect 35667 24092 36452 24120
rect 35667 24089 35679 24092
rect 35621 24083 35679 24089
rect 36446 24080 36452 24092
rect 36504 24080 36510 24132
rect 37176 24123 37234 24129
rect 37176 24089 37188 24123
rect 37222 24120 37234 24123
rect 37458 24120 37464 24132
rect 37222 24092 37464 24120
rect 37222 24089 37234 24092
rect 37176 24083 37234 24089
rect 37458 24080 37464 24092
rect 37516 24080 37522 24132
rect 35069 24055 35127 24061
rect 35069 24052 35081 24055
rect 33336 24024 35081 24052
rect 35069 24021 35081 24024
rect 35115 24052 35127 24055
rect 36630 24052 36636 24064
rect 35115 24024 36636 24052
rect 35115 24021 35127 24024
rect 35069 24015 35127 24021
rect 36630 24012 36636 24024
rect 36688 24012 36694 24064
rect 37826 24012 37832 24064
rect 37884 24052 37890 24064
rect 38289 24055 38347 24061
rect 38289 24052 38301 24055
rect 37884 24024 38301 24052
rect 37884 24012 37890 24024
rect 38289 24021 38301 24024
rect 38335 24021 38347 24055
rect 38289 24015 38347 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 10870 23808 10876 23860
rect 10928 23808 10934 23860
rect 12342 23808 12348 23860
rect 12400 23848 12406 23860
rect 12437 23851 12495 23857
rect 12437 23848 12449 23851
rect 12400 23820 12449 23848
rect 12400 23808 12406 23820
rect 12437 23817 12449 23820
rect 12483 23817 12495 23851
rect 12437 23811 12495 23817
rect 13004 23820 15516 23848
rect 9760 23783 9818 23789
rect 9760 23749 9772 23783
rect 9806 23780 9818 23783
rect 10042 23780 10048 23792
rect 9806 23752 10048 23780
rect 9806 23749 9818 23752
rect 9760 23743 9818 23749
rect 10042 23740 10048 23752
rect 10100 23740 10106 23792
rect 8202 23672 8208 23724
rect 8260 23712 8266 23724
rect 9493 23715 9551 23721
rect 9493 23712 9505 23715
rect 8260 23684 9505 23712
rect 8260 23672 8266 23684
rect 9493 23681 9505 23684
rect 9539 23681 9551 23715
rect 9493 23675 9551 23681
rect 12345 23715 12403 23721
rect 12345 23681 12357 23715
rect 12391 23712 12403 23715
rect 12802 23712 12808 23724
rect 12391 23684 12808 23712
rect 12391 23681 12403 23684
rect 12345 23675 12403 23681
rect 12802 23672 12808 23684
rect 12860 23712 12866 23724
rect 13004 23712 13032 23820
rect 13078 23740 13084 23792
rect 13136 23780 13142 23792
rect 13694 23783 13752 23789
rect 13694 23780 13706 23783
rect 13136 23752 13706 23780
rect 13136 23740 13142 23752
rect 13694 23749 13706 23752
rect 13740 23749 13752 23783
rect 13694 23743 13752 23749
rect 12860 23684 13032 23712
rect 12860 23672 12866 23684
rect 13446 23672 13452 23724
rect 13504 23672 13510 23724
rect 13998 23712 14004 23724
rect 13556 23684 14004 23712
rect 11054 23604 11060 23656
rect 11112 23644 11118 23656
rect 12250 23644 12256 23656
rect 11112 23616 12256 23644
rect 11112 23604 11118 23616
rect 12250 23604 12256 23616
rect 12308 23644 12314 23656
rect 12621 23647 12679 23653
rect 12621 23644 12633 23647
rect 12308 23616 12633 23644
rect 12308 23604 12314 23616
rect 12621 23613 12633 23616
rect 12667 23644 12679 23647
rect 13556 23644 13584 23684
rect 13998 23672 14004 23684
rect 14056 23672 14062 23724
rect 15381 23715 15439 23721
rect 15381 23681 15393 23715
rect 15427 23681 15439 23715
rect 15488 23712 15516 23820
rect 15930 23808 15936 23860
rect 15988 23808 15994 23860
rect 18141 23851 18199 23857
rect 18141 23817 18153 23851
rect 18187 23848 18199 23851
rect 18874 23848 18880 23860
rect 18187 23820 18880 23848
rect 18187 23817 18199 23820
rect 18141 23811 18199 23817
rect 18874 23808 18880 23820
rect 18932 23808 18938 23860
rect 19610 23808 19616 23860
rect 19668 23848 19674 23860
rect 19889 23851 19947 23857
rect 19889 23848 19901 23851
rect 19668 23820 19901 23848
rect 19668 23808 19674 23820
rect 19889 23817 19901 23820
rect 19935 23848 19947 23851
rect 20254 23848 20260 23860
rect 19935 23820 20260 23848
rect 19935 23817 19947 23820
rect 19889 23811 19947 23817
rect 20254 23808 20260 23820
rect 20312 23808 20318 23860
rect 20438 23808 20444 23860
rect 20496 23808 20502 23860
rect 20530 23808 20536 23860
rect 20588 23848 20594 23860
rect 20990 23848 20996 23860
rect 20588 23820 20996 23848
rect 20588 23808 20594 23820
rect 20990 23808 20996 23820
rect 21048 23848 21054 23860
rect 23290 23848 23296 23860
rect 21048 23820 23296 23848
rect 21048 23808 21054 23820
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 26326 23808 26332 23860
rect 26384 23848 26390 23860
rect 26384 23820 26556 23848
rect 26384 23808 26390 23820
rect 15565 23783 15623 23789
rect 15565 23749 15577 23783
rect 15611 23780 15623 23783
rect 16114 23780 16120 23792
rect 15611 23752 16120 23780
rect 15611 23749 15623 23752
rect 15565 23743 15623 23749
rect 16114 23740 16120 23752
rect 16172 23740 16178 23792
rect 16776 23752 21036 23780
rect 15488 23684 15608 23712
rect 15381 23675 15439 23681
rect 12667 23616 13584 23644
rect 15396 23644 15424 23675
rect 15580 23644 15608 23684
rect 15654 23672 15660 23724
rect 15712 23672 15718 23724
rect 15749 23715 15807 23721
rect 15749 23681 15761 23715
rect 15795 23712 15807 23715
rect 16390 23712 16396 23724
rect 15795 23684 16396 23712
rect 15795 23681 15807 23684
rect 15749 23675 15807 23681
rect 16390 23672 16396 23684
rect 16448 23672 16454 23724
rect 16776 23644 16804 23752
rect 17034 23672 17040 23724
rect 17092 23712 17098 23724
rect 17129 23715 17187 23721
rect 17129 23712 17141 23715
rect 17092 23684 17141 23712
rect 17092 23672 17098 23684
rect 17129 23681 17141 23684
rect 17175 23681 17187 23715
rect 17129 23675 17187 23681
rect 17310 23672 17316 23724
rect 17368 23672 17374 23724
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23712 18291 23715
rect 19426 23712 19432 23724
rect 18279 23684 19432 23712
rect 18279 23681 18291 23684
rect 18233 23675 18291 23681
rect 19426 23672 19432 23684
rect 19484 23672 19490 23724
rect 19702 23672 19708 23724
rect 19760 23672 19766 23724
rect 19981 23715 20039 23721
rect 19981 23681 19993 23715
rect 20027 23712 20039 23715
rect 20530 23712 20536 23724
rect 20027 23684 20536 23712
rect 20027 23681 20039 23684
rect 19981 23675 20039 23681
rect 20530 23672 20536 23684
rect 20588 23672 20594 23724
rect 20622 23672 20628 23724
rect 20680 23672 20686 23724
rect 20898 23672 20904 23724
rect 20956 23672 20962 23724
rect 15396 23616 15516 23644
rect 15580 23616 16804 23644
rect 18417 23647 18475 23653
rect 12667 23613 12679 23616
rect 12621 23607 12679 23613
rect 15488 23576 15516 23616
rect 18417 23613 18429 23647
rect 18463 23644 18475 23647
rect 18463 23616 18552 23644
rect 18463 23613 18475 23616
rect 18417 23607 18475 23613
rect 16666 23576 16672 23588
rect 15488 23548 16672 23576
rect 16666 23536 16672 23548
rect 16724 23536 16730 23588
rect 18524 23576 18552 23616
rect 18966 23604 18972 23656
rect 19024 23644 19030 23656
rect 19886 23644 19892 23656
rect 19024 23616 19892 23644
rect 19024 23604 19030 23616
rect 19886 23604 19892 23616
rect 19944 23604 19950 23656
rect 20070 23604 20076 23656
rect 20128 23644 20134 23656
rect 20809 23647 20867 23653
rect 20809 23644 20821 23647
rect 20128 23616 20821 23644
rect 20128 23604 20134 23616
rect 20809 23613 20821 23616
rect 20855 23613 20867 23647
rect 21008 23644 21036 23752
rect 22370 23740 22376 23792
rect 22428 23740 22434 23792
rect 24578 23740 24584 23792
rect 24636 23780 24642 23792
rect 25130 23780 25136 23792
rect 24636 23752 25136 23780
rect 24636 23740 24642 23752
rect 25130 23740 25136 23752
rect 25188 23740 25194 23792
rect 25958 23740 25964 23792
rect 26016 23780 26022 23792
rect 26528 23780 26556 23820
rect 26602 23808 26608 23860
rect 26660 23848 26666 23860
rect 27157 23851 27215 23857
rect 27157 23848 27169 23851
rect 26660 23820 27169 23848
rect 26660 23808 26666 23820
rect 27157 23817 27169 23820
rect 27203 23817 27215 23851
rect 27157 23811 27215 23817
rect 27525 23851 27583 23857
rect 27525 23817 27537 23851
rect 27571 23848 27583 23851
rect 27798 23848 27804 23860
rect 27571 23820 27804 23848
rect 27571 23817 27583 23820
rect 27525 23811 27583 23817
rect 27798 23808 27804 23820
rect 27856 23848 27862 23860
rect 28902 23848 28908 23860
rect 27856 23820 28908 23848
rect 27856 23808 27862 23820
rect 28902 23808 28908 23820
rect 28960 23808 28966 23860
rect 29454 23848 29460 23860
rect 29196 23820 29460 23848
rect 29196 23780 29224 23820
rect 29454 23808 29460 23820
rect 29512 23808 29518 23860
rect 29546 23808 29552 23860
rect 29604 23848 29610 23860
rect 29604 23820 30241 23848
rect 29604 23808 29610 23820
rect 26016 23752 26372 23780
rect 26528 23752 29224 23780
rect 26016 23740 26022 23752
rect 21082 23672 21088 23724
rect 21140 23712 21146 23724
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 21140 23684 22017 23712
rect 21140 23672 21146 23684
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 22005 23675 22063 23681
rect 22278 23672 22284 23724
rect 22336 23672 22342 23724
rect 22830 23672 22836 23724
rect 22888 23672 22894 23724
rect 23290 23672 23296 23724
rect 23348 23712 23354 23724
rect 25498 23712 25504 23724
rect 23348 23684 25504 23712
rect 23348 23672 23354 23684
rect 25498 23672 25504 23684
rect 25556 23672 25562 23724
rect 25593 23715 25651 23721
rect 25593 23681 25605 23715
rect 25639 23681 25651 23715
rect 25593 23675 25651 23681
rect 25869 23715 25927 23721
rect 25869 23681 25881 23715
rect 25915 23681 25927 23715
rect 25869 23675 25927 23681
rect 25608 23644 25636 23675
rect 21008 23616 25636 23644
rect 20809 23607 20867 23613
rect 18598 23576 18604 23588
rect 16776 23548 18368 23576
rect 18524 23548 18604 23576
rect 11974 23468 11980 23520
rect 12032 23468 12038 23520
rect 13722 23468 13728 23520
rect 13780 23508 13786 23520
rect 14829 23511 14887 23517
rect 14829 23508 14841 23511
rect 13780 23480 14841 23508
rect 13780 23468 13786 23480
rect 14829 23477 14841 23480
rect 14875 23508 14887 23511
rect 16776 23508 16804 23548
rect 14875 23480 16804 23508
rect 14875 23477 14887 23480
rect 14829 23471 14887 23477
rect 17218 23468 17224 23520
rect 17276 23468 17282 23520
rect 17770 23468 17776 23520
rect 17828 23468 17834 23520
rect 18340 23508 18368 23548
rect 18598 23536 18604 23548
rect 18656 23536 18662 23588
rect 19610 23576 19616 23588
rect 19306 23548 19616 23576
rect 19306 23508 19334 23548
rect 19610 23536 19616 23548
rect 19668 23536 19674 23588
rect 19702 23536 19708 23588
rect 19760 23576 19766 23588
rect 22186 23576 22192 23588
rect 19760 23548 22192 23576
rect 19760 23536 19766 23548
rect 22186 23536 22192 23548
rect 22244 23536 22250 23588
rect 24302 23536 24308 23588
rect 24360 23576 24366 23588
rect 25884 23576 25912 23675
rect 26142 23672 26148 23724
rect 26200 23672 26206 23724
rect 26344 23721 26372 23752
rect 29270 23740 29276 23792
rect 29328 23780 29334 23792
rect 29328 23752 30052 23780
rect 29328 23740 29334 23752
rect 26329 23715 26387 23721
rect 26329 23681 26341 23715
rect 26375 23681 26387 23715
rect 26329 23675 26387 23681
rect 27341 23715 27399 23721
rect 27341 23681 27353 23715
rect 27387 23712 27399 23715
rect 27430 23712 27436 23724
rect 27387 23684 27436 23712
rect 27387 23681 27399 23684
rect 27341 23675 27399 23681
rect 27430 23672 27436 23684
rect 27488 23672 27494 23724
rect 27617 23715 27675 23721
rect 27617 23681 27629 23715
rect 27663 23712 27675 23715
rect 28442 23712 28448 23724
rect 27663 23684 28448 23712
rect 27663 23681 27675 23684
rect 27617 23675 27675 23681
rect 26510 23604 26516 23656
rect 26568 23644 26574 23656
rect 27632 23644 27660 23675
rect 28442 23672 28448 23684
rect 28500 23672 28506 23724
rect 28534 23672 28540 23724
rect 28592 23672 28598 23724
rect 28876 23715 28934 23721
rect 28876 23712 28888 23715
rect 28644 23684 28888 23712
rect 26568 23616 27660 23644
rect 26568 23604 26574 23616
rect 28258 23604 28264 23656
rect 28316 23644 28322 23656
rect 28644 23644 28672 23684
rect 28876 23681 28888 23684
rect 28922 23681 28934 23715
rect 28876 23675 28934 23681
rect 29086 23672 29092 23724
rect 29144 23712 29150 23724
rect 30024 23721 30052 23752
rect 30098 23740 30104 23792
rect 30156 23740 30162 23792
rect 30213 23724 30241 23820
rect 33410 23808 33416 23860
rect 33468 23848 33474 23860
rect 33468 23820 34422 23848
rect 33468 23808 33474 23820
rect 31021 23783 31079 23789
rect 31021 23749 31033 23783
rect 31067 23780 31079 23783
rect 31386 23780 31392 23792
rect 31067 23752 31392 23780
rect 31067 23749 31079 23752
rect 31021 23743 31079 23749
rect 31386 23740 31392 23752
rect 31444 23740 31450 23792
rect 32950 23740 32956 23792
rect 33008 23780 33014 23792
rect 33594 23780 33600 23792
rect 33008 23752 33600 23780
rect 33008 23740 33014 23752
rect 33594 23740 33600 23752
rect 33652 23780 33658 23792
rect 34149 23783 34207 23789
rect 34149 23780 34161 23783
rect 33652 23752 34161 23780
rect 33652 23740 33658 23752
rect 34149 23749 34161 23752
rect 34195 23749 34207 23783
rect 34149 23743 34207 23749
rect 34394 23780 34422 23820
rect 34790 23808 34796 23860
rect 34848 23808 34854 23860
rect 34882 23808 34888 23860
rect 34940 23848 34946 23860
rect 35621 23851 35679 23857
rect 35621 23848 35633 23851
rect 34940 23820 35633 23848
rect 34940 23808 34946 23820
rect 35621 23817 35633 23820
rect 35667 23817 35679 23851
rect 35621 23811 35679 23817
rect 37458 23808 37464 23860
rect 37516 23808 37522 23860
rect 37826 23808 37832 23860
rect 37884 23808 37890 23860
rect 34808 23780 34836 23808
rect 35710 23780 35716 23792
rect 34394 23752 34836 23780
rect 35176 23752 35716 23780
rect 29733 23715 29791 23721
rect 29733 23712 29745 23715
rect 29144 23684 29745 23712
rect 29144 23672 29150 23684
rect 29733 23681 29745 23684
rect 29779 23681 29791 23715
rect 29733 23675 29791 23681
rect 29881 23715 29939 23721
rect 29881 23681 29893 23715
rect 29927 23681 29939 23715
rect 29881 23675 29939 23681
rect 30009 23715 30067 23721
rect 30009 23681 30021 23715
rect 30055 23681 30067 23715
rect 30009 23675 30067 23681
rect 28316 23616 28672 23644
rect 28702 23616 28948 23644
rect 28316 23604 28322 23616
rect 28702 23576 28730 23616
rect 24360 23548 25268 23576
rect 25884 23548 28730 23576
rect 28920 23576 28948 23616
rect 29270 23604 29276 23656
rect 29328 23604 29334 23656
rect 29288 23576 29316 23604
rect 28920 23548 29316 23576
rect 24360 23536 24366 23548
rect 18340 23480 19334 23508
rect 19521 23511 19579 23517
rect 19521 23477 19533 23511
rect 19567 23508 19579 23511
rect 20530 23508 20536 23520
rect 19567 23480 20536 23508
rect 19567 23477 19579 23480
rect 19521 23471 19579 23477
rect 20530 23468 20536 23480
rect 20588 23468 20594 23520
rect 20622 23468 20628 23520
rect 20680 23508 20686 23520
rect 21634 23508 21640 23520
rect 20680 23480 21640 23508
rect 20680 23468 20686 23480
rect 21634 23468 21640 23480
rect 21692 23468 21698 23520
rect 25130 23468 25136 23520
rect 25188 23468 25194 23520
rect 25240 23508 25268 23548
rect 29730 23536 29736 23588
rect 29788 23576 29794 23588
rect 29896 23576 29924 23675
rect 29788 23548 29924 23576
rect 30024 23576 30052 23675
rect 30190 23672 30196 23724
rect 30248 23721 30254 23724
rect 30248 23675 30256 23721
rect 30248 23672 30254 23675
rect 30374 23672 30380 23724
rect 30432 23712 30438 23724
rect 30837 23715 30895 23721
rect 30837 23712 30849 23715
rect 30432 23684 30849 23712
rect 30432 23672 30438 23684
rect 30837 23681 30849 23684
rect 30883 23681 30895 23715
rect 30837 23675 30895 23681
rect 30926 23672 30932 23724
rect 30984 23712 30990 23724
rect 31113 23715 31171 23721
rect 31113 23712 31125 23715
rect 30984 23684 31125 23712
rect 30984 23672 30990 23684
rect 31113 23681 31125 23684
rect 31159 23681 31171 23715
rect 31113 23675 31171 23681
rect 31205 23715 31263 23721
rect 31205 23681 31217 23715
rect 31251 23712 31263 23715
rect 31294 23712 31300 23724
rect 31251 23684 31300 23712
rect 31251 23681 31263 23684
rect 31205 23675 31263 23681
rect 31128 23644 31156 23675
rect 31294 23672 31300 23684
rect 31352 23672 31358 23724
rect 32122 23712 32128 23724
rect 31956 23684 32128 23712
rect 31956 23644 31984 23684
rect 32122 23672 32128 23684
rect 32180 23672 32186 23724
rect 32306 23672 32312 23724
rect 32364 23712 32370 23724
rect 32582 23712 32588 23724
rect 32364 23684 32588 23712
rect 32364 23672 32370 23684
rect 32582 23672 32588 23684
rect 32640 23712 32646 23724
rect 32677 23715 32735 23721
rect 32677 23712 32689 23715
rect 32640 23684 32689 23712
rect 32640 23672 32646 23684
rect 32677 23681 32689 23684
rect 32723 23681 32735 23715
rect 32677 23675 32735 23681
rect 32766 23672 32772 23724
rect 32824 23712 32830 23724
rect 33229 23715 33287 23721
rect 33229 23712 33241 23715
rect 32824 23684 33241 23712
rect 32824 23672 32830 23684
rect 33229 23681 33241 23684
rect 33275 23712 33287 23715
rect 33778 23712 33784 23724
rect 33275 23684 33784 23712
rect 33275 23681 33287 23684
rect 33229 23675 33287 23681
rect 33778 23672 33784 23684
rect 33836 23672 33842 23724
rect 33870 23672 33876 23724
rect 33928 23672 33934 23724
rect 34021 23715 34079 23721
rect 34021 23681 34033 23715
rect 34067 23712 34079 23715
rect 34067 23684 34192 23712
rect 34067 23681 34079 23684
rect 34021 23675 34079 23681
rect 34164 23656 34192 23684
rect 34238 23672 34244 23724
rect 34296 23672 34302 23724
rect 34394 23721 34422 23752
rect 34379 23715 34437 23721
rect 34379 23681 34391 23715
rect 34425 23681 34437 23715
rect 34379 23675 34437 23681
rect 34606 23672 34612 23724
rect 34664 23712 34670 23724
rect 34790 23712 34796 23724
rect 34664 23684 34796 23712
rect 34664 23672 34670 23684
rect 34790 23672 34796 23684
rect 34848 23712 34854 23724
rect 35176 23721 35204 23752
rect 35710 23740 35716 23752
rect 35768 23780 35774 23792
rect 37844 23780 37872 23808
rect 35768 23752 37872 23780
rect 35768 23740 35774 23752
rect 34977 23715 35035 23721
rect 34977 23712 34989 23715
rect 34848 23684 34989 23712
rect 34848 23672 34854 23684
rect 34977 23681 34989 23684
rect 35023 23681 35035 23715
rect 34977 23675 35035 23681
rect 35125 23715 35204 23721
rect 35125 23681 35137 23715
rect 35171 23684 35204 23715
rect 35171 23681 35183 23684
rect 35125 23675 35183 23681
rect 35250 23672 35256 23724
rect 35308 23672 35314 23724
rect 35345 23715 35403 23721
rect 35345 23681 35357 23715
rect 35391 23681 35403 23715
rect 35345 23675 35403 23681
rect 31128 23616 31984 23644
rect 32030 23604 32036 23656
rect 32088 23644 32094 23656
rect 32401 23647 32459 23653
rect 32401 23644 32413 23647
rect 32088 23616 32413 23644
rect 32088 23604 32094 23616
rect 32401 23613 32413 23616
rect 32447 23613 32459 23647
rect 32401 23607 32459 23613
rect 33413 23647 33471 23653
rect 33413 23613 33425 23647
rect 33459 23644 33471 23647
rect 33502 23644 33508 23656
rect 33459 23616 33508 23644
rect 33459 23613 33471 23616
rect 33413 23607 33471 23613
rect 33502 23604 33508 23616
rect 33560 23604 33566 23656
rect 33594 23604 33600 23656
rect 33652 23644 33658 23656
rect 34146 23644 34152 23656
rect 33652 23616 34152 23644
rect 33652 23604 33658 23616
rect 34146 23604 34152 23616
rect 34204 23644 34210 23656
rect 35360 23644 35388 23675
rect 35434 23672 35440 23724
rect 35492 23721 35498 23724
rect 35492 23712 35500 23721
rect 35492 23684 35537 23712
rect 35492 23675 35500 23684
rect 35492 23672 35498 23675
rect 35894 23672 35900 23724
rect 35952 23712 35958 23724
rect 36265 23715 36323 23721
rect 36265 23712 36277 23715
rect 35952 23684 36277 23712
rect 35952 23672 35958 23684
rect 36265 23681 36277 23684
rect 36311 23681 36323 23715
rect 36265 23675 36323 23681
rect 36354 23672 36360 23724
rect 36412 23672 36418 23724
rect 36630 23672 36636 23724
rect 36688 23712 36694 23724
rect 37458 23712 37464 23724
rect 36688 23684 37464 23712
rect 36688 23672 36694 23684
rect 37458 23672 37464 23684
rect 37516 23672 37522 23724
rect 34204 23616 35388 23644
rect 34204 23604 34210 23616
rect 35986 23604 35992 23656
rect 36044 23644 36050 23656
rect 36081 23647 36139 23653
rect 36081 23644 36093 23647
rect 36044 23616 36093 23644
rect 36044 23604 36050 23616
rect 36081 23613 36093 23616
rect 36127 23644 36139 23647
rect 37921 23647 37979 23653
rect 37921 23644 37933 23647
rect 36127 23616 37933 23644
rect 36127 23613 36139 23616
rect 36081 23607 36139 23613
rect 37921 23613 37933 23616
rect 37967 23613 37979 23647
rect 37921 23607 37979 23613
rect 38010 23604 38016 23656
rect 38068 23604 38074 23656
rect 30650 23576 30656 23588
rect 30024 23548 30656 23576
rect 29788 23536 29794 23548
rect 30650 23536 30656 23548
rect 30708 23536 30714 23588
rect 32858 23536 32864 23588
rect 32916 23576 32922 23588
rect 36262 23576 36268 23588
rect 32916 23548 36268 23576
rect 32916 23536 32922 23548
rect 36262 23536 36268 23548
rect 36320 23536 36326 23588
rect 36538 23536 36544 23588
rect 36596 23576 36602 23588
rect 36722 23576 36728 23588
rect 36596 23548 36728 23576
rect 36596 23536 36602 23548
rect 36722 23536 36728 23548
rect 36780 23536 36786 23588
rect 25774 23508 25780 23520
rect 25240 23480 25780 23508
rect 25774 23468 25780 23480
rect 25832 23508 25838 23520
rect 27338 23508 27344 23520
rect 25832 23480 27344 23508
rect 25832 23468 25838 23480
rect 27338 23468 27344 23480
rect 27396 23468 27402 23520
rect 27706 23468 27712 23520
rect 27764 23508 27770 23520
rect 28675 23511 28733 23517
rect 28675 23508 28687 23511
rect 27764 23480 28687 23508
rect 27764 23468 27770 23480
rect 28675 23477 28687 23480
rect 28721 23477 28733 23511
rect 28675 23471 28733 23477
rect 28810 23468 28816 23520
rect 28868 23508 28874 23520
rect 29638 23508 29644 23520
rect 28868 23480 29644 23508
rect 28868 23468 28874 23480
rect 29638 23468 29644 23480
rect 29696 23468 29702 23520
rect 30374 23468 30380 23520
rect 30432 23468 30438 23520
rect 31386 23468 31392 23520
rect 31444 23468 31450 23520
rect 33226 23468 33232 23520
rect 33284 23508 33290 23520
rect 34330 23508 34336 23520
rect 33284 23480 34336 23508
rect 33284 23468 33290 23480
rect 34330 23468 34336 23480
rect 34388 23468 34394 23520
rect 34514 23468 34520 23520
rect 34572 23468 34578 23520
rect 35250 23468 35256 23520
rect 35308 23508 35314 23520
rect 36078 23508 36084 23520
rect 35308 23480 36084 23508
rect 35308 23468 35314 23480
rect 36078 23468 36084 23480
rect 36136 23468 36142 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 7190 23264 7196 23316
rect 7248 23304 7254 23316
rect 11238 23304 11244 23316
rect 7248 23276 11244 23304
rect 7248 23264 7254 23276
rect 11238 23264 11244 23276
rect 11296 23264 11302 23316
rect 12802 23264 12808 23316
rect 12860 23264 12866 23316
rect 15010 23264 15016 23316
rect 15068 23264 15074 23316
rect 17310 23264 17316 23316
rect 17368 23304 17374 23316
rect 23293 23307 23351 23313
rect 17368 23276 21772 23304
rect 17368 23264 17374 23276
rect 18874 23196 18880 23248
rect 18932 23196 18938 23248
rect 19886 23196 19892 23248
rect 19944 23236 19950 23248
rect 20622 23236 20628 23248
rect 19944 23208 20628 23236
rect 19944 23196 19950 23208
rect 20622 23196 20628 23208
rect 20680 23196 20686 23248
rect 11422 23128 11428 23180
rect 11480 23128 11486 23180
rect 19334 23128 19340 23180
rect 19392 23168 19398 23180
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 19392 23140 19441 23168
rect 19392 23128 19398 23140
rect 19429 23137 19441 23140
rect 19475 23168 19487 23171
rect 20162 23168 20168 23180
rect 19475 23140 20168 23168
rect 19475 23137 19487 23140
rect 19429 23131 19487 23137
rect 20162 23128 20168 23140
rect 20220 23128 20226 23180
rect 21744 23168 21772 23276
rect 23293 23273 23305 23307
rect 23339 23304 23351 23307
rect 23566 23304 23572 23316
rect 23339 23276 23572 23304
rect 23339 23273 23351 23276
rect 23293 23267 23351 23273
rect 23566 23264 23572 23276
rect 23624 23264 23630 23316
rect 23750 23264 23756 23316
rect 23808 23304 23814 23316
rect 24762 23304 24768 23316
rect 23808 23276 24768 23304
rect 23808 23264 23814 23276
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 27982 23264 27988 23316
rect 28040 23304 28046 23316
rect 28040 23276 30788 23304
rect 28040 23264 28046 23276
rect 22097 23239 22155 23245
rect 22097 23205 22109 23239
rect 22143 23236 22155 23239
rect 22143 23208 24992 23236
rect 22143 23205 22155 23208
rect 22097 23199 22155 23205
rect 23658 23168 23664 23180
rect 21744 23140 23664 23168
rect 23658 23128 23664 23140
rect 23716 23168 23722 23180
rect 23937 23171 23995 23177
rect 23716 23140 23888 23168
rect 23716 23128 23722 23140
rect 11692 23103 11750 23109
rect 11692 23069 11704 23103
rect 11738 23100 11750 23103
rect 11974 23100 11980 23112
rect 11738 23072 11980 23100
rect 11738 23069 11750 23072
rect 11692 23063 11750 23069
rect 11974 23060 11980 23072
rect 12032 23060 12038 23112
rect 13814 23060 13820 23112
rect 13872 23100 13878 23112
rect 14829 23103 14887 23109
rect 14829 23100 14841 23103
rect 13872 23072 14841 23100
rect 13872 23060 13878 23072
rect 14829 23069 14841 23072
rect 14875 23069 14887 23103
rect 14829 23063 14887 23069
rect 15102 23060 15108 23112
rect 15160 23060 15166 23112
rect 15470 23060 15476 23112
rect 15528 23100 15534 23112
rect 15565 23103 15623 23109
rect 15565 23100 15577 23103
rect 15528 23072 15577 23100
rect 15528 23060 15534 23072
rect 15565 23069 15577 23072
rect 15611 23100 15623 23103
rect 17497 23103 17555 23109
rect 17497 23100 17509 23103
rect 15611 23072 17509 23100
rect 15611 23069 15623 23072
rect 15565 23063 15623 23069
rect 17497 23069 17509 23072
rect 17543 23100 17555 23103
rect 17696 23100 17816 23102
rect 19150 23100 19156 23112
rect 17543 23074 19156 23100
rect 17543 23072 17724 23074
rect 17788 23072 19156 23074
rect 17543 23069 17555 23072
rect 17497 23063 17555 23069
rect 19150 23060 19156 23072
rect 19208 23060 19214 23112
rect 19610 23060 19616 23112
rect 19668 23060 19674 23112
rect 19702 23060 19708 23112
rect 19760 23100 19766 23112
rect 20346 23100 20352 23112
rect 19760 23072 20352 23100
rect 19760 23060 19766 23072
rect 20346 23060 20352 23072
rect 20404 23060 20410 23112
rect 20714 23060 20720 23112
rect 20772 23100 20778 23112
rect 22002 23100 22008 23112
rect 20772 23072 22008 23100
rect 20772 23060 20778 23072
rect 22002 23060 22008 23072
rect 22060 23060 22066 23112
rect 22922 23060 22928 23112
rect 22980 23100 22986 23112
rect 23750 23100 23756 23112
rect 22980 23072 23756 23100
rect 22980 23060 22986 23072
rect 23750 23060 23756 23072
rect 23808 23060 23814 23112
rect 23860 23100 23888 23140
rect 23937 23137 23949 23171
rect 23983 23168 23995 23171
rect 24854 23168 24860 23180
rect 23983 23140 24860 23168
rect 23983 23137 23995 23140
rect 23937 23131 23995 23137
rect 24854 23128 24860 23140
rect 24912 23128 24918 23180
rect 24964 23168 24992 23208
rect 28442 23196 28448 23248
rect 28500 23196 28506 23248
rect 28534 23196 28540 23248
rect 28592 23236 28598 23248
rect 28905 23239 28963 23245
rect 28905 23236 28917 23239
rect 28592 23208 28917 23236
rect 28592 23196 28598 23208
rect 28905 23205 28917 23208
rect 28951 23205 28963 23239
rect 28905 23199 28963 23205
rect 29270 23196 29276 23248
rect 29328 23236 29334 23248
rect 29328 23208 30512 23236
rect 29328 23196 29334 23208
rect 25314 23168 25320 23180
rect 24964 23140 25320 23168
rect 25314 23128 25320 23140
rect 25372 23128 25378 23180
rect 26697 23171 26755 23177
rect 25424 23140 26464 23168
rect 24210 23100 24216 23112
rect 23860 23072 24216 23100
rect 24210 23060 24216 23072
rect 24268 23060 24274 23112
rect 24302 23060 24308 23112
rect 24360 23100 24366 23112
rect 24581 23103 24639 23109
rect 24581 23100 24593 23103
rect 24360 23072 24593 23100
rect 24360 23060 24366 23072
rect 24581 23069 24593 23072
rect 24627 23069 24639 23103
rect 24581 23063 24639 23069
rect 24762 23060 24768 23112
rect 24820 23100 24826 23112
rect 25424 23109 25452 23140
rect 25409 23103 25467 23109
rect 25409 23100 25421 23103
rect 24820 23072 25421 23100
rect 24820 23060 24826 23072
rect 25409 23069 25421 23072
rect 25455 23069 25467 23103
rect 25409 23063 25467 23069
rect 25498 23060 25504 23112
rect 25556 23100 25562 23112
rect 25593 23103 25651 23109
rect 25593 23100 25605 23103
rect 25556 23072 25605 23100
rect 25556 23060 25562 23072
rect 25593 23069 25605 23072
rect 25639 23069 25651 23103
rect 25593 23063 25651 23069
rect 25682 23060 25688 23112
rect 25740 23100 25746 23112
rect 26145 23103 26203 23109
rect 26145 23100 26157 23103
rect 25740 23072 26157 23100
rect 25740 23060 25746 23072
rect 26145 23069 26157 23072
rect 26191 23069 26203 23103
rect 26145 23063 26203 23069
rect 26329 23103 26387 23109
rect 26329 23069 26341 23103
rect 26375 23069 26387 23103
rect 26329 23063 26387 23069
rect 15832 23035 15890 23041
rect 15832 23001 15844 23035
rect 15878 23032 15890 23035
rect 16850 23032 16856 23044
rect 15878 23004 16856 23032
rect 15878 23001 15890 23004
rect 15832 22995 15890 23001
rect 16850 22992 16856 23004
rect 16908 22992 16914 23044
rect 17761 23041 17767 23044
rect 17753 23035 17767 23041
rect 17753 23001 17765 23035
rect 17819 23032 17825 23044
rect 17819 23004 17853 23032
rect 17753 22995 17767 23001
rect 17761 22992 17767 22995
rect 17819 22992 17825 23004
rect 18598 22992 18604 23044
rect 18656 23032 18662 23044
rect 20962 23035 21020 23041
rect 20962 23032 20974 23035
rect 18656 23004 20974 23032
rect 18656 22992 18662 23004
rect 20962 23001 20974 23004
rect 21008 23001 21020 23035
rect 20962 22995 21020 23001
rect 23658 22992 23664 23044
rect 23716 22992 23722 23044
rect 25222 22992 25228 23044
rect 25280 23032 25286 23044
rect 25700 23032 25728 23060
rect 26344 23032 26372 23063
rect 25280 23004 25728 23032
rect 26160 23004 26372 23032
rect 25280 22992 25286 23004
rect 26160 22976 26188 23004
rect 13078 22924 13084 22976
rect 13136 22964 13142 22976
rect 14645 22967 14703 22973
rect 14645 22964 14657 22967
rect 13136 22936 14657 22964
rect 13136 22924 13142 22936
rect 14645 22933 14657 22936
rect 14691 22933 14703 22967
rect 14645 22927 14703 22933
rect 16666 22924 16672 22976
rect 16724 22964 16730 22976
rect 16945 22967 17003 22973
rect 16945 22964 16957 22967
rect 16724 22936 16957 22964
rect 16724 22924 16730 22936
rect 16945 22933 16957 22936
rect 16991 22964 17003 22967
rect 17126 22964 17132 22976
rect 16991 22936 17132 22964
rect 16991 22933 17003 22936
rect 16945 22927 17003 22933
rect 17126 22924 17132 22936
rect 17184 22964 17190 22976
rect 17862 22964 17868 22976
rect 17184 22936 17868 22964
rect 17184 22924 17190 22936
rect 17862 22924 17868 22936
rect 17920 22924 17926 22976
rect 17954 22924 17960 22976
rect 18012 22964 18018 22976
rect 19702 22964 19708 22976
rect 18012 22936 19708 22964
rect 18012 22924 18018 22936
rect 19702 22924 19708 22936
rect 19760 22924 19766 22976
rect 19797 22967 19855 22973
rect 19797 22933 19809 22967
rect 19843 22964 19855 22967
rect 20806 22964 20812 22976
rect 19843 22936 20812 22964
rect 19843 22933 19855 22936
rect 19797 22927 19855 22933
rect 20806 22924 20812 22936
rect 20864 22924 20870 22976
rect 22738 22924 22744 22976
rect 22796 22964 22802 22976
rect 23017 22967 23075 22973
rect 23017 22964 23029 22967
rect 22796 22936 23029 22964
rect 22796 22924 22802 22936
rect 23017 22933 23029 22936
rect 23063 22964 23075 22967
rect 23753 22967 23811 22973
rect 23753 22964 23765 22967
rect 23063 22936 23765 22964
rect 23063 22933 23075 22936
rect 23017 22927 23075 22933
rect 23753 22933 23765 22936
rect 23799 22964 23811 22967
rect 23934 22964 23940 22976
rect 23799 22936 23940 22964
rect 23799 22933 23811 22936
rect 23753 22927 23811 22933
rect 23934 22924 23940 22936
rect 23992 22964 23998 22976
rect 24302 22964 24308 22976
rect 23992 22936 24308 22964
rect 23992 22924 23998 22936
rect 24302 22924 24308 22936
rect 24360 22924 24366 22976
rect 24486 22924 24492 22976
rect 24544 22964 24550 22976
rect 24673 22967 24731 22973
rect 24673 22964 24685 22967
rect 24544 22936 24685 22964
rect 24544 22924 24550 22936
rect 24673 22933 24685 22936
rect 24719 22933 24731 22967
rect 24673 22927 24731 22933
rect 26142 22924 26148 22976
rect 26200 22924 26206 22976
rect 26326 22924 26332 22976
rect 26384 22924 26390 22976
rect 26436 22964 26464 23140
rect 26697 23137 26709 23171
rect 26743 23168 26755 23171
rect 30374 23168 30380 23180
rect 26743 23140 30380 23168
rect 26743 23137 26755 23140
rect 26697 23131 26755 23137
rect 30374 23128 30380 23140
rect 30432 23128 30438 23180
rect 26786 23060 26792 23112
rect 26844 23100 26850 23112
rect 27157 23103 27215 23109
rect 27157 23100 27169 23103
rect 26844 23072 27169 23100
rect 26844 23060 26850 23072
rect 27157 23069 27169 23072
rect 27203 23069 27215 23103
rect 27157 23063 27215 23069
rect 27338 23060 27344 23112
rect 27396 23100 27402 23112
rect 28905 23103 28963 23109
rect 28905 23100 28917 23103
rect 27396 23072 28917 23100
rect 27396 23060 27402 23072
rect 28905 23069 28917 23072
rect 28951 23069 28963 23103
rect 28905 23063 28963 23069
rect 29181 23103 29239 23109
rect 29181 23069 29193 23103
rect 29227 23100 29239 23103
rect 29270 23100 29276 23112
rect 29227 23072 29276 23100
rect 29227 23069 29239 23072
rect 29181 23063 29239 23069
rect 29270 23060 29276 23072
rect 29328 23060 29334 23112
rect 29730 23060 29736 23112
rect 29788 23060 29794 23112
rect 29881 23103 29939 23109
rect 29881 23069 29893 23103
rect 29927 23100 29939 23103
rect 29927 23069 29960 23100
rect 29881 23063 29960 23069
rect 27430 22992 27436 23044
rect 27488 22992 27494 23044
rect 27982 22992 27988 23044
rect 28040 23032 28046 23044
rect 28077 23035 28135 23041
rect 28077 23032 28089 23035
rect 28040 23004 28089 23032
rect 28040 22992 28046 23004
rect 28077 23001 28089 23004
rect 28123 23001 28135 23035
rect 28077 22995 28135 23001
rect 28261 23035 28319 23041
rect 28261 23001 28273 23035
rect 28307 23032 28319 23035
rect 28350 23032 28356 23044
rect 28307 23004 28356 23032
rect 28307 23001 28319 23004
rect 28261 22995 28319 23001
rect 28350 22992 28356 23004
rect 28408 22992 28414 23044
rect 28718 22992 28724 23044
rect 28776 23032 28782 23044
rect 29932 23032 29960 23063
rect 30006 23060 30012 23112
rect 30064 23060 30070 23112
rect 30190 23060 30196 23112
rect 30248 23109 30254 23112
rect 30248 23100 30256 23109
rect 30248 23072 30293 23100
rect 30248 23063 30256 23072
rect 30248 23060 30254 23063
rect 30101 23035 30159 23041
rect 28776 23004 30052 23032
rect 28776 22992 28782 23004
rect 28000 22964 28028 22992
rect 30024 22976 30052 23004
rect 30101 23001 30113 23035
rect 30147 23001 30159 23035
rect 30484 23032 30512 23208
rect 30760 23168 30788 23276
rect 30834 23264 30840 23316
rect 30892 23264 30898 23316
rect 32766 23264 32772 23316
rect 32824 23304 32830 23316
rect 33870 23304 33876 23316
rect 32824 23276 33876 23304
rect 32824 23264 32830 23276
rect 33870 23264 33876 23276
rect 33928 23264 33934 23316
rect 34422 23264 34428 23316
rect 34480 23304 34486 23316
rect 35158 23304 35164 23316
rect 34480 23276 35164 23304
rect 34480 23264 34486 23276
rect 35158 23264 35164 23276
rect 35216 23264 35222 23316
rect 35529 23307 35587 23313
rect 35529 23273 35541 23307
rect 35575 23304 35587 23307
rect 35894 23304 35900 23316
rect 35575 23276 35900 23304
rect 35575 23273 35587 23276
rect 35529 23267 35587 23273
rect 35894 23264 35900 23276
rect 35952 23264 35958 23316
rect 36004 23276 37127 23304
rect 31570 23196 31576 23248
rect 31628 23236 31634 23248
rect 36004 23236 36032 23276
rect 31628 23208 33713 23236
rect 31628 23196 31634 23208
rect 33685 23168 33713 23208
rect 34440 23208 36032 23236
rect 37099 23236 37127 23276
rect 37458 23264 37464 23316
rect 37516 23304 37522 23316
rect 37553 23307 37611 23313
rect 37553 23304 37565 23307
rect 37516 23276 37565 23304
rect 37516 23264 37522 23276
rect 37553 23273 37565 23276
rect 37599 23273 37611 23307
rect 37553 23267 37611 23273
rect 39298 23236 39304 23248
rect 37099 23208 39304 23236
rect 30760 23140 33640 23168
rect 33685 23140 34376 23168
rect 30837 23103 30895 23109
rect 30837 23069 30849 23103
rect 30883 23100 30895 23103
rect 31018 23100 31024 23112
rect 30883 23072 31024 23100
rect 30883 23069 30895 23072
rect 30837 23063 30895 23069
rect 31018 23060 31024 23072
rect 31076 23060 31082 23112
rect 31113 23103 31171 23109
rect 31113 23069 31125 23103
rect 31159 23100 31171 23103
rect 31570 23100 31576 23112
rect 31159 23072 31576 23100
rect 31159 23069 31171 23072
rect 31113 23063 31171 23069
rect 31570 23060 31576 23072
rect 31628 23060 31634 23112
rect 31846 23060 31852 23112
rect 31904 23060 31910 23112
rect 32125 23103 32183 23109
rect 32125 23069 32137 23103
rect 32171 23100 32183 23103
rect 32214 23100 32220 23112
rect 32171 23072 32220 23100
rect 32171 23069 32183 23072
rect 32125 23063 32183 23069
rect 32214 23060 32220 23072
rect 32272 23060 32278 23112
rect 32309 23103 32367 23109
rect 32309 23069 32321 23103
rect 32355 23100 32367 23103
rect 32766 23100 32772 23112
rect 32355 23072 32772 23100
rect 32355 23069 32367 23072
rect 32309 23063 32367 23069
rect 32766 23060 32772 23072
rect 32824 23060 32830 23112
rect 32907 23103 32965 23109
rect 32907 23069 32919 23103
rect 32953 23069 32965 23103
rect 32907 23063 32965 23069
rect 33275 23103 33333 23109
rect 33275 23069 33287 23103
rect 33321 23100 33333 23103
rect 33410 23100 33416 23112
rect 33321 23072 33416 23100
rect 33321 23069 33333 23072
rect 33275 23063 33333 23069
rect 31864 23032 31892 23060
rect 30484 23004 31892 23032
rect 30101 22995 30159 23001
rect 26436 22936 28028 22964
rect 28626 22924 28632 22976
rect 28684 22964 28690 22976
rect 29089 22967 29147 22973
rect 29089 22964 29101 22967
rect 28684 22936 29101 22964
rect 28684 22924 28690 22936
rect 29089 22933 29101 22936
rect 29135 22933 29147 22967
rect 29089 22927 29147 22933
rect 30006 22924 30012 22976
rect 30064 22924 30070 22976
rect 30116 22964 30144 22995
rect 32398 22992 32404 23044
rect 32456 23032 32462 23044
rect 32932 23032 32960 23063
rect 33410 23060 33416 23072
rect 33468 23060 33474 23112
rect 32456 23004 32960 23032
rect 33045 23035 33103 23041
rect 32456 22992 32462 23004
rect 33045 23001 33057 23035
rect 33091 23001 33103 23035
rect 33045 22995 33103 23001
rect 30282 22964 30288 22976
rect 30116 22936 30288 22964
rect 30282 22924 30288 22936
rect 30340 22924 30346 22976
rect 30374 22924 30380 22976
rect 30432 22924 30438 22976
rect 30558 22924 30564 22976
rect 30616 22964 30622 22976
rect 31021 22967 31079 22973
rect 31021 22964 31033 22967
rect 30616 22936 31033 22964
rect 30616 22924 30622 22936
rect 31021 22933 31033 22936
rect 31067 22933 31079 22967
rect 31021 22927 31079 22933
rect 32950 22924 32956 22976
rect 33008 22964 33014 22976
rect 33060 22964 33088 22995
rect 33134 22992 33140 23044
rect 33192 22992 33198 23044
rect 33612 23032 33640 23140
rect 34057 23103 34115 23109
rect 34057 23069 34069 23103
rect 34103 23069 34115 23103
rect 34057 23063 34115 23069
rect 34072 23032 34100 23063
rect 34238 23060 34244 23112
rect 34296 23060 34302 23112
rect 34348 23109 34376 23140
rect 34333 23103 34391 23109
rect 34333 23069 34345 23103
rect 34379 23069 34391 23103
rect 34333 23063 34391 23069
rect 34440 23044 34468 23208
rect 39298 23196 39304 23208
rect 39356 23196 39362 23248
rect 35526 23168 35532 23180
rect 34900 23140 35532 23168
rect 34790 23060 34796 23112
rect 34848 23100 34854 23112
rect 34900 23109 34928 23140
rect 35526 23128 35532 23140
rect 35584 23128 35590 23180
rect 34885 23103 34943 23109
rect 34885 23100 34897 23103
rect 34848 23072 34897 23100
rect 34848 23060 34854 23072
rect 34885 23069 34897 23072
rect 34931 23069 34943 23103
rect 34885 23063 34943 23069
rect 34978 23103 35036 23109
rect 34978 23069 34990 23103
rect 35024 23069 35036 23103
rect 34978 23063 35036 23069
rect 34422 23032 34428 23044
rect 33612 23004 34008 23032
rect 34072 23004 34428 23032
rect 33008 22936 33088 22964
rect 33008 22924 33014 22936
rect 33226 22924 33232 22976
rect 33284 22964 33290 22976
rect 33413 22967 33471 22973
rect 33413 22964 33425 22967
rect 33284 22936 33425 22964
rect 33284 22924 33290 22936
rect 33413 22933 33425 22936
rect 33459 22933 33471 22967
rect 33413 22927 33471 22933
rect 33502 22924 33508 22976
rect 33560 22964 33566 22976
rect 33873 22967 33931 22973
rect 33873 22964 33885 22967
rect 33560 22936 33885 22964
rect 33560 22924 33566 22936
rect 33873 22933 33885 22936
rect 33919 22933 33931 22967
rect 33980 22964 34008 23004
rect 34422 22992 34428 23004
rect 34480 22992 34486 23044
rect 34606 22992 34612 23044
rect 34664 23032 34670 23044
rect 34993 23032 35021 23063
rect 35158 23060 35164 23112
rect 35216 23060 35222 23112
rect 35342 23060 35348 23112
rect 35400 23109 35406 23112
rect 35400 23100 35408 23109
rect 35802 23100 35808 23112
rect 35400 23072 35808 23100
rect 35400 23063 35408 23072
rect 35400 23060 35406 23063
rect 35802 23060 35808 23072
rect 35860 23060 35866 23112
rect 36173 23103 36231 23109
rect 36173 23069 36185 23103
rect 36219 23100 36231 23103
rect 36906 23100 36912 23112
rect 36219 23072 36912 23100
rect 36219 23069 36231 23072
rect 36173 23063 36231 23069
rect 36906 23060 36912 23072
rect 36964 23060 36970 23112
rect 36998 23060 37004 23112
rect 37056 23100 37062 23112
rect 38105 23103 38163 23109
rect 38105 23100 38117 23103
rect 37056 23072 38117 23100
rect 37056 23060 37062 23072
rect 38105 23069 38117 23072
rect 38151 23069 38163 23103
rect 38105 23063 38163 23069
rect 38286 23060 38292 23112
rect 38344 23060 38350 23112
rect 34664 23004 35021 23032
rect 35253 23035 35311 23041
rect 34664 22992 34670 23004
rect 35253 23001 35265 23035
rect 35299 23032 35311 23035
rect 35710 23032 35716 23044
rect 35299 23004 35716 23032
rect 35299 23001 35311 23004
rect 35253 22995 35311 23001
rect 35710 22992 35716 23004
rect 35768 22992 35774 23044
rect 36440 23035 36498 23041
rect 36440 23001 36452 23035
rect 36486 23032 36498 23035
rect 36722 23032 36728 23044
rect 36486 23004 36728 23032
rect 36486 23001 36498 23004
rect 36440 22995 36498 23001
rect 36722 22992 36728 23004
rect 36780 22992 36786 23044
rect 38197 22967 38255 22973
rect 38197 22964 38209 22967
rect 33980 22936 38209 22964
rect 33873 22927 33931 22933
rect 38197 22933 38209 22936
rect 38243 22933 38255 22967
rect 38197 22927 38255 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 14185 22763 14243 22769
rect 14185 22729 14197 22763
rect 14231 22760 14243 22763
rect 15102 22760 15108 22772
rect 14231 22732 15108 22760
rect 14231 22729 14243 22732
rect 14185 22723 14243 22729
rect 15102 22720 15108 22732
rect 15160 22760 15166 22772
rect 15160 22732 17540 22760
rect 15160 22720 15166 22732
rect 13078 22701 13084 22704
rect 13072 22692 13084 22701
rect 13039 22664 13084 22692
rect 13072 22655 13084 22664
rect 13078 22652 13084 22655
rect 13136 22652 13142 22704
rect 14274 22652 14280 22704
rect 14332 22692 14338 22704
rect 14737 22695 14795 22701
rect 14737 22692 14749 22695
rect 14332 22664 14749 22692
rect 14332 22652 14338 22664
rect 14737 22661 14749 22664
rect 14783 22661 14795 22695
rect 14737 22655 14795 22661
rect 16758 22652 16764 22704
rect 16816 22692 16822 22704
rect 17405 22695 17463 22701
rect 17405 22692 17417 22695
rect 16816 22664 17417 22692
rect 16816 22652 16822 22664
rect 17405 22661 17417 22664
rect 17451 22661 17463 22695
rect 17512 22692 17540 22732
rect 18598 22720 18604 22772
rect 18656 22720 18662 22772
rect 19334 22760 19340 22772
rect 18708 22732 19340 22760
rect 18708 22692 18736 22732
rect 19334 22720 19340 22732
rect 19392 22720 19398 22772
rect 20438 22720 20444 22772
rect 20496 22720 20502 22772
rect 21361 22763 21419 22769
rect 21361 22729 21373 22763
rect 21407 22760 21419 22763
rect 22554 22760 22560 22772
rect 21407 22732 22560 22760
rect 21407 22729 21419 22732
rect 21361 22723 21419 22729
rect 22554 22720 22560 22732
rect 22612 22720 22618 22772
rect 24486 22760 24492 22772
rect 22747 22732 24492 22760
rect 17512 22664 18736 22692
rect 17405 22655 17463 22661
rect 20346 22652 20352 22704
rect 20404 22692 20410 22704
rect 22747 22692 22775 22732
rect 24486 22720 24492 22732
rect 24544 22720 24550 22772
rect 27062 22760 27068 22772
rect 25056 22732 27068 22760
rect 20404 22664 21496 22692
rect 20404 22652 20410 22664
rect 12805 22627 12863 22633
rect 12805 22593 12817 22627
rect 12851 22624 12863 22627
rect 12894 22624 12900 22636
rect 12851 22596 12900 22624
rect 12851 22593 12863 22596
rect 12805 22587 12863 22593
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 15286 22584 15292 22636
rect 15344 22624 15350 22636
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 15344 22596 16129 22624
rect 15344 22584 15350 22596
rect 16117 22593 16129 22596
rect 16163 22624 16175 22627
rect 16206 22624 16212 22636
rect 16163 22596 16212 22624
rect 16163 22593 16175 22596
rect 16117 22587 16175 22593
rect 16206 22584 16212 22596
rect 16264 22584 16270 22636
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22624 16359 22627
rect 16482 22624 16488 22636
rect 16347 22596 16488 22624
rect 16347 22593 16359 22596
rect 16301 22587 16359 22593
rect 16482 22584 16488 22596
rect 16540 22584 16546 22636
rect 16574 22584 16580 22636
rect 16632 22624 16638 22636
rect 17129 22627 17187 22633
rect 17129 22624 17141 22627
rect 16632 22596 17141 22624
rect 16632 22584 16638 22596
rect 17129 22593 17141 22596
rect 17175 22593 17187 22627
rect 17129 22587 17187 22593
rect 17222 22627 17280 22633
rect 17222 22593 17234 22627
rect 17268 22593 17280 22627
rect 17222 22587 17280 22593
rect 15562 22516 15568 22568
rect 15620 22516 15626 22568
rect 15838 22516 15844 22568
rect 15896 22556 15902 22568
rect 17236 22556 17264 22587
rect 17494 22584 17500 22636
rect 17552 22584 17558 22636
rect 17594 22627 17652 22633
rect 17594 22593 17606 22627
rect 17640 22593 17652 22627
rect 17594 22587 17652 22593
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22624 18475 22627
rect 18690 22624 18696 22636
rect 18463 22596 18696 22624
rect 18463 22593 18475 22596
rect 18417 22587 18475 22593
rect 15896 22528 17264 22556
rect 15896 22516 15902 22528
rect 17310 22516 17316 22568
rect 17368 22556 17374 22568
rect 17604 22556 17632 22587
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 19061 22627 19119 22633
rect 19061 22593 19073 22627
rect 19107 22624 19119 22627
rect 19150 22624 19156 22636
rect 19107 22596 19156 22624
rect 19107 22593 19119 22596
rect 19061 22587 19119 22593
rect 19150 22584 19156 22596
rect 19208 22624 19214 22636
rect 20714 22624 20720 22636
rect 19208 22596 20720 22624
rect 19208 22584 19214 22596
rect 20714 22584 20720 22596
rect 20772 22584 20778 22636
rect 21468 22633 21496 22664
rect 22204 22664 22775 22692
rect 22204 22636 22232 22664
rect 24210 22652 24216 22704
rect 24268 22692 24274 22704
rect 25056 22692 25084 22732
rect 27062 22720 27068 22732
rect 27120 22720 27126 22772
rect 27338 22720 27344 22772
rect 27396 22760 27402 22772
rect 27522 22760 27528 22772
rect 27396 22732 27528 22760
rect 27396 22720 27402 22732
rect 27522 22720 27528 22732
rect 27580 22720 27586 22772
rect 28626 22720 28632 22772
rect 28684 22720 28690 22772
rect 29086 22720 29092 22772
rect 29144 22760 29150 22772
rect 30466 22760 30472 22772
rect 29144 22732 30472 22760
rect 29144 22720 29150 22732
rect 30466 22720 30472 22732
rect 30524 22720 30530 22772
rect 32769 22763 32827 22769
rect 32769 22729 32781 22763
rect 32815 22729 32827 22763
rect 32769 22723 32827 22729
rect 33689 22763 33747 22769
rect 33689 22729 33701 22763
rect 33735 22760 33747 22763
rect 36354 22760 36360 22772
rect 33735 22732 36360 22760
rect 33735 22729 33747 22732
rect 33689 22723 33747 22729
rect 30374 22692 30380 22704
rect 24268 22664 25084 22692
rect 25516 22664 30380 22692
rect 24268 22652 24274 22664
rect 21269 22627 21327 22633
rect 21269 22593 21281 22627
rect 21315 22593 21327 22627
rect 21269 22587 21327 22593
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22593 21511 22627
rect 21453 22587 21511 22593
rect 17368 22528 17632 22556
rect 17368 22516 17374 22528
rect 17862 22516 17868 22568
rect 17920 22556 17926 22568
rect 18233 22559 18291 22565
rect 18233 22556 18245 22559
rect 17920 22528 18245 22556
rect 17920 22516 17926 22528
rect 18233 22525 18245 22528
rect 18279 22525 18291 22559
rect 18233 22519 18291 22525
rect 18782 22516 18788 22568
rect 18840 22556 18846 22568
rect 19337 22559 19395 22565
rect 19337 22556 19349 22559
rect 18840 22528 19349 22556
rect 18840 22516 18846 22528
rect 19337 22525 19349 22528
rect 19383 22525 19395 22559
rect 19337 22519 19395 22525
rect 17402 22488 17408 22500
rect 16040 22460 17408 22488
rect 13446 22380 13452 22432
rect 13504 22420 13510 22432
rect 16040 22420 16068 22460
rect 17402 22448 17408 22460
rect 17460 22488 17466 22500
rect 17954 22488 17960 22500
rect 17460 22460 17960 22488
rect 17460 22448 17466 22460
rect 17954 22448 17960 22460
rect 18012 22448 18018 22500
rect 21284 22488 21312 22587
rect 21468 22556 21496 22587
rect 22186 22584 22192 22636
rect 22244 22584 22250 22636
rect 22278 22584 22284 22636
rect 22336 22624 22342 22636
rect 22557 22627 22615 22633
rect 22557 22624 22569 22627
rect 22336 22596 22569 22624
rect 22336 22584 22342 22596
rect 22557 22593 22569 22596
rect 22603 22593 22615 22627
rect 22557 22587 22615 22593
rect 22738 22584 22744 22636
rect 22796 22624 22802 22636
rect 23661 22627 23719 22633
rect 23661 22624 23673 22627
rect 22796 22596 23673 22624
rect 22796 22584 22802 22596
rect 23661 22593 23673 22596
rect 23707 22624 23719 22627
rect 24026 22624 24032 22636
rect 23707 22596 24032 22624
rect 23707 22593 23719 22596
rect 23661 22587 23719 22593
rect 24026 22584 24032 22596
rect 24084 22584 24090 22636
rect 25133 22627 25191 22633
rect 25133 22593 25145 22627
rect 25179 22624 25191 22627
rect 25222 22624 25228 22636
rect 25179 22596 25228 22624
rect 25179 22593 25191 22596
rect 25133 22587 25191 22593
rect 25222 22584 25228 22596
rect 25280 22584 25286 22636
rect 25516 22633 25544 22664
rect 30374 22652 30380 22664
rect 30432 22652 30438 22704
rect 31294 22692 31300 22704
rect 31220 22664 31300 22692
rect 25501 22627 25559 22633
rect 25501 22593 25513 22627
rect 25547 22593 25559 22627
rect 25501 22587 25559 22593
rect 25958 22584 25964 22636
rect 26016 22584 26022 22636
rect 26050 22584 26056 22636
rect 26108 22624 26114 22636
rect 26145 22627 26203 22633
rect 26145 22624 26157 22627
rect 26108 22596 26157 22624
rect 26108 22584 26114 22596
rect 26145 22593 26157 22596
rect 26191 22593 26203 22627
rect 26145 22587 26203 22593
rect 26237 22627 26295 22633
rect 26237 22593 26249 22627
rect 26283 22593 26295 22627
rect 26237 22587 26295 22593
rect 26381 22627 26439 22633
rect 26381 22593 26393 22627
rect 26427 22624 26439 22627
rect 26427 22593 26464 22624
rect 26381 22587 26464 22593
rect 21468 22528 22416 22556
rect 21284 22460 22232 22488
rect 13504 22392 16068 22420
rect 16117 22423 16175 22429
rect 13504 22380 13510 22392
rect 16117 22389 16129 22423
rect 16163 22420 16175 22423
rect 16666 22420 16672 22432
rect 16163 22392 16672 22420
rect 16163 22389 16175 22392
rect 16117 22383 16175 22389
rect 16666 22380 16672 22392
rect 16724 22380 16730 22432
rect 17773 22423 17831 22429
rect 17773 22389 17785 22423
rect 17819 22420 17831 22423
rect 19518 22420 19524 22432
rect 17819 22392 19524 22420
rect 17819 22389 17831 22392
rect 17773 22383 17831 22389
rect 19518 22380 19524 22392
rect 19576 22380 19582 22432
rect 22204 22420 22232 22460
rect 22278 22448 22284 22500
rect 22336 22448 22342 22500
rect 22388 22488 22416 22528
rect 22830 22516 22836 22568
rect 22888 22556 22894 22568
rect 23290 22556 23296 22568
rect 22888 22528 23296 22556
rect 22888 22516 22894 22528
rect 23290 22516 23296 22528
rect 23348 22516 23354 22568
rect 24949 22559 25007 22565
rect 24949 22525 24961 22559
rect 24995 22556 25007 22559
rect 25682 22556 25688 22568
rect 24995 22528 25688 22556
rect 24995 22525 25007 22528
rect 24949 22519 25007 22525
rect 25682 22516 25688 22528
rect 25740 22516 25746 22568
rect 26252 22556 26280 22587
rect 26436 22556 26464 22587
rect 26602 22584 26608 22636
rect 26660 22624 26666 22636
rect 27154 22624 27160 22636
rect 26660 22596 27160 22624
rect 26660 22584 26666 22596
rect 27154 22584 27160 22596
rect 27212 22624 27218 22636
rect 27525 22627 27583 22633
rect 27525 22624 27537 22627
rect 27212 22596 27537 22624
rect 27212 22584 27218 22596
rect 27525 22593 27537 22596
rect 27571 22593 27583 22627
rect 27525 22587 27583 22593
rect 27614 22584 27620 22636
rect 27672 22624 27678 22636
rect 27801 22627 27859 22633
rect 27801 22624 27813 22627
rect 27672 22596 27813 22624
rect 27672 22584 27678 22596
rect 27801 22593 27813 22596
rect 27847 22624 27859 22627
rect 28258 22624 28264 22636
rect 27847 22596 28264 22624
rect 27847 22593 27859 22596
rect 27801 22587 27859 22593
rect 28258 22584 28264 22596
rect 28316 22584 28322 22636
rect 28445 22627 28503 22633
rect 28445 22593 28457 22627
rect 28491 22624 28503 22627
rect 28718 22624 28724 22636
rect 28491 22596 28724 22624
rect 28491 22593 28503 22596
rect 28445 22587 28503 22593
rect 26878 22556 26884 22568
rect 26252 22528 26372 22556
rect 26436 22528 26884 22556
rect 24670 22488 24676 22500
rect 22388 22460 24676 22488
rect 24670 22448 24676 22460
rect 24728 22448 24734 22500
rect 25406 22448 25412 22500
rect 25464 22448 25470 22500
rect 25590 22448 25596 22500
rect 25648 22488 25654 22500
rect 26050 22488 26056 22500
rect 25648 22460 26056 22488
rect 25648 22448 25654 22460
rect 26050 22448 26056 22460
rect 26108 22448 26114 22500
rect 26344 22488 26372 22528
rect 26878 22516 26884 22528
rect 26936 22516 26942 22568
rect 27062 22516 27068 22568
rect 27120 22556 27126 22568
rect 28460 22556 28488 22587
rect 28718 22584 28724 22596
rect 28776 22584 28782 22636
rect 29089 22627 29147 22633
rect 29089 22624 29101 22627
rect 29012 22596 29101 22624
rect 27120 22528 28488 22556
rect 27120 22516 27126 22528
rect 26344 22460 28396 22488
rect 23290 22420 23296 22432
rect 22204 22392 23296 22420
rect 23290 22380 23296 22392
rect 23348 22380 23354 22432
rect 23658 22380 23664 22432
rect 23716 22420 23722 22432
rect 23753 22423 23811 22429
rect 23753 22420 23765 22423
rect 23716 22392 23765 22420
rect 23716 22380 23722 22392
rect 23753 22389 23765 22392
rect 23799 22389 23811 22423
rect 23753 22383 23811 22389
rect 24854 22380 24860 22432
rect 24912 22420 24918 22432
rect 26513 22423 26571 22429
rect 26513 22420 26525 22423
rect 24912 22392 26525 22420
rect 24912 22380 24918 22392
rect 26513 22389 26525 22392
rect 26559 22389 26571 22423
rect 26513 22383 26571 22389
rect 27062 22380 27068 22432
rect 27120 22420 27126 22432
rect 27709 22423 27767 22429
rect 27709 22420 27721 22423
rect 27120 22392 27721 22420
rect 27120 22380 27126 22392
rect 27709 22389 27721 22392
rect 27755 22389 27767 22423
rect 28368 22420 28396 22460
rect 28442 22448 28448 22500
rect 28500 22488 28506 22500
rect 29012 22488 29040 22596
rect 29089 22593 29101 22596
rect 29135 22593 29147 22627
rect 29089 22587 29147 22593
rect 29365 22627 29423 22633
rect 29365 22593 29377 22627
rect 29411 22624 29423 22627
rect 29454 22624 29460 22636
rect 29411 22596 29460 22624
rect 29411 22593 29423 22596
rect 29365 22587 29423 22593
rect 29454 22584 29460 22596
rect 29512 22584 29518 22636
rect 29638 22584 29644 22636
rect 29696 22624 29702 22636
rect 30285 22627 30343 22633
rect 30285 22624 30297 22627
rect 29696 22596 30297 22624
rect 29696 22584 29702 22596
rect 30285 22593 30297 22596
rect 30331 22593 30343 22627
rect 30285 22587 30343 22593
rect 30834 22584 30840 22636
rect 30892 22584 30898 22636
rect 31220 22633 31248 22664
rect 31294 22652 31300 22664
rect 31352 22692 31358 22704
rect 31570 22692 31576 22704
rect 31352 22664 31576 22692
rect 31352 22652 31358 22664
rect 31570 22652 31576 22664
rect 31628 22652 31634 22704
rect 32674 22692 32680 22704
rect 31680 22664 32680 22692
rect 31680 22633 31708 22664
rect 32674 22652 32680 22664
rect 32732 22652 32738 22704
rect 32784 22692 32812 22723
rect 36354 22720 36360 22732
rect 36412 22720 36418 22772
rect 32784 22664 33916 22692
rect 33888 22636 33916 22664
rect 34146 22652 34152 22704
rect 34204 22692 34210 22704
rect 34333 22695 34391 22701
rect 34333 22692 34345 22695
rect 34204 22664 34345 22692
rect 34204 22652 34210 22664
rect 34333 22661 34345 22664
rect 34379 22661 34391 22695
rect 34333 22655 34391 22661
rect 35158 22652 35164 22704
rect 35216 22692 35222 22704
rect 35526 22692 35532 22704
rect 35216 22664 35532 22692
rect 35216 22652 35222 22664
rect 35526 22652 35532 22664
rect 35584 22692 35590 22704
rect 37737 22695 37795 22701
rect 37737 22692 37749 22695
rect 35584 22664 37749 22692
rect 35584 22652 35590 22664
rect 37737 22661 37749 22664
rect 37783 22661 37795 22695
rect 37737 22655 37795 22661
rect 31205 22627 31263 22633
rect 31205 22593 31217 22627
rect 31251 22593 31263 22627
rect 31205 22587 31263 22593
rect 31665 22627 31723 22633
rect 31665 22593 31677 22627
rect 31711 22593 31723 22627
rect 32766 22624 32772 22636
rect 32727 22596 32772 22624
rect 31665 22587 31723 22593
rect 32766 22584 32772 22596
rect 32824 22584 32830 22636
rect 33134 22584 33140 22636
rect 33192 22624 33198 22636
rect 33870 22624 33876 22636
rect 33192 22596 33640 22624
rect 33832 22596 33876 22624
rect 33192 22584 33198 22596
rect 33612 22568 33640 22596
rect 33870 22584 33876 22596
rect 33928 22584 33934 22636
rect 33962 22584 33968 22636
rect 34020 22624 34026 22636
rect 34241 22627 34299 22633
rect 34020 22596 34065 22624
rect 34020 22584 34026 22596
rect 34241 22593 34253 22627
rect 34287 22593 34299 22627
rect 34241 22587 34299 22593
rect 30926 22556 30932 22568
rect 28500 22460 29040 22488
rect 29196 22528 30932 22556
rect 28500 22448 28506 22460
rect 29196 22420 29224 22528
rect 30926 22516 30932 22528
rect 30984 22516 30990 22568
rect 31294 22516 31300 22568
rect 31352 22516 31358 22568
rect 31386 22516 31392 22568
rect 31444 22556 31450 22568
rect 33229 22559 33287 22565
rect 33229 22556 33241 22559
rect 31444 22528 33241 22556
rect 31444 22516 31450 22528
rect 33229 22525 33241 22528
rect 33275 22525 33287 22559
rect 33229 22519 33287 22525
rect 33594 22516 33600 22568
rect 33652 22556 33658 22568
rect 34256 22556 34284 22587
rect 35342 22584 35348 22636
rect 35400 22584 35406 22636
rect 35437 22627 35495 22633
rect 35437 22593 35449 22627
rect 35483 22593 35495 22627
rect 35437 22587 35495 22593
rect 33652 22528 34284 22556
rect 33652 22516 33658 22528
rect 34422 22516 34428 22568
rect 34480 22556 34486 22568
rect 35452 22556 35480 22587
rect 35710 22584 35716 22636
rect 35768 22584 35774 22636
rect 36357 22627 36415 22633
rect 36357 22593 36369 22627
rect 36403 22624 36415 22627
rect 36998 22624 37004 22636
rect 36403 22596 37004 22624
rect 36403 22593 36415 22596
rect 36357 22587 36415 22593
rect 36998 22584 37004 22596
rect 37056 22584 37062 22636
rect 37458 22584 37464 22636
rect 37516 22584 37522 22636
rect 34480 22528 35480 22556
rect 34480 22516 34486 22528
rect 35618 22516 35624 22568
rect 35676 22556 35682 22568
rect 35894 22556 35900 22568
rect 35676 22528 35900 22556
rect 35676 22516 35682 22528
rect 35894 22516 35900 22528
rect 35952 22556 35958 22568
rect 36265 22559 36323 22565
rect 36265 22556 36277 22559
rect 35952 22528 36277 22556
rect 35952 22516 35958 22528
rect 36265 22525 36277 22528
rect 36311 22525 36323 22559
rect 36265 22519 36323 22525
rect 36722 22516 36728 22568
rect 36780 22516 36786 22568
rect 29365 22491 29423 22497
rect 29365 22457 29377 22491
rect 29411 22488 29423 22491
rect 29546 22488 29552 22500
rect 29411 22460 29552 22488
rect 29411 22457 29423 22460
rect 29365 22451 29423 22457
rect 29546 22448 29552 22460
rect 29604 22448 29610 22500
rect 33137 22491 33195 22497
rect 31726 22460 32996 22488
rect 28368 22392 29224 22420
rect 27709 22383 27767 22389
rect 29270 22380 29276 22432
rect 29328 22420 29334 22432
rect 31726 22420 31754 22460
rect 29328 22392 31754 22420
rect 29328 22380 29334 22392
rect 32214 22380 32220 22432
rect 32272 22420 32278 22432
rect 32585 22423 32643 22429
rect 32585 22420 32597 22423
rect 32272 22392 32597 22420
rect 32272 22380 32278 22392
rect 32585 22389 32597 22392
rect 32631 22389 32643 22423
rect 32968 22420 32996 22460
rect 33137 22457 33149 22491
rect 33183 22488 33195 22491
rect 34514 22488 34520 22500
rect 33183 22460 34520 22488
rect 33183 22457 33195 22460
rect 33137 22451 33195 22457
rect 34514 22448 34520 22460
rect 34572 22448 34578 22500
rect 35161 22491 35219 22497
rect 35161 22457 35173 22491
rect 35207 22488 35219 22491
rect 37918 22488 37924 22500
rect 35207 22460 37924 22488
rect 35207 22457 35219 22460
rect 35161 22451 35219 22457
rect 37918 22448 37924 22460
rect 37976 22448 37982 22500
rect 33318 22420 33324 22432
rect 32968 22392 33324 22420
rect 32585 22383 32643 22389
rect 33318 22380 33324 22392
rect 33376 22380 33382 22432
rect 35621 22423 35679 22429
rect 35621 22389 35633 22423
rect 35667 22420 35679 22423
rect 36170 22420 36176 22432
rect 35667 22392 36176 22420
rect 35667 22389 35679 22392
rect 35621 22383 35679 22389
rect 36170 22380 36176 22392
rect 36228 22420 36234 22432
rect 36538 22420 36544 22432
rect 36228 22392 36544 22420
rect 36228 22380 36234 22392
rect 36538 22380 36544 22392
rect 36596 22380 36602 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 17310 22176 17316 22228
rect 17368 22176 17374 22228
rect 18782 22176 18788 22228
rect 18840 22176 18846 22228
rect 19426 22176 19432 22228
rect 19484 22176 19490 22228
rect 22462 22216 22468 22228
rect 19536 22188 22468 22216
rect 17862 22108 17868 22160
rect 17920 22148 17926 22160
rect 19536 22148 19564 22188
rect 22462 22176 22468 22188
rect 22520 22176 22526 22228
rect 22554 22176 22560 22228
rect 22612 22216 22618 22228
rect 22612 22188 23796 22216
rect 22612 22176 22618 22188
rect 17920 22120 19564 22148
rect 17920 22108 17926 22120
rect 19794 22108 19800 22160
rect 19852 22108 19858 22160
rect 21361 22151 21419 22157
rect 21361 22117 21373 22151
rect 21407 22148 21419 22151
rect 21407 22120 21956 22148
rect 21407 22117 21419 22120
rect 21361 22111 21419 22117
rect 12894 22040 12900 22092
rect 12952 22080 12958 22092
rect 13541 22083 13599 22089
rect 13541 22080 13553 22083
rect 12952 22052 13553 22080
rect 12952 22040 12958 22052
rect 13541 22049 13553 22052
rect 13587 22049 13599 22083
rect 13541 22043 13599 22049
rect 14734 22040 14740 22092
rect 14792 22040 14798 22092
rect 15286 22040 15292 22092
rect 15344 22040 15350 22092
rect 15378 22040 15384 22092
rect 15436 22080 15442 22092
rect 16025 22083 16083 22089
rect 16025 22080 16037 22083
rect 15436 22052 16037 22080
rect 15436 22040 15442 22052
rect 16025 22049 16037 22052
rect 16071 22049 16083 22083
rect 16025 22043 16083 22049
rect 17218 22040 17224 22092
rect 17276 22080 17282 22092
rect 18417 22083 18475 22089
rect 18417 22080 18429 22083
rect 17276 22052 18429 22080
rect 17276 22040 17282 22052
rect 18417 22049 18429 22052
rect 18463 22049 18475 22083
rect 18417 22043 18475 22049
rect 19334 22040 19340 22092
rect 19392 22080 19398 22092
rect 19392 22052 21680 22080
rect 19392 22040 19398 22052
rect 10965 22015 11023 22021
rect 10965 21981 10977 22015
rect 11011 22012 11023 22015
rect 11054 22012 11060 22024
rect 11011 21984 11060 22012
rect 11011 21981 11023 21984
rect 10965 21975 11023 21981
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 12805 22015 12863 22021
rect 12805 21981 12817 22015
rect 12851 22012 12863 22015
rect 14274 22012 14280 22024
rect 12851 21984 14280 22012
rect 12851 21981 12863 21984
rect 12805 21975 12863 21981
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 14826 21972 14832 22024
rect 14884 21972 14890 22024
rect 15194 21972 15200 22024
rect 15252 22012 15258 22024
rect 15562 22012 15568 22024
rect 15252 21984 15568 22012
rect 15252 21972 15258 21984
rect 15562 21972 15568 21984
rect 15620 22012 15626 22024
rect 15749 22015 15807 22021
rect 15749 22012 15761 22015
rect 15620 21984 15761 22012
rect 15620 21972 15626 21984
rect 15749 21981 15761 21984
rect 15795 21981 15807 22015
rect 15749 21975 15807 21981
rect 18230 21972 18236 22024
rect 18288 22012 18294 22024
rect 18509 22015 18567 22021
rect 18509 22012 18521 22015
rect 18288 21984 18521 22012
rect 18288 21972 18294 21984
rect 18509 21981 18521 21984
rect 18555 21981 18567 22015
rect 18509 21975 18567 21981
rect 19518 21972 19524 22024
rect 19576 22012 19582 22024
rect 19613 22015 19671 22021
rect 19613 22012 19625 22015
rect 19576 21984 19625 22012
rect 19576 21972 19582 21984
rect 19613 21981 19625 21984
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 19886 21972 19892 22024
rect 19944 21972 19950 22024
rect 20162 21972 20168 22024
rect 20220 22012 20226 22024
rect 21652 22021 21680 22052
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 20220 21984 20361 22012
rect 20220 21972 20226 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 21269 22015 21327 22021
rect 21269 21981 21281 22015
rect 21315 21981 21327 22015
rect 21269 21975 21327 21981
rect 21637 22015 21695 22021
rect 21637 21981 21649 22015
rect 21683 21981 21695 22015
rect 21928 22012 21956 22120
rect 22278 22108 22284 22160
rect 22336 22148 22342 22160
rect 23198 22148 23204 22160
rect 22336 22120 23204 22148
rect 22336 22108 22342 22120
rect 23198 22108 23204 22120
rect 23256 22108 23262 22160
rect 23768 22148 23796 22188
rect 23842 22176 23848 22228
rect 23900 22216 23906 22228
rect 27338 22216 27344 22228
rect 23900 22188 27344 22216
rect 23900 22176 23906 22188
rect 27338 22176 27344 22188
rect 27396 22176 27402 22228
rect 27890 22216 27896 22228
rect 27448 22188 27896 22216
rect 24762 22148 24768 22160
rect 23768 22120 24768 22148
rect 24762 22108 24768 22120
rect 24820 22108 24826 22160
rect 24854 22108 24860 22160
rect 24912 22108 24918 22160
rect 26510 22108 26516 22160
rect 26568 22108 26574 22160
rect 22097 22083 22155 22089
rect 22097 22049 22109 22083
rect 22143 22080 22155 22083
rect 22830 22080 22836 22092
rect 22143 22052 22836 22080
rect 22143 22049 22155 22052
rect 22097 22043 22155 22049
rect 22830 22040 22836 22052
rect 22888 22040 22894 22092
rect 23293 22083 23351 22089
rect 23293 22049 23305 22083
rect 23339 22080 23351 22083
rect 25041 22083 25099 22089
rect 25041 22080 25053 22083
rect 23339 22052 25053 22080
rect 23339 22049 23351 22052
rect 23293 22043 23351 22049
rect 25041 22049 25053 22052
rect 25087 22049 25099 22083
rect 26053 22083 26111 22089
rect 26053 22080 26065 22083
rect 25041 22043 25099 22049
rect 25608 22052 26065 22080
rect 22738 22012 22744 22024
rect 21928 21984 22744 22012
rect 21637 21975 21695 21981
rect 11232 21947 11290 21953
rect 11232 21913 11244 21947
rect 11278 21944 11290 21947
rect 11790 21944 11796 21956
rect 11278 21916 11796 21944
rect 11278 21913 11290 21916
rect 11232 21907 11290 21913
rect 11790 21904 11796 21916
rect 11848 21904 11854 21956
rect 16758 21904 16764 21956
rect 16816 21944 16822 21956
rect 21082 21944 21088 21956
rect 16816 21916 21088 21944
rect 16816 21904 16822 21916
rect 21082 21904 21088 21916
rect 21140 21904 21146 21956
rect 21284 21944 21312 21975
rect 22738 21972 22744 21984
rect 22796 21972 22802 22024
rect 23017 22015 23075 22021
rect 23017 21981 23029 22015
rect 23063 22012 23075 22015
rect 23382 22012 23388 22024
rect 23063 21984 23388 22012
rect 23063 21981 23075 21984
rect 23017 21975 23075 21981
rect 23382 21972 23388 21984
rect 23440 21972 23446 22024
rect 23845 22015 23903 22021
rect 23845 21981 23857 22015
rect 23891 21981 23903 22015
rect 23845 21975 23903 21981
rect 22186 21944 22192 21956
rect 21284 21916 22192 21944
rect 22186 21904 22192 21916
rect 22244 21904 22250 21956
rect 22278 21904 22284 21956
rect 22336 21944 22342 21956
rect 23860 21944 23888 21975
rect 23934 21972 23940 22024
rect 23992 22012 23998 22024
rect 24029 22015 24087 22021
rect 24029 22012 24041 22015
rect 23992 21984 24041 22012
rect 23992 21972 23998 21984
rect 24029 21981 24041 21984
rect 24075 21981 24087 22015
rect 24029 21975 24087 21981
rect 24762 21972 24768 22024
rect 24820 22012 24826 22024
rect 25608 22012 25636 22052
rect 26053 22049 26065 22052
rect 26099 22080 26111 22083
rect 27062 22080 27068 22092
rect 26099 22052 27068 22080
rect 26099 22049 26111 22052
rect 26053 22043 26111 22049
rect 27062 22040 27068 22052
rect 27120 22040 27126 22092
rect 24820 21984 25636 22012
rect 26145 22015 26203 22021
rect 24820 21972 24826 21984
rect 26145 21981 26157 22015
rect 26191 22012 26203 22015
rect 27448 22012 27476 22188
rect 27890 22176 27896 22188
rect 27948 22176 27954 22228
rect 27982 22176 27988 22228
rect 28040 22216 28046 22228
rect 28040 22188 28764 22216
rect 28040 22176 28046 22188
rect 28626 22148 28632 22160
rect 27632 22120 28632 22148
rect 27632 22089 27660 22120
rect 28626 22108 28632 22120
rect 28684 22108 28690 22160
rect 28736 22148 28764 22188
rect 30006 22176 30012 22228
rect 30064 22216 30070 22228
rect 33134 22216 33140 22228
rect 30064 22188 33140 22216
rect 30064 22176 30070 22188
rect 33134 22176 33140 22188
rect 33192 22176 33198 22228
rect 33229 22219 33287 22225
rect 33229 22185 33241 22219
rect 33275 22216 33287 22219
rect 34422 22216 34428 22228
rect 33275 22188 34428 22216
rect 33275 22185 33287 22188
rect 33229 22179 33287 22185
rect 34422 22176 34428 22188
rect 34480 22176 34486 22228
rect 35529 22219 35587 22225
rect 35529 22185 35541 22219
rect 35575 22216 35587 22219
rect 35618 22216 35624 22228
rect 35575 22188 35624 22216
rect 35575 22185 35587 22188
rect 35529 22179 35587 22185
rect 35618 22176 35624 22188
rect 35676 22176 35682 22228
rect 38838 22216 38844 22228
rect 36372 22188 38844 22216
rect 30834 22148 30840 22160
rect 28736 22120 30840 22148
rect 30834 22108 30840 22120
rect 30892 22108 30898 22160
rect 32490 22148 32496 22160
rect 31404 22120 32496 22148
rect 27617 22083 27675 22089
rect 27617 22049 27629 22083
rect 27663 22080 27675 22083
rect 27663 22052 27697 22080
rect 27663 22049 27675 22052
rect 27617 22043 27675 22049
rect 27798 22040 27804 22092
rect 27856 22040 27862 22092
rect 28534 22089 28540 22092
rect 28517 22083 28540 22089
rect 28517 22049 28529 22083
rect 28517 22043 28540 22049
rect 28534 22040 28540 22043
rect 28592 22040 28598 22092
rect 29546 22040 29552 22092
rect 29604 22080 29610 22092
rect 30009 22083 30067 22089
rect 30009 22080 30021 22083
rect 29604 22052 30021 22080
rect 29604 22040 29610 22052
rect 30009 22049 30021 22052
rect 30055 22049 30067 22083
rect 30009 22043 30067 22049
rect 26191 21984 27476 22012
rect 26191 21981 26203 21984
rect 26145 21975 26203 21981
rect 27522 21972 27528 22024
rect 27580 21972 27586 22024
rect 28074 21972 28080 22024
rect 28132 22012 28138 22024
rect 28629 22015 28687 22021
rect 28629 22012 28641 22015
rect 28132 21984 28641 22012
rect 28132 21972 28138 21984
rect 28629 21981 28641 21984
rect 28675 21981 28687 22015
rect 28629 21975 28687 21981
rect 28994 21972 29000 22024
rect 29052 21972 29058 22024
rect 29825 22015 29883 22021
rect 29825 21981 29837 22015
rect 29871 21981 29883 22015
rect 29825 21975 29883 21981
rect 29917 22015 29975 22021
rect 29917 21981 29929 22015
rect 29963 22012 29975 22015
rect 30098 22012 30104 22024
rect 29963 21984 30104 22012
rect 29963 21981 29975 21984
rect 29917 21975 29975 21981
rect 24581 21947 24639 21953
rect 24581 21944 24593 21947
rect 22336 21916 24593 21944
rect 22336 21904 22342 21916
rect 24581 21913 24593 21916
rect 24627 21944 24639 21947
rect 25406 21944 25412 21956
rect 24627 21916 25412 21944
rect 24627 21913 24639 21916
rect 24581 21907 24639 21913
rect 25406 21904 25412 21916
rect 25464 21904 25470 21956
rect 27540 21944 27568 21972
rect 28442 21944 28448 21956
rect 27540 21916 28448 21944
rect 28442 21904 28448 21916
rect 28500 21904 28506 21956
rect 28534 21904 28540 21956
rect 28592 21944 28598 21956
rect 28902 21944 28908 21956
rect 28592 21916 28908 21944
rect 28592 21904 28598 21916
rect 28902 21904 28908 21916
rect 28960 21904 28966 21956
rect 29840 21944 29868 21975
rect 30098 21972 30104 21984
rect 30156 21972 30162 22024
rect 31018 21972 31024 22024
rect 31076 21972 31082 22024
rect 31110 21972 31116 22024
rect 31168 22012 31174 22024
rect 31297 22015 31355 22021
rect 31168 21984 31213 22012
rect 31168 21972 31174 21984
rect 31297 21981 31309 22015
rect 31343 22012 31355 22015
rect 31404 22012 31432 22120
rect 32490 22108 32496 22120
rect 32548 22148 32554 22160
rect 32950 22148 32956 22160
rect 32548 22120 32956 22148
rect 32548 22108 32554 22120
rect 32950 22108 32956 22120
rect 33008 22108 33014 22160
rect 33410 22108 33416 22160
rect 33468 22108 33474 22160
rect 34882 22148 34888 22160
rect 33796 22120 34888 22148
rect 33428 22080 33456 22108
rect 33796 22092 33824 22120
rect 34882 22108 34888 22120
rect 34940 22108 34946 22160
rect 36372 22148 36400 22188
rect 38838 22176 38844 22188
rect 38896 22176 38902 22228
rect 36280 22120 36400 22148
rect 32416 22052 33456 22080
rect 31343 21984 31432 22012
rect 31343 21981 31355 21984
rect 31297 21975 31355 21981
rect 31478 21972 31484 22024
rect 31536 22021 31542 22024
rect 32306 22021 32312 22024
rect 31536 22012 31544 22021
rect 32125 22015 32183 22021
rect 32125 22012 32137 22015
rect 31536 21984 32137 22012
rect 31536 21975 31544 21984
rect 32125 21981 32137 21984
rect 32171 21981 32183 22015
rect 32125 21975 32183 21981
rect 32273 22015 32312 22021
rect 32273 21981 32285 22015
rect 32273 21975 32312 21981
rect 31536 21972 31542 21975
rect 32306 21972 32312 21975
rect 32364 21972 32370 22024
rect 32416 22021 32444 22052
rect 33778 22040 33784 22092
rect 33836 22040 33842 22092
rect 33870 22040 33876 22092
rect 33928 22080 33934 22092
rect 34146 22080 34152 22092
rect 33928 22052 34152 22080
rect 33928 22040 33934 22052
rect 34146 22040 34152 22052
rect 34204 22040 34210 22092
rect 35526 22080 35532 22092
rect 35176 22052 35532 22080
rect 32674 22021 32680 22024
rect 32401 22015 32459 22021
rect 32401 21981 32413 22015
rect 32447 21981 32459 22015
rect 32401 21975 32459 21981
rect 32631 22015 32680 22021
rect 32631 21981 32643 22015
rect 32677 21981 32680 22015
rect 32631 21975 32680 21981
rect 32674 21972 32680 21975
rect 32732 21972 32738 22024
rect 32766 21972 32772 22024
rect 32824 22012 32830 22024
rect 33226 22012 33232 22024
rect 32824 21984 33232 22012
rect 32824 21972 32830 21984
rect 33226 21972 33232 21984
rect 33284 21972 33290 22024
rect 33410 21972 33416 22024
rect 33468 21972 33474 22024
rect 33505 22015 33563 22021
rect 33505 21981 33517 22015
rect 33551 22012 33563 22015
rect 33686 22012 33692 22024
rect 33551 21984 33692 22012
rect 33551 21981 33563 21984
rect 33505 21975 33563 21981
rect 33686 21972 33692 21984
rect 33744 22012 33750 22024
rect 33962 22012 33968 22024
rect 33744 21984 33968 22012
rect 33744 21972 33750 21984
rect 33962 21972 33968 21984
rect 34020 21972 34026 22024
rect 34790 21972 34796 22024
rect 34848 22012 34854 22024
rect 35066 22021 35072 22024
rect 34885 22015 34943 22021
rect 34885 22012 34897 22015
rect 34848 21984 34897 22012
rect 34848 21972 34854 21984
rect 34885 21981 34897 21984
rect 34931 21981 34943 22015
rect 34885 21975 34943 21981
rect 35033 22015 35072 22021
rect 35033 21981 35045 22015
rect 35033 21975 35072 21981
rect 35066 21972 35072 21975
rect 35124 21972 35130 22024
rect 35176 22021 35204 22052
rect 35526 22040 35532 22052
rect 35584 22040 35590 22092
rect 36280 22089 36308 22120
rect 36265 22083 36323 22089
rect 36265 22049 36277 22083
rect 36311 22049 36323 22083
rect 36265 22043 36323 22049
rect 36906 22040 36912 22092
rect 36964 22040 36970 22092
rect 35161 22015 35219 22021
rect 35161 21981 35173 22015
rect 35207 21981 35219 22015
rect 35161 21975 35219 21981
rect 35391 22015 35449 22021
rect 35391 21981 35403 22015
rect 35437 22012 35449 22015
rect 35802 22012 35808 22024
rect 35437 21984 35808 22012
rect 35437 21981 35449 21984
rect 35391 21975 35449 21981
rect 35802 21972 35808 21984
rect 35860 21972 35866 22024
rect 35986 21972 35992 22024
rect 36044 21972 36050 22024
rect 36525 21984 37320 22012
rect 30374 21944 30380 21956
rect 29840 21916 30380 21944
rect 30374 21904 30380 21916
rect 30432 21904 30438 21956
rect 30558 21904 30564 21956
rect 30616 21944 30622 21956
rect 31389 21947 31447 21953
rect 31389 21944 31401 21947
rect 30616 21916 31401 21944
rect 30616 21904 30622 21916
rect 31389 21913 31401 21916
rect 31435 21913 31447 21947
rect 32493 21947 32551 21953
rect 32493 21944 32505 21947
rect 31389 21907 31447 21913
rect 31496 21916 32505 21944
rect 12342 21836 12348 21888
rect 12400 21836 12406 21888
rect 13078 21836 13084 21888
rect 13136 21876 13142 21888
rect 18138 21876 18144 21888
rect 13136 21848 18144 21876
rect 13136 21836 13142 21848
rect 18138 21836 18144 21848
rect 18196 21836 18202 21888
rect 18598 21836 18604 21888
rect 18656 21876 18662 21888
rect 20441 21879 20499 21885
rect 20441 21876 20453 21879
rect 18656 21848 20453 21876
rect 18656 21836 18662 21848
rect 20441 21845 20453 21848
rect 20487 21845 20499 21879
rect 20441 21839 20499 21845
rect 22370 21836 22376 21888
rect 22428 21876 22434 21888
rect 22649 21879 22707 21885
rect 22649 21876 22661 21879
rect 22428 21848 22661 21876
rect 22428 21836 22434 21848
rect 22649 21845 22661 21848
rect 22695 21845 22707 21879
rect 22649 21839 22707 21845
rect 23109 21879 23167 21885
rect 23109 21845 23121 21879
rect 23155 21876 23167 21879
rect 23198 21876 23204 21888
rect 23155 21848 23204 21876
rect 23155 21845 23167 21848
rect 23109 21839 23167 21845
rect 23198 21836 23204 21848
rect 23256 21836 23262 21888
rect 23937 21879 23995 21885
rect 23937 21845 23949 21879
rect 23983 21876 23995 21879
rect 24118 21876 24124 21888
rect 23983 21848 24124 21876
rect 23983 21845 23995 21848
rect 23937 21839 23995 21845
rect 24118 21836 24124 21848
rect 24176 21836 24182 21888
rect 24210 21836 24216 21888
rect 24268 21876 24274 21888
rect 26418 21876 26424 21888
rect 24268 21848 26424 21876
rect 24268 21836 24274 21848
rect 26418 21836 26424 21848
rect 26476 21836 26482 21888
rect 27157 21879 27215 21885
rect 27157 21845 27169 21879
rect 27203 21876 27215 21879
rect 28258 21876 28264 21888
rect 27203 21848 28264 21876
rect 27203 21845 27215 21848
rect 27157 21839 27215 21845
rect 28258 21836 28264 21848
rect 28316 21836 28322 21888
rect 28350 21836 28356 21888
rect 28408 21836 28414 21888
rect 28994 21836 29000 21888
rect 29052 21876 29058 21888
rect 31496 21876 31524 21916
rect 32048 21888 32076 21916
rect 32493 21913 32505 21916
rect 32539 21913 32551 21947
rect 32493 21907 32551 21913
rect 32600 21916 32904 21944
rect 29052 21848 31524 21876
rect 29052 21836 29058 21848
rect 31570 21836 31576 21888
rect 31628 21876 31634 21888
rect 31665 21879 31723 21885
rect 31665 21876 31677 21879
rect 31628 21848 31677 21876
rect 31628 21836 31634 21848
rect 31665 21845 31677 21848
rect 31711 21845 31723 21879
rect 31665 21839 31723 21845
rect 32030 21836 32036 21888
rect 32088 21836 32094 21888
rect 32122 21836 32128 21888
rect 32180 21876 32186 21888
rect 32600 21876 32628 21916
rect 32180 21848 32628 21876
rect 32180 21836 32186 21848
rect 32766 21836 32772 21888
rect 32824 21836 32830 21888
rect 32876 21876 32904 21916
rect 35250 21904 35256 21956
rect 35308 21944 35314 21956
rect 36525 21944 36553 21984
rect 37182 21953 37188 21956
rect 35308 21916 36553 21944
rect 35308 21904 35314 21916
rect 37176 21907 37188 21953
rect 37182 21904 37188 21907
rect 37240 21904 37246 21956
rect 37292 21944 37320 21984
rect 37550 21972 37556 22024
rect 37608 22012 37614 22024
rect 38286 22012 38292 22024
rect 37608 21984 38292 22012
rect 37608 21972 37614 21984
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 37292 21916 38332 21944
rect 38304 21888 38332 21916
rect 38194 21876 38200 21888
rect 32876 21848 38200 21876
rect 38194 21836 38200 21848
rect 38252 21836 38258 21888
rect 38286 21836 38292 21888
rect 38344 21836 38350 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 11790 21632 11796 21684
rect 11848 21632 11854 21684
rect 12158 21632 12164 21684
rect 12216 21672 12222 21684
rect 12253 21675 12311 21681
rect 12253 21672 12265 21675
rect 12216 21644 12265 21672
rect 12216 21632 12222 21644
rect 12253 21641 12265 21644
rect 12299 21641 12311 21675
rect 12253 21635 12311 21641
rect 14737 21675 14795 21681
rect 14737 21641 14749 21675
rect 14783 21672 14795 21675
rect 15838 21672 15844 21684
rect 14783 21644 15844 21672
rect 14783 21641 14795 21644
rect 14737 21635 14795 21641
rect 15838 21632 15844 21644
rect 15896 21632 15902 21684
rect 18230 21632 18236 21684
rect 18288 21632 18294 21684
rect 19242 21672 19248 21684
rect 18708 21644 19248 21672
rect 12342 21564 12348 21616
rect 12400 21564 12406 21616
rect 13814 21604 13820 21616
rect 13372 21576 13820 21604
rect 12161 21539 12219 21545
rect 12161 21505 12173 21539
rect 12207 21536 12219 21539
rect 12360 21536 12388 21564
rect 13372 21545 13400 21576
rect 13814 21564 13820 21576
rect 13872 21564 13878 21616
rect 14274 21564 14280 21616
rect 14332 21604 14338 21616
rect 17954 21604 17960 21616
rect 14332 21576 17960 21604
rect 14332 21564 14338 21576
rect 17954 21564 17960 21576
rect 18012 21604 18018 21616
rect 18708 21613 18736 21644
rect 19242 21632 19248 21644
rect 19300 21632 19306 21684
rect 20254 21632 20260 21684
rect 20312 21672 20318 21684
rect 20622 21672 20628 21684
rect 20312 21644 20628 21672
rect 20312 21632 20318 21644
rect 20622 21632 20628 21644
rect 20680 21632 20686 21684
rect 21361 21675 21419 21681
rect 21361 21641 21373 21675
rect 21407 21672 21419 21675
rect 22186 21672 22192 21684
rect 21407 21644 22192 21672
rect 21407 21641 21419 21644
rect 21361 21635 21419 21641
rect 22186 21632 22192 21644
rect 22244 21672 22250 21684
rect 23382 21672 23388 21684
rect 22244 21644 23388 21672
rect 22244 21632 22250 21644
rect 23382 21632 23388 21644
rect 23440 21632 23446 21684
rect 23842 21632 23848 21684
rect 23900 21632 23906 21684
rect 23934 21632 23940 21684
rect 23992 21632 23998 21684
rect 24394 21632 24400 21684
rect 24452 21672 24458 21684
rect 25041 21675 25099 21681
rect 25041 21672 25053 21675
rect 24452 21644 25053 21672
rect 24452 21632 24458 21644
rect 25041 21641 25053 21644
rect 25087 21641 25099 21675
rect 25041 21635 25099 21641
rect 26602 21632 26608 21684
rect 26660 21672 26666 21684
rect 27154 21672 27160 21684
rect 26660 21644 27160 21672
rect 26660 21632 26666 21644
rect 27154 21632 27160 21644
rect 27212 21632 27218 21684
rect 28074 21632 28080 21684
rect 28132 21632 28138 21684
rect 28994 21672 29000 21684
rect 28276 21644 29000 21672
rect 18693 21607 18751 21613
rect 18693 21604 18705 21607
rect 18012 21576 18705 21604
rect 18012 21564 18018 21576
rect 18693 21573 18705 21576
rect 18739 21573 18751 21607
rect 18693 21567 18751 21573
rect 19150 21564 19156 21616
rect 19208 21604 19214 21616
rect 19429 21607 19487 21613
rect 19429 21604 19441 21607
rect 19208 21576 19441 21604
rect 19208 21564 19214 21576
rect 19429 21573 19441 21576
rect 19475 21573 19487 21607
rect 20990 21604 20996 21616
rect 19429 21567 19487 21573
rect 19536 21576 20996 21604
rect 13357 21539 13415 21545
rect 12207 21508 13216 21536
rect 12207 21505 12219 21508
rect 12161 21499 12219 21505
rect 12250 21428 12256 21480
rect 12308 21468 12314 21480
rect 12345 21471 12403 21477
rect 12345 21468 12357 21471
rect 12308 21440 12357 21468
rect 12308 21428 12314 21440
rect 12345 21437 12357 21440
rect 12391 21437 12403 21471
rect 12345 21431 12403 21437
rect 5166 21360 5172 21412
rect 5224 21400 5230 21412
rect 13078 21400 13084 21412
rect 5224 21372 13084 21400
rect 5224 21360 5230 21372
rect 13078 21360 13084 21372
rect 13136 21360 13142 21412
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 11054 21332 11060 21344
rect 6972 21304 11060 21332
rect 6972 21292 6978 21304
rect 11054 21292 11060 21304
rect 11112 21292 11118 21344
rect 13188 21332 13216 21508
rect 13357 21505 13369 21539
rect 13403 21505 13415 21539
rect 13357 21499 13415 21505
rect 13630 21496 13636 21548
rect 13688 21536 13694 21548
rect 14369 21539 14427 21545
rect 14369 21536 14381 21539
rect 13688 21508 14381 21536
rect 13688 21496 13694 21508
rect 14369 21505 14381 21508
rect 14415 21505 14427 21539
rect 14369 21499 14427 21505
rect 14826 21496 14832 21548
rect 14884 21536 14890 21548
rect 15473 21539 15531 21545
rect 15473 21536 15485 21539
rect 14884 21508 15485 21536
rect 14884 21496 14890 21508
rect 15473 21505 15485 21508
rect 15519 21505 15531 21539
rect 15473 21499 15531 21505
rect 13446 21428 13452 21480
rect 13504 21428 13510 21480
rect 14277 21471 14335 21477
rect 14277 21468 14289 21471
rect 13740 21440 14289 21468
rect 13740 21409 13768 21440
rect 14277 21437 14289 21440
rect 14323 21437 14335 21471
rect 14277 21431 14335 21437
rect 13725 21403 13783 21409
rect 13725 21369 13737 21403
rect 13771 21369 13783 21403
rect 15488 21400 15516 21499
rect 15562 21496 15568 21548
rect 15620 21536 15626 21548
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 15620 21508 16865 21536
rect 15620 21496 15626 21508
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21536 17095 21539
rect 19536 21536 19564 21576
rect 20990 21564 20996 21576
rect 21048 21564 21054 21616
rect 22738 21604 22744 21616
rect 21192 21576 22744 21604
rect 17083 21508 19564 21536
rect 17083 21505 17095 21508
rect 17037 21499 17095 21505
rect 15654 21428 15660 21480
rect 15712 21468 15718 21480
rect 15749 21471 15807 21477
rect 15749 21468 15761 21471
rect 15712 21440 15761 21468
rect 15712 21428 15718 21440
rect 15749 21437 15761 21440
rect 15795 21468 15807 21471
rect 16758 21468 16764 21480
rect 15795 21440 16764 21468
rect 15795 21437 15807 21440
rect 15749 21431 15807 21437
rect 16758 21428 16764 21440
rect 16816 21428 16822 21480
rect 17052 21400 17080 21499
rect 20070 21496 20076 21548
rect 20128 21536 20134 21548
rect 21192 21545 21220 21576
rect 22738 21564 22744 21576
rect 22796 21564 22802 21616
rect 24118 21564 24124 21616
rect 24176 21564 24182 21616
rect 25590 21564 25596 21616
rect 25648 21604 25654 21616
rect 26142 21604 26148 21616
rect 25648 21576 26148 21604
rect 25648 21564 25654 21576
rect 26142 21564 26148 21576
rect 26200 21564 26206 21616
rect 26237 21607 26295 21613
rect 26237 21573 26249 21607
rect 26283 21604 26295 21607
rect 28276 21604 28304 21644
rect 28994 21632 29000 21644
rect 29052 21632 29058 21684
rect 29822 21632 29828 21684
rect 29880 21672 29886 21684
rect 30006 21672 30012 21684
rect 29880 21644 30012 21672
rect 29880 21632 29886 21644
rect 30006 21632 30012 21644
rect 30064 21632 30070 21684
rect 31018 21632 31024 21684
rect 31076 21672 31082 21684
rect 31389 21675 31447 21681
rect 31389 21672 31401 21675
rect 31076 21644 31401 21672
rect 31076 21632 31082 21644
rect 31389 21641 31401 21644
rect 31435 21641 31447 21675
rect 31389 21635 31447 21641
rect 32232 21644 32628 21672
rect 28626 21604 28632 21616
rect 26283 21576 28304 21604
rect 28368 21576 28632 21604
rect 26283 21573 26295 21576
rect 26237 21567 26295 21573
rect 20198 21539 20256 21545
rect 20198 21536 20210 21539
rect 20128 21508 20210 21536
rect 20128 21496 20134 21508
rect 20198 21505 20210 21508
rect 20244 21505 20256 21539
rect 21177 21539 21235 21545
rect 21177 21536 21189 21539
rect 20198 21499 20256 21505
rect 20364 21508 21189 21536
rect 17773 21471 17831 21477
rect 17773 21437 17785 21471
rect 17819 21468 17831 21471
rect 18506 21468 18512 21480
rect 17819 21440 18512 21468
rect 17819 21437 17831 21440
rect 17773 21431 17831 21437
rect 18506 21428 18512 21440
rect 18564 21428 18570 21480
rect 19150 21428 19156 21480
rect 19208 21468 19214 21480
rect 20364 21468 20392 21508
rect 21177 21505 21189 21508
rect 21223 21505 21235 21539
rect 21177 21499 21235 21505
rect 21450 21496 21456 21548
rect 21508 21496 21514 21548
rect 22278 21496 22284 21548
rect 22336 21496 22342 21548
rect 22370 21496 22376 21548
rect 22428 21496 22434 21548
rect 22465 21539 22523 21545
rect 22465 21505 22477 21539
rect 22511 21536 22523 21539
rect 22554 21536 22560 21548
rect 22511 21508 22560 21536
rect 22511 21505 22523 21508
rect 22465 21499 22523 21505
rect 22554 21496 22560 21508
rect 22612 21496 22618 21548
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21536 22707 21539
rect 23566 21536 23572 21548
rect 22695 21508 23572 21536
rect 22695 21505 22707 21508
rect 22649 21499 22707 21505
rect 19208 21440 20392 21468
rect 20717 21471 20775 21477
rect 19208 21428 19214 21440
rect 20717 21437 20729 21471
rect 20763 21437 20775 21471
rect 20717 21431 20775 21437
rect 15488 21372 17080 21400
rect 18141 21403 18199 21409
rect 13725 21363 13783 21369
rect 18141 21369 18153 21403
rect 18187 21400 18199 21403
rect 18690 21400 18696 21412
rect 18187 21372 18696 21400
rect 18187 21369 18199 21372
rect 18141 21363 18199 21369
rect 18690 21360 18696 21372
rect 18748 21400 18754 21412
rect 20438 21400 20444 21412
rect 18748 21372 20444 21400
rect 18748 21360 18754 21372
rect 20438 21360 20444 21372
rect 20496 21360 20502 21412
rect 20732 21400 20760 21431
rect 21082 21428 21088 21480
rect 21140 21468 21146 21480
rect 22664 21468 22692 21499
rect 23566 21496 23572 21508
rect 23624 21496 23630 21548
rect 23750 21496 23756 21548
rect 23808 21496 23814 21548
rect 24486 21496 24492 21548
rect 24544 21536 24550 21548
rect 24581 21539 24639 21545
rect 24581 21536 24593 21539
rect 24544 21508 24593 21536
rect 24544 21496 24550 21508
rect 24581 21505 24593 21508
rect 24627 21505 24639 21539
rect 24581 21499 24639 21505
rect 24857 21539 24915 21545
rect 24857 21505 24869 21539
rect 24903 21536 24915 21539
rect 25038 21536 25044 21548
rect 24903 21508 25044 21536
rect 24903 21505 24915 21508
rect 24857 21499 24915 21505
rect 25038 21496 25044 21508
rect 25096 21536 25102 21548
rect 25406 21536 25412 21548
rect 25096 21508 25412 21536
rect 25096 21496 25102 21508
rect 25406 21496 25412 21508
rect 25464 21496 25470 21548
rect 25961 21539 26019 21545
rect 25961 21505 25973 21539
rect 26007 21505 26019 21539
rect 25961 21499 26019 21505
rect 26381 21539 26439 21545
rect 26381 21505 26393 21539
rect 26427 21536 26439 21539
rect 26878 21536 26884 21548
rect 26427 21508 26884 21536
rect 26427 21505 26439 21508
rect 26381 21499 26439 21505
rect 21140 21440 22692 21468
rect 21140 21428 21146 21440
rect 24302 21428 24308 21480
rect 24360 21468 24366 21480
rect 24673 21471 24731 21477
rect 24673 21468 24685 21471
rect 24360 21440 24685 21468
rect 24360 21428 24366 21440
rect 24673 21437 24685 21440
rect 24719 21437 24731 21471
rect 24673 21431 24731 21437
rect 25590 21428 25596 21480
rect 25648 21468 25654 21480
rect 25866 21468 25872 21480
rect 25648 21440 25872 21468
rect 25648 21428 25654 21440
rect 25866 21428 25872 21440
rect 25924 21428 25930 21480
rect 25976 21468 26004 21499
rect 26878 21496 26884 21508
rect 26936 21496 26942 21548
rect 27062 21496 27068 21548
rect 27120 21536 27126 21548
rect 28368 21545 28396 21576
rect 28626 21564 28632 21576
rect 28684 21564 28690 21616
rect 29270 21604 29276 21616
rect 28736 21576 29276 21604
rect 27249 21539 27307 21545
rect 27249 21536 27261 21539
rect 27120 21508 27261 21536
rect 27120 21496 27126 21508
rect 27249 21505 27261 21508
rect 27295 21505 27307 21539
rect 27249 21499 27307 21505
rect 28353 21539 28411 21545
rect 28353 21505 28365 21539
rect 28399 21505 28411 21539
rect 28353 21499 28411 21505
rect 28442 21496 28448 21548
rect 28500 21496 28506 21548
rect 28534 21496 28540 21548
rect 28592 21496 28598 21548
rect 26050 21468 26056 21480
rect 25976 21440 26056 21468
rect 26050 21428 26056 21440
rect 26108 21468 26114 21480
rect 26108 21440 26740 21468
rect 26108 21428 26114 21440
rect 21177 21403 21235 21409
rect 21177 21400 21189 21403
rect 20732 21372 21189 21400
rect 21177 21369 21189 21372
rect 21223 21369 21235 21403
rect 21177 21363 21235 21369
rect 21634 21360 21640 21412
rect 21692 21400 21698 21412
rect 22738 21400 22744 21412
rect 21692 21372 22744 21400
rect 21692 21360 21698 21372
rect 22738 21360 22744 21372
rect 22796 21360 22802 21412
rect 22830 21360 22836 21412
rect 22888 21400 22894 21412
rect 23569 21403 23627 21409
rect 23569 21400 23581 21403
rect 22888 21372 23581 21400
rect 22888 21360 22894 21372
rect 23569 21369 23581 21372
rect 23615 21369 23627 21403
rect 26712 21400 26740 21440
rect 27154 21428 27160 21480
rect 27212 21468 27218 21480
rect 27341 21471 27399 21477
rect 27341 21468 27353 21471
rect 27212 21440 27353 21468
rect 27212 21428 27218 21440
rect 27341 21437 27353 21440
rect 27387 21437 27399 21471
rect 27798 21468 27804 21480
rect 27341 21431 27399 21437
rect 27448 21440 27804 21468
rect 27448 21400 27476 21440
rect 27798 21428 27804 21440
rect 27856 21428 27862 21480
rect 28258 21428 28264 21480
rect 28316 21468 28322 21480
rect 28736 21468 28764 21576
rect 29270 21564 29276 21576
rect 29328 21564 29334 21616
rect 30101 21607 30159 21613
rect 30101 21573 30113 21607
rect 30147 21604 30159 21607
rect 30190 21604 30196 21616
rect 30147 21576 30196 21604
rect 30147 21573 30159 21576
rect 30101 21567 30159 21573
rect 30190 21564 30196 21576
rect 30248 21564 30254 21616
rect 30282 21564 30288 21616
rect 30340 21564 30346 21616
rect 32122 21604 32128 21616
rect 30852 21576 32128 21604
rect 28994 21496 29000 21548
rect 29052 21536 29058 21548
rect 29089 21539 29147 21545
rect 29089 21536 29101 21539
rect 29052 21508 29101 21536
rect 29052 21496 29058 21508
rect 29089 21505 29101 21508
rect 29135 21505 29147 21539
rect 29089 21499 29147 21505
rect 29178 21496 29184 21548
rect 29236 21536 29242 21548
rect 30377 21539 30435 21545
rect 29236 21508 29581 21536
rect 29236 21496 29242 21508
rect 28316 21440 28764 21468
rect 28316 21428 28322 21440
rect 28810 21428 28816 21480
rect 28868 21468 28874 21480
rect 29365 21471 29423 21477
rect 28868 21440 29316 21468
rect 28868 21428 28874 21440
rect 23569 21363 23627 21369
rect 23676 21372 26648 21400
rect 26712 21372 27476 21400
rect 27617 21403 27675 21409
rect 15562 21332 15568 21344
rect 13188 21304 15568 21332
rect 15562 21292 15568 21304
rect 15620 21292 15626 21344
rect 17221 21335 17279 21341
rect 17221 21301 17233 21335
rect 17267 21332 17279 21335
rect 17770 21332 17776 21344
rect 17267 21304 17776 21332
rect 17267 21301 17279 21304
rect 17221 21295 17279 21301
rect 17770 21292 17776 21304
rect 17828 21332 17834 21344
rect 19978 21332 19984 21344
rect 17828 21304 19984 21332
rect 17828 21292 17834 21304
rect 19978 21292 19984 21304
rect 20036 21292 20042 21344
rect 20070 21292 20076 21344
rect 20128 21292 20134 21344
rect 20162 21292 20168 21344
rect 20220 21332 20226 21344
rect 20530 21332 20536 21344
rect 20220 21304 20536 21332
rect 20220 21292 20226 21304
rect 20530 21292 20536 21304
rect 20588 21292 20594 21344
rect 20622 21292 20628 21344
rect 20680 21292 20686 21344
rect 22002 21292 22008 21344
rect 22060 21292 22066 21344
rect 22462 21292 22468 21344
rect 22520 21332 22526 21344
rect 23676 21332 23704 21372
rect 22520 21304 23704 21332
rect 22520 21292 22526 21304
rect 24578 21292 24584 21344
rect 24636 21292 24642 21344
rect 26510 21292 26516 21344
rect 26568 21292 26574 21344
rect 26620 21332 26648 21372
rect 27617 21369 27629 21403
rect 27663 21400 27675 21403
rect 28994 21400 29000 21412
rect 27663 21372 29000 21400
rect 27663 21369 27675 21372
rect 27617 21363 27675 21369
rect 28994 21360 29000 21372
rect 29052 21360 29058 21412
rect 29288 21400 29316 21440
rect 29365 21437 29377 21471
rect 29411 21468 29423 21471
rect 29454 21468 29460 21480
rect 29411 21440 29460 21468
rect 29411 21437 29423 21440
rect 29365 21431 29423 21437
rect 29454 21428 29460 21440
rect 29512 21428 29518 21480
rect 29553 21468 29581 21508
rect 30377 21505 30389 21539
rect 30423 21536 30435 21539
rect 30650 21536 30656 21548
rect 30423 21508 30656 21536
rect 30423 21505 30435 21508
rect 30377 21499 30435 21505
rect 30650 21496 30656 21508
rect 30708 21496 30714 21548
rect 30852 21545 30880 21576
rect 32122 21564 32128 21576
rect 32180 21564 32186 21616
rect 30837 21539 30895 21545
rect 30837 21505 30849 21539
rect 30883 21505 30895 21539
rect 30837 21499 30895 21505
rect 31021 21539 31079 21545
rect 31021 21505 31033 21539
rect 31067 21505 31079 21539
rect 31021 21499 31079 21505
rect 31036 21468 31064 21499
rect 31110 21496 31116 21548
rect 31168 21496 31174 21548
rect 31205 21539 31263 21545
rect 31205 21505 31217 21539
rect 31251 21505 31263 21539
rect 31205 21499 31263 21505
rect 31220 21468 31248 21499
rect 31386 21496 31392 21548
rect 31444 21536 31450 21548
rect 32232 21536 32260 21644
rect 32490 21564 32496 21616
rect 32548 21564 32554 21616
rect 32600 21613 32628 21644
rect 33318 21632 33324 21684
rect 33376 21672 33382 21684
rect 34606 21672 34612 21684
rect 33376 21644 34612 21672
rect 33376 21632 33382 21644
rect 34606 21632 34612 21644
rect 34664 21632 34670 21684
rect 37182 21632 37188 21684
rect 37240 21672 37246 21684
rect 37461 21675 37519 21681
rect 37461 21672 37473 21675
rect 37240 21644 37473 21672
rect 37240 21632 37246 21644
rect 37461 21641 37473 21644
rect 37507 21641 37519 21675
rect 37461 21635 37519 21641
rect 37829 21675 37887 21681
rect 37829 21641 37841 21675
rect 37875 21672 37887 21675
rect 38286 21672 38292 21684
rect 37875 21644 38292 21672
rect 37875 21641 37887 21644
rect 37829 21635 37887 21641
rect 38286 21632 38292 21644
rect 38344 21632 38350 21684
rect 32585 21607 32643 21613
rect 32585 21573 32597 21607
rect 32631 21573 32643 21607
rect 35250 21604 35256 21616
rect 32585 21567 32643 21573
rect 34624 21576 35256 21604
rect 31444 21508 32260 21536
rect 31444 21496 31450 21508
rect 32306 21496 32312 21548
rect 32364 21496 32370 21548
rect 32674 21496 32680 21548
rect 32732 21496 32738 21548
rect 32766 21496 32772 21548
rect 32824 21536 32830 21548
rect 33321 21539 33379 21545
rect 33321 21536 33333 21539
rect 32824 21508 33333 21536
rect 32824 21496 32830 21508
rect 33321 21505 33333 21508
rect 33367 21505 33379 21539
rect 33321 21499 33379 21505
rect 33505 21539 33563 21545
rect 33505 21505 33517 21539
rect 33551 21536 33563 21539
rect 33594 21536 33600 21548
rect 33551 21508 33600 21536
rect 33551 21505 33563 21508
rect 33505 21499 33563 21505
rect 33594 21496 33600 21508
rect 33652 21496 33658 21548
rect 34514 21496 34520 21548
rect 34572 21496 34578 21548
rect 34624 21545 34652 21576
rect 35250 21564 35256 21576
rect 35308 21564 35314 21616
rect 35434 21564 35440 21616
rect 35492 21604 35498 21616
rect 35621 21607 35679 21613
rect 35621 21604 35633 21607
rect 35492 21576 35633 21604
rect 35492 21564 35498 21576
rect 35621 21573 35633 21576
rect 35667 21573 35679 21607
rect 36078 21604 36084 21616
rect 35621 21567 35679 21573
rect 35719 21576 36084 21604
rect 34610 21539 34668 21545
rect 34610 21505 34622 21539
rect 34656 21505 34668 21539
rect 34610 21499 34668 21505
rect 34793 21539 34851 21545
rect 34793 21505 34805 21539
rect 34839 21505 34851 21539
rect 34793 21499 34851 21505
rect 32692 21468 32720 21496
rect 34422 21468 34428 21480
rect 29553 21440 31064 21468
rect 31129 21440 34428 21468
rect 29641 21403 29699 21409
rect 29641 21400 29653 21403
rect 29288 21372 29653 21400
rect 29641 21369 29653 21372
rect 29687 21369 29699 21403
rect 30466 21400 30472 21412
rect 29641 21363 29699 21369
rect 29748 21372 30472 21400
rect 26970 21332 26976 21344
rect 26620 21304 26976 21332
rect 26970 21292 26976 21304
rect 27028 21292 27034 21344
rect 27433 21335 27491 21341
rect 27433 21301 27445 21335
rect 27479 21332 27491 21335
rect 27522 21332 27528 21344
rect 27479 21304 27528 21332
rect 27479 21301 27491 21304
rect 27433 21295 27491 21301
rect 27522 21292 27528 21304
rect 27580 21292 27586 21344
rect 28442 21292 28448 21344
rect 28500 21332 28506 21344
rect 29181 21335 29239 21341
rect 29181 21332 29193 21335
rect 28500 21304 29193 21332
rect 28500 21292 28506 21304
rect 29181 21301 29193 21304
rect 29227 21301 29239 21335
rect 29181 21295 29239 21301
rect 29546 21292 29552 21344
rect 29604 21332 29610 21344
rect 29748 21332 29776 21372
rect 30466 21360 30472 21372
rect 30524 21360 30530 21412
rect 30742 21360 30748 21412
rect 30800 21400 30806 21412
rect 31129 21400 31157 21440
rect 34422 21428 34428 21440
rect 34480 21428 34486 21480
rect 34698 21428 34704 21480
rect 34756 21468 34762 21480
rect 34808 21468 34836 21499
rect 34882 21496 34888 21548
rect 34940 21496 34946 21548
rect 35023 21539 35081 21545
rect 35023 21505 35035 21539
rect 35069 21536 35081 21539
rect 35342 21536 35348 21548
rect 35069 21508 35348 21536
rect 35069 21505 35081 21508
rect 35023 21499 35081 21505
rect 35342 21496 35348 21508
rect 35400 21496 35406 21548
rect 35719 21468 35747 21576
rect 36078 21564 36084 21576
rect 36136 21564 36142 21616
rect 35805 21539 35863 21545
rect 35805 21505 35817 21539
rect 35851 21505 35863 21539
rect 35805 21499 35863 21505
rect 34756 21440 35747 21468
rect 35820 21468 35848 21499
rect 36446 21496 36452 21548
rect 36504 21496 36510 21548
rect 37642 21536 37648 21548
rect 36556 21508 37648 21536
rect 36556 21468 36584 21508
rect 37642 21496 37648 21508
rect 37700 21496 37706 21548
rect 38930 21536 38936 21548
rect 37752 21508 38936 21536
rect 35820 21440 36584 21468
rect 36725 21471 36783 21477
rect 34756 21428 34762 21440
rect 36725 21437 36737 21471
rect 36771 21468 36783 21471
rect 37752 21468 37780 21508
rect 38930 21496 38936 21508
rect 38988 21496 38994 21548
rect 36771 21440 37780 21468
rect 36771 21437 36783 21440
rect 36725 21431 36783 21437
rect 37918 21428 37924 21480
rect 37976 21428 37982 21480
rect 38102 21428 38108 21480
rect 38160 21428 38166 21480
rect 30800 21372 31157 21400
rect 30800 21360 30806 21372
rect 32582 21360 32588 21412
rect 32640 21400 32646 21412
rect 35989 21403 36047 21409
rect 35989 21400 36001 21403
rect 32640 21372 36001 21400
rect 32640 21360 32646 21372
rect 35989 21369 36001 21372
rect 36035 21369 36047 21403
rect 35989 21363 36047 21369
rect 29604 21304 29776 21332
rect 30101 21335 30159 21341
rect 29604 21292 29610 21304
rect 30101 21301 30113 21335
rect 30147 21332 30159 21335
rect 30190 21332 30196 21344
rect 30147 21304 30196 21332
rect 30147 21301 30159 21304
rect 30101 21295 30159 21301
rect 30190 21292 30196 21304
rect 30248 21292 30254 21344
rect 31202 21292 31208 21344
rect 31260 21332 31266 21344
rect 31570 21332 31576 21344
rect 31260 21304 31576 21332
rect 31260 21292 31266 21304
rect 31570 21292 31576 21304
rect 31628 21292 31634 21344
rect 32306 21292 32312 21344
rect 32364 21332 32370 21344
rect 32861 21335 32919 21341
rect 32861 21332 32873 21335
rect 32364 21304 32873 21332
rect 32364 21292 32370 21304
rect 32861 21301 32873 21304
rect 32907 21301 32919 21335
rect 32861 21295 32919 21301
rect 33502 21292 33508 21344
rect 33560 21292 33566 21344
rect 33689 21335 33747 21341
rect 33689 21301 33701 21335
rect 33735 21332 33747 21335
rect 33962 21332 33968 21344
rect 33735 21304 33968 21332
rect 33735 21301 33747 21304
rect 33689 21295 33747 21301
rect 33962 21292 33968 21304
rect 34020 21292 34026 21344
rect 34054 21292 34060 21344
rect 34112 21332 34118 21344
rect 35161 21335 35219 21341
rect 35161 21332 35173 21335
rect 34112 21304 35173 21332
rect 34112 21292 34118 21304
rect 35161 21301 35173 21304
rect 35207 21301 35219 21335
rect 35161 21295 35219 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 13630 21088 13636 21140
rect 13688 21088 13694 21140
rect 22002 21128 22008 21140
rect 17788 21100 22008 21128
rect 12621 21063 12679 21069
rect 12621 21029 12633 21063
rect 12667 21060 12679 21063
rect 12667 21032 13216 21060
rect 12667 21029 12679 21032
rect 12621 21023 12679 21029
rect 13188 21001 13216 21032
rect 16758 21020 16764 21072
rect 16816 21060 16822 21072
rect 17589 21063 17647 21069
rect 17589 21060 17601 21063
rect 16816 21032 17601 21060
rect 16816 21020 16822 21032
rect 17589 21029 17601 21032
rect 17635 21029 17647 21063
rect 17589 21023 17647 21029
rect 13173 20995 13231 21001
rect 13173 20961 13185 20995
rect 13219 20961 13231 20995
rect 15286 20992 15292 21004
rect 13173 20955 13231 20961
rect 14660 20964 15292 20992
rect 11238 20884 11244 20936
rect 11296 20884 11302 20936
rect 12618 20884 12624 20936
rect 12676 20924 12682 20936
rect 14660 20933 14688 20964
rect 15286 20952 15292 20964
rect 15344 20952 15350 21004
rect 15470 20952 15476 21004
rect 15528 20952 15534 21004
rect 13265 20927 13323 20933
rect 13265 20924 13277 20927
rect 12676 20896 13277 20924
rect 12676 20884 12682 20896
rect 13265 20893 13277 20896
rect 13311 20893 13323 20927
rect 13265 20887 13323 20893
rect 14645 20927 14703 20933
rect 14645 20893 14657 20927
rect 14691 20893 14703 20927
rect 14645 20887 14703 20893
rect 15010 20884 15016 20936
rect 15068 20884 15074 20936
rect 15194 20884 15200 20936
rect 15252 20924 15258 20936
rect 15749 20927 15807 20933
rect 15749 20924 15761 20927
rect 15252 20896 15761 20924
rect 15252 20884 15258 20896
rect 15749 20893 15761 20896
rect 15795 20893 15807 20927
rect 15749 20887 15807 20893
rect 17589 20927 17647 20933
rect 17589 20893 17601 20927
rect 17635 20924 17647 20927
rect 17788 20924 17816 21100
rect 22002 21088 22008 21100
rect 22060 21088 22066 21140
rect 22554 21088 22560 21140
rect 22612 21088 22618 21140
rect 23750 21088 23756 21140
rect 23808 21128 23814 21140
rect 24581 21131 24639 21137
rect 24581 21128 24593 21131
rect 23808 21100 24593 21128
rect 23808 21088 23814 21100
rect 24581 21097 24593 21100
rect 24627 21097 24639 21131
rect 24581 21091 24639 21097
rect 25682 21088 25688 21140
rect 25740 21128 25746 21140
rect 25866 21128 25872 21140
rect 25740 21100 25872 21128
rect 25740 21088 25746 21100
rect 25866 21088 25872 21100
rect 25924 21128 25930 21140
rect 25961 21131 26019 21137
rect 25961 21128 25973 21131
rect 25924 21100 25973 21128
rect 25924 21088 25930 21100
rect 25961 21097 25973 21100
rect 26007 21097 26019 21131
rect 25961 21091 26019 21097
rect 26050 21088 26056 21140
rect 26108 21128 26114 21140
rect 26789 21131 26847 21137
rect 26789 21128 26801 21131
rect 26108 21100 26801 21128
rect 26108 21088 26114 21100
rect 26789 21097 26801 21100
rect 26835 21097 26847 21131
rect 26789 21091 26847 21097
rect 26970 21088 26976 21140
rect 27028 21128 27034 21140
rect 30558 21128 30564 21140
rect 27028 21100 30564 21128
rect 27028 21088 27034 21100
rect 30558 21088 30564 21100
rect 30616 21088 30622 21140
rect 37274 21128 37280 21140
rect 33520 21100 37280 21128
rect 19150 21060 19156 21072
rect 17880 21032 19156 21060
rect 17880 20933 17908 21032
rect 19150 21020 19156 21032
rect 19208 21020 19214 21072
rect 19242 21020 19248 21072
rect 19300 21060 19306 21072
rect 19978 21060 19984 21072
rect 19300 21032 19984 21060
rect 19300 21020 19306 21032
rect 19978 21020 19984 21032
rect 20036 21060 20042 21072
rect 20036 21032 20392 21060
rect 20036 21020 20042 21032
rect 18877 20995 18935 21001
rect 18877 20961 18889 20995
rect 18923 20992 18935 20995
rect 18923 20964 19840 20992
rect 18923 20961 18935 20964
rect 18877 20955 18935 20961
rect 17635 20896 17816 20924
rect 17865 20927 17923 20933
rect 17635 20893 17647 20896
rect 17589 20887 17647 20893
rect 17865 20893 17877 20927
rect 17911 20893 17923 20927
rect 17865 20887 17923 20893
rect 18325 20927 18383 20933
rect 18325 20893 18337 20927
rect 18371 20893 18383 20927
rect 18325 20887 18383 20893
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20924 18567 20927
rect 19242 20924 19248 20936
rect 18555 20896 19248 20924
rect 18555 20893 18567 20896
rect 18509 20887 18567 20893
rect 11508 20859 11566 20865
rect 11508 20825 11520 20859
rect 11554 20856 11566 20859
rect 14829 20859 14887 20865
rect 11554 20828 12434 20856
rect 11554 20825 11566 20828
rect 11508 20819 11566 20825
rect 12406 20788 12434 20828
rect 14829 20825 14841 20859
rect 14875 20856 14887 20859
rect 15562 20856 15568 20868
rect 14875 20828 15568 20856
rect 14875 20825 14887 20828
rect 14829 20819 14887 20825
rect 15562 20816 15568 20828
rect 15620 20816 15626 20868
rect 17126 20816 17132 20868
rect 17184 20816 17190 20868
rect 17880 20856 17908 20887
rect 17696 20828 17908 20856
rect 18340 20856 18368 20887
rect 19242 20884 19248 20896
rect 19300 20884 19306 20936
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19812 20933 19840 20964
rect 19521 20927 19579 20933
rect 19521 20924 19533 20927
rect 19392 20896 19533 20924
rect 19392 20884 19398 20896
rect 19521 20893 19533 20896
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20924 19855 20927
rect 20162 20924 20168 20936
rect 19843 20896 20168 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 20162 20884 20168 20896
rect 20220 20884 20226 20936
rect 20257 20927 20315 20933
rect 20257 20893 20269 20927
rect 20303 20893 20315 20927
rect 20364 20924 20392 21032
rect 20622 21020 20628 21072
rect 20680 21060 20686 21072
rect 23017 21063 23075 21069
rect 23017 21060 23029 21063
rect 20680 21032 23029 21060
rect 20680 21020 20686 21032
rect 23017 21029 23029 21032
rect 23063 21029 23075 21063
rect 23017 21023 23075 21029
rect 23290 21020 23296 21072
rect 23348 21060 23354 21072
rect 26145 21063 26203 21069
rect 23348 21032 26096 21060
rect 23348 21020 23354 21032
rect 20438 20952 20444 21004
rect 20496 20992 20502 21004
rect 20901 20995 20959 21001
rect 20901 20992 20913 20995
rect 20496 20964 20913 20992
rect 20496 20952 20502 20964
rect 20901 20961 20913 20964
rect 20947 20961 20959 20995
rect 20901 20955 20959 20961
rect 21913 20995 21971 21001
rect 21913 20961 21925 20995
rect 21959 20992 21971 20995
rect 22094 20992 22100 21004
rect 21959 20964 22100 20992
rect 21959 20961 21971 20964
rect 21913 20955 21971 20961
rect 22094 20952 22100 20964
rect 22152 20952 22158 21004
rect 22186 20952 22192 21004
rect 22244 20992 22250 21004
rect 22281 20995 22339 21001
rect 22281 20992 22293 20995
rect 22244 20964 22293 20992
rect 22244 20952 22250 20964
rect 22281 20961 22293 20964
rect 22327 20961 22339 20995
rect 22281 20955 22339 20961
rect 22373 20995 22431 21001
rect 22373 20961 22385 20995
rect 22419 20992 22431 20995
rect 22922 20992 22928 21004
rect 22419 20964 22928 20992
rect 22419 20961 22431 20964
rect 22373 20955 22431 20961
rect 22922 20952 22928 20964
rect 22980 20952 22986 21004
rect 23201 20995 23259 21001
rect 23201 20961 23213 20995
rect 23247 20992 23259 20995
rect 24210 20992 24216 21004
rect 23247 20964 24216 20992
rect 23247 20961 23259 20964
rect 23201 20955 23259 20961
rect 20533 20927 20591 20933
rect 20533 20924 20545 20927
rect 20364 20896 20545 20924
rect 20257 20887 20315 20893
rect 20533 20893 20545 20896
rect 20579 20893 20591 20927
rect 20533 20887 20591 20893
rect 20272 20856 20300 20887
rect 21082 20884 21088 20936
rect 21140 20924 21146 20936
rect 21450 20924 21456 20936
rect 21140 20896 21456 20924
rect 21140 20884 21146 20896
rect 21450 20884 21456 20896
rect 21508 20924 21514 20936
rect 23216 20924 23244 20955
rect 24210 20952 24216 20964
rect 24268 20952 24274 21004
rect 25222 20952 25228 21004
rect 25280 20952 25286 21004
rect 26068 20992 26096 21032
rect 26145 21029 26157 21063
rect 26191 21060 26203 21063
rect 27614 21060 27620 21072
rect 26191 21032 27620 21060
rect 26191 21029 26203 21032
rect 26145 21023 26203 21029
rect 27614 21020 27620 21032
rect 27672 21020 27678 21072
rect 29270 21020 29276 21072
rect 29328 21060 29334 21072
rect 31113 21063 31171 21069
rect 31113 21060 31125 21063
rect 29328 21032 31125 21060
rect 29328 21020 29334 21032
rect 31113 21029 31125 21032
rect 31159 21029 31171 21063
rect 31113 21023 31171 21029
rect 31956 21032 33272 21060
rect 26234 20992 26240 21004
rect 26068 20964 26240 20992
rect 26234 20952 26240 20964
rect 26292 20992 26298 21004
rect 26292 20964 27660 20992
rect 26292 20952 26298 20964
rect 21508 20896 23244 20924
rect 23293 20927 23351 20933
rect 21508 20884 21514 20896
rect 23293 20893 23305 20927
rect 23339 20893 23351 20927
rect 23293 20887 23351 20893
rect 22094 20856 22100 20868
rect 18340 20828 22100 20856
rect 17696 20788 17724 20828
rect 22094 20816 22100 20828
rect 22152 20816 22158 20868
rect 22646 20816 22652 20868
rect 22704 20856 22710 20868
rect 23308 20856 23336 20887
rect 23382 20884 23388 20936
rect 23440 20884 23446 20936
rect 23474 20884 23480 20936
rect 23532 20884 23538 20936
rect 26694 20924 26700 20936
rect 23584 20896 26700 20924
rect 23584 20856 23612 20896
rect 26694 20884 26700 20896
rect 26752 20884 26758 20936
rect 27632 20933 27660 20964
rect 27798 20952 27804 21004
rect 27856 20992 27862 21004
rect 28997 20995 29055 21001
rect 28997 20992 29009 20995
rect 27856 20964 29009 20992
rect 27856 20952 27862 20964
rect 28997 20961 29009 20964
rect 29043 20992 29055 20995
rect 29546 20992 29552 21004
rect 29043 20964 29552 20992
rect 29043 20961 29055 20964
rect 28997 20955 29055 20961
rect 29546 20952 29552 20964
rect 29604 20952 29610 21004
rect 30006 20952 30012 21004
rect 30064 20992 30070 21004
rect 30374 20992 30380 21004
rect 30064 20964 30236 20992
rect 30064 20952 30070 20964
rect 27433 20927 27491 20933
rect 27433 20924 27445 20927
rect 26896 20896 27445 20924
rect 22704 20828 23612 20856
rect 22704 20816 22710 20828
rect 24670 20816 24676 20868
rect 24728 20856 24734 20868
rect 25777 20859 25835 20865
rect 25777 20856 25789 20859
rect 24728 20828 25789 20856
rect 24728 20816 24734 20828
rect 25777 20825 25789 20828
rect 25823 20825 25835 20859
rect 25777 20819 25835 20825
rect 25866 20816 25872 20868
rect 25924 20856 25930 20868
rect 26605 20859 26663 20865
rect 26605 20856 26617 20859
rect 25924 20828 26617 20856
rect 25924 20816 25930 20828
rect 26605 20825 26617 20828
rect 26651 20825 26663 20859
rect 26605 20819 26663 20825
rect 12406 20760 17724 20788
rect 17770 20748 17776 20800
rect 17828 20748 17834 20800
rect 18506 20748 18512 20800
rect 18564 20748 18570 20800
rect 22922 20748 22928 20800
rect 22980 20788 22986 20800
rect 24854 20788 24860 20800
rect 22980 20760 24860 20788
rect 22980 20748 22986 20760
rect 24854 20748 24860 20760
rect 24912 20748 24918 20800
rect 24946 20748 24952 20800
rect 25004 20748 25010 20800
rect 25038 20748 25044 20800
rect 25096 20748 25102 20800
rect 25314 20748 25320 20800
rect 25372 20788 25378 20800
rect 25958 20788 25964 20800
rect 26016 20797 26022 20800
rect 26016 20791 26035 20797
rect 25372 20760 25964 20788
rect 25372 20748 25378 20760
rect 25958 20748 25964 20760
rect 26023 20757 26035 20791
rect 26016 20751 26035 20757
rect 26016 20748 26022 20751
rect 26694 20748 26700 20800
rect 26752 20788 26758 20800
rect 26805 20791 26863 20797
rect 26805 20788 26817 20791
rect 26752 20760 26817 20788
rect 26752 20748 26758 20760
rect 26805 20757 26817 20760
rect 26851 20788 26863 20791
rect 26896 20788 26924 20896
rect 27433 20893 27445 20896
rect 27479 20893 27491 20927
rect 27433 20887 27491 20893
rect 27617 20927 27675 20933
rect 27617 20893 27629 20927
rect 27663 20893 27675 20927
rect 27617 20887 27675 20893
rect 28687 20927 28745 20933
rect 28687 20893 28699 20927
rect 28733 20924 28745 20927
rect 28810 20924 28816 20936
rect 28733 20896 28816 20924
rect 28733 20893 28745 20896
rect 28687 20887 28745 20893
rect 28810 20884 28816 20896
rect 28868 20884 28874 20936
rect 29089 20927 29147 20933
rect 29089 20893 29101 20927
rect 29135 20924 29147 20927
rect 29454 20924 29460 20936
rect 29135 20896 29460 20924
rect 29135 20893 29147 20896
rect 29089 20887 29147 20893
rect 29454 20884 29460 20896
rect 29512 20884 29518 20936
rect 30101 20927 30159 20933
rect 30101 20893 30113 20927
rect 30147 20893 30159 20927
rect 30101 20887 30159 20893
rect 27338 20816 27344 20868
rect 27396 20856 27402 20868
rect 30116 20856 30144 20887
rect 27396 20828 30144 20856
rect 30208 20856 30236 20964
rect 30300 20964 30380 20992
rect 30300 20933 30328 20964
rect 30374 20952 30380 20964
rect 30432 20992 30438 21004
rect 31478 20992 31484 21004
rect 30432 20964 31484 20992
rect 30432 20952 30438 20964
rect 31478 20952 31484 20964
rect 31536 20952 31542 21004
rect 30285 20927 30343 20933
rect 30285 20893 30297 20927
rect 30331 20893 30343 20927
rect 30285 20887 30343 20893
rect 30469 20927 30527 20933
rect 30469 20893 30481 20927
rect 30515 20893 30527 20927
rect 30469 20887 30527 20893
rect 30377 20859 30435 20865
rect 30377 20856 30389 20859
rect 30208 20828 30389 20856
rect 27396 20816 27402 20828
rect 30377 20825 30389 20828
rect 30423 20825 30435 20859
rect 30484 20856 30512 20887
rect 30558 20884 30564 20936
rect 30616 20924 30622 20936
rect 31294 20924 31300 20936
rect 30616 20896 31300 20924
rect 30616 20884 30622 20896
rect 31294 20884 31300 20896
rect 31352 20924 31358 20936
rect 31389 20927 31447 20933
rect 31389 20924 31401 20927
rect 31352 20896 31401 20924
rect 31352 20884 31358 20896
rect 31389 20893 31401 20896
rect 31435 20893 31447 20927
rect 31956 20924 31984 21032
rect 32030 20952 32036 21004
rect 32088 20992 32094 21004
rect 32088 20964 32812 20992
rect 32088 20952 32094 20964
rect 32125 20927 32183 20933
rect 32125 20924 32137 20927
rect 31956 20896 32137 20924
rect 31389 20887 31447 20893
rect 32125 20893 32137 20896
rect 32171 20893 32183 20927
rect 32125 20887 32183 20893
rect 32214 20884 32220 20936
rect 32272 20884 32278 20936
rect 32306 20884 32312 20936
rect 32364 20884 32370 20936
rect 32401 20927 32459 20933
rect 32401 20893 32413 20927
rect 32447 20924 32459 20927
rect 32582 20924 32588 20936
rect 32447 20896 32588 20924
rect 32447 20893 32459 20896
rect 32401 20887 32459 20893
rect 32582 20884 32588 20896
rect 32640 20884 32646 20936
rect 30742 20856 30748 20868
rect 30484 20828 30748 20856
rect 30377 20819 30435 20825
rect 30742 20816 30748 20828
rect 30800 20816 30806 20868
rect 31110 20816 31116 20868
rect 31168 20816 31174 20868
rect 32674 20856 32680 20868
rect 31220 20828 32680 20856
rect 26851 20760 26924 20788
rect 26851 20757 26863 20760
rect 26805 20751 26863 20757
rect 26970 20748 26976 20800
rect 27028 20748 27034 20800
rect 27706 20748 27712 20800
rect 27764 20748 27770 20800
rect 28537 20791 28595 20797
rect 28537 20757 28549 20791
rect 28583 20788 28595 20791
rect 28810 20788 28816 20800
rect 28583 20760 28816 20788
rect 28583 20757 28595 20760
rect 28537 20751 28595 20757
rect 28810 20748 28816 20760
rect 28868 20748 28874 20800
rect 30653 20791 30711 20797
rect 30653 20757 30665 20791
rect 30699 20788 30711 20791
rect 31220 20788 31248 20828
rect 32674 20816 32680 20828
rect 32732 20816 32738 20868
rect 32784 20856 32812 20964
rect 33244 20936 33272 21032
rect 33318 21020 33324 21072
rect 33376 21060 33382 21072
rect 33413 21063 33471 21069
rect 33413 21060 33425 21063
rect 33376 21032 33425 21060
rect 33376 21020 33382 21032
rect 33413 21029 33425 21032
rect 33459 21029 33471 21063
rect 33413 21023 33471 21029
rect 33226 20884 33232 20936
rect 33284 20884 33290 20936
rect 33318 20884 33324 20936
rect 33376 20884 33382 20936
rect 33520 20933 33548 21100
rect 37274 21088 37280 21100
rect 37332 21088 37338 21140
rect 34057 21063 34115 21069
rect 34057 21029 34069 21063
rect 34103 21060 34115 21063
rect 34103 21032 35572 21060
rect 34103 21029 34115 21032
rect 34057 21023 34115 21029
rect 35544 21004 35572 21032
rect 34422 20952 34428 21004
rect 34480 20992 34486 21004
rect 34606 20992 34612 21004
rect 34480 20964 34612 20992
rect 34480 20952 34486 20964
rect 34606 20952 34612 20964
rect 34664 20952 34670 21004
rect 35526 20952 35532 21004
rect 35584 20952 35590 21004
rect 35805 20995 35863 21001
rect 35805 20961 35817 20995
rect 35851 20961 35863 20995
rect 35805 20955 35863 20961
rect 33505 20927 33563 20933
rect 33505 20893 33517 20927
rect 33551 20893 33563 20927
rect 33505 20887 33563 20893
rect 34054 20884 34060 20936
rect 34112 20884 34118 20936
rect 34146 20884 34152 20936
rect 34204 20924 34210 20936
rect 34333 20927 34391 20933
rect 34333 20924 34345 20927
rect 34204 20896 34345 20924
rect 34204 20884 34210 20896
rect 34333 20893 34345 20896
rect 34379 20893 34391 20927
rect 34333 20887 34391 20893
rect 35250 20884 35256 20936
rect 35308 20924 35314 20936
rect 35437 20927 35495 20933
rect 35437 20924 35449 20927
rect 35308 20896 35449 20924
rect 35308 20884 35314 20896
rect 35437 20893 35449 20896
rect 35483 20893 35495 20927
rect 35437 20887 35495 20893
rect 32784 20828 34284 20856
rect 30699 20760 31248 20788
rect 30699 20757 30711 20760
rect 30653 20751 30711 20757
rect 31294 20748 31300 20800
rect 31352 20748 31358 20800
rect 31938 20748 31944 20800
rect 31996 20748 32002 20800
rect 32950 20748 32956 20800
rect 33008 20788 33014 20800
rect 34256 20797 34284 20828
rect 35710 20816 35716 20868
rect 35768 20816 35774 20868
rect 35820 20856 35848 20955
rect 36265 20927 36323 20933
rect 36265 20893 36277 20927
rect 36311 20924 36323 20927
rect 36354 20924 36360 20936
rect 36311 20896 36360 20924
rect 36311 20893 36323 20896
rect 36265 20887 36323 20893
rect 36354 20884 36360 20896
rect 36412 20884 36418 20936
rect 36510 20859 36568 20865
rect 36510 20856 36522 20859
rect 35820 20828 36522 20856
rect 36510 20825 36522 20828
rect 36556 20825 36568 20859
rect 36510 20819 36568 20825
rect 33045 20791 33103 20797
rect 33045 20788 33057 20791
rect 33008 20760 33057 20788
rect 33008 20748 33014 20760
rect 33045 20757 33057 20760
rect 33091 20757 33103 20791
rect 33045 20751 33103 20757
rect 34241 20791 34299 20797
rect 34241 20757 34253 20791
rect 34287 20788 34299 20791
rect 35728 20788 35756 20816
rect 37645 20791 37703 20797
rect 37645 20788 37657 20791
rect 34287 20760 37657 20788
rect 34287 20757 34299 20760
rect 34241 20751 34299 20757
rect 37645 20757 37657 20760
rect 37691 20757 37703 20791
rect 37645 20751 37703 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 12434 20584 12440 20596
rect 12360 20556 12440 20584
rect 12360 20457 12388 20556
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 15010 20584 15016 20596
rect 12544 20556 15016 20584
rect 12544 20457 12572 20556
rect 15010 20544 15016 20556
rect 15068 20544 15074 20596
rect 15102 20544 15108 20596
rect 15160 20544 15166 20596
rect 16206 20544 16212 20596
rect 16264 20584 16270 20596
rect 16942 20584 16948 20596
rect 16264 20556 16948 20584
rect 16264 20544 16270 20556
rect 16942 20544 16948 20556
rect 17000 20544 17006 20596
rect 17034 20544 17040 20596
rect 17092 20584 17098 20596
rect 17092 20556 18460 20584
rect 17092 20544 17098 20556
rect 15120 20516 15148 20544
rect 15746 20516 15752 20528
rect 15028 20488 15148 20516
rect 15212 20488 15752 20516
rect 12345 20451 12403 20457
rect 12345 20417 12357 20451
rect 12391 20417 12403 20451
rect 12345 20411 12403 20417
rect 12529 20451 12587 20457
rect 12529 20417 12541 20451
rect 12575 20417 12587 20451
rect 15028 20448 15056 20488
rect 12529 20411 12587 20417
rect 13004 20420 15056 20448
rect 15105 20451 15163 20457
rect 13004 20389 13032 20420
rect 15105 20417 15117 20451
rect 15151 20448 15163 20451
rect 15212 20448 15240 20488
rect 15746 20476 15752 20488
rect 15804 20476 15810 20528
rect 16040 20488 17816 20516
rect 15151 20420 15240 20448
rect 15151 20417 15163 20420
rect 15105 20411 15163 20417
rect 15286 20408 15292 20460
rect 15344 20448 15350 20460
rect 16040 20457 16068 20488
rect 17788 20460 17816 20488
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15344 20420 16037 20448
rect 15344 20408 15350 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20417 16359 20451
rect 16301 20411 16359 20417
rect 12989 20383 13047 20389
rect 12989 20380 13001 20383
rect 12406 20352 13001 20380
rect 12406 20324 12434 20352
rect 12989 20349 13001 20352
rect 13035 20349 13047 20383
rect 12989 20343 13047 20349
rect 13262 20340 13268 20392
rect 13320 20340 13326 20392
rect 13446 20340 13452 20392
rect 13504 20380 13510 20392
rect 14369 20383 14427 20389
rect 14369 20380 14381 20383
rect 13504 20352 14381 20380
rect 13504 20340 13510 20352
rect 14369 20349 14381 20352
rect 14415 20349 14427 20383
rect 14369 20343 14427 20349
rect 15010 20340 15016 20392
rect 15068 20380 15074 20392
rect 15381 20383 15439 20389
rect 15381 20380 15393 20383
rect 15068 20352 15393 20380
rect 15068 20340 15074 20352
rect 15381 20349 15393 20352
rect 15427 20349 15439 20383
rect 15381 20343 15439 20349
rect 15470 20340 15476 20392
rect 15528 20340 15534 20392
rect 15562 20340 15568 20392
rect 15620 20380 15626 20392
rect 16316 20380 16344 20411
rect 16574 20408 16580 20460
rect 16632 20448 16638 20460
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 16632 20420 16865 20448
rect 16632 20408 16638 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 16942 20408 16948 20460
rect 17000 20448 17006 20460
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 17000 20420 17049 20448
rect 17000 20408 17006 20420
rect 17037 20417 17049 20420
rect 17083 20448 17095 20451
rect 17494 20448 17500 20460
rect 17083 20420 17500 20448
rect 17083 20417 17095 20420
rect 17037 20411 17095 20417
rect 17494 20408 17500 20420
rect 17552 20448 17558 20460
rect 17681 20451 17739 20457
rect 17681 20448 17693 20451
rect 17552 20420 17693 20448
rect 17552 20408 17558 20420
rect 17681 20417 17693 20420
rect 17727 20417 17739 20451
rect 17681 20411 17739 20417
rect 17770 20408 17776 20460
rect 17828 20408 17834 20460
rect 18432 20457 18460 20556
rect 20530 20544 20536 20596
rect 20588 20584 20594 20596
rect 20625 20587 20683 20593
rect 20625 20584 20637 20587
rect 20588 20556 20637 20584
rect 20588 20544 20594 20556
rect 20625 20553 20637 20556
rect 20671 20553 20683 20587
rect 20625 20547 20683 20553
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 21361 20587 21419 20593
rect 21361 20584 21373 20587
rect 20772 20556 21373 20584
rect 20772 20544 20778 20556
rect 21361 20553 21373 20556
rect 21407 20584 21419 20587
rect 22278 20584 22284 20596
rect 21407 20556 22284 20584
rect 21407 20553 21419 20556
rect 21361 20547 21419 20553
rect 22278 20544 22284 20556
rect 22336 20544 22342 20596
rect 23842 20544 23848 20596
rect 23900 20584 23906 20596
rect 24673 20587 24731 20593
rect 24673 20584 24685 20587
rect 23900 20556 24685 20584
rect 23900 20544 23906 20556
rect 24673 20553 24685 20556
rect 24719 20553 24731 20587
rect 24673 20547 24731 20553
rect 25222 20544 25228 20596
rect 25280 20584 25286 20596
rect 25593 20587 25651 20593
rect 25593 20584 25605 20587
rect 25280 20556 25605 20584
rect 25280 20544 25286 20556
rect 25593 20553 25605 20556
rect 25639 20553 25651 20587
rect 25593 20547 25651 20553
rect 25884 20556 28488 20584
rect 18506 20476 18512 20528
rect 18564 20516 18570 20528
rect 19153 20519 19211 20525
rect 19153 20516 19165 20519
rect 18564 20488 19165 20516
rect 18564 20476 18570 20488
rect 19153 20485 19165 20488
rect 19199 20485 19211 20519
rect 19153 20479 19211 20485
rect 24029 20519 24087 20525
rect 24029 20485 24041 20519
rect 24075 20516 24087 20519
rect 24075 20488 25176 20516
rect 24075 20485 24087 20488
rect 24029 20479 24087 20485
rect 18417 20451 18475 20457
rect 18417 20417 18429 20451
rect 18463 20417 18475 20451
rect 18417 20411 18475 20417
rect 18690 20408 18696 20460
rect 18748 20408 18754 20460
rect 18785 20451 18843 20457
rect 18785 20417 18797 20451
rect 18831 20448 18843 20451
rect 20254 20448 20260 20460
rect 18831 20420 20260 20448
rect 18831 20417 18843 20420
rect 18785 20411 18843 20417
rect 20254 20408 20260 20420
rect 20312 20408 20318 20460
rect 21266 20408 21272 20460
rect 21324 20408 21330 20460
rect 21450 20408 21456 20460
rect 21508 20448 21514 20460
rect 22186 20448 22192 20460
rect 21508 20420 22192 20448
rect 21508 20408 21514 20420
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 22462 20408 22468 20460
rect 22520 20408 22526 20460
rect 22738 20408 22744 20460
rect 22796 20408 22802 20460
rect 22830 20408 22836 20460
rect 22888 20408 22894 20460
rect 23106 20408 23112 20460
rect 23164 20408 23170 20460
rect 23290 20408 23296 20460
rect 23348 20408 23354 20460
rect 23658 20408 23664 20460
rect 23716 20448 23722 20460
rect 24489 20451 24547 20457
rect 24489 20448 24501 20451
rect 23716 20420 24501 20448
rect 23716 20408 23722 20420
rect 24489 20417 24501 20420
rect 24535 20417 24547 20451
rect 24489 20411 24547 20417
rect 17957 20383 18015 20389
rect 17957 20380 17969 20383
rect 15620 20352 17969 20380
rect 15620 20340 15626 20352
rect 17957 20349 17969 20352
rect 18003 20380 18015 20383
rect 20070 20380 20076 20392
rect 18003 20352 20076 20380
rect 18003 20349 18015 20352
rect 17957 20343 18015 20349
rect 20070 20340 20076 20352
rect 20128 20340 20134 20392
rect 20533 20383 20591 20389
rect 20533 20349 20545 20383
rect 20579 20349 20591 20383
rect 20533 20343 20591 20349
rect 20717 20383 20775 20389
rect 20717 20349 20729 20383
rect 20763 20380 20775 20383
rect 20898 20380 20904 20392
rect 20763 20352 20904 20380
rect 20763 20349 20775 20352
rect 20717 20343 20775 20349
rect 12342 20272 12348 20324
rect 12400 20284 12434 20324
rect 12400 20272 12406 20284
rect 13998 20272 14004 20324
rect 14056 20312 14062 20324
rect 17865 20315 17923 20321
rect 17865 20312 17877 20315
rect 14056 20284 17877 20312
rect 14056 20272 14062 20284
rect 17865 20281 17877 20284
rect 17911 20281 17923 20315
rect 17865 20275 17923 20281
rect 19426 20272 19432 20324
rect 19484 20272 19490 20324
rect 20162 20272 20168 20324
rect 20220 20272 20226 20324
rect 20548 20312 20576 20343
rect 20898 20340 20904 20352
rect 20956 20340 20962 20392
rect 20990 20340 20996 20392
rect 21048 20380 21054 20392
rect 25148 20389 25176 20488
rect 25406 20476 25412 20528
rect 25464 20516 25470 20528
rect 25884 20516 25912 20556
rect 25464 20488 25912 20516
rect 25464 20476 25470 20488
rect 25958 20476 25964 20528
rect 26016 20516 26022 20528
rect 26016 20488 26188 20516
rect 26016 20476 26022 20488
rect 25682 20408 25688 20460
rect 25740 20448 25746 20460
rect 26160 20457 26188 20488
rect 26234 20476 26240 20528
rect 26292 20516 26298 20528
rect 26421 20519 26479 20525
rect 26421 20516 26433 20519
rect 26292 20488 26433 20516
rect 26292 20476 26298 20488
rect 26421 20485 26433 20488
rect 26467 20485 26479 20519
rect 26421 20479 26479 20485
rect 28350 20476 28356 20528
rect 28408 20476 28414 20528
rect 28460 20516 28488 20556
rect 28534 20544 28540 20596
rect 28592 20544 28598 20596
rect 30742 20584 30748 20596
rect 28828 20556 30748 20584
rect 28828 20516 28856 20556
rect 30742 20544 30748 20556
rect 30800 20544 30806 20596
rect 30837 20587 30895 20593
rect 30837 20553 30849 20587
rect 30883 20584 30895 20587
rect 33318 20584 33324 20596
rect 30883 20556 33324 20584
rect 30883 20553 30895 20556
rect 30837 20547 30895 20553
rect 33318 20544 33324 20556
rect 33376 20544 33382 20596
rect 33778 20544 33784 20596
rect 33836 20584 33842 20596
rect 35802 20584 35808 20596
rect 33836 20556 35808 20584
rect 33836 20544 33842 20556
rect 35802 20544 35808 20556
rect 35860 20544 35866 20596
rect 36262 20544 36268 20596
rect 36320 20584 36326 20596
rect 36817 20587 36875 20593
rect 36817 20584 36829 20587
rect 36320 20556 36829 20584
rect 36320 20544 36326 20556
rect 36817 20553 36829 20556
rect 36863 20553 36875 20587
rect 36817 20547 36875 20553
rect 28460 20488 28856 20516
rect 28902 20476 28908 20528
rect 28960 20516 28966 20528
rect 28960 20488 30328 20516
rect 28960 20476 28966 20488
rect 26053 20451 26111 20457
rect 26053 20448 26065 20451
rect 25740 20420 26065 20448
rect 25740 20408 25746 20420
rect 26053 20417 26065 20420
rect 26099 20417 26111 20451
rect 26053 20411 26111 20417
rect 26146 20451 26204 20457
rect 26146 20417 26158 20451
rect 26192 20417 26204 20451
rect 26146 20411 26204 20417
rect 27062 20408 27068 20460
rect 27120 20448 27126 20460
rect 27893 20451 27951 20457
rect 27893 20448 27905 20451
rect 27120 20420 27905 20448
rect 27120 20408 27126 20420
rect 27893 20417 27905 20420
rect 27939 20448 27951 20451
rect 28629 20451 28687 20457
rect 27939 20420 28212 20448
rect 27939 20417 27951 20420
rect 27893 20411 27951 20417
rect 24397 20383 24455 20389
rect 21048 20352 23980 20380
rect 21048 20340 21054 20352
rect 20364 20284 20576 20312
rect 12437 20247 12495 20253
rect 12437 20213 12449 20247
rect 12483 20244 12495 20247
rect 14642 20244 14648 20256
rect 12483 20216 14648 20244
rect 12483 20213 12495 20216
rect 12437 20207 12495 20213
rect 14642 20204 14648 20216
rect 14700 20204 14706 20256
rect 15102 20204 15108 20256
rect 15160 20244 15166 20256
rect 15197 20247 15255 20253
rect 15197 20244 15209 20247
rect 15160 20216 15209 20244
rect 15160 20204 15166 20216
rect 15197 20213 15209 20216
rect 15243 20213 15255 20247
rect 15197 20207 15255 20213
rect 15286 20204 15292 20256
rect 15344 20204 15350 20256
rect 16022 20204 16028 20256
rect 16080 20204 16086 20256
rect 17218 20204 17224 20256
rect 17276 20204 17282 20256
rect 17494 20204 17500 20256
rect 17552 20244 17558 20256
rect 19334 20244 19340 20256
rect 17552 20216 19340 20244
rect 17552 20204 17558 20216
rect 19334 20204 19340 20216
rect 19392 20204 19398 20256
rect 20070 20204 20076 20256
rect 20128 20244 20134 20256
rect 20364 20244 20392 20284
rect 22094 20272 22100 20324
rect 22152 20272 22158 20324
rect 23952 20312 23980 20352
rect 24397 20349 24409 20383
rect 24443 20349 24455 20383
rect 24397 20343 24455 20349
rect 25133 20383 25191 20389
rect 25133 20349 25145 20383
rect 25179 20380 25191 20383
rect 25222 20380 25228 20392
rect 25179 20352 25228 20380
rect 25179 20349 25191 20352
rect 25133 20343 25191 20349
rect 24412 20312 24440 20343
rect 25222 20340 25228 20352
rect 25280 20380 25286 20392
rect 26326 20380 26332 20392
rect 25280 20352 26332 20380
rect 25280 20340 25286 20352
rect 26326 20340 26332 20352
rect 26384 20340 26390 20392
rect 26602 20340 26608 20392
rect 26660 20380 26666 20392
rect 27430 20380 27436 20392
rect 26660 20352 27436 20380
rect 26660 20340 26666 20352
rect 27430 20340 27436 20352
rect 27488 20340 27494 20392
rect 27617 20383 27675 20389
rect 27617 20349 27629 20383
rect 27663 20380 27675 20383
rect 27982 20380 27988 20392
rect 27663 20352 27988 20380
rect 27663 20349 27675 20352
rect 27617 20343 27675 20349
rect 27982 20340 27988 20352
rect 28040 20340 28046 20392
rect 28184 20380 28212 20420
rect 28629 20417 28641 20451
rect 28675 20448 28687 20451
rect 28718 20448 28724 20460
rect 28675 20420 28724 20448
rect 28675 20417 28687 20420
rect 28629 20411 28687 20417
rect 28718 20408 28724 20420
rect 28776 20408 28782 20460
rect 29270 20408 29276 20460
rect 29328 20408 29334 20460
rect 30300 20457 30328 20488
rect 30374 20476 30380 20528
rect 30432 20516 30438 20528
rect 30469 20519 30527 20525
rect 30469 20516 30481 20519
rect 30432 20488 30481 20516
rect 30432 20476 30438 20488
rect 30469 20485 30481 20488
rect 30515 20485 30527 20519
rect 36633 20519 36691 20525
rect 30469 20479 30527 20485
rect 33336 20488 34008 20516
rect 33336 20460 33364 20488
rect 30285 20451 30343 20457
rect 30285 20417 30297 20451
rect 30331 20417 30343 20451
rect 30285 20411 30343 20417
rect 30561 20451 30619 20457
rect 30561 20417 30573 20451
rect 30607 20417 30619 20451
rect 30561 20411 30619 20417
rect 28534 20380 28540 20392
rect 28184 20352 28540 20380
rect 28534 20340 28540 20352
rect 28592 20340 28598 20392
rect 29362 20340 29368 20392
rect 29420 20380 29426 20392
rect 29730 20380 29736 20392
rect 29420 20352 29736 20380
rect 29420 20340 29426 20352
rect 29730 20340 29736 20352
rect 29788 20340 29794 20392
rect 30576 20380 30604 20411
rect 30650 20408 30656 20460
rect 30708 20408 30714 20460
rect 30852 20420 32628 20448
rect 30742 20380 30748 20392
rect 30576 20352 30748 20380
rect 30742 20340 30748 20352
rect 30800 20340 30806 20392
rect 25501 20315 25559 20321
rect 25501 20312 25513 20315
rect 23952 20284 25513 20312
rect 25501 20281 25513 20284
rect 25547 20312 25559 20315
rect 26510 20312 26516 20324
rect 25547 20284 26516 20312
rect 25547 20281 25559 20284
rect 25501 20275 25559 20281
rect 26510 20272 26516 20284
rect 26568 20272 26574 20324
rect 27801 20315 27859 20321
rect 27801 20281 27813 20315
rect 27847 20312 27859 20315
rect 27890 20312 27896 20324
rect 27847 20284 27896 20312
rect 27847 20281 27859 20284
rect 27801 20275 27859 20281
rect 27890 20272 27896 20284
rect 27948 20272 27954 20324
rect 28350 20272 28356 20324
rect 28408 20272 28414 20324
rect 30852 20312 30880 20420
rect 31297 20383 31355 20389
rect 31297 20349 31309 20383
rect 31343 20380 31355 20383
rect 31386 20380 31392 20392
rect 31343 20352 31392 20380
rect 31343 20349 31355 20352
rect 31297 20343 31355 20349
rect 31386 20340 31392 20352
rect 31444 20340 31450 20392
rect 31846 20340 31852 20392
rect 31904 20380 31910 20392
rect 32493 20383 32551 20389
rect 32493 20380 32505 20383
rect 31904 20352 32505 20380
rect 31904 20340 31910 20352
rect 32493 20349 32505 20352
rect 32539 20349 32551 20383
rect 32493 20343 32551 20349
rect 29564 20284 30880 20312
rect 20128 20216 20392 20244
rect 20128 20204 20134 20216
rect 21266 20204 21272 20256
rect 21324 20244 21330 20256
rect 22186 20244 22192 20256
rect 21324 20216 22192 20244
rect 21324 20204 21330 20216
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 22462 20204 22468 20256
rect 22520 20244 22526 20256
rect 27433 20247 27491 20253
rect 27433 20244 27445 20247
rect 22520 20216 27445 20244
rect 22520 20204 22526 20216
rect 27433 20213 27445 20216
rect 27479 20213 27491 20247
rect 27433 20207 27491 20213
rect 27522 20204 27528 20256
rect 27580 20244 27586 20256
rect 29564 20244 29592 20284
rect 31478 20272 31484 20324
rect 31536 20312 31542 20324
rect 31573 20315 31631 20321
rect 31573 20312 31585 20315
rect 31536 20284 31585 20312
rect 31536 20272 31542 20284
rect 31573 20281 31585 20284
rect 31619 20281 31631 20315
rect 32398 20312 32404 20324
rect 31573 20275 31631 20281
rect 31680 20284 32404 20312
rect 27580 20216 29592 20244
rect 27580 20204 27586 20216
rect 29638 20204 29644 20256
rect 29696 20204 29702 20256
rect 30834 20204 30840 20256
rect 30892 20244 30898 20256
rect 31680 20244 31708 20284
rect 32398 20272 32404 20284
rect 32456 20272 32462 20324
rect 30892 20216 31708 20244
rect 31757 20247 31815 20253
rect 30892 20204 30898 20216
rect 31757 20213 31769 20247
rect 31803 20244 31815 20247
rect 31846 20244 31852 20256
rect 31803 20216 31852 20244
rect 31803 20213 31815 20216
rect 31757 20207 31815 20213
rect 31846 20204 31852 20216
rect 31904 20204 31910 20256
rect 32600 20244 32628 20420
rect 32674 20408 32680 20460
rect 32732 20408 32738 20460
rect 32769 20451 32827 20457
rect 32769 20417 32781 20451
rect 32815 20448 32827 20451
rect 33134 20448 33140 20460
rect 32815 20420 33140 20448
rect 32815 20417 32827 20420
rect 32769 20411 32827 20417
rect 33134 20408 33140 20420
rect 33192 20408 33198 20460
rect 33318 20408 33324 20460
rect 33376 20408 33382 20460
rect 33778 20408 33784 20460
rect 33836 20448 33842 20460
rect 33980 20457 34008 20488
rect 34072 20488 36584 20516
rect 34072 20460 34100 20488
rect 33873 20451 33931 20457
rect 33873 20448 33885 20451
rect 33836 20420 33885 20448
rect 33836 20408 33842 20420
rect 33873 20417 33885 20420
rect 33919 20417 33931 20451
rect 33873 20411 33931 20417
rect 33965 20451 34023 20457
rect 33965 20417 33977 20451
rect 34011 20417 34023 20451
rect 33965 20411 34023 20417
rect 34054 20408 34060 20460
rect 34112 20408 34118 20460
rect 34146 20408 34152 20460
rect 34204 20408 34210 20460
rect 34241 20451 34299 20457
rect 34241 20417 34253 20451
rect 34287 20417 34299 20451
rect 34241 20411 34299 20417
rect 32950 20340 32956 20392
rect 33008 20380 33014 20392
rect 33045 20383 33103 20389
rect 33045 20380 33057 20383
rect 33008 20352 33057 20380
rect 33008 20340 33014 20352
rect 33045 20349 33057 20352
rect 33091 20349 33103 20383
rect 33045 20343 33103 20349
rect 33226 20340 33232 20392
rect 33284 20380 33290 20392
rect 34256 20380 34284 20411
rect 34422 20408 34428 20460
rect 34480 20448 34486 20460
rect 34701 20451 34759 20457
rect 34701 20448 34713 20451
rect 34480 20420 34713 20448
rect 34480 20408 34486 20420
rect 34701 20417 34713 20420
rect 34747 20417 34759 20451
rect 34701 20411 34759 20417
rect 34974 20408 34980 20460
rect 35032 20408 35038 20460
rect 35618 20408 35624 20460
rect 35676 20448 35682 20460
rect 35805 20451 35863 20457
rect 35805 20448 35817 20451
rect 35676 20420 35817 20448
rect 35676 20408 35682 20420
rect 35805 20417 35817 20420
rect 35851 20417 35863 20451
rect 35805 20411 35863 20417
rect 35897 20451 35955 20457
rect 35897 20417 35909 20451
rect 35943 20417 35955 20451
rect 35897 20411 35955 20417
rect 33284 20352 34284 20380
rect 33284 20340 33290 20352
rect 35250 20340 35256 20392
rect 35308 20380 35314 20392
rect 35710 20380 35716 20392
rect 35308 20352 35716 20380
rect 35308 20340 35314 20352
rect 35710 20340 35716 20352
rect 35768 20340 35774 20392
rect 32858 20272 32864 20324
rect 32916 20312 32922 20324
rect 35912 20312 35940 20411
rect 35986 20408 35992 20460
rect 36044 20448 36050 20460
rect 36173 20451 36231 20457
rect 36173 20448 36185 20451
rect 36044 20420 36185 20448
rect 36044 20408 36050 20420
rect 36173 20417 36185 20420
rect 36219 20448 36231 20451
rect 36446 20448 36452 20460
rect 36219 20420 36452 20448
rect 36219 20417 36231 20420
rect 36173 20411 36231 20417
rect 36446 20408 36452 20420
rect 36504 20408 36510 20460
rect 36556 20448 36584 20488
rect 36633 20485 36645 20519
rect 36679 20516 36691 20519
rect 37366 20516 37372 20528
rect 36679 20488 37372 20516
rect 36679 20485 36691 20488
rect 36633 20479 36691 20485
rect 37366 20476 37372 20488
rect 37424 20476 37430 20528
rect 37921 20519 37979 20525
rect 37921 20485 37933 20519
rect 37967 20516 37979 20519
rect 38010 20516 38016 20528
rect 37967 20488 38016 20516
rect 37967 20485 37979 20488
rect 37921 20479 37979 20485
rect 36909 20451 36967 20457
rect 36909 20448 36921 20451
rect 36556 20420 36921 20448
rect 36909 20417 36921 20420
rect 36955 20417 36967 20451
rect 36909 20411 36967 20417
rect 37826 20408 37832 20460
rect 37884 20408 37890 20460
rect 36078 20340 36084 20392
rect 36136 20340 36142 20392
rect 37936 20312 37964 20479
rect 38010 20476 38016 20488
rect 38068 20476 38074 20528
rect 38102 20340 38108 20392
rect 38160 20340 38166 20392
rect 32916 20284 35940 20312
rect 36004 20284 37964 20312
rect 32916 20272 32922 20284
rect 32950 20244 32956 20256
rect 32600 20216 32956 20244
rect 32950 20204 32956 20216
rect 33008 20204 33014 20256
rect 33134 20204 33140 20256
rect 33192 20244 33198 20256
rect 33410 20244 33416 20256
rect 33192 20216 33416 20244
rect 33192 20204 33198 20216
rect 33410 20204 33416 20216
rect 33468 20204 33474 20256
rect 33689 20247 33747 20253
rect 33689 20213 33701 20247
rect 33735 20244 33747 20247
rect 34422 20244 34428 20256
rect 33735 20216 34428 20244
rect 33735 20213 33747 20216
rect 33689 20207 33747 20213
rect 34422 20204 34428 20216
rect 34480 20204 34486 20256
rect 35621 20247 35679 20253
rect 35621 20213 35633 20247
rect 35667 20244 35679 20247
rect 36004 20244 36032 20284
rect 35667 20216 36032 20244
rect 35667 20213 35679 20216
rect 35621 20207 35679 20213
rect 36170 20204 36176 20256
rect 36228 20244 36234 20256
rect 36633 20247 36691 20253
rect 36633 20244 36645 20247
rect 36228 20216 36645 20244
rect 36228 20204 36234 20216
rect 36633 20213 36645 20216
rect 36679 20213 36691 20247
rect 36633 20207 36691 20213
rect 37458 20204 37464 20256
rect 37516 20204 37522 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 12618 20000 12624 20052
rect 12676 20000 12682 20052
rect 13262 20000 13268 20052
rect 13320 20000 13326 20052
rect 14734 20000 14740 20052
rect 14792 20040 14798 20052
rect 15470 20040 15476 20052
rect 14792 20012 15476 20040
rect 14792 20000 14798 20012
rect 15470 20000 15476 20012
rect 15528 20000 15534 20052
rect 16574 20000 16580 20052
rect 16632 20000 16638 20052
rect 20438 20000 20444 20052
rect 20496 20000 20502 20052
rect 21913 20043 21971 20049
rect 21913 20009 21925 20043
rect 21959 20040 21971 20043
rect 23290 20040 23296 20052
rect 21959 20012 23296 20040
rect 21959 20009 21971 20012
rect 21913 20003 21971 20009
rect 23290 20000 23296 20012
rect 23348 20000 23354 20052
rect 23474 20000 23480 20052
rect 23532 20040 23538 20052
rect 23937 20043 23995 20049
rect 23937 20040 23949 20043
rect 23532 20012 23949 20040
rect 23532 20000 23538 20012
rect 23937 20009 23949 20012
rect 23983 20009 23995 20043
rect 23937 20003 23995 20009
rect 24026 20000 24032 20052
rect 24084 20040 24090 20052
rect 26602 20040 26608 20052
rect 24084 20012 26608 20040
rect 24084 20000 24090 20012
rect 26602 20000 26608 20012
rect 26660 20000 26666 20052
rect 31113 20043 31171 20049
rect 31113 20040 31125 20043
rect 26804 20012 31125 20040
rect 16022 19972 16028 19984
rect 13372 19944 16028 19972
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 12342 19836 12348 19848
rect 11296 19808 12348 19836
rect 11296 19796 11302 19808
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 11508 19771 11566 19777
rect 11508 19737 11520 19771
rect 11554 19768 11566 19771
rect 13372 19768 13400 19944
rect 16022 19932 16028 19944
rect 16080 19932 16086 19984
rect 16132 19944 18184 19972
rect 15286 19904 15292 19916
rect 13740 19876 15292 19904
rect 13740 19845 13768 19876
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 16132 19904 16160 19944
rect 15488 19876 16160 19904
rect 17221 19907 17279 19913
rect 13449 19839 13507 19845
rect 13449 19805 13461 19839
rect 13495 19805 13507 19839
rect 13449 19799 13507 19805
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19805 13783 19839
rect 13725 19799 13783 19805
rect 11554 19740 13400 19768
rect 13464 19768 13492 19799
rect 14734 19796 14740 19848
rect 14792 19796 14798 19848
rect 14829 19839 14887 19845
rect 14829 19805 14841 19839
rect 14875 19836 14887 19839
rect 14918 19836 14924 19848
rect 14875 19808 14924 19836
rect 14875 19805 14887 19808
rect 14829 19799 14887 19805
rect 14918 19796 14924 19808
rect 14976 19796 14982 19848
rect 15013 19839 15071 19845
rect 15013 19805 15025 19839
rect 15059 19805 15071 19839
rect 15013 19799 15071 19805
rect 14458 19768 14464 19780
rect 13464 19740 14464 19768
rect 11554 19737 11566 19740
rect 11508 19731 11566 19737
rect 14458 19728 14464 19740
rect 14516 19728 14522 19780
rect 15028 19768 15056 19799
rect 15102 19796 15108 19848
rect 15160 19836 15166 19848
rect 15488 19836 15516 19876
rect 17221 19873 17233 19907
rect 17267 19904 17279 19907
rect 18046 19904 18052 19916
rect 17267 19876 18052 19904
rect 17267 19873 17279 19876
rect 17221 19867 17279 19873
rect 18046 19864 18052 19876
rect 18104 19864 18110 19916
rect 18156 19904 18184 19944
rect 19978 19932 19984 19984
rect 20036 19932 20042 19984
rect 20254 19932 20260 19984
rect 20312 19972 20318 19984
rect 20806 19972 20812 19984
rect 20312 19944 20812 19972
rect 20312 19932 20318 19944
rect 20806 19932 20812 19944
rect 20864 19932 20870 19984
rect 20898 19932 20904 19984
rect 20956 19972 20962 19984
rect 21634 19972 21640 19984
rect 20956 19944 21640 19972
rect 20956 19932 20962 19944
rect 21634 19932 21640 19944
rect 21692 19972 21698 19984
rect 22738 19972 22744 19984
rect 21692 19944 22744 19972
rect 21692 19932 21698 19944
rect 21726 19904 21732 19916
rect 18156 19876 21732 19904
rect 21726 19864 21732 19876
rect 21784 19864 21790 19916
rect 15160 19808 15516 19836
rect 15565 19839 15623 19845
rect 15160 19796 15166 19808
rect 15565 19805 15577 19839
rect 15611 19836 15623 19839
rect 15654 19836 15660 19848
rect 15611 19808 15660 19836
rect 15611 19805 15623 19808
rect 15565 19799 15623 19805
rect 15654 19796 15660 19808
rect 15712 19796 15718 19848
rect 16666 19796 16672 19848
rect 16724 19836 16730 19848
rect 16945 19839 17003 19845
rect 16945 19836 16957 19839
rect 16724 19808 16957 19836
rect 16724 19796 16730 19808
rect 16945 19805 16957 19808
rect 16991 19805 17003 19839
rect 16945 19799 17003 19805
rect 17954 19796 17960 19848
rect 18012 19796 18018 19848
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19836 19671 19839
rect 20530 19836 20536 19848
rect 19659 19808 20536 19836
rect 19659 19805 19671 19808
rect 19613 19799 19671 19805
rect 20530 19796 20536 19808
rect 20588 19796 20594 19848
rect 20714 19796 20720 19848
rect 20772 19796 20778 19848
rect 20806 19796 20812 19848
rect 20864 19796 20870 19848
rect 20898 19796 20904 19848
rect 20956 19796 20962 19848
rect 21085 19839 21143 19845
rect 21085 19805 21097 19839
rect 21131 19805 21143 19839
rect 21928 19836 21956 19944
rect 22738 19932 22744 19944
rect 22796 19972 22802 19984
rect 22796 19944 24164 19972
rect 22796 19932 22802 19944
rect 22002 19864 22008 19916
rect 22060 19904 22066 19916
rect 22925 19907 22983 19913
rect 22060 19876 22416 19904
rect 22060 19864 22066 19876
rect 22388 19848 22416 19876
rect 22925 19873 22937 19907
rect 22971 19904 22983 19907
rect 22971 19876 23520 19904
rect 22971 19873 22983 19876
rect 22925 19867 22983 19873
rect 22097 19839 22155 19845
rect 22097 19836 22109 19839
rect 21928 19808 22109 19836
rect 21085 19799 21143 19805
rect 22097 19805 22109 19808
rect 22143 19805 22155 19839
rect 22097 19799 22155 19805
rect 15746 19768 15752 19780
rect 15028 19740 15752 19768
rect 15746 19728 15752 19740
rect 15804 19768 15810 19780
rect 15841 19771 15899 19777
rect 15841 19768 15853 19771
rect 15804 19740 15853 19768
rect 15804 19728 15810 19740
rect 15841 19737 15853 19740
rect 15887 19768 15899 19771
rect 15887 19740 18276 19768
rect 15887 19737 15899 19740
rect 15841 19731 15899 19737
rect 13633 19703 13691 19709
rect 13633 19669 13645 19703
rect 13679 19700 13691 19703
rect 14553 19703 14611 19709
rect 14553 19700 14565 19703
rect 13679 19672 14565 19700
rect 13679 19669 13691 19672
rect 13633 19663 13691 19669
rect 14553 19669 14565 19672
rect 14599 19669 14611 19703
rect 14553 19663 14611 19669
rect 15930 19660 15936 19712
rect 15988 19700 15994 19712
rect 16482 19700 16488 19712
rect 15988 19672 16488 19700
rect 15988 19660 15994 19672
rect 16482 19660 16488 19672
rect 16540 19700 16546 19712
rect 17037 19703 17095 19709
rect 17037 19700 17049 19703
rect 16540 19672 17049 19700
rect 16540 19660 16546 19672
rect 17037 19669 17049 19672
rect 17083 19700 17095 19703
rect 18046 19700 18052 19712
rect 17083 19672 18052 19700
rect 17083 19669 17095 19672
rect 17037 19663 17095 19669
rect 18046 19660 18052 19672
rect 18104 19660 18110 19712
rect 18248 19700 18276 19740
rect 18690 19728 18696 19780
rect 18748 19728 18754 19780
rect 18874 19728 18880 19780
rect 18932 19768 18938 19780
rect 19797 19771 19855 19777
rect 19797 19768 19809 19771
rect 18932 19740 19809 19768
rect 18932 19728 18938 19740
rect 19797 19737 19809 19740
rect 19843 19768 19855 19771
rect 21100 19768 21128 19799
rect 22186 19796 22192 19848
rect 22244 19796 22250 19848
rect 22370 19796 22376 19848
rect 22428 19796 22434 19848
rect 22465 19839 22523 19845
rect 22465 19805 22477 19839
rect 22511 19805 22523 19839
rect 22465 19799 22523 19805
rect 22278 19768 22284 19780
rect 19843 19740 22284 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 22278 19728 22284 19740
rect 22336 19728 22342 19780
rect 22480 19768 22508 19799
rect 23014 19796 23020 19848
rect 23072 19836 23078 19848
rect 23109 19839 23167 19845
rect 23109 19836 23121 19839
rect 23072 19808 23121 19836
rect 23072 19796 23078 19808
rect 23109 19805 23121 19808
rect 23155 19805 23167 19839
rect 23492 19836 23520 19876
rect 23566 19864 23572 19916
rect 23624 19904 23630 19916
rect 24029 19907 24087 19913
rect 24029 19904 24041 19907
rect 23624 19876 24041 19904
rect 23624 19864 23630 19876
rect 24029 19873 24041 19876
rect 24075 19873 24087 19907
rect 24136 19904 24164 19944
rect 24854 19932 24860 19984
rect 24912 19972 24918 19984
rect 25041 19975 25099 19981
rect 25041 19972 25053 19975
rect 24912 19944 25053 19972
rect 24912 19932 24918 19944
rect 25041 19941 25053 19944
rect 25087 19941 25099 19975
rect 25041 19935 25099 19941
rect 26237 19907 26295 19913
rect 26237 19904 26249 19907
rect 24136 19876 26249 19904
rect 24029 19867 24087 19873
rect 26237 19873 26249 19876
rect 26283 19873 26295 19907
rect 26237 19867 26295 19873
rect 23658 19836 23664 19848
rect 23492 19808 23664 19836
rect 23109 19799 23167 19805
rect 23658 19796 23664 19808
rect 23716 19796 23722 19848
rect 23753 19839 23811 19845
rect 23753 19805 23765 19839
rect 23799 19805 23811 19839
rect 23753 19799 23811 19805
rect 23845 19839 23903 19845
rect 23845 19805 23857 19839
rect 23891 19836 23903 19839
rect 24210 19836 24216 19848
rect 23891 19808 24216 19836
rect 23891 19805 23903 19808
rect 23845 19799 23903 19805
rect 22480 19740 23336 19768
rect 18892 19700 18920 19728
rect 18248 19672 18920 19700
rect 20346 19660 20352 19712
rect 20404 19700 20410 19712
rect 23014 19700 23020 19712
rect 20404 19672 23020 19700
rect 20404 19660 20410 19672
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 23308 19709 23336 19740
rect 23474 19728 23480 19780
rect 23532 19768 23538 19780
rect 23768 19768 23796 19799
rect 24210 19796 24216 19808
rect 24268 19796 24274 19848
rect 25317 19839 25375 19845
rect 25317 19805 25329 19839
rect 25363 19836 25375 19839
rect 25406 19836 25412 19848
rect 25363 19808 25412 19836
rect 25363 19805 25375 19808
rect 25317 19799 25375 19805
rect 25406 19796 25412 19808
rect 25464 19796 25470 19848
rect 26050 19836 26056 19848
rect 25516 19808 26056 19836
rect 25516 19777 25544 19808
rect 26050 19796 26056 19808
rect 26108 19836 26114 19848
rect 26145 19839 26203 19845
rect 26145 19836 26157 19839
rect 26108 19808 26157 19836
rect 26108 19796 26114 19808
rect 26145 19805 26157 19808
rect 26191 19805 26203 19839
rect 26145 19799 26203 19805
rect 26326 19796 26332 19848
rect 26384 19836 26390 19848
rect 26697 19839 26755 19845
rect 26697 19836 26709 19839
rect 26384 19808 26709 19836
rect 26384 19796 26390 19808
rect 26697 19805 26709 19808
rect 26743 19805 26755 19839
rect 26804 19836 26832 20012
rect 31113 20009 31125 20012
rect 31159 20040 31171 20043
rect 31294 20040 31300 20052
rect 31159 20012 31300 20040
rect 31159 20009 31171 20012
rect 31113 20003 31171 20009
rect 31294 20000 31300 20012
rect 31352 20040 31358 20052
rect 32030 20040 32036 20052
rect 31352 20012 32036 20040
rect 31352 20000 31358 20012
rect 32030 20000 32036 20012
rect 32088 20000 32094 20052
rect 32125 20043 32183 20049
rect 32125 20009 32137 20043
rect 32171 20040 32183 20043
rect 33226 20040 33232 20052
rect 32171 20012 33232 20040
rect 32171 20009 32183 20012
rect 32125 20003 32183 20009
rect 33226 20000 33232 20012
rect 33284 20000 33290 20052
rect 33965 20043 34023 20049
rect 33965 20009 33977 20043
rect 34011 20040 34023 20043
rect 34146 20040 34152 20052
rect 34011 20012 34152 20040
rect 34011 20009 34023 20012
rect 33965 20003 34023 20009
rect 34146 20000 34152 20012
rect 34204 20000 34210 20052
rect 34698 20000 34704 20052
rect 34756 20040 34762 20052
rect 34974 20040 34980 20052
rect 34756 20012 34980 20040
rect 34756 20000 34762 20012
rect 34974 20000 34980 20012
rect 35032 20000 35038 20052
rect 35250 20000 35256 20052
rect 35308 20040 35314 20052
rect 35526 20040 35532 20052
rect 35308 20012 35532 20040
rect 35308 20000 35314 20012
rect 35526 20000 35532 20012
rect 35584 20000 35590 20052
rect 27338 19932 27344 19984
rect 27396 19972 27402 19984
rect 28718 19972 28724 19984
rect 27396 19944 28724 19972
rect 27396 19932 27402 19944
rect 28718 19932 28724 19944
rect 28776 19972 28782 19984
rect 28994 19972 29000 19984
rect 28776 19944 29000 19972
rect 28776 19932 28782 19944
rect 28994 19932 29000 19944
rect 29052 19932 29058 19984
rect 31018 19932 31024 19984
rect 31076 19972 31082 19984
rect 31076 19944 33824 19972
rect 31076 19932 31082 19944
rect 26878 19864 26884 19916
rect 26936 19904 26942 19916
rect 26936 19876 27108 19904
rect 26936 19864 26942 19876
rect 26973 19839 27031 19845
rect 26973 19836 26985 19839
rect 26804 19808 26985 19836
rect 26697 19799 26755 19805
rect 26973 19805 26985 19808
rect 27019 19805 27031 19839
rect 27080 19836 27108 19876
rect 27246 19864 27252 19916
rect 27304 19904 27310 19916
rect 28629 19907 28687 19913
rect 28629 19904 28641 19907
rect 27304 19876 28641 19904
rect 27304 19864 27310 19876
rect 28629 19873 28641 19876
rect 28675 19873 28687 19907
rect 33042 19904 33048 19916
rect 28629 19867 28687 19873
rect 30760 19876 33048 19904
rect 27341 19839 27399 19845
rect 27341 19836 27353 19839
rect 27080 19808 27353 19836
rect 26973 19799 27031 19805
rect 27341 19805 27353 19808
rect 27387 19805 27399 19839
rect 27341 19799 27399 19805
rect 23532 19740 23796 19768
rect 25501 19771 25559 19777
rect 23532 19728 23538 19740
rect 25501 19737 25513 19771
rect 25547 19737 25559 19771
rect 25501 19731 25559 19737
rect 25593 19771 25651 19777
rect 25593 19737 25605 19771
rect 25639 19737 25651 19771
rect 26510 19768 26516 19780
rect 25593 19731 25651 19737
rect 26068 19740 26516 19768
rect 23293 19703 23351 19709
rect 23293 19669 23305 19703
rect 23339 19700 23351 19703
rect 23382 19700 23388 19712
rect 23339 19672 23388 19700
rect 23339 19669 23351 19672
rect 23293 19663 23351 19669
rect 23382 19660 23388 19672
rect 23440 19700 23446 19712
rect 24762 19700 24768 19712
rect 23440 19672 24768 19700
rect 23440 19660 23446 19672
rect 24762 19660 24768 19672
rect 24820 19660 24826 19712
rect 25608 19700 25636 19731
rect 26068 19712 26096 19740
rect 26510 19728 26516 19740
rect 26568 19728 26574 19780
rect 26712 19768 26740 19799
rect 27430 19796 27436 19848
rect 27488 19836 27494 19848
rect 28077 19839 28135 19845
rect 28077 19836 28089 19839
rect 27488 19808 28089 19836
rect 27488 19796 27494 19808
rect 28077 19805 28089 19808
rect 28123 19805 28135 19839
rect 28077 19799 28135 19805
rect 28261 19839 28319 19845
rect 28261 19805 28273 19839
rect 28307 19836 28319 19839
rect 28902 19836 28908 19848
rect 28307 19808 28908 19836
rect 28307 19805 28319 19808
rect 28261 19799 28319 19805
rect 28902 19796 28908 19808
rect 28960 19796 28966 19848
rect 29733 19839 29791 19845
rect 29733 19805 29745 19839
rect 29779 19836 29791 19839
rect 30760 19836 30788 19876
rect 33042 19864 33048 19876
rect 33100 19864 33106 19916
rect 33686 19904 33692 19916
rect 33152 19876 33692 19904
rect 32309 19839 32367 19845
rect 32309 19836 32321 19839
rect 29779 19808 30788 19836
rect 30852 19808 32321 19836
rect 29779 19805 29791 19808
rect 29733 19799 29791 19805
rect 26786 19768 26792 19780
rect 26712 19740 26792 19768
rect 26786 19728 26792 19740
rect 26844 19768 26850 19780
rect 27246 19768 27252 19780
rect 26844 19740 27252 19768
rect 26844 19728 26850 19740
rect 27246 19728 27252 19740
rect 27304 19728 27310 19780
rect 29454 19768 29460 19780
rect 28184 19740 29460 19768
rect 26050 19700 26056 19712
rect 25608 19672 26056 19700
rect 26050 19660 26056 19672
rect 26108 19660 26114 19712
rect 26234 19660 26240 19712
rect 26292 19700 26298 19712
rect 28184 19700 28212 19740
rect 29454 19728 29460 19740
rect 29512 19728 29518 19780
rect 29638 19728 29644 19780
rect 29696 19768 29702 19780
rect 29978 19771 30036 19777
rect 29978 19768 29990 19771
rect 29696 19740 29990 19768
rect 29696 19728 29702 19740
rect 29978 19737 29990 19740
rect 30024 19737 30036 19771
rect 29978 19731 30036 19737
rect 30466 19728 30472 19780
rect 30524 19768 30530 19780
rect 30852 19768 30880 19808
rect 32309 19805 32321 19808
rect 32355 19805 32367 19839
rect 32309 19799 32367 19805
rect 32401 19839 32459 19845
rect 32401 19805 32413 19839
rect 32447 19836 32459 19839
rect 33152 19836 33180 19876
rect 33686 19864 33692 19876
rect 33744 19864 33750 19916
rect 33796 19904 33824 19944
rect 34624 19944 35388 19972
rect 34624 19904 34652 19944
rect 33796 19876 34652 19904
rect 35360 19904 35388 19944
rect 35618 19932 35624 19984
rect 35676 19932 35682 19984
rect 36354 19904 36360 19916
rect 35360 19876 36360 19904
rect 36354 19864 36360 19876
rect 36412 19864 36418 19916
rect 32447 19808 33180 19836
rect 32447 19805 32459 19808
rect 32401 19799 32459 19805
rect 33226 19796 33232 19848
rect 33284 19836 33290 19848
rect 33413 19839 33471 19845
rect 33413 19836 33425 19839
rect 33284 19808 33425 19836
rect 33284 19796 33290 19808
rect 33413 19805 33425 19808
rect 33459 19805 33471 19839
rect 33413 19799 33471 19805
rect 33781 19839 33839 19845
rect 33781 19805 33793 19839
rect 33827 19836 33839 19839
rect 33870 19836 33876 19848
rect 33827 19808 33876 19836
rect 33827 19805 33839 19808
rect 33781 19799 33839 19805
rect 33870 19796 33876 19808
rect 33928 19796 33934 19848
rect 34790 19796 34796 19848
rect 34848 19836 34854 19848
rect 34977 19839 35035 19845
rect 34977 19836 34989 19839
rect 34848 19808 34989 19836
rect 34848 19796 34854 19808
rect 34977 19805 34989 19808
rect 35023 19805 35035 19839
rect 34977 19799 35035 19805
rect 35066 19796 35072 19848
rect 35124 19836 35130 19848
rect 35124 19808 35169 19836
rect 35124 19796 35130 19808
rect 35250 19796 35256 19848
rect 35308 19796 35314 19848
rect 35526 19845 35532 19848
rect 35483 19839 35532 19845
rect 35483 19805 35495 19839
rect 35529 19805 35532 19839
rect 35483 19799 35532 19805
rect 35526 19796 35532 19799
rect 35584 19836 35590 19848
rect 35802 19836 35808 19848
rect 35584 19808 35808 19836
rect 35584 19796 35590 19808
rect 35802 19796 35808 19808
rect 35860 19796 35866 19848
rect 35986 19796 35992 19848
rect 36044 19836 36050 19848
rect 36081 19839 36139 19845
rect 36081 19836 36093 19839
rect 36044 19808 36093 19836
rect 36044 19796 36050 19808
rect 36081 19805 36093 19808
rect 36127 19805 36139 19839
rect 36081 19799 36139 19805
rect 36170 19796 36176 19848
rect 36228 19836 36234 19848
rect 36265 19839 36323 19845
rect 36265 19836 36277 19839
rect 36228 19808 36277 19836
rect 36228 19796 36234 19808
rect 36265 19805 36277 19808
rect 36311 19805 36323 19839
rect 36265 19799 36323 19805
rect 36538 19796 36544 19848
rect 36596 19836 36602 19848
rect 36909 19839 36967 19845
rect 36909 19836 36921 19839
rect 36596 19808 36921 19836
rect 36596 19796 36602 19808
rect 36909 19805 36921 19808
rect 36955 19805 36967 19839
rect 36909 19799 36967 19805
rect 37176 19839 37234 19845
rect 37176 19805 37188 19839
rect 37222 19836 37234 19839
rect 37458 19836 37464 19848
rect 37222 19808 37464 19836
rect 37222 19805 37234 19808
rect 37176 19799 37234 19805
rect 37458 19796 37464 19808
rect 37516 19796 37522 19848
rect 30524 19740 30880 19768
rect 30524 19728 30530 19740
rect 32030 19728 32036 19780
rect 32088 19768 32094 19780
rect 32677 19771 32735 19777
rect 32677 19768 32689 19771
rect 32088 19740 32689 19768
rect 32088 19728 32094 19740
rect 32677 19737 32689 19740
rect 32723 19737 32735 19771
rect 32677 19731 32735 19737
rect 32769 19771 32827 19777
rect 32769 19737 32781 19771
rect 32815 19768 32827 19771
rect 33502 19768 33508 19780
rect 32815 19740 33508 19768
rect 32815 19737 32827 19740
rect 32769 19731 32827 19737
rect 33502 19728 33508 19740
rect 33560 19728 33566 19780
rect 33594 19728 33600 19780
rect 33652 19728 33658 19780
rect 33689 19771 33747 19777
rect 33689 19737 33701 19771
rect 33735 19737 33747 19771
rect 33689 19731 33747 19737
rect 35345 19771 35403 19777
rect 35345 19737 35357 19771
rect 35391 19768 35403 19771
rect 37826 19768 37832 19780
rect 35391 19740 37832 19768
rect 35391 19737 35403 19740
rect 35345 19731 35403 19737
rect 26292 19672 28212 19700
rect 26292 19660 26298 19672
rect 28258 19660 28264 19712
rect 28316 19660 28322 19712
rect 31294 19660 31300 19712
rect 31352 19700 31358 19712
rect 31662 19700 31668 19712
rect 31352 19672 31668 19700
rect 31352 19660 31358 19672
rect 31662 19660 31668 19672
rect 31720 19660 31726 19712
rect 32398 19660 32404 19712
rect 32456 19700 32462 19712
rect 33704 19700 33732 19731
rect 32456 19672 33732 19700
rect 32456 19660 32462 19672
rect 34882 19660 34888 19712
rect 34940 19700 34946 19712
rect 35360 19700 35388 19731
rect 37826 19728 37832 19740
rect 37884 19768 37890 19780
rect 37884 19740 38332 19768
rect 37884 19728 37890 19740
rect 34940 19672 35388 19700
rect 36357 19703 36415 19709
rect 34940 19660 34946 19672
rect 36357 19669 36369 19703
rect 36403 19700 36415 19703
rect 36630 19700 36636 19712
rect 36403 19672 36636 19700
rect 36403 19669 36415 19672
rect 36357 19663 36415 19669
rect 36630 19660 36636 19672
rect 36688 19660 36694 19712
rect 38304 19709 38332 19740
rect 38289 19703 38347 19709
rect 38289 19669 38301 19703
rect 38335 19669 38347 19703
rect 38289 19663 38347 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 13814 19456 13820 19508
rect 13872 19456 13878 19508
rect 14734 19456 14740 19508
rect 14792 19496 14798 19508
rect 15013 19499 15071 19505
rect 15013 19496 15025 19499
rect 14792 19468 15025 19496
rect 14792 19456 14798 19468
rect 15013 19465 15025 19468
rect 15059 19465 15071 19499
rect 20254 19496 20260 19508
rect 15013 19459 15071 19465
rect 16592 19468 20260 19496
rect 14921 19431 14979 19437
rect 14921 19397 14933 19431
rect 14967 19428 14979 19431
rect 16592 19428 16620 19468
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 20717 19499 20775 19505
rect 20717 19465 20729 19499
rect 20763 19496 20775 19499
rect 20806 19496 20812 19508
rect 20763 19468 20812 19496
rect 20763 19465 20775 19468
rect 20717 19459 20775 19465
rect 20806 19456 20812 19468
rect 20864 19456 20870 19508
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 21266 19496 21272 19508
rect 21223 19468 21272 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 23198 19456 23204 19508
rect 23256 19496 23262 19508
rect 24670 19496 24676 19508
rect 23256 19468 24676 19496
rect 23256 19456 23262 19468
rect 24670 19456 24676 19468
rect 24728 19456 24734 19508
rect 25038 19456 25044 19508
rect 25096 19496 25102 19508
rect 25409 19499 25467 19505
rect 25409 19496 25421 19499
rect 25096 19468 25421 19496
rect 25096 19456 25102 19468
rect 25409 19465 25421 19468
rect 25455 19465 25467 19499
rect 25409 19459 25467 19465
rect 26418 19456 26424 19508
rect 26476 19456 26482 19508
rect 27154 19456 27160 19508
rect 27212 19496 27218 19508
rect 27338 19496 27344 19508
rect 27212 19468 27344 19496
rect 27212 19456 27218 19468
rect 27338 19456 27344 19468
rect 27396 19456 27402 19508
rect 30006 19496 30012 19508
rect 27448 19468 30012 19496
rect 14967 19400 16620 19428
rect 14967 19397 14979 19400
rect 14921 19391 14979 19397
rect 16666 19388 16672 19440
rect 16724 19428 16730 19440
rect 19337 19431 19395 19437
rect 19337 19428 19349 19431
rect 16724 19400 19349 19428
rect 16724 19388 16730 19400
rect 19337 19397 19349 19400
rect 19383 19428 19395 19431
rect 19610 19428 19616 19440
rect 19383 19400 19616 19428
rect 19383 19397 19395 19400
rect 19337 19391 19395 19397
rect 19610 19388 19616 19400
rect 19668 19388 19674 19440
rect 20530 19388 20536 19440
rect 20588 19428 20594 19440
rect 22005 19431 22063 19437
rect 22005 19428 22017 19431
rect 20588 19400 22017 19428
rect 20588 19388 20594 19400
rect 22005 19397 22017 19400
rect 22051 19428 22063 19431
rect 22094 19428 22100 19440
rect 22051 19400 22100 19428
rect 22051 19397 22063 19400
rect 22005 19391 22063 19397
rect 22094 19388 22100 19400
rect 22152 19388 22158 19440
rect 24394 19388 24400 19440
rect 24452 19428 24458 19440
rect 26436 19428 26464 19456
rect 24452 19400 27200 19428
rect 24452 19388 24458 19400
rect 12342 19320 12348 19372
rect 12400 19360 12406 19372
rect 12437 19363 12495 19369
rect 12437 19360 12449 19363
rect 12400 19332 12449 19360
rect 12400 19320 12406 19332
rect 12437 19329 12449 19332
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 14826 19320 14832 19372
rect 14884 19320 14890 19372
rect 15841 19363 15899 19369
rect 15841 19329 15853 19363
rect 15887 19360 15899 19363
rect 16574 19360 16580 19372
rect 15887 19332 16580 19360
rect 15887 19329 15899 19332
rect 15841 19323 15899 19329
rect 16574 19320 16580 19332
rect 16632 19320 16638 19372
rect 17126 19320 17132 19372
rect 17184 19320 17190 19372
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19360 17371 19363
rect 17678 19360 17684 19372
rect 17359 19332 17684 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 17770 19320 17776 19372
rect 17828 19320 17834 19372
rect 18046 19320 18052 19372
rect 18104 19320 18110 19372
rect 18141 19363 18199 19369
rect 18141 19329 18153 19363
rect 18187 19360 18199 19363
rect 20622 19360 20628 19372
rect 18187 19332 20628 19360
rect 18187 19329 18199 19332
rect 18141 19323 18199 19329
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 21085 19363 21143 19369
rect 21085 19329 21097 19363
rect 21131 19360 21143 19363
rect 21450 19360 21456 19372
rect 21131 19332 21456 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 21450 19320 21456 19332
rect 21508 19320 21514 19372
rect 23293 19363 23351 19369
rect 23293 19329 23305 19363
rect 23339 19360 23351 19363
rect 23474 19360 23480 19372
rect 23339 19332 23480 19360
rect 23339 19329 23351 19332
rect 23293 19323 23351 19329
rect 23474 19320 23480 19332
rect 23532 19360 23538 19372
rect 23750 19360 23756 19372
rect 23532 19332 23756 19360
rect 23532 19320 23538 19332
rect 23750 19320 23756 19332
rect 23808 19320 23814 19372
rect 24302 19320 24308 19372
rect 24360 19320 24366 19372
rect 24486 19320 24492 19372
rect 24544 19320 24550 19372
rect 24581 19363 24639 19369
rect 24581 19329 24593 19363
rect 24627 19329 24639 19363
rect 24581 19323 24639 19329
rect 12713 19295 12771 19301
rect 12713 19261 12725 19295
rect 12759 19292 12771 19295
rect 14366 19292 14372 19304
rect 12759 19264 14372 19292
rect 12759 19261 12771 19264
rect 12713 19255 12771 19261
rect 14366 19252 14372 19264
rect 14424 19252 14430 19304
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 14553 19295 14611 19301
rect 14553 19292 14565 19295
rect 14516 19264 14565 19292
rect 14516 19252 14522 19264
rect 14553 19261 14565 19264
rect 14599 19261 14611 19295
rect 14553 19255 14611 19261
rect 15194 19252 15200 19304
rect 15252 19252 15258 19304
rect 15289 19295 15347 19301
rect 15289 19261 15301 19295
rect 15335 19292 15347 19295
rect 15378 19292 15384 19304
rect 15335 19264 15384 19292
rect 15335 19261 15347 19264
rect 15289 19255 15347 19261
rect 15378 19252 15384 19264
rect 15436 19252 15442 19304
rect 15933 19295 15991 19301
rect 15933 19261 15945 19295
rect 15979 19292 15991 19295
rect 17144 19292 17172 19320
rect 15979 19264 17172 19292
rect 15979 19261 15991 19264
rect 15933 19255 15991 19261
rect 13538 19184 13544 19236
rect 13596 19224 13602 19236
rect 15948 19224 15976 19255
rect 16758 19224 16764 19236
rect 13596 19196 15976 19224
rect 16040 19196 16764 19224
rect 13596 19184 13602 19196
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 15930 19156 15936 19168
rect 14516 19128 15936 19156
rect 14516 19116 14522 19128
rect 15930 19116 15936 19128
rect 15988 19116 15994 19168
rect 16040 19165 16068 19196
rect 16758 19184 16764 19196
rect 16816 19184 16822 19236
rect 17034 19184 17040 19236
rect 17092 19224 17098 19236
rect 17788 19233 17816 19320
rect 18064 19292 18092 19320
rect 18233 19295 18291 19301
rect 18233 19292 18245 19295
rect 18064 19264 18245 19292
rect 17129 19227 17187 19233
rect 17129 19224 17141 19227
rect 17092 19196 17141 19224
rect 17092 19184 17098 19196
rect 17129 19193 17141 19196
rect 17175 19193 17187 19227
rect 17129 19187 17187 19193
rect 17773 19227 17831 19233
rect 17773 19193 17785 19227
rect 17819 19193 17831 19227
rect 17773 19187 17831 19193
rect 16025 19159 16083 19165
rect 16025 19125 16037 19159
rect 16071 19125 16083 19159
rect 16025 19119 16083 19125
rect 16206 19116 16212 19168
rect 16264 19116 16270 19168
rect 18064 19156 18092 19264
rect 18233 19261 18245 19264
rect 18279 19261 18291 19295
rect 18233 19255 18291 19261
rect 18417 19295 18475 19301
rect 18417 19261 18429 19295
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 18432 19224 18460 19255
rect 18506 19252 18512 19304
rect 18564 19292 18570 19304
rect 19334 19292 19340 19304
rect 18564 19264 19340 19292
rect 18564 19252 18570 19264
rect 19334 19252 19340 19264
rect 19392 19292 19398 19304
rect 19429 19295 19487 19301
rect 19429 19292 19441 19295
rect 19392 19264 19441 19292
rect 19392 19252 19398 19264
rect 19429 19261 19441 19264
rect 19475 19261 19487 19295
rect 19429 19255 19487 19261
rect 19613 19295 19671 19301
rect 19613 19261 19625 19295
rect 19659 19292 19671 19295
rect 20990 19292 20996 19304
rect 19659 19264 20996 19292
rect 19659 19261 19671 19264
rect 19613 19255 19671 19261
rect 20990 19252 20996 19264
rect 21048 19252 21054 19304
rect 21361 19295 21419 19301
rect 21361 19261 21373 19295
rect 21407 19261 21419 19295
rect 21361 19255 21419 19261
rect 21082 19224 21088 19236
rect 18432 19196 21088 19224
rect 21082 19184 21088 19196
rect 21140 19184 21146 19236
rect 18506 19156 18512 19168
rect 18064 19128 18512 19156
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 18966 19116 18972 19168
rect 19024 19116 19030 19168
rect 21376 19156 21404 19255
rect 21726 19252 21732 19304
rect 21784 19292 21790 19304
rect 22002 19292 22008 19304
rect 21784 19264 22008 19292
rect 21784 19252 21790 19264
rect 22002 19252 22008 19264
rect 22060 19252 22066 19304
rect 23109 19295 23167 19301
rect 23109 19292 23121 19295
rect 22204 19264 23121 19292
rect 21910 19184 21916 19236
rect 21968 19224 21974 19236
rect 22204 19224 22232 19264
rect 23109 19261 23121 19264
rect 23155 19261 23167 19295
rect 23109 19255 23167 19261
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19292 23627 19295
rect 23934 19292 23940 19304
rect 23615 19264 23940 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 23934 19252 23940 19264
rect 23992 19252 23998 19304
rect 24210 19252 24216 19304
rect 24268 19292 24274 19304
rect 24596 19292 24624 19323
rect 24670 19320 24676 19372
rect 24728 19320 24734 19372
rect 24762 19320 24768 19372
rect 24820 19360 24826 19372
rect 25317 19363 25375 19369
rect 25317 19360 25329 19363
rect 24820 19332 25329 19360
rect 24820 19320 24826 19332
rect 25317 19329 25329 19332
rect 25363 19329 25375 19363
rect 25317 19323 25375 19329
rect 25958 19320 25964 19372
rect 26016 19320 26022 19372
rect 26142 19320 26148 19372
rect 26200 19320 26206 19372
rect 26234 19320 26240 19372
rect 26292 19320 26298 19372
rect 26381 19363 26439 19369
rect 26381 19329 26393 19363
rect 26427 19360 26439 19363
rect 26878 19360 26884 19372
rect 26427 19332 26884 19360
rect 26427 19329 26439 19332
rect 26381 19323 26439 19329
rect 26878 19320 26884 19332
rect 26936 19320 26942 19372
rect 27172 19369 27200 19400
rect 27157 19363 27215 19369
rect 27157 19329 27169 19363
rect 27203 19329 27215 19363
rect 27157 19323 27215 19329
rect 27246 19320 27252 19372
rect 27304 19360 27310 19372
rect 27448 19369 27476 19468
rect 30006 19456 30012 19468
rect 30064 19456 30070 19508
rect 31018 19496 31024 19508
rect 30208 19468 31024 19496
rect 28718 19388 28724 19440
rect 28776 19428 28782 19440
rect 28813 19431 28871 19437
rect 28813 19428 28825 19431
rect 28776 19400 28825 19428
rect 28776 19388 28782 19400
rect 28813 19397 28825 19400
rect 28859 19397 28871 19431
rect 28813 19391 28871 19397
rect 28994 19388 29000 19440
rect 29052 19388 29058 19440
rect 29454 19388 29460 19440
rect 29512 19428 29518 19440
rect 30208 19428 30236 19468
rect 31018 19456 31024 19468
rect 31076 19456 31082 19508
rect 31110 19456 31116 19508
rect 31168 19496 31174 19508
rect 31481 19499 31539 19505
rect 31481 19496 31493 19499
rect 31168 19468 31493 19496
rect 31168 19456 31174 19468
rect 31481 19465 31493 19468
rect 31527 19465 31539 19499
rect 31481 19459 31539 19465
rect 32858 19456 32864 19508
rect 32916 19456 32922 19508
rect 33318 19496 33324 19508
rect 33152 19468 33324 19496
rect 33152 19428 33180 19468
rect 33318 19456 33324 19468
rect 33376 19456 33382 19508
rect 35345 19499 35403 19505
rect 35345 19496 35357 19499
rect 33980 19468 35357 19496
rect 29512 19400 30236 19428
rect 29512 19388 29518 19400
rect 27341 19363 27399 19369
rect 27341 19360 27353 19363
rect 27304 19332 27353 19360
rect 27304 19320 27310 19332
rect 27341 19329 27353 19332
rect 27387 19329 27399 19363
rect 27341 19323 27399 19329
rect 27433 19363 27491 19369
rect 27433 19329 27445 19363
rect 27479 19329 27491 19363
rect 27433 19323 27491 19329
rect 27553 19363 27611 19369
rect 27553 19329 27565 19363
rect 27599 19360 27611 19363
rect 27599 19329 27614 19360
rect 27553 19323 27614 19329
rect 26896 19292 26924 19320
rect 27586 19304 27614 19323
rect 27890 19320 27896 19372
rect 27948 19360 27954 19372
rect 27948 19332 29868 19360
rect 27948 19320 27954 19332
rect 27062 19292 27068 19304
rect 24268 19264 26832 19292
rect 26896 19264 27068 19292
rect 24268 19252 24274 19264
rect 21968 19196 22232 19224
rect 21968 19184 21974 19196
rect 22370 19184 22376 19236
rect 22428 19224 22434 19236
rect 25866 19224 25872 19236
rect 22428 19196 25872 19224
rect 22428 19184 22434 19196
rect 25866 19184 25872 19196
rect 25924 19184 25930 19236
rect 22465 19159 22523 19165
rect 22465 19156 22477 19159
rect 21376 19128 22477 19156
rect 22465 19125 22477 19128
rect 22511 19125 22523 19159
rect 22465 19119 22523 19125
rect 23474 19116 23480 19168
rect 23532 19116 23538 19168
rect 24857 19159 24915 19165
rect 24857 19125 24869 19159
rect 24903 19156 24915 19159
rect 25130 19156 25136 19168
rect 24903 19128 25136 19156
rect 24903 19125 24915 19128
rect 24857 19119 24915 19125
rect 25130 19116 25136 19128
rect 25188 19116 25194 19168
rect 26418 19116 26424 19168
rect 26476 19156 26482 19168
rect 26513 19159 26571 19165
rect 26513 19156 26525 19159
rect 26476 19128 26525 19156
rect 26476 19116 26482 19128
rect 26513 19125 26525 19128
rect 26559 19125 26571 19159
rect 26804 19156 26832 19264
rect 27062 19252 27068 19264
rect 27120 19252 27126 19304
rect 27586 19264 27620 19304
rect 27614 19252 27620 19264
rect 27672 19252 27678 19304
rect 29089 19295 29147 19301
rect 29089 19261 29101 19295
rect 29135 19292 29147 19295
rect 29362 19292 29368 19304
rect 29135 19264 29368 19292
rect 29135 19261 29147 19264
rect 29089 19255 29147 19261
rect 29362 19252 29368 19264
rect 29420 19292 29426 19304
rect 29638 19292 29644 19304
rect 29420 19264 29644 19292
rect 29420 19252 29426 19264
rect 29638 19252 29644 19264
rect 29696 19252 29702 19304
rect 26878 19184 26884 19236
rect 26936 19224 26942 19236
rect 27709 19227 27767 19233
rect 27709 19224 27721 19227
rect 26936 19196 27721 19224
rect 26936 19184 26942 19196
rect 27709 19193 27721 19196
rect 27755 19193 27767 19227
rect 29733 19227 29791 19233
rect 29733 19224 29745 19227
rect 27709 19187 27767 19193
rect 27816 19196 29745 19224
rect 27816 19156 27844 19196
rect 29733 19193 29745 19196
rect 29779 19193 29791 19227
rect 29840 19224 29868 19332
rect 29914 19320 29920 19372
rect 29972 19320 29978 19372
rect 30208 19369 30236 19400
rect 30944 19400 33180 19428
rect 30193 19363 30251 19369
rect 30193 19329 30205 19363
rect 30239 19329 30251 19363
rect 30193 19323 30251 19329
rect 30834 19320 30840 19372
rect 30892 19320 30898 19372
rect 30944 19369 30972 19400
rect 33226 19388 33232 19440
rect 33284 19428 33290 19440
rect 33980 19437 34008 19468
rect 35345 19465 35357 19468
rect 35391 19465 35403 19499
rect 35345 19459 35403 19465
rect 33505 19431 33563 19437
rect 33505 19428 33517 19431
rect 33284 19400 33517 19428
rect 33284 19388 33290 19400
rect 33505 19397 33517 19400
rect 33551 19397 33563 19431
rect 33505 19391 33563 19397
rect 33965 19431 34023 19437
rect 33965 19397 33977 19431
rect 34011 19397 34023 19431
rect 33965 19391 34023 19397
rect 34054 19388 34060 19440
rect 34112 19428 34118 19440
rect 34112 19400 34284 19428
rect 34112 19388 34118 19400
rect 30929 19363 30987 19369
rect 30929 19329 30941 19363
rect 30975 19329 30987 19363
rect 30929 19323 30987 19329
rect 31018 19320 31024 19372
rect 31076 19360 31082 19372
rect 31113 19363 31171 19369
rect 31113 19360 31125 19363
rect 31076 19332 31125 19360
rect 31076 19320 31082 19332
rect 31113 19329 31125 19332
rect 31159 19329 31171 19363
rect 31113 19323 31171 19329
rect 31201 19363 31259 19369
rect 31201 19329 31213 19363
rect 31247 19329 31259 19363
rect 31201 19323 31259 19329
rect 31343 19363 31401 19369
rect 31343 19329 31355 19363
rect 31389 19360 31401 19363
rect 31662 19360 31668 19372
rect 31389 19332 31668 19360
rect 31389 19329 31401 19332
rect 31343 19323 31401 19329
rect 30101 19295 30159 19301
rect 30101 19261 30113 19295
rect 30147 19292 30159 19295
rect 30282 19292 30288 19304
rect 30147 19264 30288 19292
rect 30147 19261 30159 19264
rect 30101 19255 30159 19261
rect 30282 19252 30288 19264
rect 30340 19252 30346 19304
rect 30852 19292 30880 19320
rect 31220 19292 31248 19323
rect 31662 19320 31668 19332
rect 31720 19320 31726 19372
rect 32858 19320 32864 19372
rect 32916 19360 32922 19372
rect 33137 19363 33195 19369
rect 33137 19360 33149 19363
rect 32916 19332 33149 19360
rect 32916 19320 32922 19332
rect 33137 19329 33149 19332
rect 33183 19360 33195 19363
rect 33686 19360 33692 19372
rect 33183 19332 33692 19360
rect 33183 19329 33195 19332
rect 33137 19323 33195 19329
rect 33686 19320 33692 19332
rect 33744 19320 33750 19372
rect 33870 19320 33876 19372
rect 33928 19360 33934 19372
rect 34256 19369 34284 19400
rect 34606 19388 34612 19440
rect 34664 19428 34670 19440
rect 35069 19431 35127 19437
rect 35069 19428 35081 19431
rect 34664 19400 35081 19428
rect 34664 19388 34670 19400
rect 35069 19397 35081 19400
rect 35115 19397 35127 19431
rect 35069 19391 35127 19397
rect 36354 19388 36360 19440
rect 36412 19428 36418 19440
rect 38105 19431 38163 19437
rect 36412 19400 36952 19428
rect 36412 19388 36418 19400
rect 34149 19363 34207 19369
rect 34149 19360 34161 19363
rect 33928 19332 34161 19360
rect 33928 19320 33934 19332
rect 34149 19329 34161 19332
rect 34195 19329 34207 19363
rect 34149 19323 34207 19329
rect 34241 19363 34299 19369
rect 34241 19329 34253 19363
rect 34287 19329 34299 19363
rect 34241 19323 34299 19329
rect 34514 19320 34520 19372
rect 34572 19360 34578 19372
rect 34882 19369 34888 19372
rect 34701 19363 34759 19369
rect 34701 19360 34713 19363
rect 34572 19332 34713 19360
rect 34572 19320 34578 19332
rect 34701 19329 34713 19332
rect 34747 19329 34759 19363
rect 34701 19323 34759 19329
rect 34849 19363 34888 19369
rect 34849 19329 34861 19363
rect 34849 19323 34888 19329
rect 34882 19320 34888 19323
rect 34940 19320 34946 19372
rect 34975 19320 34981 19372
rect 35033 19360 35039 19372
rect 35207 19363 35265 19369
rect 35033 19332 35077 19360
rect 35033 19320 35039 19332
rect 35207 19329 35219 19363
rect 35253 19360 35265 19363
rect 35342 19360 35348 19372
rect 35253 19332 35348 19360
rect 35253 19329 35265 19332
rect 35207 19323 35265 19329
rect 35342 19320 35348 19332
rect 35400 19320 35406 19372
rect 35802 19320 35808 19372
rect 35860 19320 35866 19372
rect 36081 19363 36139 19369
rect 36081 19360 36093 19363
rect 35912 19332 36093 19360
rect 30852 19264 31248 19292
rect 33042 19252 33048 19304
rect 33100 19252 33106 19304
rect 33413 19295 33471 19301
rect 33413 19261 33425 19295
rect 33459 19261 33471 19295
rect 33413 19255 33471 19261
rect 30466 19224 30472 19236
rect 29840 19196 30472 19224
rect 29733 19187 29791 19193
rect 30466 19184 30472 19196
rect 30524 19184 30530 19236
rect 31754 19184 31760 19236
rect 31812 19224 31818 19236
rect 32214 19224 32220 19236
rect 31812 19196 32220 19224
rect 31812 19184 31818 19196
rect 32214 19184 32220 19196
rect 32272 19184 32278 19236
rect 32490 19184 32496 19236
rect 32548 19224 32554 19236
rect 33428 19224 33456 19255
rect 33502 19252 33508 19304
rect 33560 19292 33566 19304
rect 35912 19292 35940 19332
rect 36081 19329 36093 19332
rect 36127 19329 36139 19363
rect 36081 19323 36139 19329
rect 36722 19320 36728 19372
rect 36780 19320 36786 19372
rect 36924 19369 36952 19400
rect 38105 19397 38117 19431
rect 38151 19428 38163 19431
rect 39022 19428 39028 19440
rect 38151 19400 39028 19428
rect 38151 19397 38163 19400
rect 38105 19391 38163 19397
rect 39022 19388 39028 19400
rect 39080 19388 39086 19440
rect 36909 19363 36967 19369
rect 36909 19329 36921 19363
rect 36955 19360 36967 19363
rect 37550 19360 37556 19372
rect 36955 19332 37556 19360
rect 36955 19329 36967 19332
rect 36909 19323 36967 19329
rect 37550 19320 37556 19332
rect 37608 19320 37614 19372
rect 37829 19363 37887 19369
rect 37829 19329 37841 19363
rect 37875 19360 37887 19363
rect 37918 19360 37924 19372
rect 37875 19332 37924 19360
rect 37875 19329 37887 19332
rect 37829 19323 37887 19329
rect 37918 19320 37924 19332
rect 37976 19320 37982 19372
rect 33560 19264 35940 19292
rect 33560 19252 33566 19264
rect 34808 19236 34836 19264
rect 36814 19252 36820 19304
rect 36872 19252 36878 19304
rect 32548 19196 33456 19224
rect 33965 19227 34023 19233
rect 32548 19184 32554 19196
rect 33965 19193 33977 19227
rect 34011 19224 34023 19227
rect 34054 19224 34060 19236
rect 34011 19196 34060 19224
rect 34011 19193 34023 19196
rect 33965 19187 34023 19193
rect 34054 19184 34060 19196
rect 34112 19184 34118 19236
rect 34790 19184 34796 19236
rect 34848 19184 34854 19236
rect 26804 19128 27844 19156
rect 28537 19159 28595 19165
rect 26513 19119 26571 19125
rect 28537 19125 28549 19159
rect 28583 19156 28595 19159
rect 28718 19156 28724 19168
rect 28583 19128 28724 19156
rect 28583 19125 28595 19128
rect 28537 19119 28595 19125
rect 28718 19116 28724 19128
rect 28776 19116 28782 19168
rect 30006 19116 30012 19168
rect 30064 19156 30070 19168
rect 30742 19156 30748 19168
rect 30064 19128 30748 19156
rect 30064 19116 30070 19128
rect 30742 19116 30748 19128
rect 30800 19116 30806 19168
rect 31018 19116 31024 19168
rect 31076 19156 31082 19168
rect 31662 19156 31668 19168
rect 31076 19128 31668 19156
rect 31076 19116 31082 19128
rect 31662 19116 31668 19128
rect 31720 19156 31726 19168
rect 34974 19156 34980 19168
rect 31720 19128 34980 19156
rect 31720 19116 31726 19128
rect 34974 19116 34980 19128
rect 35032 19116 35038 19168
rect 35158 19116 35164 19168
rect 35216 19156 35222 19168
rect 35618 19156 35624 19168
rect 35216 19128 35624 19156
rect 35216 19116 35222 19128
rect 35618 19116 35624 19128
rect 35676 19116 35682 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 12897 18955 12955 18961
rect 12897 18921 12909 18955
rect 12943 18952 12955 18955
rect 13538 18952 13544 18964
rect 12943 18924 13544 18952
rect 12943 18921 12955 18924
rect 12897 18915 12955 18921
rect 13538 18912 13544 18924
rect 13596 18912 13602 18964
rect 13633 18955 13691 18961
rect 13633 18921 13645 18955
rect 13679 18952 13691 18955
rect 13679 18924 18644 18952
rect 13679 18921 13691 18924
rect 13633 18915 13691 18921
rect 13648 18816 13676 18915
rect 14734 18884 14740 18896
rect 14568 18856 14740 18884
rect 13096 18788 13676 18816
rect 12894 18708 12900 18760
rect 12952 18708 12958 18760
rect 13096 18757 13124 18788
rect 14090 18776 14096 18828
rect 14148 18816 14154 18828
rect 14568 18825 14596 18856
rect 14734 18844 14740 18856
rect 14792 18844 14798 18896
rect 14826 18844 14832 18896
rect 14884 18884 14890 18896
rect 15565 18887 15623 18893
rect 15565 18884 15577 18887
rect 14884 18856 15577 18884
rect 14884 18844 14890 18856
rect 15565 18853 15577 18856
rect 15611 18853 15623 18887
rect 15565 18847 15623 18853
rect 14553 18819 14611 18825
rect 14553 18816 14565 18819
rect 14148 18788 14565 18816
rect 14148 18776 14154 18788
rect 14553 18785 14565 18788
rect 14599 18785 14611 18819
rect 15470 18816 15476 18828
rect 14553 18779 14611 18785
rect 14752 18788 15476 18816
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18717 13139 18751
rect 13081 18711 13139 18717
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18748 13599 18751
rect 14458 18748 14464 18760
rect 13587 18720 14464 18748
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 14642 18708 14648 18760
rect 14700 18748 14706 18760
rect 14752 18757 14780 18788
rect 15470 18776 15476 18788
rect 15528 18776 15534 18828
rect 16206 18776 16212 18828
rect 16264 18776 16270 18828
rect 16669 18819 16727 18825
rect 16669 18785 16681 18819
rect 16715 18816 16727 18819
rect 17218 18816 17224 18828
rect 16715 18788 17224 18816
rect 16715 18785 16727 18788
rect 16669 18779 16727 18785
rect 17218 18776 17224 18788
rect 17276 18776 17282 18828
rect 18616 18825 18644 18924
rect 20898 18912 20904 18964
rect 20956 18952 20962 18964
rect 21177 18955 21235 18961
rect 21177 18952 21189 18955
rect 20956 18924 21189 18952
rect 20956 18912 20962 18924
rect 21177 18921 21189 18924
rect 21223 18921 21235 18955
rect 21177 18915 21235 18921
rect 21726 18912 21732 18964
rect 21784 18912 21790 18964
rect 21821 18955 21879 18961
rect 21821 18921 21833 18955
rect 21867 18952 21879 18955
rect 23106 18952 23112 18964
rect 21867 18924 23112 18952
rect 21867 18921 21879 18924
rect 21821 18915 21879 18921
rect 23106 18912 23112 18924
rect 23164 18912 23170 18964
rect 23750 18912 23756 18964
rect 23808 18952 23814 18964
rect 23937 18955 23995 18961
rect 23937 18952 23949 18955
rect 23808 18924 23949 18952
rect 23808 18912 23814 18924
rect 23937 18921 23949 18924
rect 23983 18952 23995 18955
rect 24762 18952 24768 18964
rect 23983 18924 24768 18952
rect 23983 18921 23995 18924
rect 23937 18915 23995 18921
rect 24762 18912 24768 18924
rect 24820 18912 24826 18964
rect 25866 18912 25872 18964
rect 25924 18912 25930 18964
rect 27985 18955 28043 18961
rect 27985 18952 27997 18955
rect 25976 18924 27997 18952
rect 22370 18884 22376 18896
rect 21008 18856 22376 18884
rect 21008 18825 21036 18856
rect 22370 18844 22376 18856
rect 22428 18844 22434 18896
rect 23842 18844 23848 18896
rect 23900 18884 23906 18896
rect 24578 18884 24584 18896
rect 23900 18856 24584 18884
rect 23900 18844 23906 18856
rect 24578 18844 24584 18856
rect 24636 18844 24642 18896
rect 24673 18887 24731 18893
rect 24673 18853 24685 18887
rect 24719 18853 24731 18887
rect 25976 18884 26004 18924
rect 27985 18921 27997 18924
rect 28031 18921 28043 18955
rect 27985 18915 28043 18921
rect 28626 18912 28632 18964
rect 28684 18952 28690 18964
rect 29914 18952 29920 18964
rect 28684 18924 29920 18952
rect 28684 18912 28690 18924
rect 29914 18912 29920 18924
rect 29972 18912 29978 18964
rect 32214 18912 32220 18964
rect 32272 18952 32278 18964
rect 32858 18952 32864 18964
rect 32272 18924 32864 18952
rect 32272 18912 32278 18924
rect 32858 18912 32864 18924
rect 32916 18912 32922 18964
rect 33134 18912 33140 18964
rect 33192 18952 33198 18964
rect 33502 18952 33508 18964
rect 33192 18924 33508 18952
rect 33192 18912 33198 18924
rect 33502 18912 33508 18924
rect 33560 18912 33566 18964
rect 33594 18912 33600 18964
rect 33652 18952 33658 18964
rect 35066 18952 35072 18964
rect 33652 18924 35072 18952
rect 33652 18912 33658 18924
rect 35066 18912 35072 18924
rect 35124 18952 35130 18964
rect 35618 18952 35624 18964
rect 35124 18924 35624 18952
rect 35124 18912 35130 18924
rect 35618 18912 35624 18924
rect 35676 18912 35682 18964
rect 36446 18912 36452 18964
rect 36504 18952 36510 18964
rect 37921 18955 37979 18961
rect 37921 18952 37933 18955
rect 36504 18924 37933 18952
rect 36504 18912 36510 18924
rect 37921 18921 37933 18924
rect 37967 18921 37979 18955
rect 37921 18915 37979 18921
rect 24673 18847 24731 18853
rect 24780 18856 26004 18884
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18785 18659 18819
rect 18601 18779 18659 18785
rect 18785 18819 18843 18825
rect 18785 18785 18797 18819
rect 18831 18816 18843 18819
rect 20993 18819 21051 18825
rect 20993 18816 21005 18819
rect 18831 18788 21005 18816
rect 18831 18785 18843 18788
rect 18785 18779 18843 18785
rect 20993 18785 21005 18788
rect 21039 18785 21051 18819
rect 20993 18779 21051 18785
rect 21450 18776 21456 18828
rect 21508 18816 21514 18828
rect 21913 18819 21971 18825
rect 21913 18816 21925 18819
rect 21508 18788 21925 18816
rect 21508 18776 21514 18788
rect 21913 18785 21925 18788
rect 21959 18785 21971 18819
rect 21913 18779 21971 18785
rect 22002 18776 22008 18828
rect 22060 18816 22066 18828
rect 24688 18816 24716 18847
rect 22060 18788 24716 18816
rect 22060 18776 22066 18788
rect 14737 18751 14795 18757
rect 14737 18748 14749 18751
rect 14700 18720 14749 18748
rect 14700 18708 14706 18720
rect 14737 18717 14749 18720
rect 14783 18717 14795 18751
rect 14737 18711 14795 18717
rect 15010 18708 15016 18760
rect 15068 18708 15074 18760
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 15396 18720 15761 18748
rect 14921 18683 14979 18689
rect 14921 18649 14933 18683
rect 14967 18680 14979 18683
rect 15396 18680 15424 18720
rect 15749 18717 15761 18720
rect 15795 18748 15807 18751
rect 16224 18748 16252 18776
rect 15795 18720 16252 18748
rect 16577 18751 16635 18757
rect 15795 18717 15807 18720
rect 15749 18711 15807 18717
rect 16577 18717 16589 18751
rect 16623 18748 16635 18751
rect 16758 18748 16764 18760
rect 16623 18720 16764 18748
rect 16623 18717 16635 18720
rect 16577 18711 16635 18717
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 17126 18708 17132 18760
rect 17184 18748 17190 18760
rect 17313 18751 17371 18757
rect 17313 18748 17325 18751
rect 17184 18720 17325 18748
rect 17184 18708 17190 18720
rect 17313 18717 17325 18720
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18748 17555 18751
rect 18966 18748 18972 18760
rect 17543 18720 18972 18748
rect 17543 18717 17555 18720
rect 17497 18711 17555 18717
rect 14967 18652 15424 18680
rect 14967 18649 14979 18652
rect 14921 18643 14979 18649
rect 15470 18640 15476 18692
rect 15528 18640 15534 18692
rect 15657 18683 15715 18689
rect 15657 18649 15669 18683
rect 15703 18649 15715 18683
rect 15657 18643 15715 18649
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 14734 18612 14740 18624
rect 11112 18584 14740 18612
rect 11112 18572 11118 18584
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 15010 18572 15016 18624
rect 15068 18612 15074 18624
rect 15672 18612 15700 18643
rect 15068 18584 15700 18612
rect 15068 18572 15074 18584
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 16853 18615 16911 18621
rect 16853 18612 16865 18615
rect 16080 18584 16865 18612
rect 16080 18572 16086 18584
rect 16853 18581 16865 18584
rect 16899 18581 16911 18615
rect 17328 18612 17356 18711
rect 18966 18708 18972 18720
rect 19024 18708 19030 18760
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 20530 18708 20536 18760
rect 20588 18708 20594 18760
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18748 20959 18751
rect 21468 18748 21496 18776
rect 20947 18720 21496 18748
rect 20947 18717 20959 18720
rect 20901 18711 20959 18717
rect 21634 18708 21640 18760
rect 21692 18708 21698 18760
rect 22830 18708 22836 18760
rect 22888 18748 22894 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 22888 18720 22937 18748
rect 22888 18708 22894 18720
rect 22925 18717 22937 18720
rect 22971 18717 22983 18751
rect 22925 18711 22983 18717
rect 23201 18751 23259 18757
rect 23201 18717 23213 18751
rect 23247 18748 23259 18751
rect 23290 18748 23296 18760
rect 23247 18720 23296 18748
rect 23247 18717 23259 18720
rect 23201 18711 23259 18717
rect 23290 18708 23296 18720
rect 23348 18708 23354 18760
rect 23750 18708 23756 18760
rect 23808 18748 23814 18760
rect 23845 18751 23903 18757
rect 23845 18748 23857 18751
rect 23808 18720 23857 18748
rect 23808 18708 23814 18720
rect 23845 18717 23857 18720
rect 23891 18717 23903 18751
rect 23845 18711 23903 18717
rect 23934 18708 23940 18760
rect 23992 18748 23998 18760
rect 24780 18748 24808 18856
rect 26050 18844 26056 18896
rect 26108 18884 26114 18896
rect 26970 18884 26976 18896
rect 26108 18856 26976 18884
rect 26108 18844 26114 18856
rect 26970 18844 26976 18856
rect 27028 18844 27034 18896
rect 27249 18887 27307 18893
rect 27249 18853 27261 18887
rect 27295 18884 27307 18887
rect 27338 18884 27344 18896
rect 27295 18856 27344 18884
rect 27295 18853 27307 18856
rect 27249 18847 27307 18853
rect 27338 18844 27344 18856
rect 27396 18844 27402 18896
rect 29362 18884 29368 18896
rect 28092 18856 29368 18884
rect 25133 18819 25191 18825
rect 25133 18785 25145 18819
rect 25179 18816 25191 18819
rect 25222 18816 25228 18828
rect 25179 18788 25228 18816
rect 25179 18785 25191 18788
rect 25133 18779 25191 18785
rect 25222 18776 25228 18788
rect 25280 18776 25286 18828
rect 27706 18816 27712 18828
rect 25884 18788 27712 18816
rect 25884 18760 25912 18788
rect 27706 18776 27712 18788
rect 27764 18776 27770 18828
rect 23992 18720 24808 18748
rect 23992 18708 23998 18720
rect 25866 18708 25872 18760
rect 25924 18708 25930 18760
rect 26050 18708 26056 18760
rect 26108 18708 26114 18760
rect 26510 18708 26516 18760
rect 26568 18748 26574 18760
rect 26697 18751 26755 18757
rect 26697 18748 26709 18751
rect 26568 18720 26709 18748
rect 26568 18708 26574 18720
rect 26697 18717 26709 18720
rect 26743 18717 26755 18751
rect 26697 18711 26755 18717
rect 26786 18708 26792 18760
rect 26844 18748 26850 18760
rect 26881 18751 26939 18757
rect 26881 18748 26893 18751
rect 26844 18720 26893 18748
rect 26844 18708 26850 18720
rect 26881 18717 26893 18720
rect 26927 18717 26939 18751
rect 26881 18711 26939 18717
rect 27062 18708 27068 18760
rect 27120 18757 27126 18760
rect 27120 18748 27128 18757
rect 27522 18748 27528 18760
rect 27120 18720 27528 18748
rect 27120 18711 27128 18720
rect 27120 18708 27126 18711
rect 27522 18708 27528 18720
rect 27580 18708 27586 18760
rect 28092 18748 28120 18856
rect 29362 18844 29368 18856
rect 29420 18844 29426 18896
rect 30006 18884 30012 18896
rect 29932 18856 30012 18884
rect 28534 18816 28540 18828
rect 28460 18788 28540 18816
rect 27632 18720 28120 18748
rect 17681 18683 17739 18689
rect 17681 18649 17693 18683
rect 17727 18680 17739 18683
rect 17770 18680 17776 18692
rect 17727 18652 17776 18680
rect 17727 18649 17739 18652
rect 17681 18643 17739 18649
rect 17770 18640 17776 18652
rect 17828 18640 17834 18692
rect 18509 18683 18567 18689
rect 17880 18652 18460 18680
rect 17880 18612 17908 18652
rect 17328 18584 17908 18612
rect 18141 18615 18199 18621
rect 16853 18575 16911 18581
rect 18141 18581 18153 18615
rect 18187 18612 18199 18615
rect 18322 18612 18328 18624
rect 18187 18584 18328 18612
rect 18187 18581 18199 18584
rect 18141 18575 18199 18581
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 18432 18612 18460 18652
rect 18509 18649 18521 18683
rect 18555 18680 18567 18683
rect 18598 18680 18604 18692
rect 18555 18652 18604 18680
rect 18555 18649 18567 18652
rect 18509 18643 18567 18649
rect 18598 18640 18604 18652
rect 18656 18640 18662 18692
rect 19429 18683 19487 18689
rect 19429 18649 19441 18683
rect 19475 18649 19487 18683
rect 19429 18643 19487 18649
rect 19981 18683 20039 18689
rect 19981 18649 19993 18683
rect 20027 18680 20039 18683
rect 20622 18680 20628 18692
rect 20027 18652 20628 18680
rect 20027 18649 20039 18652
rect 19981 18643 20039 18649
rect 19444 18612 19472 18643
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 23014 18640 23020 18692
rect 23072 18680 23078 18692
rect 23661 18683 23719 18689
rect 23661 18680 23673 18683
rect 23072 18652 23673 18680
rect 23072 18640 23078 18652
rect 23661 18649 23673 18652
rect 23707 18680 23719 18683
rect 24394 18680 24400 18692
rect 23707 18652 24400 18680
rect 23707 18649 23719 18652
rect 23661 18643 23719 18649
rect 24394 18640 24400 18652
rect 24452 18640 24458 18692
rect 25130 18640 25136 18692
rect 25188 18640 25194 18692
rect 25222 18640 25228 18692
rect 25280 18640 25286 18692
rect 26973 18683 27031 18689
rect 26973 18649 26985 18683
rect 27019 18680 27031 18683
rect 27632 18680 27660 18720
rect 28166 18708 28172 18760
rect 28224 18708 28230 18760
rect 28350 18708 28356 18760
rect 28408 18708 28414 18760
rect 28460 18757 28488 18788
rect 28534 18776 28540 18788
rect 28592 18816 28598 18828
rect 29454 18816 29460 18828
rect 28592 18788 29460 18816
rect 28592 18776 28598 18788
rect 29454 18776 29460 18788
rect 29512 18776 29518 18828
rect 28445 18751 28503 18757
rect 28445 18717 28457 18751
rect 28491 18717 28503 18751
rect 29089 18751 29147 18757
rect 29089 18748 29101 18751
rect 28445 18711 28503 18717
rect 28552 18720 29101 18748
rect 27019 18652 27660 18680
rect 27019 18649 27031 18652
rect 26973 18643 27031 18649
rect 27706 18640 27712 18692
rect 27764 18680 27770 18692
rect 28552 18680 28580 18720
rect 29089 18717 29101 18720
rect 29135 18717 29147 18751
rect 29089 18711 29147 18717
rect 29181 18751 29239 18757
rect 29181 18717 29193 18751
rect 29227 18748 29239 18751
rect 29822 18748 29828 18760
rect 29227 18720 29828 18748
rect 29227 18717 29239 18720
rect 29181 18711 29239 18717
rect 29822 18708 29828 18720
rect 29880 18708 29886 18760
rect 29932 18757 29960 18856
rect 30006 18844 30012 18856
rect 30064 18844 30070 18896
rect 30469 18887 30527 18893
rect 30469 18853 30481 18887
rect 30515 18853 30527 18887
rect 30469 18847 30527 18853
rect 30484 18816 30512 18847
rect 30834 18844 30840 18896
rect 30892 18884 30898 18896
rect 30892 18856 31064 18884
rect 30892 18844 30898 18856
rect 31036 18825 31064 18856
rect 31570 18844 31576 18896
rect 31628 18884 31634 18896
rect 31628 18856 33732 18884
rect 31628 18844 31634 18856
rect 30920 18819 30978 18825
rect 30920 18816 30932 18819
rect 30484 18788 30932 18816
rect 30920 18785 30932 18788
rect 30966 18785 30978 18819
rect 30920 18779 30978 18785
rect 31021 18819 31079 18825
rect 31021 18785 31033 18819
rect 31067 18785 31079 18819
rect 31294 18816 31300 18828
rect 31021 18779 31079 18785
rect 31119 18788 31300 18816
rect 29917 18751 29975 18757
rect 29917 18717 29929 18751
rect 29963 18717 29975 18751
rect 29917 18711 29975 18717
rect 30006 18708 30012 18760
rect 30064 18747 30070 18760
rect 30101 18751 30159 18757
rect 30101 18747 30113 18751
rect 30064 18719 30113 18747
rect 30064 18708 30070 18719
rect 30101 18717 30113 18719
rect 30147 18717 30159 18751
rect 30101 18711 30159 18717
rect 30331 18751 30389 18757
rect 30331 18717 30343 18751
rect 30377 18748 30389 18751
rect 31119 18748 31147 18788
rect 31294 18776 31300 18788
rect 31352 18776 31358 18828
rect 31496 18788 33088 18816
rect 30377 18720 31147 18748
rect 30377 18717 30389 18720
rect 30331 18711 30389 18717
rect 31202 18708 31208 18760
rect 31260 18708 31266 18760
rect 31496 18757 31524 18788
rect 31481 18751 31539 18757
rect 31481 18717 31493 18751
rect 31527 18717 31539 18751
rect 31481 18711 31539 18717
rect 31662 18708 31668 18760
rect 31720 18708 31726 18760
rect 32398 18708 32404 18760
rect 32456 18748 32462 18760
rect 32769 18751 32827 18757
rect 32769 18748 32781 18751
rect 32456 18720 32781 18748
rect 32456 18708 32462 18720
rect 32769 18717 32781 18720
rect 32815 18717 32827 18751
rect 32769 18711 32827 18717
rect 32858 18708 32864 18760
rect 32916 18708 32922 18760
rect 27764 18652 28580 18680
rect 28905 18683 28963 18689
rect 27764 18640 27770 18652
rect 28905 18649 28917 18683
rect 28951 18680 28963 18683
rect 29362 18680 29368 18692
rect 28951 18652 29368 18680
rect 28951 18649 28963 18652
rect 28905 18643 28963 18649
rect 18432 18584 19472 18612
rect 22738 18572 22744 18624
rect 22796 18572 22802 18624
rect 23109 18615 23167 18621
rect 23109 18581 23121 18615
rect 23155 18612 23167 18615
rect 23382 18612 23388 18624
rect 23155 18584 23388 18612
rect 23155 18581 23167 18584
rect 23109 18575 23167 18581
rect 23382 18572 23388 18584
rect 23440 18612 23446 18624
rect 24578 18612 24584 18624
rect 23440 18584 24584 18612
rect 23440 18572 23446 18584
rect 24578 18572 24584 18584
rect 24636 18572 24642 18624
rect 26237 18615 26295 18621
rect 26237 18581 26249 18615
rect 26283 18612 26295 18615
rect 27338 18612 27344 18624
rect 26283 18584 27344 18612
rect 26283 18581 26295 18584
rect 26237 18575 26295 18581
rect 27338 18572 27344 18584
rect 27396 18572 27402 18624
rect 27522 18572 27528 18624
rect 27580 18612 27586 18624
rect 28920 18612 28948 18643
rect 29362 18640 29368 18652
rect 29420 18640 29426 18692
rect 30193 18683 30251 18689
rect 30193 18649 30205 18683
rect 30239 18680 30251 18683
rect 30466 18680 30472 18692
rect 30239 18652 30472 18680
rect 30239 18649 30251 18652
rect 30193 18643 30251 18649
rect 30466 18640 30472 18652
rect 30524 18680 30530 18692
rect 32306 18680 32312 18692
rect 30524 18652 32312 18680
rect 30524 18640 30530 18652
rect 32306 18640 32312 18652
rect 32364 18640 32370 18692
rect 27580 18584 28948 18612
rect 27580 18572 27586 18584
rect 28994 18572 29000 18624
rect 29052 18621 29058 18624
rect 29052 18575 29061 18621
rect 29052 18572 29058 18575
rect 30558 18572 30564 18624
rect 30616 18612 30622 18624
rect 31202 18612 31208 18624
rect 30616 18584 31208 18612
rect 30616 18572 30622 18584
rect 31202 18572 31208 18584
rect 31260 18572 31266 18624
rect 31294 18572 31300 18624
rect 31352 18612 31358 18624
rect 32490 18612 32496 18624
rect 31352 18584 32496 18612
rect 31352 18572 31358 18584
rect 32490 18572 32496 18584
rect 32548 18572 32554 18624
rect 32582 18572 32588 18624
rect 32640 18572 32646 18624
rect 33060 18612 33088 18788
rect 33226 18776 33232 18828
rect 33284 18776 33290 18828
rect 33704 18748 33732 18856
rect 33962 18844 33968 18896
rect 34020 18844 34026 18896
rect 35529 18887 35587 18893
rect 35529 18884 35541 18887
rect 34348 18856 35541 18884
rect 33781 18819 33839 18825
rect 33781 18785 33793 18819
rect 33827 18816 33839 18819
rect 33980 18816 34008 18844
rect 34348 18825 34376 18856
rect 35529 18853 35541 18856
rect 35575 18853 35587 18887
rect 35529 18847 35587 18853
rect 33827 18788 34008 18816
rect 34333 18819 34391 18825
rect 33827 18785 33839 18788
rect 33781 18779 33839 18785
rect 34333 18785 34345 18819
rect 34379 18785 34391 18819
rect 36262 18816 36268 18828
rect 34333 18779 34391 18785
rect 34440 18788 36268 18816
rect 33965 18751 34023 18757
rect 33965 18748 33977 18751
rect 33152 18720 33456 18748
rect 33704 18720 33977 18748
rect 33152 18692 33180 18720
rect 33134 18640 33140 18692
rect 33192 18640 33198 18692
rect 33428 18680 33456 18720
rect 33965 18717 33977 18720
rect 34011 18748 34023 18751
rect 34440 18748 34468 18788
rect 36262 18776 36268 18788
rect 36320 18776 36326 18828
rect 34011 18720 34468 18748
rect 34011 18717 34023 18720
rect 33965 18711 34023 18717
rect 34514 18708 34520 18760
rect 34572 18748 34578 18760
rect 34885 18751 34943 18757
rect 34885 18748 34897 18751
rect 34572 18720 34897 18748
rect 34572 18708 34578 18720
rect 34885 18717 34897 18720
rect 34931 18717 34943 18751
rect 34885 18711 34943 18717
rect 34974 18708 34980 18760
rect 35032 18748 35038 18760
rect 35032 18720 35077 18748
rect 35032 18708 35038 18720
rect 35158 18708 35164 18760
rect 35216 18708 35222 18760
rect 35342 18708 35348 18760
rect 35400 18757 35406 18760
rect 35400 18748 35408 18757
rect 35400 18720 35445 18748
rect 35400 18711 35408 18720
rect 35400 18708 35406 18711
rect 36538 18708 36544 18760
rect 36596 18708 36602 18760
rect 35253 18683 35311 18689
rect 33428 18652 35112 18680
rect 33686 18612 33692 18624
rect 33060 18584 33692 18612
rect 33686 18572 33692 18584
rect 33744 18572 33750 18624
rect 33962 18572 33968 18624
rect 34020 18572 34026 18624
rect 35084 18612 35112 18652
rect 35253 18649 35265 18683
rect 35299 18649 35311 18683
rect 35253 18643 35311 18649
rect 35268 18612 35296 18643
rect 36446 18640 36452 18692
rect 36504 18680 36510 18692
rect 36786 18683 36844 18689
rect 36786 18680 36798 18683
rect 36504 18652 36798 18680
rect 36504 18640 36510 18652
rect 36786 18649 36798 18652
rect 36832 18649 36844 18683
rect 36786 18643 36844 18649
rect 35084 18584 35296 18612
rect 35342 18572 35348 18624
rect 35400 18612 35406 18624
rect 37826 18612 37832 18624
rect 35400 18584 37832 18612
rect 35400 18572 35406 18584
rect 37826 18572 37832 18584
rect 37884 18572 37890 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 14366 18368 14372 18420
rect 14424 18368 14430 18420
rect 15378 18368 15384 18420
rect 15436 18408 15442 18420
rect 15565 18411 15623 18417
rect 15565 18408 15577 18411
rect 15436 18380 15577 18408
rect 15436 18368 15442 18380
rect 15565 18377 15577 18380
rect 15611 18377 15623 18411
rect 16942 18408 16948 18420
rect 15565 18371 15623 18377
rect 15948 18380 16948 18408
rect 12894 18300 12900 18352
rect 12952 18340 12958 18352
rect 15948 18340 15976 18380
rect 16942 18368 16948 18380
rect 17000 18408 17006 18420
rect 17000 18380 18460 18408
rect 17000 18368 17006 18380
rect 12952 18312 15976 18340
rect 12952 18300 12958 18312
rect 16022 18300 16028 18352
rect 16080 18300 16086 18352
rect 14090 18232 14096 18284
rect 14148 18232 14154 18284
rect 14185 18275 14243 18281
rect 14185 18241 14197 18275
rect 14231 18272 14243 18275
rect 14826 18272 14832 18284
rect 14231 18244 14832 18272
rect 14231 18241 14243 18244
rect 14185 18235 14243 18241
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 15010 18164 15016 18216
rect 15068 18204 15074 18216
rect 15197 18207 15255 18213
rect 15197 18204 15209 18207
rect 15068 18176 15209 18204
rect 15068 18164 15074 18176
rect 15197 18173 15209 18176
rect 15243 18173 15255 18207
rect 15396 18204 15424 18235
rect 16206 18232 16212 18284
rect 16264 18232 16270 18284
rect 16298 18232 16304 18284
rect 16356 18232 16362 18284
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18272 17371 18275
rect 18322 18272 18328 18284
rect 17359 18244 18328 18272
rect 17359 18241 17371 18244
rect 17313 18235 17371 18241
rect 18322 18232 18328 18244
rect 18380 18232 18386 18284
rect 18432 18281 18460 18380
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 19613 18411 19671 18417
rect 19613 18408 19625 18411
rect 19392 18380 19625 18408
rect 19392 18368 19398 18380
rect 19613 18377 19625 18380
rect 19659 18408 19671 18411
rect 20070 18408 20076 18420
rect 19659 18380 20076 18408
rect 19659 18377 19671 18380
rect 19613 18371 19671 18377
rect 20070 18368 20076 18380
rect 20128 18368 20134 18420
rect 20162 18368 20168 18420
rect 20220 18408 20226 18420
rect 23109 18411 23167 18417
rect 23109 18408 23121 18411
rect 20220 18380 23121 18408
rect 20220 18368 20226 18380
rect 23109 18377 23121 18380
rect 23155 18377 23167 18411
rect 23109 18371 23167 18377
rect 23198 18368 23204 18420
rect 23256 18408 23262 18420
rect 23474 18408 23480 18420
rect 23256 18380 23480 18408
rect 23256 18368 23262 18380
rect 23474 18368 23480 18380
rect 23532 18368 23538 18420
rect 24302 18368 24308 18420
rect 24360 18408 24366 18420
rect 24673 18411 24731 18417
rect 24673 18408 24685 18411
rect 24360 18380 24685 18408
rect 24360 18368 24366 18380
rect 24673 18377 24685 18380
rect 24719 18377 24731 18411
rect 29914 18408 29920 18420
rect 24673 18371 24731 18377
rect 26988 18380 29920 18408
rect 20438 18340 20444 18352
rect 18616 18312 20444 18340
rect 18616 18281 18644 18312
rect 18417 18275 18475 18281
rect 18417 18241 18429 18275
rect 18463 18241 18475 18275
rect 18417 18235 18475 18241
rect 18601 18275 18659 18281
rect 18601 18241 18613 18275
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 18693 18275 18751 18281
rect 18693 18241 18705 18275
rect 18739 18241 18751 18275
rect 18693 18235 18751 18241
rect 17589 18207 17647 18213
rect 15396 18176 16160 18204
rect 15197 18167 15255 18173
rect 16132 18145 16160 18176
rect 17589 18173 17601 18207
rect 17635 18204 17647 18207
rect 18506 18204 18512 18216
rect 17635 18176 18512 18204
rect 17635 18173 17647 18176
rect 17589 18167 17647 18173
rect 18506 18164 18512 18176
rect 18564 18204 18570 18216
rect 18708 18204 18736 18235
rect 18564 18176 18736 18204
rect 18564 18164 18570 18176
rect 16117 18139 16175 18145
rect 16117 18105 16129 18139
rect 16163 18105 16175 18139
rect 16117 18099 16175 18105
rect 17497 18139 17555 18145
rect 17497 18105 17509 18139
rect 17543 18136 17555 18139
rect 18800 18136 18828 18312
rect 20438 18300 20444 18312
rect 20496 18300 20502 18352
rect 20622 18300 20628 18352
rect 20680 18340 20686 18352
rect 20717 18343 20775 18349
rect 20717 18340 20729 18343
rect 20680 18312 20729 18340
rect 20680 18300 20686 18312
rect 20717 18309 20729 18312
rect 20763 18309 20775 18343
rect 20717 18303 20775 18309
rect 22738 18300 22744 18352
rect 22796 18340 22802 18352
rect 25222 18340 25228 18352
rect 22796 18312 23429 18340
rect 22796 18300 22802 18312
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18272 19579 18275
rect 20640 18272 20668 18300
rect 19567 18244 20668 18272
rect 19567 18241 19579 18244
rect 19521 18235 19579 18241
rect 22278 18232 22284 18284
rect 22336 18232 22342 18284
rect 22370 18232 22376 18284
rect 22428 18232 22434 18284
rect 22462 18232 22468 18284
rect 22520 18272 22526 18284
rect 23401 18281 23429 18312
rect 24044 18312 25228 18340
rect 24044 18284 24072 18312
rect 25222 18300 25228 18312
rect 25280 18300 25286 18352
rect 22649 18275 22707 18281
rect 22649 18272 22661 18275
rect 22520 18244 22661 18272
rect 22520 18232 22526 18244
rect 22649 18241 22661 18244
rect 22695 18241 22707 18275
rect 22649 18235 22707 18241
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18241 23351 18275
rect 23293 18235 23351 18241
rect 23385 18275 23443 18281
rect 23385 18241 23397 18275
rect 23431 18241 23443 18275
rect 23385 18235 23443 18241
rect 23661 18275 23719 18281
rect 23661 18241 23673 18275
rect 23707 18272 23719 18275
rect 24026 18272 24032 18284
rect 23707 18244 24032 18272
rect 23707 18241 23719 18244
rect 23661 18235 23719 18241
rect 19794 18164 19800 18216
rect 19852 18164 19858 18216
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 20806 18204 20812 18216
rect 20128 18176 20812 18204
rect 20128 18164 20134 18176
rect 20806 18164 20812 18176
rect 20864 18164 20870 18216
rect 20993 18207 21051 18213
rect 20993 18173 21005 18207
rect 21039 18204 21051 18207
rect 22186 18204 22192 18216
rect 21039 18176 22192 18204
rect 21039 18173 21051 18176
rect 20993 18167 21051 18173
rect 22186 18164 22192 18176
rect 22244 18164 22250 18216
rect 23309 18204 23337 18235
rect 24026 18232 24032 18244
rect 24084 18232 24090 18284
rect 24121 18275 24179 18281
rect 24121 18241 24133 18275
rect 24167 18272 24179 18275
rect 24302 18272 24308 18284
rect 24167 18244 24308 18272
rect 24167 18241 24179 18244
rect 24121 18235 24179 18241
rect 24302 18232 24308 18244
rect 24360 18232 24366 18284
rect 25682 18232 25688 18284
rect 25740 18232 25746 18284
rect 25866 18232 25872 18284
rect 25924 18232 25930 18284
rect 26234 18232 26240 18284
rect 26292 18272 26298 18284
rect 26421 18275 26479 18281
rect 26421 18272 26433 18275
rect 26292 18244 26433 18272
rect 26292 18232 26298 18244
rect 26421 18241 26433 18244
rect 26467 18241 26479 18275
rect 26421 18235 26479 18241
rect 26602 18232 26608 18284
rect 26660 18232 26666 18284
rect 26988 18272 27016 18380
rect 29914 18368 29920 18380
rect 29972 18408 29978 18420
rect 30834 18408 30840 18420
rect 29972 18380 30840 18408
rect 29972 18368 29978 18380
rect 30834 18368 30840 18380
rect 30892 18368 30898 18420
rect 32214 18368 32220 18420
rect 32272 18408 32278 18420
rect 32272 18380 32536 18408
rect 32272 18368 32278 18380
rect 27341 18343 27399 18349
rect 27341 18340 27353 18343
rect 27264 18312 27353 18340
rect 27264 18284 27292 18312
rect 27341 18309 27353 18312
rect 27387 18309 27399 18343
rect 27614 18340 27620 18352
rect 27341 18303 27399 18309
rect 27586 18300 27620 18340
rect 27672 18300 27678 18352
rect 32398 18340 32404 18352
rect 29288 18312 32404 18340
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 26988 18244 27169 18272
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 23566 18204 23572 18216
rect 23309 18176 23572 18204
rect 23566 18164 23572 18176
rect 23624 18164 23630 18216
rect 24394 18164 24400 18216
rect 24452 18164 24458 18216
rect 25958 18164 25964 18216
rect 26016 18164 26022 18216
rect 26050 18164 26056 18216
rect 26108 18204 26114 18216
rect 27172 18204 27200 18235
rect 27246 18232 27252 18284
rect 27304 18232 27310 18284
rect 27586 18281 27614 18300
rect 27434 18275 27492 18281
rect 27434 18241 27446 18275
rect 27480 18241 27492 18275
rect 27434 18235 27492 18241
rect 27553 18275 27614 18281
rect 27553 18241 27565 18275
rect 27599 18241 27614 18275
rect 27553 18235 27614 18241
rect 26108 18176 27200 18204
rect 27448 18204 27476 18235
rect 27568 18234 27614 18235
rect 29086 18232 29092 18284
rect 29144 18232 29150 18284
rect 29288 18281 29316 18312
rect 32398 18300 32404 18312
rect 32456 18300 32462 18352
rect 32508 18340 32536 18380
rect 35250 18368 35256 18420
rect 35308 18408 35314 18420
rect 35526 18408 35532 18420
rect 35308 18380 35532 18408
rect 35308 18368 35314 18380
rect 35526 18368 35532 18380
rect 35584 18368 35590 18420
rect 32508 18312 32608 18340
rect 32580 18303 32608 18312
rect 32692 18312 34928 18340
rect 32580 18297 32643 18303
rect 29273 18275 29331 18281
rect 29273 18241 29285 18275
rect 29319 18241 29331 18275
rect 29273 18235 29331 18241
rect 29365 18275 29423 18281
rect 29365 18241 29377 18275
rect 29411 18272 29423 18275
rect 29454 18272 29460 18284
rect 29411 18244 29460 18272
rect 29411 18241 29423 18244
rect 29365 18235 29423 18241
rect 29454 18232 29460 18244
rect 29512 18232 29518 18284
rect 30009 18275 30067 18281
rect 30009 18241 30021 18275
rect 30055 18272 30067 18275
rect 30282 18272 30288 18284
rect 30055 18244 30288 18272
rect 30055 18241 30067 18244
rect 30009 18235 30067 18241
rect 30282 18232 30288 18244
rect 30340 18232 30346 18284
rect 30374 18232 30380 18284
rect 30432 18232 30438 18284
rect 30558 18232 30564 18284
rect 30616 18272 30622 18284
rect 30837 18275 30895 18281
rect 30837 18272 30849 18275
rect 30616 18244 30849 18272
rect 30616 18232 30622 18244
rect 30837 18241 30849 18244
rect 30883 18241 30895 18275
rect 31754 18272 31760 18284
rect 30837 18235 30895 18241
rect 30944 18244 31760 18272
rect 30193 18207 30251 18213
rect 27448 18176 30144 18204
rect 26108 18164 26114 18176
rect 17543 18108 18828 18136
rect 22557 18139 22615 18145
rect 17543 18105 17555 18108
rect 17497 18099 17555 18105
rect 22557 18105 22569 18139
rect 22603 18136 22615 18139
rect 23382 18136 23388 18148
rect 22603 18108 23388 18136
rect 22603 18105 22615 18108
rect 22557 18099 22615 18105
rect 23382 18096 23388 18108
rect 23440 18096 23446 18148
rect 24578 18096 24584 18148
rect 24636 18136 24642 18148
rect 28905 18139 28963 18145
rect 28905 18136 28917 18139
rect 24636 18108 28917 18136
rect 24636 18096 24642 18108
rect 28905 18105 28917 18108
rect 28951 18105 28963 18139
rect 28905 18099 28963 18105
rect 30006 18096 30012 18148
rect 30064 18096 30070 18148
rect 30116 18136 30144 18176
rect 30193 18173 30205 18207
rect 30239 18204 30251 18207
rect 30944 18204 30972 18244
rect 31754 18232 31760 18244
rect 31812 18232 31818 18284
rect 32580 18266 32597 18297
rect 32585 18263 32597 18266
rect 32631 18263 32643 18297
rect 32585 18257 32643 18263
rect 30239 18176 30972 18204
rect 30239 18173 30251 18176
rect 30193 18167 30251 18173
rect 31570 18164 31576 18216
rect 31628 18164 31634 18216
rect 32214 18164 32220 18216
rect 32272 18204 32278 18216
rect 32490 18204 32496 18216
rect 32272 18176 32496 18204
rect 32272 18164 32278 18176
rect 32490 18164 32496 18176
rect 32548 18164 32554 18216
rect 32582 18164 32588 18216
rect 32640 18204 32646 18216
rect 32692 18204 32720 18312
rect 32953 18275 33011 18281
rect 32953 18241 32965 18275
rect 32999 18272 33011 18275
rect 33226 18272 33232 18284
rect 32999 18244 33232 18272
rect 32999 18241 33011 18244
rect 32953 18235 33011 18241
rect 33226 18232 33232 18244
rect 33284 18232 33290 18284
rect 33410 18232 33416 18284
rect 33468 18232 33474 18284
rect 33506 18275 33564 18281
rect 33506 18241 33518 18275
rect 33552 18241 33564 18275
rect 33506 18235 33564 18241
rect 32640 18176 32720 18204
rect 32640 18164 32646 18176
rect 32858 18164 32864 18216
rect 32916 18164 32922 18216
rect 30742 18136 30748 18148
rect 30116 18108 30748 18136
rect 30742 18096 30748 18108
rect 30800 18096 30806 18148
rect 30834 18096 30840 18148
rect 30892 18136 30898 18148
rect 33520 18136 33548 18235
rect 33594 18232 33600 18284
rect 33652 18272 33658 18284
rect 33689 18275 33747 18281
rect 33689 18272 33701 18275
rect 33652 18244 33701 18272
rect 33652 18232 33658 18244
rect 33689 18241 33701 18244
rect 33735 18241 33747 18275
rect 33689 18235 33747 18241
rect 33781 18275 33839 18281
rect 33781 18241 33793 18275
rect 33827 18241 33839 18275
rect 33781 18235 33839 18241
rect 33796 18204 33824 18235
rect 33870 18232 33876 18284
rect 33928 18281 33934 18284
rect 33928 18272 33936 18281
rect 33928 18244 33973 18272
rect 33928 18235 33936 18244
rect 33928 18232 33934 18235
rect 34790 18232 34796 18284
rect 34848 18232 34854 18284
rect 34900 18281 34928 18312
rect 34974 18300 34980 18352
rect 35032 18340 35038 18352
rect 35161 18343 35219 18349
rect 35161 18340 35173 18343
rect 35032 18312 35173 18340
rect 35032 18300 35038 18312
rect 35161 18309 35173 18312
rect 35207 18340 35219 18343
rect 35342 18340 35348 18352
rect 35207 18312 35348 18340
rect 35207 18309 35219 18312
rect 35161 18303 35219 18309
rect 35342 18300 35348 18312
rect 35400 18300 35406 18352
rect 35802 18300 35808 18352
rect 35860 18340 35866 18352
rect 35860 18312 36216 18340
rect 35860 18300 35866 18312
rect 34886 18275 34944 18281
rect 34886 18241 34898 18275
rect 34932 18241 34944 18275
rect 34886 18235 34944 18241
rect 35066 18232 35072 18284
rect 35124 18232 35130 18284
rect 35250 18232 35256 18284
rect 35308 18281 35314 18284
rect 36188 18281 36216 18312
rect 35308 18235 35316 18281
rect 36081 18275 36139 18281
rect 36081 18273 36093 18275
rect 36079 18272 36093 18273
rect 35820 18244 36093 18272
rect 35308 18232 35314 18235
rect 33704 18176 33824 18204
rect 33704 18148 33732 18176
rect 30892 18108 33548 18136
rect 30892 18096 30898 18108
rect 33686 18096 33692 18148
rect 33744 18096 33750 18148
rect 34606 18136 34612 18148
rect 33980 18108 34612 18136
rect 17129 18071 17187 18077
rect 17129 18037 17141 18071
rect 17175 18068 17187 18071
rect 17402 18068 17408 18080
rect 17175 18040 17408 18068
rect 17175 18037 17187 18040
rect 17129 18031 17187 18037
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 18138 18028 18144 18080
rect 18196 18028 18202 18080
rect 19150 18028 19156 18080
rect 19208 18028 19214 18080
rect 20349 18071 20407 18077
rect 20349 18037 20361 18071
rect 20395 18068 20407 18071
rect 20530 18068 20536 18080
rect 20395 18040 20536 18068
rect 20395 18037 20407 18040
rect 20349 18031 20407 18037
rect 20530 18028 20536 18040
rect 20588 18028 20594 18080
rect 21634 18028 21640 18080
rect 21692 18068 21698 18080
rect 22097 18071 22155 18077
rect 22097 18068 22109 18071
rect 21692 18040 22109 18068
rect 21692 18028 21698 18040
rect 22097 18037 22109 18040
rect 22143 18037 22155 18071
rect 22097 18031 22155 18037
rect 23474 18028 23480 18080
rect 23532 18068 23538 18080
rect 23569 18071 23627 18077
rect 23569 18068 23581 18071
rect 23532 18040 23581 18068
rect 23532 18028 23538 18040
rect 23569 18037 23581 18040
rect 23615 18068 23627 18071
rect 24210 18068 24216 18080
rect 23615 18040 24216 18068
rect 23615 18037 23627 18040
rect 23569 18031 23627 18037
rect 24210 18028 24216 18040
rect 24268 18028 24274 18080
rect 25498 18028 25504 18080
rect 25556 18028 25562 18080
rect 26510 18028 26516 18080
rect 26568 18028 26574 18080
rect 27709 18071 27767 18077
rect 27709 18037 27721 18071
rect 27755 18068 27767 18071
rect 28258 18068 28264 18080
rect 27755 18040 28264 18068
rect 27755 18037 27767 18040
rect 27709 18031 27767 18037
rect 28258 18028 28264 18040
rect 28316 18028 28322 18080
rect 29086 18028 29092 18080
rect 29144 18068 29150 18080
rect 31294 18068 31300 18080
rect 29144 18040 31300 18068
rect 29144 18028 29150 18040
rect 31294 18028 31300 18040
rect 31352 18028 31358 18080
rect 32309 18071 32367 18077
rect 32309 18037 32321 18071
rect 32355 18068 32367 18071
rect 33980 18068 34008 18108
rect 34606 18096 34612 18108
rect 34664 18096 34670 18148
rect 35437 18139 35495 18145
rect 35437 18105 35449 18139
rect 35483 18136 35495 18139
rect 35820 18136 35848 18244
rect 36081 18241 36093 18244
rect 36127 18241 36139 18275
rect 36081 18235 36139 18241
rect 36173 18275 36231 18281
rect 36173 18241 36185 18275
rect 36219 18241 36231 18275
rect 36173 18235 36231 18241
rect 36262 18232 36268 18284
rect 36320 18272 36326 18284
rect 36449 18275 36507 18281
rect 36449 18272 36461 18275
rect 36320 18244 36461 18272
rect 36320 18232 36326 18244
rect 36449 18241 36461 18244
rect 36495 18241 36507 18275
rect 36449 18235 36507 18241
rect 37826 18232 37832 18284
rect 37884 18232 37890 18284
rect 35897 18207 35955 18213
rect 35897 18173 35909 18207
rect 35943 18204 35955 18207
rect 36354 18204 36360 18216
rect 35943 18176 36360 18204
rect 35943 18173 35955 18176
rect 35897 18167 35955 18173
rect 36354 18164 36360 18176
rect 36412 18204 36418 18216
rect 37921 18207 37979 18213
rect 37921 18204 37933 18207
rect 36412 18176 37933 18204
rect 36412 18164 36418 18176
rect 37921 18173 37933 18176
rect 37967 18173 37979 18207
rect 37921 18167 37979 18173
rect 38102 18164 38108 18216
rect 38160 18164 38166 18216
rect 35483 18108 35848 18136
rect 35483 18105 35495 18108
rect 35437 18099 35495 18105
rect 32355 18040 34008 18068
rect 34057 18071 34115 18077
rect 32355 18037 32367 18040
rect 32309 18031 32367 18037
rect 34057 18037 34069 18071
rect 34103 18068 34115 18071
rect 34514 18068 34520 18080
rect 34103 18040 34520 18068
rect 34103 18037 34115 18040
rect 34057 18031 34115 18037
rect 34514 18028 34520 18040
rect 34572 18028 34578 18080
rect 35342 18028 35348 18080
rect 35400 18068 35406 18080
rect 36078 18068 36084 18080
rect 35400 18040 36084 18068
rect 35400 18028 35406 18040
rect 36078 18028 36084 18040
rect 36136 18068 36142 18080
rect 36357 18071 36415 18077
rect 36357 18068 36369 18071
rect 36136 18040 36369 18068
rect 36136 18028 36142 18040
rect 36357 18037 36369 18040
rect 36403 18037 36415 18071
rect 36357 18031 36415 18037
rect 37458 18028 37464 18080
rect 37516 18028 37522 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 15010 17824 15016 17876
rect 15068 17824 15074 17876
rect 15378 17824 15384 17876
rect 15436 17864 15442 17876
rect 15930 17864 15936 17876
rect 15436 17836 15936 17864
rect 15436 17824 15442 17836
rect 15930 17824 15936 17836
rect 15988 17864 15994 17876
rect 16298 17864 16304 17876
rect 15988 17836 16304 17864
rect 15988 17824 15994 17836
rect 16298 17824 16304 17836
rect 16356 17864 16362 17876
rect 16482 17864 16488 17876
rect 16356 17836 16488 17864
rect 16356 17824 16362 17836
rect 16482 17824 16488 17836
rect 16540 17864 16546 17876
rect 17865 17867 17923 17873
rect 17865 17864 17877 17867
rect 16540 17836 17877 17864
rect 16540 17824 16546 17836
rect 17865 17833 17877 17836
rect 17911 17833 17923 17867
rect 17865 17827 17923 17833
rect 18506 17824 18512 17876
rect 18564 17864 18570 17876
rect 18693 17867 18751 17873
rect 18693 17864 18705 17867
rect 18564 17836 18705 17864
rect 18564 17824 18570 17836
rect 18693 17833 18705 17836
rect 18739 17833 18751 17867
rect 18693 17827 18751 17833
rect 19518 17824 19524 17876
rect 19576 17864 19582 17876
rect 22002 17864 22008 17876
rect 19576 17836 22008 17864
rect 19576 17824 19582 17836
rect 22002 17824 22008 17836
rect 22060 17824 22066 17876
rect 22370 17824 22376 17876
rect 22428 17864 22434 17876
rect 22649 17867 22707 17873
rect 22649 17864 22661 17867
rect 22428 17836 22661 17864
rect 22428 17824 22434 17836
rect 22649 17833 22661 17836
rect 22695 17833 22707 17867
rect 22649 17827 22707 17833
rect 23566 17824 23572 17876
rect 23624 17824 23630 17876
rect 23937 17867 23995 17873
rect 23937 17833 23949 17867
rect 23983 17864 23995 17867
rect 26510 17864 26516 17876
rect 23983 17836 26516 17864
rect 23983 17833 23995 17836
rect 23937 17827 23995 17833
rect 26510 17824 26516 17836
rect 26568 17824 26574 17876
rect 27522 17864 27528 17876
rect 26620 17836 27528 17864
rect 20349 17799 20407 17805
rect 18708 17768 19334 17796
rect 16022 17728 16028 17740
rect 15212 17700 16028 17728
rect 15212 17669 15240 17700
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 16684 17700 18276 17728
rect 15197 17663 15255 17669
rect 15197 17629 15209 17663
rect 15243 17629 15255 17663
rect 15197 17623 15255 17629
rect 15378 17620 15384 17672
rect 15436 17620 15442 17672
rect 15473 17663 15531 17669
rect 15473 17629 15485 17663
rect 15519 17629 15531 17663
rect 15473 17623 15531 17629
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17660 15991 17663
rect 16684 17660 16712 17700
rect 18248 17672 18276 17700
rect 15979 17632 16712 17660
rect 16761 17663 16819 17669
rect 15979 17629 15991 17632
rect 15933 17623 15991 17629
rect 16761 17629 16773 17663
rect 16807 17629 16819 17663
rect 16761 17623 16819 17629
rect 17221 17663 17279 17669
rect 17221 17629 17233 17663
rect 17267 17660 17279 17663
rect 17494 17660 17500 17672
rect 17267 17632 17500 17660
rect 17267 17629 17279 17632
rect 17221 17623 17279 17629
rect 15488 17536 15516 17623
rect 15838 17552 15844 17604
rect 15896 17592 15902 17604
rect 16393 17595 16451 17601
rect 16393 17592 16405 17595
rect 15896 17564 16405 17592
rect 15896 17552 15902 17564
rect 16393 17561 16405 17564
rect 16439 17561 16451 17595
rect 16776 17592 16804 17623
rect 17494 17620 17500 17632
rect 17552 17620 17558 17672
rect 17770 17620 17776 17672
rect 17828 17620 17834 17672
rect 18230 17620 18236 17672
rect 18288 17620 18294 17672
rect 18708 17669 18736 17768
rect 19306 17728 19334 17768
rect 20349 17765 20361 17799
rect 20395 17796 20407 17799
rect 21266 17796 21272 17808
rect 20395 17768 21272 17796
rect 20395 17765 20407 17768
rect 20349 17759 20407 17765
rect 21266 17756 21272 17768
rect 21324 17756 21330 17808
rect 23290 17756 23296 17808
rect 23348 17796 23354 17808
rect 24670 17796 24676 17808
rect 23348 17768 24676 17796
rect 23348 17756 23354 17768
rect 24670 17756 24676 17768
rect 24728 17756 24734 17808
rect 24765 17799 24823 17805
rect 24765 17765 24777 17799
rect 24811 17765 24823 17799
rect 24765 17759 24823 17765
rect 24780 17728 24808 17759
rect 25498 17756 25504 17808
rect 25556 17796 25562 17808
rect 26620 17796 26648 17836
rect 27522 17824 27528 17836
rect 27580 17824 27586 17876
rect 30101 17867 30159 17873
rect 30101 17833 30113 17867
rect 30147 17864 30159 17867
rect 31386 17864 31392 17876
rect 30147 17836 31392 17864
rect 30147 17833 30159 17836
rect 30101 17827 30159 17833
rect 31386 17824 31392 17836
rect 31444 17864 31450 17876
rect 31938 17864 31944 17876
rect 31444 17836 31944 17864
rect 31444 17824 31450 17836
rect 31938 17824 31944 17836
rect 31996 17864 32002 17876
rect 32309 17867 32367 17873
rect 32309 17864 32321 17867
rect 31996 17836 32321 17864
rect 31996 17824 32002 17836
rect 32309 17833 32321 17836
rect 32355 17833 32367 17867
rect 32309 17827 32367 17833
rect 32490 17824 32496 17876
rect 32548 17864 32554 17876
rect 34146 17864 34152 17876
rect 32548 17836 34152 17864
rect 32548 17824 32554 17836
rect 34146 17824 34152 17836
rect 34204 17824 34210 17876
rect 35342 17824 35348 17876
rect 35400 17824 35406 17876
rect 36446 17824 36452 17876
rect 36504 17824 36510 17876
rect 37826 17824 37832 17876
rect 37884 17864 37890 17876
rect 38289 17867 38347 17873
rect 38289 17864 38301 17867
rect 37884 17836 38301 17864
rect 37884 17824 37890 17836
rect 38289 17833 38301 17836
rect 38335 17833 38347 17867
rect 38289 17827 38347 17833
rect 25556 17768 26648 17796
rect 25556 17756 25562 17768
rect 27154 17756 27160 17808
rect 27212 17796 27218 17808
rect 27709 17799 27767 17805
rect 27709 17796 27721 17799
rect 27212 17768 27721 17796
rect 27212 17756 27218 17768
rect 27709 17765 27721 17768
rect 27755 17765 27767 17799
rect 27709 17759 27767 17765
rect 28166 17756 28172 17808
rect 28224 17796 28230 17808
rect 28353 17799 28411 17805
rect 28353 17796 28365 17799
rect 28224 17768 28365 17796
rect 28224 17756 28230 17768
rect 28353 17765 28365 17768
rect 28399 17765 28411 17799
rect 28353 17759 28411 17765
rect 30742 17756 30748 17808
rect 30800 17796 30806 17808
rect 32582 17796 32588 17808
rect 30800 17768 32588 17796
rect 30800 17756 30806 17768
rect 32582 17756 32588 17768
rect 32640 17756 32646 17808
rect 33965 17799 34023 17805
rect 33965 17765 33977 17799
rect 34011 17765 34023 17799
rect 33965 17759 34023 17765
rect 19306 17700 21036 17728
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17629 18751 17663
rect 18693 17623 18751 17629
rect 18874 17620 18880 17672
rect 18932 17620 18938 17672
rect 19058 17620 19064 17672
rect 19116 17660 19122 17672
rect 19518 17660 19524 17672
rect 19116 17632 19524 17660
rect 19116 17620 19122 17632
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 20625 17663 20683 17669
rect 20625 17629 20637 17663
rect 20671 17660 20683 17663
rect 20714 17660 20720 17672
rect 20671 17632 20720 17660
rect 20671 17629 20683 17632
rect 20625 17623 20683 17629
rect 17788 17592 17816 17620
rect 16776 17564 17816 17592
rect 16393 17555 16451 17561
rect 19150 17552 19156 17604
rect 19208 17592 19214 17604
rect 19628 17592 19656 17623
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 20898 17620 20904 17672
rect 20956 17620 20962 17672
rect 21008 17660 21036 17700
rect 23952 17700 24808 17728
rect 24857 17731 24915 17737
rect 21008 17632 22146 17660
rect 19208 17564 19656 17592
rect 19208 17552 19214 17564
rect 20806 17552 20812 17604
rect 20864 17552 20870 17604
rect 21266 17552 21272 17604
rect 21324 17592 21330 17604
rect 21453 17595 21511 17601
rect 21453 17592 21465 17595
rect 21324 17564 21465 17592
rect 21324 17552 21330 17564
rect 21453 17561 21465 17564
rect 21499 17561 21511 17595
rect 21453 17555 21511 17561
rect 21637 17595 21695 17601
rect 21637 17561 21649 17595
rect 21683 17592 21695 17595
rect 22002 17592 22008 17604
rect 21683 17564 22008 17592
rect 21683 17561 21695 17564
rect 21637 17555 21695 17561
rect 22002 17552 22008 17564
rect 22060 17552 22066 17604
rect 22118 17592 22146 17632
rect 22830 17620 22836 17672
rect 22888 17620 22894 17672
rect 23109 17663 23167 17669
rect 23109 17629 23121 17663
rect 23155 17660 23167 17663
rect 23198 17660 23204 17672
rect 23155 17632 23204 17660
rect 23155 17629 23167 17632
rect 23109 17623 23167 17629
rect 23198 17620 23204 17632
rect 23256 17620 23262 17672
rect 23753 17663 23811 17669
rect 23753 17629 23765 17663
rect 23799 17654 23811 17663
rect 23952 17660 23980 17700
rect 24857 17697 24869 17731
rect 24903 17697 24915 17731
rect 30834 17728 30840 17740
rect 24857 17691 24915 17697
rect 27172 17700 30840 17728
rect 24044 17669 24164 17670
rect 23860 17654 23980 17660
rect 23799 17632 23980 17654
rect 24029 17663 24164 17669
rect 23799 17629 23888 17632
rect 23753 17626 23888 17629
rect 24029 17629 24041 17663
rect 24075 17660 24164 17663
rect 24578 17660 24584 17672
rect 24075 17642 24584 17660
rect 24075 17629 24087 17642
rect 24136 17632 24584 17642
rect 23753 17623 23811 17626
rect 24029 17623 24087 17629
rect 24578 17620 24584 17632
rect 24636 17620 24642 17672
rect 24670 17620 24676 17672
rect 24728 17620 24734 17672
rect 24762 17620 24768 17672
rect 24820 17660 24826 17672
rect 24872 17660 24900 17691
rect 24820 17632 24900 17660
rect 24820 17620 24826 17632
rect 25774 17620 25780 17672
rect 25832 17620 25838 17672
rect 26326 17620 26332 17672
rect 26384 17660 26390 17672
rect 27172 17669 27200 17700
rect 30834 17688 30840 17700
rect 30892 17688 30898 17740
rect 30926 17688 30932 17740
rect 30984 17728 30990 17740
rect 31662 17728 31668 17740
rect 30984 17700 31668 17728
rect 30984 17688 30990 17700
rect 31662 17688 31668 17700
rect 31720 17728 31726 17740
rect 32309 17731 32367 17737
rect 32309 17728 32321 17731
rect 31720 17700 32321 17728
rect 31720 17688 31726 17700
rect 32309 17697 32321 17700
rect 32355 17697 32367 17731
rect 32309 17691 32367 17697
rect 32950 17688 32956 17740
rect 33008 17728 33014 17740
rect 33594 17728 33600 17740
rect 33008 17700 33600 17728
rect 33008 17688 33014 17700
rect 33594 17688 33600 17700
rect 33652 17688 33658 17740
rect 27614 17669 27620 17672
rect 27157 17663 27215 17669
rect 26384 17632 26740 17660
rect 26384 17620 26390 17632
rect 23017 17595 23075 17601
rect 23017 17592 23029 17595
rect 22118 17564 23029 17592
rect 23017 17561 23029 17564
rect 23063 17592 23075 17595
rect 23934 17592 23940 17604
rect 23063 17564 23940 17592
rect 23063 17561 23075 17564
rect 23017 17555 23075 17561
rect 23934 17552 23940 17564
rect 23992 17552 23998 17604
rect 26602 17552 26608 17604
rect 26660 17552 26666 17604
rect 26712 17592 26740 17632
rect 27157 17629 27169 17663
rect 27203 17629 27215 17663
rect 27577 17663 27620 17669
rect 27157 17623 27215 17629
rect 27264 17632 27476 17660
rect 27264 17592 27292 17632
rect 26712 17564 27292 17592
rect 27338 17552 27344 17604
rect 27396 17552 27402 17604
rect 27448 17601 27476 17632
rect 27577 17629 27589 17663
rect 27672 17660 27678 17672
rect 27672 17632 28948 17660
rect 27577 17623 27620 17629
rect 27614 17620 27620 17623
rect 27672 17620 27678 17632
rect 27433 17595 27491 17601
rect 27433 17561 27445 17595
rect 27479 17592 27491 17595
rect 27982 17592 27988 17604
rect 27479 17564 27988 17592
rect 27479 17561 27491 17564
rect 27433 17555 27491 17561
rect 27982 17552 27988 17564
rect 28040 17552 28046 17604
rect 28626 17552 28632 17604
rect 28684 17552 28690 17604
rect 28920 17601 28948 17632
rect 29730 17620 29736 17672
rect 29788 17620 29794 17672
rect 30558 17620 30564 17672
rect 30616 17620 30622 17672
rect 31386 17620 31392 17672
rect 31444 17620 31450 17672
rect 31478 17620 31484 17672
rect 31536 17660 31542 17672
rect 31941 17663 31999 17669
rect 31941 17660 31953 17663
rect 31536 17632 31953 17660
rect 31536 17620 31542 17632
rect 31941 17629 31953 17632
rect 31987 17629 31999 17663
rect 31941 17623 31999 17629
rect 32030 17620 32036 17672
rect 32088 17660 32094 17672
rect 32214 17660 32220 17672
rect 32088 17632 32220 17660
rect 32088 17620 32094 17632
rect 32214 17620 32220 17632
rect 32272 17660 32278 17672
rect 32858 17660 32864 17672
rect 32272 17632 32864 17660
rect 32272 17620 32278 17632
rect 32858 17620 32864 17632
rect 32916 17620 32922 17672
rect 33318 17620 33324 17672
rect 33376 17620 33382 17672
rect 33410 17620 33416 17672
rect 33468 17620 33474 17672
rect 33502 17620 33508 17672
rect 33560 17660 33566 17672
rect 33560 17632 33640 17660
rect 33560 17620 33566 17632
rect 28905 17595 28963 17601
rect 28905 17561 28917 17595
rect 28951 17592 28963 17595
rect 28951 17564 29224 17592
rect 28951 17561 28963 17564
rect 28905 17555 28963 17561
rect 15470 17484 15476 17536
rect 15528 17524 15534 17536
rect 16206 17524 16212 17536
rect 15528 17496 16212 17524
rect 15528 17484 15534 17496
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 16298 17484 16304 17536
rect 16356 17524 16362 17536
rect 19521 17527 19579 17533
rect 19521 17524 19533 17527
rect 16356 17496 19533 17524
rect 16356 17484 16362 17496
rect 19521 17493 19533 17496
rect 19567 17493 19579 17527
rect 19521 17487 19579 17493
rect 20898 17484 20904 17536
rect 20956 17524 20962 17536
rect 21821 17527 21879 17533
rect 21821 17524 21833 17527
rect 20956 17496 21833 17524
rect 20956 17484 20962 17496
rect 21821 17493 21833 17496
rect 21867 17493 21879 17527
rect 21821 17487 21879 17493
rect 26970 17484 26976 17536
rect 27028 17524 27034 17536
rect 28350 17524 28356 17536
rect 27028 17496 28356 17524
rect 27028 17484 27034 17496
rect 28350 17484 28356 17496
rect 28408 17484 28414 17536
rect 28534 17484 28540 17536
rect 28592 17524 28598 17536
rect 28813 17527 28871 17533
rect 28813 17524 28825 17527
rect 28592 17496 28825 17524
rect 28592 17484 28598 17496
rect 28813 17493 28825 17496
rect 28859 17493 28871 17527
rect 29196 17524 29224 17564
rect 29270 17552 29276 17604
rect 29328 17592 29334 17604
rect 29917 17595 29975 17601
rect 29917 17592 29929 17595
rect 29328 17564 29929 17592
rect 29328 17552 29334 17564
rect 29917 17561 29929 17564
rect 29963 17561 29975 17595
rect 29917 17555 29975 17561
rect 31294 17552 31300 17604
rect 31352 17592 31358 17604
rect 33612 17601 33640 17632
rect 33778 17620 33784 17672
rect 33836 17669 33842 17672
rect 33836 17660 33844 17669
rect 33980 17660 34008 17759
rect 34054 17756 34060 17808
rect 34112 17796 34118 17808
rect 34112 17768 36032 17796
rect 34112 17756 34118 17768
rect 34698 17688 34704 17740
rect 34756 17728 34762 17740
rect 36004 17737 36032 17768
rect 34885 17731 34943 17737
rect 34885 17728 34897 17731
rect 34756 17700 34897 17728
rect 34756 17688 34762 17700
rect 34885 17697 34897 17700
rect 34931 17697 34943 17731
rect 34885 17691 34943 17697
rect 35989 17731 36047 17737
rect 35989 17697 36001 17731
rect 36035 17728 36047 17731
rect 36722 17728 36728 17740
rect 36035 17700 36728 17728
rect 36035 17697 36047 17700
rect 35989 17691 36047 17697
rect 36722 17688 36728 17700
rect 36780 17688 36786 17740
rect 35069 17663 35127 17669
rect 35069 17660 35081 17663
rect 33836 17632 33881 17660
rect 33980 17632 35081 17660
rect 33836 17623 33844 17632
rect 35069 17629 35081 17632
rect 35115 17629 35127 17663
rect 35069 17623 35127 17629
rect 33836 17620 33842 17623
rect 35158 17620 35164 17672
rect 35216 17620 35222 17672
rect 35437 17663 35495 17669
rect 35437 17629 35449 17663
rect 35483 17629 35495 17663
rect 35437 17623 35495 17629
rect 33597 17595 33655 17601
rect 31352 17564 33548 17592
rect 31352 17552 31358 17564
rect 29638 17524 29644 17536
rect 29196 17496 29644 17524
rect 28813 17487 28871 17493
rect 29638 17484 29644 17496
rect 29696 17524 29702 17536
rect 30558 17524 30564 17536
rect 29696 17496 30564 17524
rect 29696 17484 29702 17496
rect 30558 17484 30564 17496
rect 30616 17484 30622 17536
rect 32125 17527 32183 17533
rect 32125 17493 32137 17527
rect 32171 17524 32183 17527
rect 33410 17524 33416 17536
rect 32171 17496 33416 17524
rect 32171 17493 32183 17496
rect 32125 17487 32183 17493
rect 33410 17484 33416 17496
rect 33468 17484 33474 17536
rect 33520 17524 33548 17564
rect 33597 17561 33609 17595
rect 33643 17561 33655 17595
rect 33597 17555 33655 17561
rect 33686 17552 33692 17604
rect 33744 17552 33750 17604
rect 35452 17592 35480 17623
rect 36078 17620 36084 17672
rect 36136 17620 36142 17672
rect 36538 17620 36544 17672
rect 36596 17660 36602 17672
rect 36814 17660 36820 17672
rect 36596 17632 36820 17660
rect 36596 17620 36602 17632
rect 36814 17620 36820 17632
rect 36872 17660 36878 17672
rect 36909 17663 36967 17669
rect 36909 17660 36921 17663
rect 36872 17632 36921 17660
rect 36872 17620 36878 17632
rect 36909 17629 36921 17632
rect 36955 17629 36967 17663
rect 36909 17623 36967 17629
rect 37176 17663 37234 17669
rect 37176 17629 37188 17663
rect 37222 17660 37234 17663
rect 37458 17660 37464 17672
rect 37222 17632 37464 17660
rect 37222 17629 37234 17632
rect 37176 17623 37234 17629
rect 37458 17620 37464 17632
rect 37516 17620 37522 17672
rect 34808 17564 35480 17592
rect 34808 17524 34836 17564
rect 33520 17496 34836 17524
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 15194 17280 15200 17332
rect 15252 17280 15258 17332
rect 19058 17320 19064 17332
rect 17236 17292 19064 17320
rect 15470 17252 15476 17264
rect 14936 17224 15476 17252
rect 14936 17193 14964 17224
rect 15470 17212 15476 17224
rect 15528 17212 15534 17264
rect 14921 17187 14979 17193
rect 14921 17153 14933 17187
rect 14967 17153 14979 17187
rect 14921 17147 14979 17153
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17184 15071 17187
rect 15657 17187 15715 17193
rect 15657 17184 15669 17187
rect 15059 17156 15669 17184
rect 15059 17153 15071 17156
rect 15013 17147 15071 17153
rect 15657 17153 15669 17156
rect 15703 17153 15715 17187
rect 15657 17147 15715 17153
rect 15838 17144 15844 17196
rect 15896 17144 15902 17196
rect 15930 17144 15936 17196
rect 15988 17144 15994 17196
rect 16114 17144 16120 17196
rect 16172 17144 16178 17196
rect 16209 17187 16267 17193
rect 16209 17153 16221 17187
rect 16255 17184 16267 17187
rect 16298 17184 16304 17196
rect 16255 17156 16304 17184
rect 16255 17153 16267 17156
rect 16209 17147 16267 17153
rect 16022 17076 16028 17128
rect 16080 17116 16086 17128
rect 16224 17116 16252 17147
rect 16298 17144 16304 17156
rect 16356 17144 16362 17196
rect 17236 17193 17264 17292
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 22103 17323 22161 17329
rect 22103 17289 22115 17323
rect 22149 17320 22161 17323
rect 22278 17320 22284 17332
rect 22149 17292 22284 17320
rect 22149 17289 22161 17292
rect 22103 17283 22161 17289
rect 22278 17280 22284 17292
rect 22336 17280 22342 17332
rect 23017 17323 23075 17329
rect 23017 17289 23029 17323
rect 23063 17320 23075 17323
rect 24486 17320 24492 17332
rect 23063 17292 24492 17320
rect 23063 17289 23075 17292
rect 23017 17283 23075 17289
rect 24486 17280 24492 17292
rect 24544 17280 24550 17332
rect 24857 17323 24915 17329
rect 24857 17289 24869 17323
rect 24903 17320 24915 17323
rect 26694 17320 26700 17332
rect 24903 17292 26700 17320
rect 24903 17289 24915 17292
rect 24857 17283 24915 17289
rect 26694 17280 26700 17292
rect 26752 17280 26758 17332
rect 29914 17320 29920 17332
rect 27356 17292 29920 17320
rect 18046 17212 18052 17264
rect 18104 17252 18110 17264
rect 18966 17252 18972 17264
rect 18104 17224 18972 17252
rect 18104 17212 18110 17224
rect 18966 17212 18972 17224
rect 19024 17252 19030 17264
rect 19613 17255 19671 17261
rect 19613 17252 19625 17255
rect 19024 17224 19625 17252
rect 19024 17212 19030 17224
rect 19613 17221 19625 17224
rect 19659 17221 19671 17255
rect 20254 17252 20260 17264
rect 19613 17215 19671 17221
rect 19812 17224 20260 17252
rect 17221 17187 17279 17193
rect 17221 17153 17233 17187
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 17402 17144 17408 17196
rect 17460 17184 17466 17196
rect 17957 17187 18015 17193
rect 17957 17184 17969 17187
rect 17460 17156 17969 17184
rect 17460 17144 17466 17156
rect 17957 17153 17969 17156
rect 18003 17153 18015 17187
rect 17957 17147 18015 17153
rect 18506 17144 18512 17196
rect 18564 17184 18570 17196
rect 18693 17187 18751 17193
rect 18693 17184 18705 17187
rect 18564 17156 18705 17184
rect 18564 17144 18570 17156
rect 18693 17153 18705 17156
rect 18739 17184 18751 17187
rect 19426 17184 19432 17196
rect 18739 17156 19432 17184
rect 18739 17153 18751 17156
rect 18693 17147 18751 17153
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 19812 17193 19840 17224
rect 20254 17212 20260 17224
rect 20312 17212 20318 17264
rect 21910 17212 21916 17264
rect 21968 17252 21974 17264
rect 22005 17255 22063 17261
rect 22005 17252 22017 17255
rect 21968 17224 22017 17252
rect 21968 17212 21974 17224
rect 22005 17221 22017 17224
rect 22051 17221 22063 17255
rect 22005 17215 22063 17221
rect 22186 17212 22192 17264
rect 22244 17212 22250 17264
rect 22370 17212 22376 17264
rect 22428 17252 22434 17264
rect 26602 17252 26608 17264
rect 22428 17224 26608 17252
rect 22428 17212 22434 17224
rect 19797 17187 19855 17193
rect 19797 17153 19809 17187
rect 19843 17153 19855 17187
rect 19797 17147 19855 17153
rect 19889 17187 19947 17193
rect 19889 17153 19901 17187
rect 19935 17153 19947 17187
rect 19889 17147 19947 17153
rect 16080 17088 16252 17116
rect 16080 17076 16086 17088
rect 17494 17076 17500 17128
rect 17552 17076 17558 17128
rect 18138 17076 18144 17128
rect 18196 17116 18202 17128
rect 18785 17119 18843 17125
rect 18785 17116 18797 17119
rect 18196 17088 18797 17116
rect 18196 17076 18202 17088
rect 18785 17085 18797 17088
rect 18831 17085 18843 17119
rect 18785 17079 18843 17085
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 19904 17116 19932 17147
rect 20162 17144 20168 17196
rect 20220 17184 20226 17196
rect 20438 17184 20444 17196
rect 20220 17156 20444 17184
rect 20220 17144 20226 17156
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 20530 17144 20536 17196
rect 20588 17184 20594 17196
rect 20625 17187 20683 17193
rect 20625 17184 20637 17187
rect 20588 17156 20637 17184
rect 20588 17144 20594 17156
rect 20625 17153 20637 17156
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17184 20867 17187
rect 21634 17184 21640 17196
rect 20855 17156 21640 17184
rect 20855 17153 20867 17156
rect 20809 17147 20867 17153
rect 21634 17144 21640 17156
rect 21692 17144 21698 17196
rect 22281 17187 22339 17193
rect 22281 17153 22293 17187
rect 22327 17184 22339 17187
rect 22646 17184 22652 17196
rect 22327 17156 22652 17184
rect 22327 17153 22339 17156
rect 22281 17147 22339 17153
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 22741 17187 22799 17193
rect 22741 17153 22753 17187
rect 22787 17184 22799 17187
rect 23382 17184 23388 17196
rect 22787 17156 23388 17184
rect 22787 17153 22799 17156
rect 22741 17147 22799 17153
rect 23382 17144 23388 17156
rect 23440 17144 23446 17196
rect 23492 17193 23520 17224
rect 26602 17212 26608 17224
rect 26660 17212 26666 17264
rect 27356 17196 27384 17292
rect 29914 17280 29920 17292
rect 29972 17280 29978 17332
rect 30009 17323 30067 17329
rect 30009 17289 30021 17323
rect 30055 17320 30067 17323
rect 30098 17320 30104 17332
rect 30055 17292 30104 17320
rect 30055 17289 30067 17292
rect 30009 17283 30067 17289
rect 30098 17280 30104 17292
rect 30156 17280 30162 17332
rect 33873 17323 33931 17329
rect 33873 17289 33885 17323
rect 33919 17320 33931 17323
rect 35158 17320 35164 17332
rect 33919 17292 35164 17320
rect 33919 17289 33931 17292
rect 33873 17283 33931 17289
rect 35158 17280 35164 17292
rect 35216 17280 35222 17332
rect 37826 17280 37832 17332
rect 37884 17280 37890 17332
rect 29178 17212 29184 17264
rect 29236 17252 29242 17264
rect 29730 17252 29736 17264
rect 29236 17224 29736 17252
rect 29236 17212 29242 17224
rect 29730 17212 29736 17224
rect 29788 17212 29794 17264
rect 30116 17252 30144 17280
rect 31294 17252 31300 17264
rect 30116 17224 31300 17252
rect 23477 17187 23535 17193
rect 23477 17153 23489 17187
rect 23523 17153 23535 17187
rect 23733 17187 23791 17193
rect 23733 17184 23745 17187
rect 23477 17147 23535 17153
rect 23584 17156 23745 17184
rect 19392 17088 19932 17116
rect 23017 17119 23075 17125
rect 19392 17076 19398 17088
rect 23017 17085 23029 17119
rect 23063 17116 23075 17119
rect 23106 17116 23112 17128
rect 23063 17088 23112 17116
rect 23063 17085 23075 17088
rect 23017 17079 23075 17085
rect 23106 17076 23112 17088
rect 23164 17076 23170 17128
rect 23198 17076 23204 17128
rect 23256 17116 23262 17128
rect 23584 17116 23612 17156
rect 23733 17153 23745 17156
rect 23779 17153 23791 17187
rect 23733 17147 23791 17153
rect 25685 17187 25743 17193
rect 25685 17153 25697 17187
rect 25731 17184 25743 17187
rect 25731 17156 27200 17184
rect 25731 17153 25743 17156
rect 25685 17147 25743 17153
rect 23256 17088 23612 17116
rect 25573 17119 25631 17125
rect 23256 17076 23262 17088
rect 25573 17085 25585 17119
rect 25619 17116 25631 17119
rect 25961 17119 26019 17125
rect 25619 17088 25912 17116
rect 25619 17085 25631 17088
rect 25573 17079 25631 17085
rect 15010 17008 15016 17060
rect 15068 17048 15074 17060
rect 18046 17048 18052 17060
rect 15068 17020 18052 17048
rect 15068 17008 15074 17020
rect 18046 17008 18052 17020
rect 18104 17008 18110 17060
rect 18233 17051 18291 17057
rect 18233 17017 18245 17051
rect 18279 17048 18291 17051
rect 18874 17048 18880 17060
rect 18279 17020 18880 17048
rect 18279 17017 18291 17020
rect 18233 17011 18291 17017
rect 18874 17008 18880 17020
rect 18932 17008 18938 17060
rect 20073 17051 20131 17057
rect 20073 17017 20085 17051
rect 20119 17048 20131 17051
rect 21266 17048 21272 17060
rect 20119 17020 21272 17048
rect 20119 17017 20131 17020
rect 20073 17011 20131 17017
rect 21266 17008 21272 17020
rect 21324 17008 21330 17060
rect 25409 17051 25467 17057
rect 25409 17048 25421 17051
rect 24412 17020 25421 17048
rect 17034 16940 17040 16992
rect 17092 16940 17098 16992
rect 17405 16983 17463 16989
rect 17405 16949 17417 16983
rect 17451 16980 17463 16983
rect 19150 16980 19156 16992
rect 17451 16952 19156 16980
rect 17451 16949 17463 16952
rect 17405 16943 17463 16949
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 20806 16940 20812 16992
rect 20864 16980 20870 16992
rect 20901 16983 20959 16989
rect 20901 16980 20913 16983
rect 20864 16952 20913 16980
rect 20864 16940 20870 16952
rect 20901 16949 20913 16952
rect 20947 16949 20959 16983
rect 20901 16943 20959 16949
rect 22833 16983 22891 16989
rect 22833 16949 22845 16983
rect 22879 16980 22891 16983
rect 23014 16980 23020 16992
rect 22879 16952 23020 16980
rect 22879 16949 22891 16952
rect 22833 16943 22891 16949
rect 23014 16940 23020 16952
rect 23072 16940 23078 16992
rect 23842 16940 23848 16992
rect 23900 16980 23906 16992
rect 24412 16980 24440 17020
rect 25409 17017 25421 17020
rect 25455 17017 25467 17051
rect 25409 17011 25467 17017
rect 23900 16952 24440 16980
rect 25884 16980 25912 17088
rect 25961 17085 25973 17119
rect 26007 17085 26019 17119
rect 25961 17079 26019 17085
rect 25976 17048 26004 17079
rect 26050 17076 26056 17128
rect 26108 17076 26114 17128
rect 27172 17125 27200 17156
rect 27338 17144 27344 17196
rect 27396 17144 27402 17196
rect 27433 17187 27491 17193
rect 27433 17153 27445 17187
rect 27479 17184 27491 17187
rect 27706 17184 27712 17196
rect 27479 17156 27712 17184
rect 27479 17153 27491 17156
rect 27433 17147 27491 17153
rect 27706 17144 27712 17156
rect 27764 17144 27770 17196
rect 28534 17144 28540 17196
rect 28592 17184 28598 17196
rect 28629 17187 28687 17193
rect 28629 17184 28641 17187
rect 28592 17156 28641 17184
rect 28592 17144 28598 17156
rect 28629 17153 28641 17156
rect 28675 17153 28687 17187
rect 28629 17147 28687 17153
rect 28896 17187 28954 17193
rect 28896 17153 28908 17187
rect 28942 17184 28954 17187
rect 28942 17156 30604 17184
rect 28942 17153 28954 17156
rect 28896 17147 28954 17153
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17085 27215 17119
rect 27157 17079 27215 17085
rect 27522 17076 27528 17128
rect 27580 17076 27586 17128
rect 27614 17076 27620 17128
rect 27672 17076 27678 17128
rect 26142 17048 26148 17060
rect 25976 17020 26148 17048
rect 26142 17008 26148 17020
rect 26200 17048 26206 17060
rect 27632 17048 27660 17076
rect 26200 17020 27660 17048
rect 30576 17048 30604 17156
rect 30650 17144 30656 17196
rect 30708 17144 30714 17196
rect 30742 17144 30748 17196
rect 30800 17144 30806 17196
rect 30926 17144 30932 17196
rect 30984 17144 30990 17196
rect 31036 17193 31064 17224
rect 31294 17212 31300 17224
rect 31352 17212 31358 17264
rect 32674 17212 32680 17264
rect 32732 17252 32738 17264
rect 32732 17224 32904 17252
rect 32732 17212 32738 17224
rect 31202 17193 31208 17196
rect 31021 17187 31079 17193
rect 31021 17153 31033 17187
rect 31067 17153 31079 17187
rect 31021 17147 31079 17153
rect 31159 17187 31208 17193
rect 31159 17153 31171 17187
rect 31205 17153 31208 17187
rect 31159 17147 31208 17153
rect 31202 17144 31208 17147
rect 31260 17144 31266 17196
rect 31846 17144 31852 17196
rect 31904 17184 31910 17196
rect 32306 17184 32312 17196
rect 31904 17156 32312 17184
rect 31904 17144 31910 17156
rect 32306 17144 32312 17156
rect 32364 17184 32370 17196
rect 32493 17187 32551 17193
rect 32493 17184 32505 17187
rect 32364 17156 32505 17184
rect 32364 17144 32370 17156
rect 32493 17153 32505 17156
rect 32539 17153 32551 17187
rect 32876 17184 32904 17224
rect 33226 17212 33232 17264
rect 33284 17252 33290 17264
rect 33505 17255 33563 17261
rect 33505 17252 33517 17255
rect 33284 17224 33517 17252
rect 33284 17212 33290 17224
rect 33505 17221 33517 17224
rect 33551 17221 33563 17255
rect 33505 17215 33563 17221
rect 33594 17212 33600 17264
rect 33652 17212 33658 17264
rect 34333 17255 34391 17261
rect 34333 17221 34345 17255
rect 34379 17252 34391 17255
rect 37921 17255 37979 17261
rect 37921 17252 37933 17255
rect 34379 17224 37933 17252
rect 34379 17221 34391 17224
rect 34333 17215 34391 17221
rect 33321 17187 33379 17193
rect 33321 17184 33333 17187
rect 32876 17156 33333 17184
rect 32493 17147 32551 17153
rect 33321 17153 33333 17156
rect 33367 17153 33379 17187
rect 33321 17147 33379 17153
rect 33689 17187 33747 17193
rect 33689 17153 33701 17187
rect 33735 17184 33747 17187
rect 34238 17184 34244 17196
rect 33735 17156 34244 17184
rect 33735 17153 33747 17156
rect 33689 17147 33747 17153
rect 34238 17144 34244 17156
rect 34296 17144 34302 17196
rect 34514 17144 34520 17196
rect 34572 17144 34578 17196
rect 34606 17144 34612 17196
rect 34664 17144 34670 17196
rect 35544 17193 35572 17224
rect 37921 17221 37933 17224
rect 37967 17221 37979 17255
rect 37921 17215 37979 17221
rect 34885 17187 34943 17193
rect 34885 17153 34897 17187
rect 34931 17153 34943 17187
rect 34885 17147 34943 17153
rect 35529 17187 35587 17193
rect 35529 17153 35541 17187
rect 35575 17153 35587 17187
rect 35529 17147 35587 17153
rect 31662 17076 31668 17128
rect 31720 17116 31726 17128
rect 32401 17119 32459 17125
rect 32401 17116 32413 17119
rect 31720 17088 32413 17116
rect 31720 17076 31726 17088
rect 32401 17085 32413 17088
rect 32447 17085 32459 17119
rect 32401 17079 32459 17085
rect 32582 17076 32588 17128
rect 32640 17116 32646 17128
rect 34900 17116 34928 17147
rect 36354 17144 36360 17196
rect 36412 17184 36418 17196
rect 36449 17187 36507 17193
rect 36449 17184 36461 17187
rect 36412 17156 36461 17184
rect 36412 17144 36418 17156
rect 36449 17153 36461 17156
rect 36495 17153 36507 17187
rect 38838 17184 38844 17196
rect 36449 17147 36507 17153
rect 37936 17156 38844 17184
rect 32640 17088 34928 17116
rect 35805 17119 35863 17125
rect 32640 17076 32646 17088
rect 35805 17085 35817 17119
rect 35851 17085 35863 17119
rect 35805 17079 35863 17085
rect 36725 17119 36783 17125
rect 36725 17085 36737 17119
rect 36771 17116 36783 17119
rect 37936 17116 37964 17156
rect 38838 17144 38844 17156
rect 38896 17144 38902 17196
rect 36771 17088 37964 17116
rect 36771 17085 36783 17088
rect 36725 17079 36783 17085
rect 31846 17048 31852 17060
rect 30576 17020 31852 17048
rect 26200 17008 26206 17020
rect 31846 17008 31852 17020
rect 31904 17008 31910 17060
rect 34793 17051 34851 17057
rect 34793 17017 34805 17051
rect 34839 17048 34851 17051
rect 35342 17048 35348 17060
rect 34839 17020 35348 17048
rect 34839 17017 34851 17020
rect 34793 17011 34851 17017
rect 35342 17008 35348 17020
rect 35400 17008 35406 17060
rect 35820 17048 35848 17079
rect 38102 17076 38108 17128
rect 38160 17076 38166 17128
rect 39022 17048 39028 17060
rect 35820 17020 39028 17048
rect 39022 17008 39028 17020
rect 39080 17008 39086 17060
rect 29000 16980 29006 16992
rect 25884 16952 29006 16980
rect 23900 16940 23906 16952
rect 29000 16940 29006 16952
rect 29058 16940 29064 16992
rect 31297 16983 31355 16989
rect 31297 16949 31309 16983
rect 31343 16980 31355 16983
rect 31478 16980 31484 16992
rect 31343 16952 31484 16980
rect 31343 16949 31355 16952
rect 31297 16943 31355 16949
rect 31478 16940 31484 16952
rect 31536 16940 31542 16992
rect 31662 16940 31668 16992
rect 31720 16980 31726 16992
rect 32769 16983 32827 16989
rect 32769 16980 32781 16983
rect 31720 16952 32781 16980
rect 31720 16940 31726 16952
rect 32769 16949 32781 16952
rect 32815 16949 32827 16983
rect 32769 16943 32827 16949
rect 37090 16940 37096 16992
rect 37148 16980 37154 16992
rect 37461 16983 37519 16989
rect 37461 16980 37473 16983
rect 37148 16952 37473 16980
rect 37148 16940 37154 16952
rect 37461 16949 37473 16952
rect 37507 16949 37519 16983
rect 37461 16943 37519 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 15010 16736 15016 16788
rect 15068 16736 15074 16788
rect 16206 16736 16212 16788
rect 16264 16776 16270 16788
rect 16264 16748 16436 16776
rect 16264 16736 16270 16748
rect 15838 16668 15844 16720
rect 15896 16708 15902 16720
rect 16408 16717 16436 16748
rect 16850 16736 16856 16788
rect 16908 16776 16914 16788
rect 17494 16776 17500 16788
rect 16908 16748 17500 16776
rect 16908 16736 16914 16748
rect 17494 16736 17500 16748
rect 17552 16776 17558 16788
rect 22002 16776 22008 16788
rect 17552 16748 22008 16776
rect 17552 16736 17558 16748
rect 22002 16736 22008 16748
rect 22060 16736 22066 16788
rect 22646 16736 22652 16788
rect 22704 16776 22710 16788
rect 23845 16779 23903 16785
rect 23845 16776 23857 16779
rect 22704 16748 23857 16776
rect 22704 16736 22710 16748
rect 23845 16745 23857 16748
rect 23891 16745 23903 16779
rect 23845 16739 23903 16745
rect 24949 16779 25007 16785
rect 24949 16745 24961 16779
rect 24995 16776 25007 16779
rect 27706 16776 27712 16788
rect 24995 16748 27712 16776
rect 24995 16745 25007 16748
rect 24949 16739 25007 16745
rect 16393 16711 16451 16717
rect 15896 16680 16344 16708
rect 15896 16668 15902 16680
rect 16316 16640 16344 16680
rect 16393 16677 16405 16711
rect 16439 16677 16451 16711
rect 17681 16711 17739 16717
rect 17681 16708 17693 16711
rect 16393 16671 16451 16677
rect 16592 16680 17693 16708
rect 16485 16643 16543 16649
rect 16485 16640 16497 16643
rect 16316 16612 16497 16640
rect 16485 16609 16497 16612
rect 16531 16609 16543 16643
rect 16485 16603 16543 16609
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16572 15899 16575
rect 16022 16572 16028 16584
rect 15887 16544 16028 16572
rect 15887 16541 15899 16544
rect 15841 16535 15899 16541
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 16114 16532 16120 16584
rect 16172 16572 16178 16584
rect 16209 16575 16267 16581
rect 16209 16572 16221 16575
rect 16172 16544 16221 16572
rect 16172 16532 16178 16544
rect 16209 16541 16221 16544
rect 16255 16572 16267 16575
rect 16592 16572 16620 16680
rect 17681 16677 17693 16680
rect 17727 16677 17739 16711
rect 17681 16671 17739 16677
rect 19426 16668 19432 16720
rect 19484 16708 19490 16720
rect 19484 16680 21496 16708
rect 19484 16668 19490 16680
rect 16666 16600 16672 16652
rect 16724 16640 16730 16652
rect 16724 16612 16804 16640
rect 16724 16600 16730 16612
rect 16776 16581 16804 16612
rect 18414 16600 18420 16652
rect 18472 16600 18478 16652
rect 20257 16643 20315 16649
rect 20257 16609 20269 16643
rect 20303 16640 20315 16643
rect 21358 16640 21364 16652
rect 20303 16612 21364 16640
rect 20303 16609 20315 16612
rect 20257 16603 20315 16609
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 21468 16640 21496 16680
rect 22005 16643 22063 16649
rect 22005 16640 22017 16643
rect 21468 16612 22017 16640
rect 22005 16609 22017 16612
rect 22051 16609 22063 16643
rect 22005 16603 22063 16609
rect 25498 16600 25504 16652
rect 25556 16640 25562 16652
rect 25556 16612 25820 16640
rect 25556 16600 25562 16612
rect 16255 16544 16620 16572
rect 16761 16575 16819 16581
rect 16255 16541 16267 16544
rect 16209 16535 16267 16541
rect 16761 16541 16773 16575
rect 16807 16541 16819 16575
rect 16761 16535 16819 16541
rect 17586 16532 17592 16584
rect 17644 16532 17650 16584
rect 18046 16532 18052 16584
rect 18104 16572 18110 16584
rect 18141 16575 18199 16581
rect 18141 16572 18153 16575
rect 18104 16544 18153 16572
rect 18104 16532 18110 16544
rect 18141 16541 18153 16544
rect 18187 16541 18199 16575
rect 18141 16535 18199 16541
rect 20349 16575 20407 16581
rect 20349 16541 20361 16575
rect 20395 16541 20407 16575
rect 20349 16535 20407 16541
rect 14829 16507 14887 16513
rect 14829 16473 14841 16507
rect 14875 16504 14887 16507
rect 16574 16504 16580 16516
rect 14875 16476 16580 16504
rect 14875 16473 14887 16476
rect 14829 16467 14887 16473
rect 16574 16464 16580 16476
rect 16632 16464 16638 16516
rect 20364 16504 20392 16535
rect 20438 16532 20444 16584
rect 20496 16572 20502 16584
rect 20533 16575 20591 16581
rect 20533 16572 20545 16575
rect 20496 16544 20545 16572
rect 20496 16532 20502 16544
rect 20533 16541 20545 16544
rect 20579 16541 20591 16575
rect 20533 16535 20591 16541
rect 21726 16532 21732 16584
rect 21784 16572 21790 16584
rect 22370 16572 22376 16584
rect 21784 16544 22376 16572
rect 21784 16532 21790 16544
rect 22370 16532 22376 16544
rect 22428 16532 22434 16584
rect 23845 16575 23903 16581
rect 23845 16541 23857 16575
rect 23891 16572 23903 16575
rect 23934 16572 23940 16584
rect 23891 16544 23940 16572
rect 23891 16541 23903 16544
rect 23845 16535 23903 16541
rect 23934 16532 23940 16544
rect 23992 16532 23998 16584
rect 24029 16575 24087 16581
rect 24029 16541 24041 16575
rect 24075 16572 24087 16575
rect 24394 16572 24400 16584
rect 24075 16544 24400 16572
rect 24075 16541 24087 16544
rect 24029 16535 24087 16541
rect 24394 16532 24400 16544
rect 24452 16532 24458 16584
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16572 24639 16575
rect 25682 16572 25688 16584
rect 24627 16544 25688 16572
rect 24627 16541 24639 16544
rect 24581 16535 24639 16541
rect 25682 16532 25688 16544
rect 25740 16532 25746 16584
rect 25792 16581 25820 16612
rect 25884 16581 25912 16748
rect 27706 16736 27712 16748
rect 27764 16736 27770 16788
rect 28626 16736 28632 16788
rect 28684 16776 28690 16788
rect 29086 16776 29092 16788
rect 28684 16748 29092 16776
rect 28684 16736 28690 16748
rect 29086 16736 29092 16748
rect 29144 16736 29150 16788
rect 30098 16736 30104 16788
rect 30156 16776 30162 16788
rect 30193 16779 30251 16785
rect 30193 16776 30205 16779
rect 30156 16748 30205 16776
rect 30156 16736 30162 16748
rect 30193 16745 30205 16748
rect 30239 16745 30251 16779
rect 31570 16776 31576 16788
rect 30193 16739 30251 16745
rect 30852 16748 31576 16776
rect 26053 16711 26111 16717
rect 26053 16677 26065 16711
rect 26099 16708 26111 16711
rect 28445 16711 28503 16717
rect 26099 16680 28396 16708
rect 26099 16677 26111 16680
rect 26053 16671 26111 16677
rect 27341 16643 27399 16649
rect 27341 16609 27353 16643
rect 27387 16640 27399 16643
rect 27522 16640 27528 16652
rect 27387 16612 27528 16640
rect 27387 16609 27399 16612
rect 27341 16603 27399 16609
rect 27522 16600 27528 16612
rect 27580 16600 27586 16652
rect 27798 16600 27804 16652
rect 27856 16640 27862 16652
rect 27985 16643 28043 16649
rect 27985 16640 27997 16643
rect 27856 16612 27997 16640
rect 27856 16600 27862 16612
rect 27985 16609 27997 16612
rect 28031 16609 28043 16643
rect 28368 16640 28396 16680
rect 28445 16677 28457 16711
rect 28491 16708 28503 16711
rect 28491 16680 29868 16708
rect 28491 16677 28503 16680
rect 28445 16671 28503 16677
rect 29840 16649 29868 16680
rect 30852 16649 30880 16748
rect 31570 16736 31576 16748
rect 31628 16776 31634 16788
rect 31628 16748 32996 16776
rect 31628 16736 31634 16748
rect 32217 16711 32275 16717
rect 32217 16677 32229 16711
rect 32263 16708 32275 16711
rect 32582 16708 32588 16720
rect 32263 16680 32588 16708
rect 32263 16677 32275 16680
rect 32217 16671 32275 16677
rect 32582 16668 32588 16680
rect 32640 16668 32646 16720
rect 32968 16652 32996 16748
rect 33686 16736 33692 16788
rect 33744 16776 33750 16788
rect 34333 16779 34391 16785
rect 34333 16776 34345 16779
rect 33744 16748 34345 16776
rect 33744 16736 33750 16748
rect 34333 16745 34345 16748
rect 34379 16745 34391 16779
rect 34333 16739 34391 16745
rect 34790 16736 34796 16788
rect 34848 16776 34854 16788
rect 36081 16779 36139 16785
rect 34848 16748 36032 16776
rect 34848 16736 34854 16748
rect 29825 16643 29883 16649
rect 28368 16612 29500 16640
rect 27985 16603 28043 16609
rect 25777 16575 25835 16581
rect 25777 16541 25789 16575
rect 25823 16541 25835 16575
rect 25777 16535 25835 16541
rect 25869 16575 25927 16581
rect 25869 16541 25881 16575
rect 25915 16541 25927 16575
rect 25869 16535 25927 16541
rect 26142 16532 26148 16584
rect 26200 16572 26206 16584
rect 26513 16575 26571 16581
rect 26513 16572 26525 16575
rect 26200 16544 26525 16572
rect 26200 16532 26206 16544
rect 26513 16541 26525 16544
rect 26559 16541 26571 16575
rect 26513 16535 26571 16541
rect 27246 16532 27252 16584
rect 27304 16572 27310 16584
rect 28077 16575 28135 16581
rect 28077 16572 28089 16575
rect 27304 16544 28089 16572
rect 27304 16532 27310 16544
rect 28077 16541 28089 16544
rect 28123 16541 28135 16575
rect 28077 16535 28135 16541
rect 20898 16504 20904 16516
rect 20364 16476 20904 16504
rect 20898 16464 20904 16476
rect 20956 16464 20962 16516
rect 20993 16507 21051 16513
rect 20993 16473 21005 16507
rect 21039 16473 21051 16507
rect 20993 16467 21051 16473
rect 15010 16396 15016 16448
rect 15068 16445 15074 16448
rect 15068 16439 15087 16445
rect 15075 16405 15087 16439
rect 15068 16399 15087 16405
rect 15197 16439 15255 16445
rect 15197 16405 15209 16439
rect 15243 16436 15255 16439
rect 15286 16436 15292 16448
rect 15243 16408 15292 16436
rect 15243 16405 15255 16408
rect 15197 16399 15255 16405
rect 15068 16396 15074 16399
rect 15286 16396 15292 16408
rect 15344 16396 15350 16448
rect 20254 16396 20260 16448
rect 20312 16436 20318 16448
rect 21008 16436 21036 16467
rect 23474 16464 23480 16516
rect 23532 16504 23538 16516
rect 24118 16504 24124 16516
rect 23532 16476 24124 16504
rect 23532 16464 23538 16476
rect 24118 16464 24124 16476
rect 24176 16504 24182 16516
rect 24765 16507 24823 16513
rect 24765 16504 24777 16507
rect 24176 16476 24777 16504
rect 24176 16464 24182 16476
rect 24765 16473 24777 16476
rect 24811 16473 24823 16507
rect 24765 16467 24823 16473
rect 20312 16408 21036 16436
rect 20312 16396 20318 16408
rect 22738 16396 22744 16448
rect 22796 16436 22802 16448
rect 23109 16439 23167 16445
rect 23109 16436 23121 16439
rect 22796 16408 23121 16436
rect 22796 16396 22802 16408
rect 23109 16405 23121 16408
rect 23155 16405 23167 16439
rect 23109 16399 23167 16405
rect 25409 16439 25467 16445
rect 25409 16405 25421 16439
rect 25455 16436 25467 16439
rect 27338 16436 27344 16448
rect 25455 16408 27344 16436
rect 25455 16405 25467 16408
rect 25409 16399 25467 16405
rect 27338 16396 27344 16408
rect 27396 16396 27402 16448
rect 28092 16436 28120 16535
rect 28258 16532 28264 16584
rect 28316 16572 28322 16584
rect 28905 16575 28963 16581
rect 28905 16572 28917 16575
rect 28316 16544 28917 16572
rect 28316 16532 28322 16544
rect 28905 16541 28917 16544
rect 28951 16541 28963 16575
rect 28905 16535 28963 16541
rect 29089 16575 29147 16581
rect 29089 16541 29101 16575
rect 29135 16541 29147 16575
rect 29472 16572 29500 16612
rect 29825 16609 29837 16643
rect 29871 16609 29883 16643
rect 29825 16603 29883 16609
rect 30837 16643 30895 16649
rect 30837 16609 30849 16643
rect 30883 16609 30895 16643
rect 30837 16603 30895 16609
rect 32950 16600 32956 16652
rect 33008 16600 33014 16652
rect 33962 16600 33968 16652
rect 34020 16640 34026 16652
rect 34793 16643 34851 16649
rect 34793 16640 34805 16643
rect 34020 16612 34805 16640
rect 34020 16600 34026 16612
rect 34793 16609 34805 16612
rect 34839 16609 34851 16643
rect 34793 16603 34851 16609
rect 35250 16600 35256 16652
rect 35308 16600 35314 16652
rect 29917 16575 29975 16581
rect 29917 16572 29929 16575
rect 29472 16544 29929 16572
rect 29089 16535 29147 16541
rect 29917 16541 29929 16544
rect 29963 16541 29975 16575
rect 29917 16535 29975 16541
rect 31104 16575 31162 16581
rect 31104 16541 31116 16575
rect 31150 16572 31162 16575
rect 31662 16572 31668 16584
rect 31150 16544 31668 16572
rect 31150 16541 31162 16544
rect 31104 16535 31162 16541
rect 28350 16464 28356 16516
rect 28408 16504 28414 16516
rect 28997 16507 29055 16513
rect 28997 16504 29009 16507
rect 28408 16476 29009 16504
rect 28408 16464 28414 16476
rect 28997 16473 29009 16476
rect 29043 16473 29055 16507
rect 29104 16504 29132 16535
rect 31662 16532 31668 16544
rect 31720 16532 31726 16584
rect 33502 16532 33508 16584
rect 33560 16572 33566 16584
rect 34146 16572 34152 16584
rect 33560 16544 34152 16572
rect 33560 16532 33566 16544
rect 34146 16532 34152 16544
rect 34204 16572 34210 16584
rect 34885 16575 34943 16581
rect 34885 16572 34897 16575
rect 34204 16544 34897 16572
rect 34204 16532 34210 16544
rect 34885 16541 34897 16544
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 35621 16575 35679 16581
rect 35621 16541 35633 16575
rect 35667 16572 35679 16575
rect 35802 16572 35808 16584
rect 35667 16544 35808 16572
rect 35667 16541 35679 16544
rect 35621 16535 35679 16541
rect 35802 16532 35808 16544
rect 35860 16572 35866 16584
rect 36004 16581 36032 16748
rect 36081 16745 36093 16779
rect 36127 16776 36139 16779
rect 36998 16776 37004 16788
rect 36127 16748 37004 16776
rect 36127 16745 36139 16748
rect 36081 16739 36139 16745
rect 36998 16736 37004 16748
rect 37056 16736 37062 16788
rect 37826 16736 37832 16788
rect 37884 16776 37890 16788
rect 38197 16779 38255 16785
rect 38197 16776 38209 16779
rect 37884 16748 38209 16776
rect 37884 16736 37890 16748
rect 38197 16745 38209 16748
rect 38243 16745 38255 16779
rect 38197 16739 38255 16745
rect 36814 16640 36820 16652
rect 36096 16612 36820 16640
rect 35897 16575 35955 16581
rect 35897 16572 35909 16575
rect 35860 16544 35909 16572
rect 35860 16532 35866 16544
rect 35897 16541 35909 16544
rect 35943 16541 35955 16575
rect 35897 16535 35955 16541
rect 35989 16575 36047 16581
rect 35989 16541 36001 16575
rect 36035 16541 36047 16575
rect 35989 16535 36047 16541
rect 29546 16504 29552 16516
rect 29104 16476 29552 16504
rect 28997 16467 29055 16473
rect 29546 16464 29552 16476
rect 29604 16464 29610 16516
rect 33220 16507 33278 16513
rect 33220 16473 33232 16507
rect 33266 16504 33278 16507
rect 33594 16504 33600 16516
rect 33266 16476 33600 16504
rect 33266 16473 33278 16476
rect 33220 16467 33278 16473
rect 33594 16464 33600 16476
rect 33652 16464 33658 16516
rect 34790 16464 34796 16516
rect 34848 16504 34854 16516
rect 36096 16504 36124 16612
rect 36814 16600 36820 16612
rect 36872 16600 36878 16652
rect 37090 16581 37096 16584
rect 37084 16572 37096 16581
rect 37051 16544 37096 16572
rect 37084 16535 37096 16544
rect 37090 16532 37096 16535
rect 37148 16532 37154 16584
rect 34848 16476 36124 16504
rect 34848 16464 34854 16476
rect 30282 16436 30288 16448
rect 28092 16408 30288 16436
rect 30282 16396 30288 16408
rect 30340 16396 30346 16448
rect 32122 16396 32128 16448
rect 32180 16436 32186 16448
rect 34330 16436 34336 16448
rect 32180 16408 34336 16436
rect 32180 16396 32186 16408
rect 34330 16396 34336 16408
rect 34388 16396 34394 16448
rect 36262 16396 36268 16448
rect 36320 16396 36326 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 15381 16235 15439 16241
rect 15381 16201 15393 16235
rect 15427 16232 15439 16235
rect 19426 16232 19432 16244
rect 15427 16204 19432 16232
rect 15427 16201 15439 16204
rect 15381 16195 15439 16201
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 21358 16192 21364 16244
rect 21416 16192 21422 16244
rect 21542 16192 21548 16244
rect 21600 16232 21606 16244
rect 24026 16232 24032 16244
rect 21600 16204 24032 16232
rect 21600 16192 21606 16204
rect 24026 16192 24032 16204
rect 24084 16232 24090 16244
rect 24084 16204 24624 16232
rect 24084 16192 24090 16204
rect 15933 16167 15991 16173
rect 15933 16133 15945 16167
rect 15979 16164 15991 16167
rect 17034 16164 17040 16176
rect 15979 16136 17040 16164
rect 15979 16133 15991 16136
rect 15933 16127 15991 16133
rect 17034 16124 17040 16136
rect 17092 16124 17098 16176
rect 21818 16124 21824 16176
rect 21876 16164 21882 16176
rect 23661 16167 23719 16173
rect 21876 16136 22146 16164
rect 21876 16124 21882 16136
rect 15286 16056 15292 16108
rect 15344 16056 15350 16108
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16096 15531 16099
rect 16022 16096 16028 16108
rect 15519 16068 16028 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16065 16175 16099
rect 16117 16059 16175 16065
rect 15930 15988 15936 16040
rect 15988 16028 15994 16040
rect 16132 16028 16160 16059
rect 16850 16056 16856 16108
rect 16908 16056 16914 16108
rect 16942 16056 16948 16108
rect 17000 16056 17006 16108
rect 18506 16056 18512 16108
rect 18564 16056 18570 16108
rect 18598 16056 18604 16108
rect 18656 16056 18662 16108
rect 20346 16056 20352 16108
rect 20404 16056 20410 16108
rect 20806 16056 20812 16108
rect 20864 16056 20870 16108
rect 21266 16056 21272 16108
rect 21324 16056 21330 16108
rect 21726 16056 21732 16108
rect 21784 16096 21790 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21784 16068 22017 16096
rect 21784 16056 21790 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22118 16096 22146 16136
rect 23661 16133 23673 16167
rect 23707 16164 23719 16167
rect 23750 16164 23756 16176
rect 23707 16136 23756 16164
rect 23707 16133 23719 16136
rect 23661 16127 23719 16133
rect 23750 16124 23756 16136
rect 23808 16124 23814 16176
rect 23934 16164 23940 16176
rect 23860 16136 23940 16164
rect 23860 16096 23888 16136
rect 23934 16124 23940 16136
rect 23992 16164 23998 16176
rect 24489 16167 24547 16173
rect 24489 16164 24501 16167
rect 23992 16136 24501 16164
rect 23992 16124 23998 16136
rect 24489 16133 24501 16136
rect 24535 16133 24547 16167
rect 24489 16127 24547 16133
rect 22118 16068 23888 16096
rect 22005 16059 22063 16065
rect 24302 16056 24308 16108
rect 24360 16056 24366 16108
rect 24596 16105 24624 16204
rect 25590 16192 25596 16244
rect 25648 16232 25654 16244
rect 25869 16235 25927 16241
rect 25869 16232 25881 16235
rect 25648 16204 25881 16232
rect 25648 16192 25654 16204
rect 25869 16201 25881 16204
rect 25915 16232 25927 16235
rect 27706 16232 27712 16244
rect 25915 16204 27712 16232
rect 25915 16201 25927 16204
rect 25869 16195 25927 16201
rect 27706 16192 27712 16204
rect 27764 16192 27770 16244
rect 30742 16192 30748 16244
rect 30800 16232 30806 16244
rect 30837 16235 30895 16241
rect 30837 16232 30849 16235
rect 30800 16204 30849 16232
rect 30800 16192 30806 16204
rect 30837 16201 30849 16204
rect 30883 16201 30895 16235
rect 30837 16195 30895 16201
rect 31754 16192 31760 16244
rect 31812 16232 31818 16244
rect 31812 16204 32996 16232
rect 31812 16192 31818 16204
rect 26418 16124 26424 16176
rect 26476 16164 26482 16176
rect 26476 16136 30880 16164
rect 26476 16124 26482 16136
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16065 24639 16099
rect 24581 16059 24639 16065
rect 25777 16099 25835 16105
rect 25777 16065 25789 16099
rect 25823 16096 25835 16099
rect 26050 16096 26056 16108
rect 25823 16068 26056 16096
rect 25823 16065 25835 16068
rect 25777 16059 25835 16065
rect 26050 16056 26056 16068
rect 26108 16056 26114 16108
rect 26510 16056 26516 16108
rect 26568 16096 26574 16108
rect 27617 16099 27675 16105
rect 26568 16068 27568 16096
rect 26568 16056 26574 16068
rect 15988 16000 16160 16028
rect 16301 16031 16359 16037
rect 15988 15988 15994 16000
rect 16301 15997 16313 16031
rect 16347 16028 16359 16031
rect 16574 16028 16580 16040
rect 16347 16000 16580 16028
rect 16347 15997 16359 16000
rect 16301 15991 16359 15997
rect 16574 15988 16580 16000
rect 16632 16028 16638 16040
rect 17586 16028 17592 16040
rect 16632 16000 17592 16028
rect 16632 15988 16638 16000
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 19150 15988 19156 16040
rect 19208 16028 19214 16040
rect 19245 16031 19303 16037
rect 19245 16028 19257 16031
rect 19208 16000 19257 16028
rect 19208 15988 19214 16000
rect 19245 15997 19257 16000
rect 19291 16028 19303 16031
rect 22281 16031 22339 16037
rect 22281 16028 22293 16031
rect 19291 16000 22293 16028
rect 19291 15997 19303 16000
rect 19245 15991 19303 15997
rect 22281 15997 22293 16000
rect 22327 15997 22339 16031
rect 22281 15991 22339 15997
rect 23014 15988 23020 16040
rect 23072 16028 23078 16040
rect 23072 16000 24256 16028
rect 23072 15988 23078 16000
rect 15010 15920 15016 15972
rect 15068 15960 15074 15972
rect 18414 15960 18420 15972
rect 15068 15932 18420 15960
rect 15068 15920 15074 15932
rect 18414 15920 18420 15932
rect 18472 15920 18478 15972
rect 23106 15920 23112 15972
rect 23164 15960 23170 15972
rect 24121 15963 24179 15969
rect 24121 15960 24133 15963
rect 23164 15932 24133 15960
rect 23164 15920 23170 15932
rect 24121 15929 24133 15932
rect 24167 15929 24179 15963
rect 24228 15960 24256 16000
rect 25958 15988 25964 16040
rect 26016 15988 26022 16040
rect 27540 16028 27568 16068
rect 27617 16065 27629 16099
rect 27663 16096 27675 16099
rect 28442 16096 28448 16108
rect 27663 16068 28448 16096
rect 27663 16065 27675 16068
rect 27617 16059 27675 16065
rect 28442 16056 28448 16068
rect 28500 16056 28506 16108
rect 28534 16056 28540 16108
rect 28592 16056 28598 16108
rect 28810 16105 28816 16108
rect 28804 16059 28816 16105
rect 28810 16056 28816 16059
rect 28868 16056 28874 16108
rect 30742 16056 30748 16108
rect 30800 16056 30806 16108
rect 30852 16096 30880 16136
rect 31110 16124 31116 16176
rect 31168 16164 31174 16176
rect 31168 16136 32352 16164
rect 31168 16124 31174 16136
rect 32324 16105 32352 16136
rect 32968 16108 32996 16204
rect 33594 16192 33600 16244
rect 33652 16192 33658 16244
rect 33686 16192 33692 16244
rect 33744 16232 33750 16244
rect 33965 16235 34023 16241
rect 33965 16232 33977 16235
rect 33744 16204 33977 16232
rect 33744 16192 33750 16204
rect 33965 16201 33977 16204
rect 34011 16201 34023 16235
rect 33965 16195 34023 16201
rect 34514 16192 34520 16244
rect 34572 16232 34578 16244
rect 34572 16204 36308 16232
rect 34572 16192 34578 16204
rect 35250 16173 35256 16176
rect 35244 16164 35256 16173
rect 35211 16136 35256 16164
rect 35244 16127 35256 16136
rect 35250 16124 35256 16127
rect 35308 16124 35314 16176
rect 36280 16164 36308 16204
rect 36354 16192 36360 16244
rect 36412 16192 36418 16244
rect 37918 16164 37924 16176
rect 36280 16136 37924 16164
rect 37918 16124 37924 16136
rect 37976 16124 37982 16176
rect 31573 16099 31631 16105
rect 31573 16096 31585 16099
rect 30852 16068 31585 16096
rect 31573 16065 31585 16068
rect 31619 16065 31631 16099
rect 31573 16059 31631 16065
rect 31757 16099 31815 16105
rect 31757 16065 31769 16099
rect 31803 16065 31815 16099
rect 31757 16059 31815 16065
rect 32309 16099 32367 16105
rect 32309 16065 32321 16099
rect 32355 16065 32367 16099
rect 32309 16059 32367 16065
rect 27801 16031 27859 16037
rect 27801 16028 27813 16031
rect 27540 16000 27813 16028
rect 27801 15997 27813 16000
rect 27847 15997 27859 16031
rect 27801 15991 27859 15997
rect 29546 15988 29552 16040
rect 29604 16028 29610 16040
rect 31021 16031 31079 16037
rect 29604 16000 30972 16028
rect 29604 15988 29610 16000
rect 30944 15960 30972 16000
rect 31021 15997 31033 16031
rect 31067 16028 31079 16031
rect 31110 16028 31116 16040
rect 31067 16000 31116 16028
rect 31067 15997 31079 16000
rect 31021 15991 31079 15997
rect 31110 15988 31116 16000
rect 31168 15988 31174 16040
rect 31772 15960 31800 16059
rect 32398 16056 32404 16108
rect 32456 16096 32462 16108
rect 32674 16096 32680 16108
rect 32456 16068 32680 16096
rect 32456 16056 32462 16068
rect 32674 16056 32680 16068
rect 32732 16056 32738 16108
rect 32950 16056 32956 16108
rect 33008 16056 33014 16108
rect 34057 16099 34115 16105
rect 34057 16065 34069 16099
rect 34103 16096 34115 16099
rect 34698 16096 34704 16108
rect 34103 16068 34704 16096
rect 34103 16065 34115 16068
rect 34057 16059 34115 16065
rect 34698 16056 34704 16068
rect 34756 16096 34762 16108
rect 36354 16096 36360 16108
rect 34756 16068 36360 16096
rect 34756 16056 34762 16068
rect 36354 16056 36360 16068
rect 36412 16056 36418 16108
rect 37826 16056 37832 16108
rect 37884 16056 37890 16108
rect 32582 15988 32588 16040
rect 32640 15988 32646 16040
rect 34241 16031 34299 16037
rect 34241 15997 34253 16031
rect 34287 15997 34299 16031
rect 34241 15991 34299 15997
rect 24228 15932 27476 15960
rect 24121 15923 24179 15929
rect 20070 15852 20076 15904
rect 20128 15892 20134 15904
rect 20165 15895 20223 15901
rect 20165 15892 20177 15895
rect 20128 15864 20177 15892
rect 20128 15852 20134 15864
rect 20165 15861 20177 15864
rect 20211 15861 20223 15895
rect 20165 15855 20223 15861
rect 25406 15852 25412 15904
rect 25464 15852 25470 15904
rect 27249 15895 27307 15901
rect 27249 15861 27261 15895
rect 27295 15892 27307 15895
rect 27338 15892 27344 15904
rect 27295 15864 27344 15892
rect 27295 15861 27307 15864
rect 27249 15855 27307 15861
rect 27338 15852 27344 15864
rect 27396 15852 27402 15904
rect 27448 15892 27476 15932
rect 29472 15932 30512 15960
rect 30944 15932 31800 15960
rect 29472 15892 29500 15932
rect 27448 15864 29500 15892
rect 29914 15852 29920 15904
rect 29972 15852 29978 15904
rect 30374 15852 30380 15904
rect 30432 15852 30438 15904
rect 30484 15892 30512 15932
rect 31665 15895 31723 15901
rect 31665 15892 31677 15895
rect 30484 15864 31677 15892
rect 31665 15861 31677 15864
rect 31711 15861 31723 15895
rect 34256 15892 34284 15991
rect 34790 15988 34796 16040
rect 34848 16028 34854 16040
rect 34977 16031 35035 16037
rect 34977 16028 34989 16031
rect 34848 16000 34989 16028
rect 34848 15988 34854 16000
rect 34977 15997 34989 16000
rect 35023 15997 35035 16031
rect 38013 16031 38071 16037
rect 38013 16028 38025 16031
rect 34977 15991 35035 15997
rect 37384 16000 38025 16028
rect 37384 15892 37412 16000
rect 38013 15997 38025 16000
rect 38059 16028 38071 16031
rect 38102 16028 38108 16040
rect 38059 16000 38108 16028
rect 38059 15997 38071 16000
rect 38013 15991 38071 15997
rect 38102 15988 38108 16000
rect 38160 15988 38166 16040
rect 34256 15864 37412 15892
rect 31665 15855 31723 15861
rect 37458 15852 37464 15904
rect 37516 15852 37522 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 16758 15648 16764 15700
rect 16816 15688 16822 15700
rect 17681 15691 17739 15697
rect 17681 15688 17693 15691
rect 16816 15660 17693 15688
rect 16816 15648 16822 15660
rect 17681 15657 17693 15660
rect 17727 15657 17739 15691
rect 17681 15651 17739 15657
rect 18417 15691 18475 15697
rect 18417 15657 18429 15691
rect 18463 15688 18475 15691
rect 19334 15688 19340 15700
rect 18463 15660 19340 15688
rect 18463 15657 18475 15660
rect 18417 15651 18475 15657
rect 17696 15620 17724 15651
rect 19334 15648 19340 15660
rect 19392 15688 19398 15700
rect 19978 15688 19984 15700
rect 19392 15660 19984 15688
rect 19392 15648 19398 15660
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 22554 15688 22560 15700
rect 20088 15660 22560 15688
rect 20088 15620 20116 15660
rect 22554 15648 22560 15660
rect 22612 15688 22618 15700
rect 27246 15688 27252 15700
rect 22612 15660 27252 15688
rect 22612 15648 22618 15660
rect 27246 15648 27252 15660
rect 27304 15648 27310 15700
rect 28442 15648 28448 15700
rect 28500 15648 28506 15700
rect 28994 15648 29000 15700
rect 29052 15648 29058 15700
rect 33134 15648 33140 15700
rect 33192 15688 33198 15700
rect 37369 15691 37427 15697
rect 37369 15688 37381 15691
rect 33192 15660 37381 15688
rect 33192 15648 33198 15660
rect 37369 15657 37381 15660
rect 37415 15688 37427 15691
rect 37826 15688 37832 15700
rect 37415 15660 37832 15688
rect 37415 15657 37427 15660
rect 37369 15651 37427 15657
rect 37826 15648 37832 15660
rect 37884 15648 37890 15700
rect 17696 15592 20116 15620
rect 20162 15580 20168 15632
rect 20220 15580 20226 15632
rect 20346 15580 20352 15632
rect 20404 15620 20410 15632
rect 21545 15623 21603 15629
rect 21545 15620 21557 15623
rect 20404 15592 21557 15620
rect 20404 15580 20410 15592
rect 21545 15589 21557 15592
rect 21591 15589 21603 15623
rect 21545 15583 21603 15589
rect 31938 15580 31944 15632
rect 31996 15580 32002 15632
rect 16301 15555 16359 15561
rect 16301 15521 16313 15555
rect 16347 15552 16359 15555
rect 18690 15552 18696 15564
rect 16347 15524 18696 15552
rect 16347 15521 16359 15524
rect 16301 15515 16359 15521
rect 18690 15512 18696 15524
rect 18748 15512 18754 15564
rect 18785 15555 18843 15561
rect 18785 15521 18797 15555
rect 18831 15552 18843 15555
rect 18831 15524 20024 15552
rect 18831 15521 18843 15524
rect 18785 15515 18843 15521
rect 16577 15487 16635 15493
rect 16577 15453 16589 15487
rect 16623 15484 16635 15487
rect 18506 15484 18512 15496
rect 16623 15456 18512 15484
rect 16623 15453 16635 15456
rect 16577 15447 16635 15453
rect 18506 15444 18512 15456
rect 18564 15444 18570 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15453 18659 15487
rect 18601 15447 18659 15453
rect 18616 15416 18644 15447
rect 18874 15444 18880 15496
rect 18932 15484 18938 15496
rect 19426 15484 19432 15496
rect 18932 15456 19432 15484
rect 18932 15444 18938 15456
rect 19426 15444 19432 15456
rect 19484 15484 19490 15496
rect 19996 15493 20024 15524
rect 20530 15512 20536 15564
rect 20588 15552 20594 15564
rect 21729 15555 21787 15561
rect 20588 15524 21588 15552
rect 20588 15512 20594 15524
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 19484 15456 19533 15484
rect 19484 15444 19490 15456
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19981 15487 20039 15493
rect 19981 15453 19993 15487
rect 20027 15484 20039 15487
rect 20070 15484 20076 15496
rect 20027 15456 20076 15484
rect 20027 15453 20039 15456
rect 19981 15447 20039 15453
rect 20070 15444 20076 15456
rect 20128 15444 20134 15496
rect 20254 15444 20260 15496
rect 20312 15444 20318 15496
rect 20625 15487 20683 15493
rect 20625 15453 20637 15487
rect 20671 15484 20683 15487
rect 20806 15484 20812 15496
rect 20671 15456 20812 15484
rect 20671 15453 20683 15456
rect 20625 15447 20683 15453
rect 20640 15416 20668 15447
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 21560 15493 21588 15524
rect 21729 15521 21741 15555
rect 21775 15552 21787 15555
rect 22002 15552 22008 15564
rect 21775 15524 22008 15552
rect 21775 15521 21787 15524
rect 21729 15515 21787 15521
rect 22002 15512 22008 15524
rect 22060 15512 22066 15564
rect 23569 15555 23627 15561
rect 23569 15521 23581 15555
rect 23615 15552 23627 15555
rect 26510 15552 26516 15564
rect 23615 15524 26516 15552
rect 23615 15521 23627 15524
rect 23569 15515 23627 15521
rect 26510 15512 26516 15524
rect 26568 15512 26574 15564
rect 26602 15512 26608 15564
rect 26660 15552 26666 15564
rect 27065 15555 27123 15561
rect 27065 15552 27077 15555
rect 26660 15524 27077 15552
rect 26660 15512 26666 15524
rect 27065 15521 27077 15524
rect 27111 15521 27123 15555
rect 27065 15515 27123 15521
rect 28534 15512 28540 15564
rect 28592 15552 28598 15564
rect 28592 15524 29776 15552
rect 28592 15512 28598 15524
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 21634 15444 21640 15496
rect 21692 15484 21698 15496
rect 21913 15487 21971 15493
rect 21913 15484 21925 15487
rect 21692 15456 21925 15484
rect 21692 15444 21698 15456
rect 21913 15453 21925 15456
rect 21959 15453 21971 15487
rect 21913 15447 21971 15453
rect 23382 15444 23388 15496
rect 23440 15484 23446 15496
rect 24946 15484 24952 15496
rect 23440 15456 24952 15484
rect 23440 15444 23446 15456
rect 24946 15444 24952 15456
rect 25004 15444 25010 15496
rect 27338 15493 27344 15496
rect 27332 15484 27344 15493
rect 27299 15456 27344 15484
rect 27332 15447 27344 15456
rect 27338 15444 27344 15447
rect 27396 15444 27402 15496
rect 28905 15487 28963 15493
rect 28905 15484 28917 15487
rect 27448 15456 28917 15484
rect 27448 15428 27476 15456
rect 28905 15453 28917 15456
rect 28951 15453 28963 15487
rect 28905 15447 28963 15453
rect 29089 15487 29147 15493
rect 29089 15453 29101 15487
rect 29135 15484 29147 15487
rect 29546 15484 29552 15496
rect 29135 15456 29552 15484
rect 29135 15453 29147 15456
rect 29089 15447 29147 15453
rect 29546 15444 29552 15456
rect 29604 15444 29610 15496
rect 29748 15493 29776 15524
rect 31478 15512 31484 15564
rect 31536 15552 31542 15564
rect 31573 15555 31631 15561
rect 31573 15552 31585 15555
rect 31536 15524 31585 15552
rect 31536 15512 31542 15524
rect 31573 15521 31585 15524
rect 31619 15521 31631 15555
rect 31573 15515 31631 15521
rect 38105 15555 38163 15561
rect 38105 15521 38117 15555
rect 38151 15552 38163 15555
rect 38930 15552 38936 15564
rect 38151 15524 38936 15552
rect 38151 15521 38163 15524
rect 38105 15515 38163 15521
rect 38930 15512 38936 15524
rect 38988 15512 38994 15564
rect 29733 15487 29791 15493
rect 29733 15453 29745 15487
rect 29779 15484 29791 15487
rect 29822 15484 29828 15496
rect 29779 15456 29828 15484
rect 29779 15453 29791 15456
rect 29733 15447 29791 15453
rect 29822 15444 29828 15456
rect 29880 15484 29886 15496
rect 31386 15484 31392 15496
rect 29880 15456 31392 15484
rect 29880 15444 29886 15456
rect 31386 15444 31392 15456
rect 31444 15484 31450 15496
rect 32493 15487 32551 15493
rect 32493 15484 32505 15487
rect 31444 15456 32505 15484
rect 31444 15444 31450 15456
rect 32493 15453 32505 15456
rect 32539 15484 32551 15487
rect 34698 15484 34704 15496
rect 32539 15456 34704 15484
rect 32539 15453 32551 15456
rect 32493 15447 32551 15453
rect 34698 15444 34704 15456
rect 34756 15484 34762 15496
rect 35989 15487 36047 15493
rect 35989 15484 36001 15487
rect 34756 15456 36001 15484
rect 34756 15444 34762 15456
rect 35989 15453 36001 15456
rect 36035 15453 36047 15487
rect 35989 15447 36047 15453
rect 36256 15487 36314 15493
rect 36256 15453 36268 15487
rect 36302 15484 36314 15487
rect 37458 15484 37464 15496
rect 36302 15456 37464 15484
rect 36302 15453 36314 15456
rect 36256 15447 36314 15453
rect 37458 15444 37464 15456
rect 37516 15444 37522 15496
rect 37829 15487 37887 15493
rect 37829 15453 37841 15487
rect 37875 15484 37887 15487
rect 38010 15484 38016 15496
rect 37875 15456 38016 15484
rect 37875 15453 37887 15456
rect 37829 15447 37887 15453
rect 38010 15444 38016 15456
rect 38068 15444 38074 15496
rect 18616 15388 20668 15416
rect 23293 15419 23351 15425
rect 23293 15385 23305 15419
rect 23339 15416 23351 15419
rect 23750 15416 23756 15428
rect 23339 15388 23756 15416
rect 23339 15385 23351 15388
rect 23293 15379 23351 15385
rect 23750 15376 23756 15388
rect 23808 15376 23814 15428
rect 24578 15376 24584 15428
rect 24636 15416 24642 15428
rect 24636 15388 26096 15416
rect 24636 15376 24642 15388
rect 22922 15308 22928 15360
rect 22980 15308 22986 15360
rect 25498 15308 25504 15360
rect 25556 15348 25562 15360
rect 25869 15351 25927 15357
rect 25869 15348 25881 15351
rect 25556 15320 25881 15348
rect 25556 15308 25562 15320
rect 25869 15317 25881 15320
rect 25915 15317 25927 15351
rect 26068 15348 26096 15388
rect 27430 15376 27436 15428
rect 27488 15376 27494 15428
rect 30000 15419 30058 15425
rect 30000 15385 30012 15419
rect 30046 15416 30058 15419
rect 30374 15416 30380 15428
rect 30046 15388 30380 15416
rect 30046 15385 30058 15388
rect 30000 15379 30058 15385
rect 30374 15376 30380 15388
rect 30432 15376 30438 15428
rect 32214 15376 32220 15428
rect 32272 15416 32278 15428
rect 32738 15419 32796 15425
rect 32738 15416 32750 15419
rect 32272 15388 32750 15416
rect 32272 15376 32278 15388
rect 32738 15385 32750 15388
rect 32784 15385 32796 15419
rect 32738 15379 32796 15385
rect 35161 15419 35219 15425
rect 35161 15385 35173 15419
rect 35207 15385 35219 15419
rect 35161 15379 35219 15385
rect 35345 15419 35403 15425
rect 35345 15385 35357 15419
rect 35391 15416 35403 15419
rect 35710 15416 35716 15428
rect 35391 15388 35716 15416
rect 35391 15385 35403 15388
rect 35345 15379 35403 15385
rect 29546 15348 29552 15360
rect 26068 15320 29552 15348
rect 25869 15311 25927 15317
rect 29546 15308 29552 15320
rect 29604 15308 29610 15360
rect 30742 15308 30748 15360
rect 30800 15348 30806 15360
rect 31113 15351 31171 15357
rect 31113 15348 31125 15351
rect 30800 15320 31125 15348
rect 30800 15308 30806 15320
rect 31113 15317 31125 15320
rect 31159 15317 31171 15351
rect 31113 15311 31171 15317
rect 32033 15351 32091 15357
rect 32033 15317 32045 15351
rect 32079 15348 32091 15351
rect 33594 15348 33600 15360
rect 32079 15320 33600 15348
rect 32079 15317 32091 15320
rect 32033 15311 32091 15317
rect 33594 15308 33600 15320
rect 33652 15308 33658 15360
rect 33870 15308 33876 15360
rect 33928 15308 33934 15360
rect 35176 15348 35204 15379
rect 35710 15376 35716 15388
rect 35768 15376 35774 15428
rect 35434 15348 35440 15360
rect 35176 15320 35440 15348
rect 35434 15308 35440 15320
rect 35492 15308 35498 15360
rect 35529 15351 35587 15357
rect 35529 15317 35541 15351
rect 35575 15348 35587 15351
rect 36262 15348 36268 15360
rect 35575 15320 36268 15348
rect 35575 15317 35587 15320
rect 35529 15311 35587 15317
rect 36262 15308 36268 15320
rect 36320 15308 36326 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 21177 15147 21235 15153
rect 21177 15113 21189 15147
rect 21223 15144 21235 15147
rect 22462 15144 22468 15156
rect 21223 15116 22468 15144
rect 21223 15113 21235 15116
rect 21177 15107 21235 15113
rect 22462 15104 22468 15116
rect 22520 15144 22526 15156
rect 23382 15144 23388 15156
rect 22520 15116 23388 15144
rect 22520 15104 22526 15116
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 23658 15104 23664 15156
rect 23716 15144 23722 15156
rect 27617 15147 27675 15153
rect 23716 15116 27568 15144
rect 23716 15104 23722 15116
rect 17865 15079 17923 15085
rect 17865 15045 17877 15079
rect 17911 15076 17923 15079
rect 18598 15076 18604 15088
rect 17911 15048 18604 15076
rect 17911 15045 17923 15048
rect 17865 15039 17923 15045
rect 18598 15036 18604 15048
rect 18656 15036 18662 15088
rect 17402 14968 17408 15020
rect 17460 15008 17466 15020
rect 17681 15011 17739 15017
rect 17681 15008 17693 15011
rect 17460 14980 17693 15008
rect 17460 14968 17466 14980
rect 17681 14977 17693 14980
rect 17727 14977 17739 15011
rect 17681 14971 17739 14977
rect 18138 14968 18144 15020
rect 18196 14968 18202 15020
rect 19150 14968 19156 15020
rect 19208 14968 19214 15020
rect 19797 15011 19855 15017
rect 19797 14977 19809 15011
rect 19843 15008 19855 15011
rect 20438 15008 20444 15020
rect 19843 14980 20444 15008
rect 19843 14977 19855 14980
rect 19797 14971 19855 14977
rect 20438 14968 20444 14980
rect 20496 14968 20502 15020
rect 21082 14968 21088 15020
rect 21140 14968 21146 15020
rect 22370 14968 22376 15020
rect 22428 14968 22434 15020
rect 22640 15011 22698 15017
rect 22640 14977 22652 15011
rect 22686 15008 22698 15011
rect 22922 15008 22928 15020
rect 22686 14980 22928 15008
rect 22686 14977 22698 14980
rect 22640 14971 22698 14977
rect 22922 14968 22928 14980
rect 22980 14968 22986 15020
rect 25032 15011 25090 15017
rect 25032 14977 25044 15011
rect 25078 15008 25090 15011
rect 25406 15008 25412 15020
rect 25078 14980 25412 15008
rect 25078 14977 25090 14980
rect 25032 14971 25090 14977
rect 25406 14968 25412 14980
rect 25464 14968 25470 15020
rect 27338 14968 27344 15020
rect 27396 14968 27402 15020
rect 27430 14968 27436 15020
rect 27488 14968 27494 15020
rect 27540 15008 27568 15116
rect 27617 15113 27629 15147
rect 27663 15144 27675 15147
rect 27663 15116 28764 15144
rect 27663 15113 27675 15116
rect 27617 15107 27675 15113
rect 28736 15076 28764 15116
rect 28810 15104 28816 15156
rect 28868 15144 28874 15156
rect 29641 15147 29699 15153
rect 29641 15144 29653 15147
rect 28868 15116 29653 15144
rect 28868 15104 28874 15116
rect 29641 15113 29653 15116
rect 29687 15113 29699 15147
rect 29641 15107 29699 15113
rect 29914 15104 29920 15156
rect 29972 15144 29978 15156
rect 30009 15147 30067 15153
rect 30009 15144 30021 15147
rect 29972 15116 30021 15144
rect 29972 15104 29978 15116
rect 30009 15113 30021 15116
rect 30055 15113 30067 15147
rect 30009 15107 30067 15113
rect 30098 15104 30104 15156
rect 30156 15104 30162 15156
rect 31021 15147 31079 15153
rect 31021 15113 31033 15147
rect 31067 15144 31079 15147
rect 32214 15144 32220 15156
rect 31067 15116 32220 15144
rect 31067 15113 31079 15116
rect 31021 15107 31079 15113
rect 32214 15104 32220 15116
rect 32272 15104 32278 15156
rect 32585 15147 32643 15153
rect 32585 15113 32597 15147
rect 32631 15144 32643 15147
rect 33778 15144 33784 15156
rect 32631 15116 33784 15144
rect 32631 15113 32643 15116
rect 32585 15107 32643 15113
rect 33778 15104 33784 15116
rect 33836 15144 33842 15156
rect 33836 15116 34192 15144
rect 33836 15104 33842 15116
rect 29730 15076 29736 15088
rect 28736 15048 29736 15076
rect 29730 15036 29736 15048
rect 29788 15036 29794 15088
rect 27982 15008 27988 15020
rect 27540 14980 27988 15008
rect 27982 14968 27988 14980
rect 28040 15008 28046 15020
rect 28169 15011 28227 15017
rect 28169 15008 28181 15011
rect 28040 14980 28181 15008
rect 28040 14968 28046 14980
rect 28169 14977 28181 14980
rect 28215 14977 28227 15011
rect 28169 14971 28227 14977
rect 28442 14968 28448 15020
rect 28500 15008 28506 15020
rect 28629 15011 28687 15017
rect 28629 15008 28641 15011
rect 28500 14980 28641 15008
rect 28500 14968 28506 14980
rect 28629 14977 28641 14980
rect 28675 14977 28687 15011
rect 30116 15008 30144 15104
rect 31389 15079 31447 15085
rect 31389 15045 31401 15079
rect 31435 15076 31447 15079
rect 33870 15076 33876 15088
rect 31435 15048 33876 15076
rect 31435 15045 31447 15048
rect 31389 15039 31447 15045
rect 30116 14980 30420 15008
rect 28629 14971 28687 14977
rect 19242 14900 19248 14952
rect 19300 14900 19306 14952
rect 19518 14900 19524 14952
rect 19576 14940 19582 14952
rect 20162 14940 20168 14952
rect 19576 14912 20168 14940
rect 19576 14900 19582 14912
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 21361 14943 21419 14949
rect 21361 14909 21373 14943
rect 21407 14940 21419 14943
rect 22278 14940 22284 14952
rect 21407 14912 22284 14940
rect 21407 14909 21419 14912
rect 21361 14903 21419 14909
rect 22278 14900 22284 14912
rect 22336 14900 22342 14952
rect 23382 14900 23388 14952
rect 23440 14940 23446 14952
rect 24765 14943 24823 14949
rect 24765 14940 24777 14943
rect 23440 14912 24777 14940
rect 23440 14900 23446 14912
rect 24765 14909 24777 14912
rect 24811 14909 24823 14943
rect 27448 14940 27476 14968
rect 27448 14912 28304 14940
rect 24765 14903 24823 14909
rect 18414 14832 18420 14884
rect 18472 14872 18478 14884
rect 18782 14872 18788 14884
rect 18472 14844 18788 14872
rect 18472 14832 18478 14844
rect 18782 14832 18788 14844
rect 18840 14872 18846 14884
rect 19337 14875 19395 14881
rect 19337 14872 19349 14875
rect 18840 14844 19349 14872
rect 18840 14832 18846 14844
rect 19337 14841 19349 14844
rect 19383 14841 19395 14875
rect 28276 14872 28304 14912
rect 28350 14900 28356 14952
rect 28408 14900 28414 14952
rect 28537 14943 28595 14949
rect 28537 14909 28549 14943
rect 28583 14909 28595 14943
rect 28537 14903 28595 14909
rect 28552 14872 28580 14903
rect 30190 14900 30196 14952
rect 30248 14900 30254 14952
rect 30392 14940 30420 14980
rect 30466 14968 30472 15020
rect 30524 15008 30530 15020
rect 32309 15011 32367 15017
rect 32309 15008 32321 15011
rect 30524 14980 32321 15008
rect 30524 14968 30530 14980
rect 32309 14977 32321 14980
rect 32355 14977 32367 15011
rect 32309 14971 32367 14977
rect 32490 14968 32496 15020
rect 32548 15008 32554 15020
rect 33137 15011 33195 15017
rect 33137 15008 33149 15011
rect 32548 14980 33149 15008
rect 32548 14968 32554 14980
rect 33137 14977 33149 14980
rect 33183 14977 33195 15011
rect 33502 15008 33508 15020
rect 33137 14971 33195 14977
rect 33244 14980 33508 15008
rect 31478 14940 31484 14952
rect 30392 14912 31484 14940
rect 31478 14900 31484 14912
rect 31536 14900 31542 14952
rect 31662 14900 31668 14952
rect 31720 14900 31726 14952
rect 33244 14940 33272 14980
rect 33502 14968 33508 14980
rect 33560 14968 33566 15020
rect 33612 15017 33640 15048
rect 33870 15036 33876 15048
rect 33928 15036 33934 15088
rect 33597 15011 33655 15017
rect 33597 14977 33609 15011
rect 33643 14977 33655 15011
rect 34164 15008 34192 15116
rect 34606 15104 34612 15156
rect 34664 15144 34670 15156
rect 34701 15147 34759 15153
rect 34701 15144 34713 15147
rect 34664 15116 34713 15144
rect 34664 15104 34670 15116
rect 34701 15113 34713 15116
rect 34747 15113 34759 15147
rect 35986 15144 35992 15156
rect 34701 15107 34759 15113
rect 35452 15116 35992 15144
rect 35452 15076 35480 15116
rect 35986 15104 35992 15116
rect 36044 15144 36050 15156
rect 36449 15147 36507 15153
rect 36449 15144 36461 15147
rect 36044 15116 36461 15144
rect 36044 15104 36050 15116
rect 36449 15113 36461 15116
rect 36495 15113 36507 15147
rect 36449 15107 36507 15113
rect 34624 15048 35296 15076
rect 34624 15017 34652 15048
rect 34609 15011 34667 15017
rect 34609 15008 34621 15011
rect 34164 14980 34621 15008
rect 33597 14971 33655 14977
rect 34609 14977 34621 14980
rect 34655 14977 34667 15011
rect 34609 14971 34667 14977
rect 34793 15011 34851 15017
rect 34793 14977 34805 15011
rect 34839 14977 34851 15011
rect 34793 14971 34851 14977
rect 32324 14912 33272 14940
rect 32324 14872 32352 14912
rect 33318 14900 33324 14952
rect 33376 14900 33382 14952
rect 28276 14844 32352 14872
rect 19337 14835 19395 14841
rect 20717 14807 20775 14813
rect 20717 14773 20729 14807
rect 20763 14804 20775 14807
rect 22094 14804 22100 14816
rect 20763 14776 22100 14804
rect 20763 14773 20775 14776
rect 20717 14767 20775 14773
rect 22094 14764 22100 14776
rect 22152 14764 22158 14816
rect 23750 14764 23756 14816
rect 23808 14804 23814 14816
rect 24762 14804 24768 14816
rect 23808 14776 24768 14804
rect 23808 14764 23814 14776
rect 24762 14764 24768 14776
rect 24820 14764 24826 14816
rect 26050 14764 26056 14816
rect 26108 14804 26114 14816
rect 26145 14807 26203 14813
rect 26145 14804 26157 14807
rect 26108 14776 26157 14804
rect 26108 14764 26114 14776
rect 26145 14773 26157 14776
rect 26191 14773 26203 14807
rect 26145 14767 26203 14773
rect 29454 14764 29460 14816
rect 29512 14804 29518 14816
rect 31570 14804 31576 14816
rect 29512 14776 31576 14804
rect 29512 14764 29518 14776
rect 31570 14764 31576 14776
rect 31628 14804 31634 14816
rect 34808 14804 34836 14971
rect 35268 14940 35296 15048
rect 35360 15048 35480 15076
rect 35360 15017 35388 15048
rect 35894 15036 35900 15088
rect 35952 15076 35958 15088
rect 36081 15079 36139 15085
rect 36081 15076 36093 15079
rect 35952 15048 36093 15076
rect 35952 15036 35958 15048
rect 36081 15045 36093 15048
rect 36127 15045 36139 15079
rect 36081 15039 36139 15045
rect 36262 15036 36268 15088
rect 36320 15076 36326 15088
rect 36906 15076 36912 15088
rect 36320 15048 36912 15076
rect 36320 15036 36326 15048
rect 36906 15036 36912 15048
rect 36964 15036 36970 15088
rect 38105 15079 38163 15085
rect 38105 15045 38117 15079
rect 38151 15076 38163 15079
rect 39022 15076 39028 15088
rect 38151 15048 39028 15076
rect 38151 15045 38163 15048
rect 38105 15039 38163 15045
rect 39022 15036 39028 15048
rect 39080 15036 39086 15088
rect 35345 15011 35403 15017
rect 35345 14977 35357 15011
rect 35391 14977 35403 15011
rect 35345 14971 35403 14977
rect 35437 15011 35495 15017
rect 35437 14977 35449 15011
rect 35483 15008 35495 15011
rect 36170 15008 36176 15020
rect 35483 14980 36176 15008
rect 35483 14977 35495 14980
rect 35437 14971 35495 14977
rect 36170 14968 36176 14980
rect 36228 14968 36234 15020
rect 36354 14968 36360 15020
rect 36412 15008 36418 15020
rect 37829 15011 37887 15017
rect 37829 15008 37841 15011
rect 36412 14980 37841 15008
rect 36412 14968 36418 14980
rect 37829 14977 37841 14980
rect 37875 14977 37887 15011
rect 37829 14971 37887 14977
rect 35986 14940 35992 14952
rect 35268 14912 35992 14940
rect 35986 14900 35992 14912
rect 36044 14900 36050 14952
rect 31628 14776 34836 14804
rect 35621 14807 35679 14813
rect 31628 14764 31634 14776
rect 35621 14773 35633 14807
rect 35667 14804 35679 14807
rect 36354 14804 36360 14816
rect 35667 14776 36360 14804
rect 35667 14773 35679 14776
rect 35621 14767 35679 14773
rect 36354 14764 36360 14776
rect 36412 14764 36418 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 18506 14560 18512 14612
rect 18564 14600 18570 14612
rect 18877 14603 18935 14609
rect 18877 14600 18889 14603
rect 18564 14572 18889 14600
rect 18564 14560 18570 14572
rect 18877 14569 18889 14572
rect 18923 14569 18935 14603
rect 18877 14563 18935 14569
rect 21082 14560 21088 14612
rect 21140 14600 21146 14612
rect 23201 14603 23259 14609
rect 23201 14600 23213 14603
rect 21140 14572 23213 14600
rect 21140 14560 21146 14572
rect 23201 14569 23213 14572
rect 23247 14569 23259 14603
rect 23201 14563 23259 14569
rect 23845 14603 23903 14609
rect 23845 14569 23857 14603
rect 23891 14600 23903 14603
rect 23934 14600 23940 14612
rect 23891 14572 23940 14600
rect 23891 14569 23903 14572
rect 23845 14563 23903 14569
rect 18785 14535 18843 14541
rect 18785 14501 18797 14535
rect 18831 14532 18843 14535
rect 19518 14532 19524 14544
rect 18831 14504 19524 14532
rect 18831 14501 18843 14504
rect 18785 14495 18843 14501
rect 19518 14492 19524 14504
rect 19576 14492 19582 14544
rect 19426 14356 19432 14408
rect 19484 14396 19490 14408
rect 19521 14399 19579 14405
rect 19521 14396 19533 14399
rect 19484 14368 19533 14396
rect 19484 14356 19490 14368
rect 19521 14365 19533 14368
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 20070 14356 20076 14408
rect 20128 14356 20134 14408
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14396 21879 14399
rect 22370 14396 22376 14408
rect 21867 14368 22376 14396
rect 21867 14365 21879 14368
rect 21821 14359 21879 14365
rect 22370 14356 22376 14368
rect 22428 14396 22434 14408
rect 22646 14396 22652 14408
rect 22428 14368 22652 14396
rect 22428 14356 22434 14368
rect 22646 14356 22652 14368
rect 22704 14356 22710 14408
rect 18417 14331 18475 14337
rect 18417 14297 18429 14331
rect 18463 14328 18475 14331
rect 19334 14328 19340 14340
rect 18463 14300 19340 14328
rect 18463 14297 18475 14300
rect 18417 14291 18475 14297
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 22094 14337 22100 14340
rect 19720 14300 20470 14328
rect 19242 14220 19248 14272
rect 19300 14260 19306 14272
rect 19720 14260 19748 14300
rect 22088 14291 22100 14337
rect 22094 14288 22100 14291
rect 22152 14288 22158 14340
rect 23216 14328 23244 14563
rect 23934 14560 23940 14572
rect 23992 14600 23998 14612
rect 24670 14600 24676 14612
rect 23992 14572 24676 14600
rect 23992 14560 23998 14572
rect 24670 14560 24676 14572
rect 24728 14560 24734 14612
rect 25041 14603 25099 14609
rect 25041 14569 25053 14603
rect 25087 14600 25099 14603
rect 27338 14600 27344 14612
rect 25087 14572 27344 14600
rect 25087 14569 25099 14572
rect 25041 14563 25099 14569
rect 27338 14560 27344 14572
rect 27396 14560 27402 14612
rect 32306 14560 32312 14612
rect 32364 14600 32370 14612
rect 33778 14600 33784 14612
rect 32364 14572 33784 14600
rect 32364 14560 32370 14572
rect 33778 14560 33784 14572
rect 33836 14560 33842 14612
rect 35802 14560 35808 14612
rect 35860 14600 35866 14612
rect 37093 14603 37151 14609
rect 37093 14600 37105 14603
rect 35860 14572 37105 14600
rect 35860 14560 35866 14572
rect 37093 14569 37105 14572
rect 37139 14569 37151 14603
rect 37093 14563 37151 14569
rect 27525 14535 27583 14541
rect 27525 14501 27537 14535
rect 27571 14532 27583 14535
rect 28350 14532 28356 14544
rect 27571 14504 28356 14532
rect 27571 14501 27583 14504
rect 27525 14495 27583 14501
rect 28350 14492 28356 14504
rect 28408 14492 28414 14544
rect 26050 14464 26056 14476
rect 25332 14436 26056 14464
rect 24026 14396 24032 14408
rect 23892 14371 24032 14396
rect 23891 14368 24032 14371
rect 23891 14365 23949 14368
rect 23661 14331 23719 14337
rect 23661 14328 23673 14331
rect 23216 14300 23673 14328
rect 23661 14297 23673 14300
rect 23707 14297 23719 14331
rect 23891 14331 23903 14365
rect 23937 14331 23949 14365
rect 24026 14356 24032 14368
rect 24084 14396 24090 14408
rect 24946 14396 24952 14408
rect 24084 14368 24952 14396
rect 24084 14356 24090 14368
rect 24946 14356 24952 14368
rect 25004 14356 25010 14408
rect 25332 14405 25360 14436
rect 26050 14424 26056 14436
rect 26108 14424 26114 14476
rect 27706 14424 27712 14476
rect 27764 14464 27770 14476
rect 28445 14467 28503 14473
rect 28445 14464 28457 14467
rect 27764 14436 28457 14464
rect 27764 14424 27770 14436
rect 28445 14433 28457 14436
rect 28491 14433 28503 14467
rect 28445 14427 28503 14433
rect 28534 14424 28540 14476
rect 28592 14424 28598 14476
rect 30650 14424 30656 14476
rect 30708 14464 30714 14476
rect 30708 14436 30880 14464
rect 30708 14424 30714 14436
rect 25317 14399 25375 14405
rect 25317 14365 25329 14399
rect 25363 14365 25375 14399
rect 25317 14359 25375 14365
rect 25409 14399 25467 14405
rect 25409 14365 25421 14399
rect 25455 14365 25467 14399
rect 25409 14359 25467 14365
rect 23891 14325 23949 14331
rect 23661 14291 23719 14297
rect 24854 14288 24860 14340
rect 24912 14328 24918 14340
rect 25424 14328 25452 14359
rect 25498 14356 25504 14408
rect 25556 14356 25562 14408
rect 25685 14399 25743 14405
rect 25685 14365 25697 14399
rect 25731 14365 25743 14399
rect 25685 14359 25743 14365
rect 26145 14399 26203 14405
rect 26145 14365 26157 14399
rect 26191 14396 26203 14399
rect 26191 14368 26648 14396
rect 26191 14365 26203 14368
rect 26145 14359 26203 14365
rect 24912 14300 25452 14328
rect 24912 14288 24918 14300
rect 19300 14232 19748 14260
rect 19300 14220 19306 14232
rect 22370 14220 22376 14272
rect 22428 14260 22434 14272
rect 23474 14260 23480 14272
rect 22428 14232 23480 14260
rect 22428 14220 22434 14232
rect 23474 14220 23480 14232
rect 23532 14220 23538 14272
rect 24026 14220 24032 14272
rect 24084 14220 24090 14272
rect 25700 14260 25728 14359
rect 26620 14340 26648 14368
rect 27982 14356 27988 14408
rect 28040 14396 28046 14408
rect 28040 14368 28111 14396
rect 28040 14356 28046 14368
rect 26412 14331 26470 14337
rect 26412 14297 26424 14331
rect 26458 14328 26470 14331
rect 26458 14300 26556 14328
rect 26458 14297 26470 14300
rect 26412 14291 26470 14297
rect 26326 14260 26332 14272
rect 25700 14232 26332 14260
rect 26326 14220 26332 14232
rect 26384 14220 26390 14272
rect 26528 14260 26556 14300
rect 26602 14288 26608 14340
rect 26660 14288 26666 14340
rect 26712 14300 28028 14328
rect 26712 14260 26740 14300
rect 28000 14269 28028 14300
rect 26528 14232 26740 14260
rect 27985 14263 28043 14269
rect 27985 14229 27997 14263
rect 28031 14229 28043 14263
rect 28083 14260 28111 14368
rect 28350 14356 28356 14408
rect 28408 14356 28414 14408
rect 30852 14405 30880 14436
rect 38102 14424 38108 14476
rect 38160 14424 38166 14476
rect 30745 14399 30803 14405
rect 30745 14365 30757 14399
rect 30791 14365 30803 14399
rect 30745 14359 30803 14365
rect 30837 14399 30895 14405
rect 30837 14365 30849 14399
rect 30883 14396 30895 14399
rect 31018 14396 31024 14408
rect 30883 14368 31024 14396
rect 30883 14365 30895 14368
rect 30837 14359 30895 14365
rect 30760 14328 30788 14359
rect 31018 14356 31024 14368
rect 31076 14356 31082 14408
rect 31941 14399 31999 14405
rect 31941 14365 31953 14399
rect 31987 14396 31999 14399
rect 33042 14396 33048 14408
rect 31987 14368 33048 14396
rect 31987 14365 31999 14368
rect 31941 14359 31999 14365
rect 33042 14356 33048 14368
rect 33100 14396 33106 14408
rect 34790 14396 34796 14408
rect 33100 14368 34796 14396
rect 33100 14356 33106 14368
rect 34790 14356 34796 14368
rect 34848 14396 34854 14408
rect 34885 14399 34943 14405
rect 34885 14396 34897 14399
rect 34848 14368 34897 14396
rect 34848 14356 34854 14368
rect 34885 14365 34897 14368
rect 34931 14365 34943 14399
rect 36078 14396 36084 14408
rect 34885 14359 34943 14365
rect 34992 14368 36084 14396
rect 30926 14328 30932 14340
rect 30760 14300 30932 14328
rect 30926 14288 30932 14300
rect 30984 14288 30990 14340
rect 32030 14288 32036 14340
rect 32088 14328 32094 14340
rect 32186 14331 32244 14337
rect 32186 14328 32198 14331
rect 32088 14300 32198 14328
rect 32088 14288 32094 14300
rect 32186 14297 32198 14300
rect 32232 14297 32244 14331
rect 32186 14291 32244 14297
rect 33962 14288 33968 14340
rect 34020 14288 34026 14340
rect 34146 14288 34152 14340
rect 34204 14288 34210 14340
rect 34333 14331 34391 14337
rect 34333 14297 34345 14331
rect 34379 14328 34391 14331
rect 34992 14328 35020 14368
rect 36078 14356 36084 14368
rect 36136 14396 36142 14408
rect 36909 14399 36967 14405
rect 36909 14396 36921 14399
rect 36136 14368 36921 14396
rect 36136 14356 36142 14368
rect 36909 14365 36921 14368
rect 36955 14365 36967 14399
rect 36909 14359 36967 14365
rect 37829 14399 37887 14405
rect 37829 14365 37841 14399
rect 37875 14396 37887 14399
rect 37918 14396 37924 14408
rect 37875 14368 37924 14396
rect 37875 14365 37887 14368
rect 37829 14359 37887 14365
rect 37918 14356 37924 14368
rect 37976 14356 37982 14408
rect 34379 14300 35020 14328
rect 35130 14331 35188 14337
rect 34379 14297 34391 14300
rect 34333 14291 34391 14297
rect 35130 14297 35142 14331
rect 35176 14297 35188 14331
rect 35130 14291 35188 14297
rect 30377 14263 30435 14269
rect 30377 14260 30389 14263
rect 28083 14232 30389 14260
rect 27985 14223 28043 14229
rect 30377 14229 30389 14232
rect 30423 14260 30435 14263
rect 32490 14260 32496 14272
rect 30423 14232 32496 14260
rect 30423 14229 30435 14232
rect 30377 14223 30435 14229
rect 32490 14220 32496 14232
rect 32548 14260 32554 14272
rect 33226 14260 33232 14272
rect 32548 14232 33232 14260
rect 32548 14220 32554 14232
rect 33226 14220 33232 14232
rect 33284 14220 33290 14272
rect 33318 14220 33324 14272
rect 33376 14220 33382 14272
rect 34790 14220 34796 14272
rect 34848 14260 34854 14272
rect 35145 14260 35173 14291
rect 36722 14288 36728 14340
rect 36780 14288 36786 14340
rect 37550 14288 37556 14340
rect 37608 14288 37614 14340
rect 34848 14232 35173 14260
rect 34848 14220 34854 14232
rect 35342 14220 35348 14272
rect 35400 14260 35406 14272
rect 36265 14263 36323 14269
rect 36265 14260 36277 14263
rect 35400 14232 36277 14260
rect 35400 14220 35406 14232
rect 36265 14229 36277 14232
rect 36311 14229 36323 14263
rect 36265 14223 36323 14229
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 18969 14059 19027 14065
rect 18969 14025 18981 14059
rect 19015 14056 19027 14059
rect 21269 14059 21327 14065
rect 19015 14028 20668 14056
rect 19015 14025 19027 14028
rect 18969 14019 19027 14025
rect 20640 13988 20668 14028
rect 21269 14025 21281 14059
rect 21315 14056 21327 14059
rect 22370 14056 22376 14068
rect 21315 14028 22376 14056
rect 21315 14025 21327 14028
rect 21269 14019 21327 14025
rect 22370 14016 22376 14028
rect 22428 14016 22434 14068
rect 22462 14016 22468 14068
rect 22520 14056 22526 14068
rect 22922 14056 22928 14068
rect 22520 14028 22928 14056
rect 22520 14016 22526 14028
rect 22922 14016 22928 14028
rect 22980 14016 22986 14068
rect 23014 14016 23020 14068
rect 23072 14056 23078 14068
rect 25498 14056 25504 14068
rect 23072 14028 25504 14056
rect 23072 14016 23078 14028
rect 23198 13988 23204 14000
rect 20640 13960 23204 13988
rect 23198 13948 23204 13960
rect 23256 13948 23262 14000
rect 23566 13948 23572 14000
rect 23624 13988 23630 14000
rect 24044 13997 24072 14028
rect 25498 14016 25504 14028
rect 25556 14056 25562 14068
rect 26142 14056 26148 14068
rect 25556 14028 26148 14056
rect 25556 14016 25562 14028
rect 26142 14016 26148 14028
rect 26200 14016 26206 14068
rect 27430 14016 27436 14068
rect 27488 14056 27494 14068
rect 27801 14059 27859 14065
rect 27801 14056 27813 14059
rect 27488 14028 27813 14056
rect 27488 14016 27494 14028
rect 27801 14025 27813 14028
rect 27847 14025 27859 14059
rect 27801 14019 27859 14025
rect 28902 14016 28908 14068
rect 28960 14056 28966 14068
rect 31665 14059 31723 14065
rect 31665 14056 31677 14059
rect 28960 14028 31677 14056
rect 28960 14016 28966 14028
rect 31665 14025 31677 14028
rect 31711 14025 31723 14059
rect 31665 14019 31723 14025
rect 32677 14059 32735 14065
rect 32677 14025 32689 14059
rect 32723 14056 32735 14059
rect 32766 14056 32772 14068
rect 32723 14028 32772 14056
rect 32723 14025 32735 14028
rect 32677 14019 32735 14025
rect 32766 14016 32772 14028
rect 32824 14016 32830 14068
rect 33962 14016 33968 14068
rect 34020 14056 34026 14068
rect 36081 14059 36139 14065
rect 36081 14056 36093 14059
rect 34020 14028 36093 14056
rect 34020 14016 34026 14028
rect 36081 14025 36093 14028
rect 36127 14025 36139 14059
rect 36081 14019 36139 14025
rect 36449 14059 36507 14065
rect 36449 14025 36461 14059
rect 36495 14025 36507 14059
rect 36449 14019 36507 14025
rect 23937 13991 23995 13997
rect 23937 13988 23949 13991
rect 23624 13960 23949 13988
rect 23624 13948 23630 13960
rect 23937 13957 23949 13960
rect 23983 13957 23995 13991
rect 23937 13951 23995 13957
rect 24029 13991 24087 13997
rect 24029 13957 24041 13991
rect 24075 13957 24087 13991
rect 27522 13988 27528 14000
rect 24029 13951 24087 13957
rect 24780 13960 27528 13988
rect 18782 13880 18788 13932
rect 18840 13880 18846 13932
rect 18966 13880 18972 13932
rect 19024 13880 19030 13932
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 19981 13923 20039 13929
rect 19981 13920 19993 13923
rect 19300 13892 19993 13920
rect 19300 13880 19306 13892
rect 19981 13889 19993 13892
rect 20027 13889 20039 13923
rect 19981 13883 20039 13889
rect 22370 13880 22376 13932
rect 22428 13880 22434 13932
rect 23382 13880 23388 13932
rect 23440 13920 23446 13932
rect 24780 13929 24808 13960
rect 27522 13948 27528 13960
rect 27580 13948 27586 14000
rect 29638 13988 29644 14000
rect 28368 13960 29644 13988
rect 28368 13932 28396 13960
rect 29638 13948 29644 13960
rect 29696 13948 29702 14000
rect 29825 13991 29883 13997
rect 29825 13957 29837 13991
rect 29871 13988 29883 13991
rect 29914 13988 29920 14000
rect 29871 13960 29920 13988
rect 29871 13957 29883 13960
rect 29825 13951 29883 13957
rect 29914 13948 29920 13960
rect 29972 13948 29978 14000
rect 30009 13991 30067 13997
rect 30009 13957 30021 13991
rect 30055 13988 30067 13991
rect 30055 13960 31156 13988
rect 30055 13957 30067 13960
rect 30009 13951 30067 13957
rect 24765 13923 24823 13929
rect 24765 13920 24777 13923
rect 23440 13892 24777 13920
rect 23440 13880 23446 13892
rect 24765 13889 24777 13892
rect 24811 13889 24823 13923
rect 24765 13883 24823 13889
rect 25032 13923 25090 13929
rect 25032 13889 25044 13923
rect 25078 13920 25090 13923
rect 25314 13920 25320 13932
rect 25078 13892 25320 13920
rect 25078 13889 25090 13892
rect 25032 13883 25090 13889
rect 25314 13880 25320 13892
rect 25372 13880 25378 13932
rect 28350 13880 28356 13932
rect 28408 13880 28414 13932
rect 28445 13923 28503 13929
rect 28445 13889 28457 13923
rect 28491 13920 28503 13923
rect 30650 13920 30656 13932
rect 28491 13892 30656 13920
rect 28491 13889 28503 13892
rect 28445 13883 28503 13889
rect 18690 13812 18696 13864
rect 18748 13852 18754 13864
rect 19426 13852 19432 13864
rect 18748 13824 19432 13852
rect 18748 13812 18754 13824
rect 19426 13812 19432 13824
rect 19484 13852 19490 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19484 13824 19717 13852
rect 19484 13812 19490 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 22649 13855 22707 13861
rect 22649 13821 22661 13855
rect 22695 13852 22707 13855
rect 22738 13852 22744 13864
rect 22695 13824 22744 13852
rect 22695 13821 22707 13824
rect 22649 13815 22707 13821
rect 22738 13812 22744 13824
rect 22796 13812 22802 13864
rect 23934 13812 23940 13864
rect 23992 13812 23998 13864
rect 24044 13824 24808 13852
rect 20714 13744 20720 13796
rect 20772 13784 20778 13796
rect 23106 13784 23112 13796
rect 20772 13756 23112 13784
rect 20772 13744 20778 13756
rect 23106 13744 23112 13756
rect 23164 13744 23170 13796
rect 23477 13787 23535 13793
rect 23477 13753 23489 13787
rect 23523 13784 23535 13787
rect 24044 13784 24072 13824
rect 23523 13756 24072 13784
rect 23523 13753 23535 13756
rect 23477 13747 23535 13753
rect 22002 13676 22008 13728
rect 22060 13676 22066 13728
rect 22830 13676 22836 13728
rect 22888 13716 22894 13728
rect 23198 13716 23204 13728
rect 22888 13688 23204 13716
rect 22888 13676 22894 13688
rect 23198 13676 23204 13688
rect 23256 13676 23262 13728
rect 24780 13716 24808 13824
rect 25792 13824 27568 13852
rect 25792 13716 25820 13824
rect 27540 13784 27568 13824
rect 27614 13812 27620 13864
rect 27672 13852 27678 13864
rect 28460 13852 28488 13883
rect 30650 13880 30656 13892
rect 30708 13880 30714 13932
rect 30742 13880 30748 13932
rect 30800 13880 30806 13932
rect 30837 13923 30895 13929
rect 30837 13889 30849 13923
rect 30883 13889 30895 13923
rect 30837 13883 30895 13889
rect 30929 13923 30987 13929
rect 30929 13889 30941 13923
rect 30975 13920 30987 13923
rect 31018 13920 31024 13932
rect 30975 13892 31024 13920
rect 30975 13889 30987 13892
rect 30929 13883 30987 13889
rect 27672 13824 28488 13852
rect 27672 13812 27678 13824
rect 28994 13812 29000 13864
rect 29052 13852 29058 13864
rect 30852 13852 30880 13883
rect 31018 13880 31024 13892
rect 31076 13880 31082 13932
rect 31128 13929 31156 13960
rect 34514 13948 34520 14000
rect 34572 13988 34578 14000
rect 34946 13991 35004 13997
rect 34946 13988 34958 13991
rect 34572 13960 34958 13988
rect 34572 13948 34578 13960
rect 34946 13957 34958 13960
rect 34992 13957 35004 13991
rect 36464 13988 36492 14019
rect 36814 14016 36820 14068
rect 36872 14016 36878 14068
rect 37550 14016 37556 14068
rect 37608 14056 37614 14068
rect 38121 14059 38179 14065
rect 38121 14056 38133 14059
rect 37608 14028 38133 14056
rect 37608 14016 37614 14028
rect 38121 14025 38133 14028
rect 38167 14025 38179 14059
rect 38121 14019 38179 14025
rect 38289 14059 38347 14065
rect 38289 14025 38301 14059
rect 38335 14056 38347 14059
rect 39482 14056 39488 14068
rect 38335 14028 39488 14056
rect 38335 14025 38347 14028
rect 38289 14019 38347 14025
rect 39482 14016 39488 14028
rect 39540 14016 39546 14068
rect 37734 13988 37740 14000
rect 36464 13960 37740 13988
rect 34946 13951 35004 13957
rect 37734 13948 37740 13960
rect 37792 13948 37798 14000
rect 37921 13991 37979 13997
rect 37921 13957 37933 13991
rect 37967 13988 37979 13991
rect 39390 13988 39396 14000
rect 37967 13960 39396 13988
rect 37967 13957 37979 13960
rect 37921 13951 37979 13957
rect 31113 13923 31171 13929
rect 31113 13889 31125 13923
rect 31159 13889 31171 13923
rect 31113 13883 31171 13889
rect 31570 13880 31576 13932
rect 31628 13880 31634 13932
rect 31662 13880 31668 13932
rect 31720 13920 31726 13932
rect 32401 13923 32459 13929
rect 32401 13920 32413 13923
rect 31720 13892 32413 13920
rect 31720 13880 31726 13892
rect 32401 13889 32413 13892
rect 32447 13889 32459 13923
rect 32401 13883 32459 13889
rect 33226 13880 33232 13932
rect 33284 13880 33290 13932
rect 33502 13880 33508 13932
rect 33560 13920 33566 13932
rect 33597 13923 33655 13929
rect 33597 13920 33609 13923
rect 33560 13892 33609 13920
rect 33560 13880 33566 13892
rect 33597 13889 33609 13892
rect 33643 13889 33655 13923
rect 33597 13883 33655 13889
rect 33873 13923 33931 13929
rect 33873 13889 33885 13923
rect 33919 13889 33931 13923
rect 33873 13883 33931 13889
rect 29052 13824 30880 13852
rect 33413 13855 33471 13861
rect 29052 13812 29058 13824
rect 33413 13821 33425 13855
rect 33459 13821 33471 13855
rect 33888 13852 33916 13883
rect 34698 13880 34704 13932
rect 34756 13880 34762 13932
rect 35342 13920 35348 13932
rect 34808 13892 35348 13920
rect 34808 13852 34836 13892
rect 35342 13880 35348 13892
rect 35400 13880 35406 13932
rect 35526 13880 35532 13932
rect 35584 13920 35590 13932
rect 36265 13923 36323 13929
rect 36265 13920 36277 13923
rect 35584 13892 36277 13920
rect 35584 13880 35590 13892
rect 36265 13889 36277 13892
rect 36311 13889 36323 13923
rect 36265 13883 36323 13889
rect 37645 13923 37703 13929
rect 37645 13889 37657 13923
rect 37691 13920 37703 13923
rect 37936 13920 37964 13951
rect 39390 13948 39396 13960
rect 39448 13948 39454 14000
rect 37691 13892 37964 13920
rect 37691 13889 37703 13892
rect 37645 13883 37703 13889
rect 33888 13824 34836 13852
rect 33413 13815 33471 13821
rect 27890 13784 27896 13796
rect 27540 13756 27896 13784
rect 27890 13744 27896 13756
rect 27948 13784 27954 13796
rect 28810 13784 28816 13796
rect 27948 13756 28816 13784
rect 27948 13744 27954 13756
rect 28810 13744 28816 13756
rect 28868 13744 28874 13796
rect 30466 13744 30472 13796
rect 30524 13744 30530 13796
rect 33428 13784 33456 13815
rect 33962 13784 33968 13796
rect 33428 13756 33968 13784
rect 33962 13744 33968 13756
rect 34020 13744 34026 13796
rect 36814 13744 36820 13796
rect 36872 13784 36878 13796
rect 36872 13756 38148 13784
rect 36872 13744 36878 13756
rect 24780 13688 25820 13716
rect 26142 13676 26148 13728
rect 26200 13676 26206 13728
rect 32950 13676 32956 13728
rect 33008 13716 33014 13728
rect 36262 13716 36268 13728
rect 33008 13688 36268 13716
rect 33008 13676 33014 13688
rect 36262 13676 36268 13688
rect 36320 13676 36326 13728
rect 38120 13725 38148 13756
rect 38105 13719 38163 13725
rect 38105 13685 38117 13719
rect 38151 13685 38163 13719
rect 38105 13679 38163 13685
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 19392 13484 19441 13512
rect 19392 13472 19398 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 19429 13475 19487 13481
rect 20257 13515 20315 13521
rect 20257 13481 20269 13515
rect 20303 13512 20315 13515
rect 22189 13515 22247 13521
rect 20303 13484 22094 13512
rect 20303 13481 20315 13484
rect 20257 13475 20315 13481
rect 22066 13444 22094 13484
rect 22189 13481 22201 13515
rect 22235 13512 22247 13515
rect 22370 13512 22376 13524
rect 22235 13484 22376 13512
rect 22235 13481 22247 13484
rect 22189 13475 22247 13481
rect 22370 13472 22376 13484
rect 22428 13472 22434 13524
rect 23566 13512 23572 13524
rect 22480 13484 23572 13512
rect 22480 13444 22508 13484
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 23934 13472 23940 13524
rect 23992 13512 23998 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 23992 13484 24593 13512
rect 23992 13472 23998 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 25314 13472 25320 13524
rect 25372 13472 25378 13524
rect 27338 13512 27344 13524
rect 25976 13484 27344 13512
rect 22066 13416 22508 13444
rect 24029 13447 24087 13453
rect 24029 13413 24041 13447
rect 24075 13444 24087 13447
rect 24302 13444 24308 13456
rect 24075 13416 24308 13444
rect 24075 13413 24087 13416
rect 24029 13407 24087 13413
rect 24302 13404 24308 13416
rect 24360 13404 24366 13456
rect 19978 13376 19984 13388
rect 19444 13348 19984 13376
rect 19444 13317 19472 13348
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 20349 13379 20407 13385
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 20714 13376 20720 13388
rect 20395 13348 20720 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 20714 13336 20720 13348
rect 20772 13336 20778 13388
rect 22646 13336 22652 13388
rect 22704 13336 22710 13388
rect 24210 13336 24216 13388
rect 24268 13376 24274 13388
rect 25976 13385 26004 13484
rect 27338 13472 27344 13484
rect 27396 13472 27402 13524
rect 31941 13515 31999 13521
rect 31941 13481 31953 13515
rect 31987 13512 31999 13515
rect 32030 13512 32036 13524
rect 31987 13484 32036 13512
rect 31987 13481 31999 13484
rect 31941 13475 31999 13481
rect 32030 13472 32036 13484
rect 32088 13472 32094 13524
rect 33597 13515 33655 13521
rect 33597 13481 33609 13515
rect 33643 13512 33655 13515
rect 34514 13512 34520 13524
rect 33643 13484 34520 13512
rect 33643 13481 33655 13484
rect 33597 13475 33655 13481
rect 34514 13472 34520 13484
rect 34572 13472 34578 13524
rect 34790 13472 34796 13524
rect 34848 13512 34854 13524
rect 34885 13515 34943 13521
rect 34885 13512 34897 13515
rect 34848 13484 34897 13512
rect 34848 13472 34854 13484
rect 34885 13481 34897 13484
rect 34931 13481 34943 13515
rect 34885 13475 34943 13481
rect 36817 13515 36875 13521
rect 36817 13481 36829 13515
rect 36863 13512 36875 13515
rect 37274 13512 37280 13524
rect 36863 13484 37280 13512
rect 36863 13481 36875 13484
rect 36817 13475 36875 13481
rect 37274 13472 37280 13484
rect 37332 13472 37338 13524
rect 38289 13515 38347 13521
rect 38289 13481 38301 13515
rect 38335 13512 38347 13515
rect 39022 13512 39028 13524
rect 38335 13484 39028 13512
rect 38335 13481 38347 13484
rect 38289 13475 38347 13481
rect 39022 13472 39028 13484
rect 39080 13472 39086 13524
rect 31478 13404 31484 13456
rect 31536 13444 31542 13456
rect 31536 13416 32444 13444
rect 31536 13404 31542 13416
rect 25961 13379 26019 13385
rect 25961 13376 25973 13379
rect 24268 13348 25973 13376
rect 24268 13336 24274 13348
rect 25961 13345 25973 13348
rect 26007 13345 26019 13379
rect 25961 13339 26019 13345
rect 26344 13348 26924 13376
rect 26344 13320 26372 13348
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 20073 13311 20131 13317
rect 20073 13277 20085 13311
rect 20119 13277 20131 13311
rect 20073 13271 20131 13277
rect 20165 13311 20223 13317
rect 20165 13277 20177 13311
rect 20211 13308 20223 13311
rect 20530 13308 20536 13320
rect 20211 13280 20536 13308
rect 20211 13277 20223 13280
rect 20165 13271 20223 13277
rect 19628 13172 19656 13271
rect 20088 13240 20116 13271
rect 20530 13268 20536 13280
rect 20588 13268 20594 13320
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 23382 13308 23388 13320
rect 20855 13280 23388 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 24026 13268 24032 13320
rect 24084 13308 24090 13320
rect 24581 13311 24639 13317
rect 24581 13308 24593 13311
rect 24084 13280 24593 13308
rect 24084 13268 24090 13280
rect 24581 13277 24593 13280
rect 24627 13277 24639 13311
rect 24581 13271 24639 13277
rect 24762 13268 24768 13320
rect 24820 13268 24826 13320
rect 24854 13268 24860 13320
rect 24912 13268 24918 13320
rect 25682 13268 25688 13320
rect 25740 13308 25746 13320
rect 26142 13308 26148 13320
rect 25740 13280 26148 13308
rect 25740 13268 25746 13280
rect 26142 13268 26148 13280
rect 26200 13268 26206 13320
rect 26326 13268 26332 13320
rect 26384 13268 26390 13320
rect 26896 13317 26924 13348
rect 27522 13336 27528 13388
rect 27580 13376 27586 13388
rect 27798 13376 27804 13388
rect 27580 13348 27804 13376
rect 27580 13336 27586 13348
rect 27798 13336 27804 13348
rect 27856 13336 27862 13388
rect 29822 13336 29828 13388
rect 29880 13336 29886 13388
rect 32416 13385 32444 13416
rect 34238 13404 34244 13456
rect 34296 13444 34302 13456
rect 34296 13416 35572 13444
rect 34296 13404 34302 13416
rect 32401 13379 32459 13385
rect 32401 13345 32413 13379
rect 32447 13345 32459 13379
rect 32401 13339 32459 13345
rect 32490 13336 32496 13388
rect 32548 13376 32554 13388
rect 34149 13379 34207 13385
rect 34149 13376 34161 13379
rect 32548 13348 34161 13376
rect 32548 13336 32554 13348
rect 34149 13345 34161 13348
rect 34195 13376 34207 13379
rect 35158 13376 35164 13388
rect 34195 13348 35164 13376
rect 34195 13345 34207 13348
rect 34149 13339 34207 13345
rect 35158 13336 35164 13348
rect 35216 13336 35222 13388
rect 35434 13336 35440 13388
rect 35492 13336 35498 13388
rect 35544 13376 35572 13416
rect 36078 13404 36084 13456
rect 36136 13404 36142 13456
rect 37461 13379 37519 13385
rect 35544 13348 36768 13376
rect 26605 13311 26663 13317
rect 26605 13277 26617 13311
rect 26651 13277 26663 13311
rect 26605 13271 26663 13277
rect 26881 13311 26939 13317
rect 26881 13277 26893 13311
rect 26927 13308 26939 13311
rect 27890 13308 27896 13320
rect 26927 13280 27896 13308
rect 26927 13277 26939 13280
rect 26881 13271 26939 13277
rect 21076 13243 21134 13249
rect 20088 13212 21036 13240
rect 20254 13172 20260 13184
rect 19628 13144 20260 13172
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 21008 13172 21036 13212
rect 21076 13209 21088 13243
rect 21122 13240 21134 13243
rect 22002 13240 22008 13252
rect 21122 13212 22008 13240
rect 21122 13209 21134 13212
rect 21076 13203 21134 13209
rect 22002 13200 22008 13212
rect 22060 13200 22066 13252
rect 22916 13243 22974 13249
rect 22916 13209 22928 13243
rect 22962 13240 22974 13243
rect 23566 13240 23572 13252
rect 22962 13212 23572 13240
rect 22962 13209 22974 13212
rect 22916 13203 22974 13209
rect 23566 13200 23572 13212
rect 23624 13200 23630 13252
rect 24872 13240 24900 13268
rect 26620 13240 26648 13271
rect 27890 13268 27896 13280
rect 27948 13268 27954 13320
rect 28810 13268 28816 13320
rect 28868 13308 28874 13320
rect 32122 13308 32128 13320
rect 28868 13280 32128 13308
rect 28868 13268 28874 13280
rect 32122 13268 32128 13280
rect 32180 13268 32186 13320
rect 34057 13311 34115 13317
rect 34057 13277 34069 13311
rect 34103 13308 34115 13311
rect 35345 13311 35403 13317
rect 35345 13308 35357 13311
rect 34103 13280 35357 13308
rect 34103 13277 34115 13280
rect 34057 13271 34115 13277
rect 35345 13277 35357 13280
rect 35391 13277 35403 13311
rect 35345 13271 35403 13277
rect 24872 13212 26648 13240
rect 26789 13243 26847 13249
rect 26789 13209 26801 13243
rect 26835 13209 26847 13243
rect 26789 13203 26847 13209
rect 22370 13172 22376 13184
rect 21008 13144 22376 13172
rect 22370 13132 22376 13144
rect 22428 13132 22434 13184
rect 25590 13132 25596 13184
rect 25648 13172 25654 13184
rect 25777 13175 25835 13181
rect 25777 13172 25789 13175
rect 25648 13144 25789 13172
rect 25648 13132 25654 13144
rect 25777 13141 25789 13144
rect 25823 13141 25835 13175
rect 25777 13135 25835 13141
rect 26234 13132 26240 13184
rect 26292 13172 26298 13184
rect 26804 13172 26832 13203
rect 27338 13200 27344 13252
rect 27396 13200 27402 13252
rect 28068 13243 28126 13249
rect 28068 13209 28080 13243
rect 28114 13240 28126 13243
rect 28626 13240 28632 13252
rect 28114 13212 28632 13240
rect 28114 13209 28126 13212
rect 28068 13203 28126 13209
rect 28626 13200 28632 13212
rect 28684 13200 28690 13252
rect 30092 13243 30150 13249
rect 30092 13209 30104 13243
rect 30138 13240 30150 13243
rect 30282 13240 30288 13252
rect 30138 13212 30288 13240
rect 30138 13209 30150 13212
rect 30092 13203 30150 13209
rect 30282 13200 30288 13212
rect 30340 13200 30346 13252
rect 30742 13240 30748 13252
rect 30392 13212 30748 13240
rect 26878 13172 26884 13184
rect 26292 13144 26884 13172
rect 26292 13132 26298 13144
rect 26878 13132 26884 13144
rect 26936 13172 26942 13184
rect 27614 13172 27620 13184
rect 26936 13144 27620 13172
rect 26936 13132 26942 13144
rect 27614 13132 27620 13144
rect 27672 13132 27678 13184
rect 29181 13175 29239 13181
rect 29181 13141 29193 13175
rect 29227 13172 29239 13175
rect 29270 13172 29276 13184
rect 29227 13144 29276 13172
rect 29227 13141 29239 13144
rect 29181 13135 29239 13141
rect 29270 13132 29276 13144
rect 29328 13132 29334 13184
rect 29454 13132 29460 13184
rect 29512 13172 29518 13184
rect 30392 13172 30420 13212
rect 30742 13200 30748 13212
rect 30800 13240 30806 13252
rect 34072 13240 34100 13271
rect 35986 13268 35992 13320
rect 36044 13308 36050 13320
rect 36081 13311 36139 13317
rect 36081 13308 36093 13311
rect 36044 13280 36093 13308
rect 36044 13268 36050 13280
rect 36081 13277 36093 13280
rect 36127 13277 36139 13311
rect 36081 13271 36139 13277
rect 36262 13268 36268 13320
rect 36320 13268 36326 13320
rect 36740 13317 36768 13348
rect 37461 13345 37473 13379
rect 37507 13376 37519 13379
rect 38654 13376 38660 13388
rect 37507 13348 38660 13376
rect 37507 13345 37519 13348
rect 37461 13339 37519 13345
rect 38654 13336 38660 13348
rect 38712 13336 38718 13388
rect 36725 13311 36783 13317
rect 36725 13277 36737 13311
rect 36771 13277 36783 13311
rect 36725 13271 36783 13277
rect 36906 13268 36912 13320
rect 36964 13268 36970 13320
rect 37366 13268 37372 13320
rect 37424 13268 37430 13320
rect 37553 13311 37611 13317
rect 37553 13277 37565 13311
rect 37599 13308 37611 13311
rect 37642 13308 37648 13320
rect 37599 13280 37648 13308
rect 37599 13277 37611 13280
rect 37553 13271 37611 13277
rect 37642 13268 37648 13280
rect 37700 13268 37706 13320
rect 30800 13212 34100 13240
rect 30800 13200 30806 13212
rect 29512 13144 30420 13172
rect 29512 13132 29518 13144
rect 30650 13132 30656 13184
rect 30708 13172 30714 13184
rect 31205 13175 31263 13181
rect 31205 13172 31217 13175
rect 30708 13144 31217 13172
rect 30708 13132 30714 13144
rect 31205 13141 31217 13144
rect 31251 13141 31263 13175
rect 31205 13135 31263 13141
rect 32309 13175 32367 13181
rect 32309 13141 32321 13175
rect 32355 13172 32367 13175
rect 33318 13172 33324 13184
rect 32355 13144 33324 13172
rect 32355 13141 32367 13144
rect 32309 13135 32367 13141
rect 33318 13132 33324 13144
rect 33376 13132 33382 13184
rect 33962 13132 33968 13184
rect 34020 13132 34026 13184
rect 35253 13175 35311 13181
rect 35253 13141 35265 13175
rect 35299 13172 35311 13175
rect 35342 13172 35348 13184
rect 35299 13144 35348 13172
rect 35299 13141 35311 13144
rect 35253 13135 35311 13141
rect 35342 13132 35348 13144
rect 35400 13132 35406 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 23198 12968 23204 12980
rect 21284 12940 23204 12968
rect 20441 12903 20499 12909
rect 20441 12869 20453 12903
rect 20487 12900 20499 12903
rect 20898 12900 20904 12912
rect 20487 12872 20904 12900
rect 20487 12869 20499 12872
rect 20441 12863 20499 12869
rect 20898 12860 20904 12872
rect 20956 12860 20962 12912
rect 21284 12909 21312 12940
rect 23198 12928 23204 12940
rect 23256 12928 23262 12980
rect 23566 12928 23572 12980
rect 23624 12928 23630 12980
rect 23937 12971 23995 12977
rect 23937 12937 23949 12971
rect 23983 12968 23995 12971
rect 24302 12968 24308 12980
rect 23983 12940 24308 12968
rect 23983 12937 23995 12940
rect 23937 12931 23995 12937
rect 24302 12928 24308 12940
rect 24360 12928 24366 12980
rect 24670 12928 24676 12980
rect 24728 12928 24734 12980
rect 25958 12968 25964 12980
rect 25240 12940 25964 12968
rect 21269 12903 21327 12909
rect 21269 12869 21281 12903
rect 21315 12869 21327 12903
rect 21269 12863 21327 12869
rect 22922 12860 22928 12912
rect 22980 12900 22986 12912
rect 24029 12903 24087 12909
rect 24029 12900 24041 12903
rect 22980 12872 24041 12900
rect 22980 12860 22986 12872
rect 24029 12869 24041 12872
rect 24075 12869 24087 12903
rect 24029 12863 24087 12869
rect 20257 12835 20315 12841
rect 20257 12801 20269 12835
rect 20303 12832 20315 12835
rect 20346 12832 20352 12844
rect 20303 12804 20352 12832
rect 20303 12801 20315 12804
rect 20257 12795 20315 12801
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 20530 12792 20536 12844
rect 20588 12792 20594 12844
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12832 21051 12835
rect 22094 12832 22100 12844
rect 21039 12804 22100 12832
rect 21039 12801 21051 12804
rect 20993 12795 21051 12801
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 22649 12835 22707 12841
rect 22649 12801 22661 12835
rect 22695 12801 22707 12835
rect 22649 12795 22707 12801
rect 22557 12767 22615 12773
rect 22557 12733 22569 12767
rect 22603 12733 22615 12767
rect 22664 12764 22692 12795
rect 22738 12792 22744 12844
rect 22796 12832 22802 12844
rect 24688 12832 24716 12928
rect 24765 12835 24823 12841
rect 24765 12832 24777 12835
rect 22796 12804 24624 12832
rect 24688 12804 24777 12832
rect 22796 12792 22802 12804
rect 22664 12736 23796 12764
rect 22557 12727 22615 12733
rect 22572 12696 22600 12727
rect 23658 12696 23664 12708
rect 22572 12668 23664 12696
rect 23658 12656 23664 12668
rect 23716 12656 23722 12708
rect 23768 12696 23796 12736
rect 24210 12724 24216 12776
rect 24268 12724 24274 12776
rect 24596 12764 24624 12804
rect 24765 12801 24777 12804
rect 24811 12801 24823 12835
rect 24765 12795 24823 12801
rect 24857 12835 24915 12841
rect 24857 12801 24869 12835
rect 24903 12832 24915 12835
rect 24946 12832 24952 12844
rect 24903 12804 24952 12832
rect 24903 12801 24915 12804
rect 24857 12795 24915 12801
rect 24946 12792 24952 12804
rect 25004 12792 25010 12844
rect 25240 12764 25268 12940
rect 25958 12928 25964 12940
rect 26016 12968 26022 12980
rect 27890 12968 27896 12980
rect 26016 12940 27896 12968
rect 26016 12928 26022 12940
rect 27890 12928 27896 12940
rect 27948 12928 27954 12980
rect 28626 12928 28632 12980
rect 28684 12928 28690 12980
rect 29086 12928 29092 12980
rect 29144 12968 29150 12980
rect 29454 12968 29460 12980
rect 29144 12940 29460 12968
rect 29144 12928 29150 12940
rect 29454 12928 29460 12940
rect 29512 12928 29518 12980
rect 30282 12928 30288 12980
rect 30340 12928 30346 12980
rect 30650 12928 30656 12980
rect 30708 12928 30714 12980
rect 30742 12928 30748 12980
rect 30800 12928 30806 12980
rect 30834 12928 30840 12980
rect 30892 12968 30898 12980
rect 31665 12971 31723 12977
rect 31665 12968 31677 12971
rect 30892 12940 31677 12968
rect 30892 12928 30898 12940
rect 31665 12937 31677 12940
rect 31711 12937 31723 12971
rect 31665 12931 31723 12937
rect 35618 12928 35624 12980
rect 35676 12968 35682 12980
rect 35897 12971 35955 12977
rect 35897 12968 35909 12971
rect 35676 12940 35909 12968
rect 35676 12928 35682 12940
rect 35897 12937 35909 12940
rect 35943 12937 35955 12971
rect 35897 12931 35955 12937
rect 36541 12971 36599 12977
rect 36541 12937 36553 12971
rect 36587 12968 36599 12971
rect 38562 12968 38568 12980
rect 36587 12940 38568 12968
rect 36587 12937 36599 12940
rect 36541 12931 36599 12937
rect 38562 12928 38568 12940
rect 38620 12928 38626 12980
rect 25317 12903 25375 12909
rect 25317 12869 25329 12903
rect 25363 12900 25375 12903
rect 26050 12900 26056 12912
rect 25363 12872 26056 12900
rect 25363 12869 25375 12872
rect 25317 12863 25375 12869
rect 26050 12860 26056 12872
rect 26108 12900 26114 12912
rect 28350 12900 28356 12912
rect 26108 12872 28356 12900
rect 26108 12860 26114 12872
rect 26145 12835 26203 12841
rect 26145 12832 26157 12835
rect 24596 12736 25268 12764
rect 25332 12804 26157 12832
rect 25332 12696 25360 12804
rect 26145 12801 26157 12804
rect 26191 12832 26203 12835
rect 26326 12832 26332 12844
rect 26191 12804 26332 12832
rect 26191 12801 26203 12804
rect 26145 12795 26203 12801
rect 26326 12792 26332 12804
rect 26384 12792 26390 12844
rect 26602 12792 26608 12844
rect 26660 12832 26666 12844
rect 27062 12832 27068 12844
rect 26660 12804 27068 12832
rect 26660 12792 26666 12804
rect 27062 12792 27068 12804
rect 27120 12792 27126 12844
rect 27540 12841 27568 12872
rect 28350 12860 28356 12872
rect 28408 12860 28414 12912
rect 29362 12860 29368 12912
rect 29420 12900 29426 12912
rect 29420 12872 31616 12900
rect 29420 12860 29426 12872
rect 27525 12835 27583 12841
rect 27525 12801 27537 12835
rect 27571 12801 27583 12835
rect 27525 12795 27583 12801
rect 27614 12792 27620 12844
rect 27672 12792 27678 12844
rect 27709 12835 27767 12841
rect 27709 12801 27721 12835
rect 27755 12832 27767 12835
rect 28074 12832 28080 12844
rect 27755 12804 28080 12832
rect 27755 12801 27767 12804
rect 27709 12795 27767 12801
rect 28074 12792 28080 12804
rect 28132 12792 28138 12844
rect 28997 12835 29055 12841
rect 28997 12801 29009 12835
rect 29043 12832 29055 12835
rect 29270 12832 29276 12844
rect 29043 12804 29276 12832
rect 29043 12801 29055 12804
rect 28997 12795 29055 12801
rect 29270 12792 29276 12804
rect 29328 12832 29334 12844
rect 29914 12832 29920 12844
rect 29328 12804 29920 12832
rect 29328 12792 29334 12804
rect 29914 12792 29920 12804
rect 29972 12792 29978 12844
rect 30558 12792 30564 12844
rect 30616 12832 30622 12844
rect 31588 12841 31616 12872
rect 32122 12860 32128 12912
rect 32180 12900 32186 12912
rect 32180 12872 35848 12900
rect 32180 12860 32186 12872
rect 31573 12835 31631 12841
rect 30616 12804 31244 12832
rect 30616 12792 30622 12804
rect 26053 12767 26111 12773
rect 26053 12733 26065 12767
rect 26099 12764 26111 12767
rect 27430 12764 27436 12776
rect 26099 12736 27436 12764
rect 26099 12733 26111 12736
rect 26053 12727 26111 12733
rect 27430 12724 27436 12736
rect 27488 12724 27494 12776
rect 28258 12724 28264 12776
rect 28316 12764 28322 12776
rect 29086 12764 29092 12776
rect 28316 12736 29092 12764
rect 28316 12724 28322 12736
rect 29086 12724 29092 12736
rect 29144 12724 29150 12776
rect 29181 12767 29239 12773
rect 29181 12733 29193 12767
rect 29227 12764 29239 12767
rect 30190 12764 30196 12776
rect 29227 12736 30196 12764
rect 29227 12733 29239 12736
rect 29181 12727 29239 12733
rect 29196 12696 29224 12727
rect 30190 12724 30196 12736
rect 30248 12724 30254 12776
rect 30837 12767 30895 12773
rect 30837 12733 30849 12767
rect 30883 12764 30895 12767
rect 31110 12764 31116 12776
rect 30883 12736 31116 12764
rect 30883 12733 30895 12736
rect 30837 12727 30895 12733
rect 23768 12668 25360 12696
rect 27448 12668 29224 12696
rect 27448 12640 27476 12668
rect 20257 12631 20315 12637
rect 20257 12597 20269 12631
rect 20303 12628 20315 12631
rect 22002 12628 22008 12640
rect 20303 12600 22008 12628
rect 20303 12597 20315 12600
rect 20257 12591 20315 12597
rect 22002 12588 22008 12600
rect 22060 12588 22066 12640
rect 22278 12588 22284 12640
rect 22336 12628 22342 12640
rect 22833 12631 22891 12637
rect 22833 12628 22845 12631
rect 22336 12600 22845 12628
rect 22336 12588 22342 12600
rect 22833 12597 22845 12600
rect 22879 12628 22891 12631
rect 23842 12628 23848 12640
rect 22879 12600 23848 12628
rect 22879 12597 22891 12600
rect 22833 12591 22891 12597
rect 23842 12588 23848 12600
rect 23900 12588 23906 12640
rect 26326 12588 26332 12640
rect 26384 12628 26390 12640
rect 26786 12628 26792 12640
rect 26384 12600 26792 12628
rect 26384 12588 26390 12600
rect 26786 12588 26792 12600
rect 26844 12588 26850 12640
rect 27430 12588 27436 12640
rect 27488 12588 27494 12640
rect 27890 12588 27896 12640
rect 27948 12628 27954 12640
rect 30852 12628 30880 12727
rect 31110 12724 31116 12736
rect 31168 12724 31174 12776
rect 31216 12764 31244 12804
rect 31573 12801 31585 12835
rect 31619 12801 31631 12835
rect 31573 12795 31631 12801
rect 31757 12835 31815 12841
rect 31757 12801 31769 12835
rect 31803 12801 31815 12835
rect 31757 12795 31815 12801
rect 31772 12764 31800 12795
rect 32306 12792 32312 12844
rect 32364 12792 32370 12844
rect 32858 12792 32864 12844
rect 32916 12792 32922 12844
rect 33137 12835 33195 12841
rect 33137 12801 33149 12835
rect 33183 12832 33195 12835
rect 33318 12832 33324 12844
rect 33183 12804 33324 12832
rect 33183 12801 33195 12804
rect 33137 12795 33195 12801
rect 33318 12792 33324 12804
rect 33376 12792 33382 12844
rect 33502 12792 33508 12844
rect 33560 12792 33566 12844
rect 33686 12792 33692 12844
rect 33744 12792 33750 12844
rect 34790 12792 34796 12844
rect 34848 12832 34854 12844
rect 35820 12841 35848 12872
rect 34977 12835 35035 12841
rect 34977 12832 34989 12835
rect 34848 12804 34989 12832
rect 34848 12792 34854 12804
rect 34977 12801 34989 12804
rect 35023 12801 35035 12835
rect 34977 12795 35035 12801
rect 35805 12835 35863 12841
rect 35805 12801 35817 12835
rect 35851 12801 35863 12835
rect 35805 12795 35863 12801
rect 35989 12835 36047 12841
rect 35989 12801 36001 12835
rect 36035 12801 36047 12835
rect 35989 12795 36047 12801
rect 33229 12767 33287 12773
rect 33229 12764 33241 12767
rect 31216 12736 31800 12764
rect 33152 12736 33241 12764
rect 33152 12708 33180 12736
rect 33229 12733 33241 12736
rect 33275 12733 33287 12767
rect 33229 12727 33287 12733
rect 34514 12724 34520 12776
rect 34572 12764 34578 12776
rect 35069 12767 35127 12773
rect 35069 12764 35081 12767
rect 34572 12736 35081 12764
rect 34572 12724 34578 12736
rect 35069 12733 35081 12736
rect 35115 12733 35127 12767
rect 35069 12727 35127 12733
rect 35158 12724 35164 12776
rect 35216 12724 35222 12776
rect 35526 12724 35532 12776
rect 35584 12764 35590 12776
rect 36004 12764 36032 12795
rect 36354 12792 36360 12844
rect 36412 12832 36418 12844
rect 36449 12835 36507 12841
rect 36449 12832 36461 12835
rect 36412 12804 36461 12832
rect 36412 12792 36418 12804
rect 36449 12801 36461 12804
rect 36495 12801 36507 12835
rect 36449 12795 36507 12801
rect 36630 12792 36636 12844
rect 36688 12792 36694 12844
rect 36906 12764 36912 12776
rect 35584 12736 36912 12764
rect 35584 12724 35590 12736
rect 36906 12724 36912 12736
rect 36964 12724 36970 12776
rect 33134 12656 33140 12708
rect 33192 12656 33198 12708
rect 27948 12600 30880 12628
rect 27948 12588 27954 12600
rect 34606 12588 34612 12640
rect 34664 12588 34670 12640
rect 38286 12588 38292 12640
rect 38344 12588 38350 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 20346 12384 20352 12436
rect 20404 12424 20410 12436
rect 20404 12396 23051 12424
rect 20404 12384 20410 12396
rect 20809 12359 20867 12365
rect 20809 12325 20821 12359
rect 20855 12356 20867 12359
rect 22278 12356 22284 12368
rect 20855 12328 21680 12356
rect 20855 12325 20867 12328
rect 20809 12319 20867 12325
rect 19426 12248 19432 12300
rect 19484 12248 19490 12300
rect 21652 12161 21680 12328
rect 21836 12328 22284 12356
rect 21836 12297 21864 12328
rect 22278 12316 22284 12328
rect 22336 12316 22342 12368
rect 22557 12359 22615 12365
rect 22557 12325 22569 12359
rect 22603 12356 22615 12359
rect 23023 12356 23051 12396
rect 23106 12384 23112 12436
rect 23164 12424 23170 12436
rect 23845 12427 23903 12433
rect 23845 12424 23857 12427
rect 23164 12396 23857 12424
rect 23164 12384 23170 12396
rect 23845 12393 23857 12396
rect 23891 12424 23903 12427
rect 24578 12424 24584 12436
rect 23891 12396 24584 12424
rect 23891 12393 23903 12396
rect 23845 12387 23903 12393
rect 24578 12384 24584 12396
rect 24636 12384 24642 12436
rect 26602 12424 26608 12436
rect 26160 12396 26608 12424
rect 24029 12359 24087 12365
rect 24029 12356 24041 12359
rect 22603 12328 22968 12356
rect 23023 12328 24041 12356
rect 22603 12325 22615 12328
rect 22557 12319 22615 12325
rect 21821 12291 21879 12297
rect 21821 12257 21833 12291
rect 21867 12257 21879 12291
rect 21821 12251 21879 12257
rect 22002 12180 22008 12232
rect 22060 12220 22066 12232
rect 22833 12223 22891 12229
rect 22833 12220 22845 12223
rect 22060 12192 22845 12220
rect 22060 12180 22066 12192
rect 22833 12189 22845 12192
rect 22879 12189 22891 12223
rect 22940 12220 22968 12328
rect 24029 12325 24041 12328
rect 24075 12325 24087 12359
rect 24029 12319 24087 12325
rect 23014 12248 23020 12300
rect 23072 12288 23078 12300
rect 23109 12291 23167 12297
rect 23109 12288 23121 12291
rect 23072 12260 23121 12288
rect 23072 12248 23078 12260
rect 23109 12257 23121 12260
rect 23155 12257 23167 12291
rect 23109 12251 23167 12257
rect 23842 12248 23848 12300
rect 23900 12288 23906 12300
rect 25593 12291 25651 12297
rect 25593 12288 25605 12291
rect 23900 12260 25605 12288
rect 23900 12248 23906 12260
rect 25593 12257 25605 12260
rect 25639 12288 25651 12291
rect 26160 12288 26188 12396
rect 26602 12384 26608 12396
rect 26660 12384 26666 12436
rect 28537 12427 28595 12433
rect 28537 12393 28549 12427
rect 28583 12424 28595 12427
rect 32306 12424 32312 12436
rect 28583 12396 32312 12424
rect 28583 12393 28595 12396
rect 28537 12387 28595 12393
rect 32306 12384 32312 12396
rect 32364 12384 32370 12436
rect 34790 12384 34796 12436
rect 34848 12424 34854 12436
rect 36265 12427 36323 12433
rect 36265 12424 36277 12427
rect 34848 12396 36277 12424
rect 34848 12384 34854 12396
rect 36265 12393 36277 12396
rect 36311 12393 36323 12427
rect 36265 12387 36323 12393
rect 26970 12356 26976 12368
rect 25639 12260 26188 12288
rect 26252 12328 26976 12356
rect 25639 12257 25651 12260
rect 25593 12251 25651 12257
rect 26252 12220 26280 12328
rect 26970 12316 26976 12328
rect 27028 12316 27034 12368
rect 28994 12356 29000 12368
rect 28920 12328 29000 12356
rect 26326 12248 26332 12300
rect 26384 12288 26390 12300
rect 27341 12291 27399 12297
rect 27341 12288 27353 12291
rect 26384 12260 27353 12288
rect 26384 12248 26390 12260
rect 27341 12257 27353 12260
rect 27387 12257 27399 12291
rect 27341 12251 27399 12257
rect 28626 12248 28632 12300
rect 28684 12288 28690 12300
rect 28920 12288 28948 12328
rect 28994 12316 29000 12328
rect 29052 12316 29058 12368
rect 30561 12359 30619 12365
rect 30561 12325 30573 12359
rect 30607 12356 30619 12359
rect 31662 12356 31668 12368
rect 30607 12328 31668 12356
rect 30607 12325 30619 12328
rect 30561 12319 30619 12325
rect 31662 12316 31668 12328
rect 31720 12316 31726 12368
rect 32674 12316 32680 12368
rect 32732 12316 32738 12368
rect 34808 12356 34836 12384
rect 33428 12328 34836 12356
rect 29546 12288 29552 12300
rect 28684 12260 28948 12288
rect 28684 12248 28690 12260
rect 22940 12192 26280 12220
rect 22833 12183 22891 12189
rect 26602 12180 26608 12232
rect 26660 12180 26666 12232
rect 26697 12223 26755 12229
rect 26697 12189 26709 12223
rect 26743 12189 26755 12223
rect 26697 12183 26755 12189
rect 19696 12155 19754 12161
rect 19696 12121 19708 12155
rect 19742 12152 19754 12155
rect 21637 12155 21695 12161
rect 19742 12124 21312 12152
rect 19742 12121 19754 12124
rect 19696 12115 19754 12121
rect 21284 12093 21312 12124
rect 21637 12121 21649 12155
rect 21683 12152 21695 12155
rect 23661 12155 23719 12161
rect 23661 12152 23673 12155
rect 21683 12124 23673 12152
rect 21683 12121 21695 12124
rect 21637 12115 21695 12121
rect 23661 12121 23673 12124
rect 23707 12121 23719 12155
rect 23661 12115 23719 12121
rect 23842 12112 23848 12164
rect 23900 12161 23906 12164
rect 23900 12155 23935 12161
rect 23923 12152 23935 12155
rect 25038 12152 25044 12164
rect 23923 12124 25044 12152
rect 23923 12121 23935 12124
rect 23900 12115 23935 12121
rect 23900 12112 23906 12115
rect 25038 12112 25044 12124
rect 25096 12112 25102 12164
rect 25409 12155 25467 12161
rect 25409 12121 25421 12155
rect 25455 12152 25467 12155
rect 26418 12152 26424 12164
rect 25455 12124 26424 12152
rect 25455 12121 25467 12124
rect 25409 12115 25467 12121
rect 26418 12112 26424 12124
rect 26476 12112 26482 12164
rect 26712 12152 26740 12183
rect 26878 12180 26884 12232
rect 26936 12180 26942 12232
rect 26970 12180 26976 12232
rect 27028 12220 27034 12232
rect 28534 12220 28540 12232
rect 27028 12192 28540 12220
rect 27028 12180 27034 12192
rect 28534 12180 28540 12192
rect 28592 12180 28598 12232
rect 28920 12229 28948 12260
rect 29012 12260 29552 12288
rect 29012 12232 29040 12260
rect 29546 12248 29552 12260
rect 29604 12248 29610 12300
rect 30101 12291 30159 12297
rect 30101 12257 30113 12291
rect 30147 12288 30159 12291
rect 30147 12260 31248 12288
rect 30147 12257 30159 12260
rect 30101 12251 30159 12257
rect 28813 12223 28871 12229
rect 28813 12189 28825 12223
rect 28859 12189 28871 12223
rect 28813 12183 28871 12189
rect 28905 12223 28963 12229
rect 28905 12189 28917 12223
rect 28951 12189 28963 12223
rect 28905 12183 28963 12189
rect 27246 12152 27252 12164
rect 26712 12124 27252 12152
rect 27246 12112 27252 12124
rect 27304 12112 27310 12164
rect 28828 12152 28856 12183
rect 28994 12180 29000 12232
rect 29052 12180 29058 12232
rect 29178 12180 29184 12232
rect 29236 12180 29242 12232
rect 29914 12180 29920 12232
rect 29972 12180 29978 12232
rect 30650 12180 30656 12232
rect 30708 12220 30714 12232
rect 30837 12223 30895 12229
rect 30837 12220 30849 12223
rect 30708 12192 30849 12220
rect 30708 12180 30714 12192
rect 30837 12189 30849 12192
rect 30883 12189 30895 12223
rect 30837 12183 30895 12189
rect 30926 12180 30932 12232
rect 30984 12180 30990 12232
rect 31018 12180 31024 12232
rect 31076 12180 31082 12232
rect 31220 12229 31248 12260
rect 31754 12248 31760 12300
rect 31812 12288 31818 12300
rect 32950 12288 32956 12300
rect 31812 12260 32956 12288
rect 31812 12248 31818 12260
rect 32950 12248 32956 12260
rect 33008 12248 33014 12300
rect 33428 12297 33456 12328
rect 33413 12291 33471 12297
rect 33413 12257 33425 12291
rect 33459 12257 33471 12291
rect 33413 12251 33471 12257
rect 33502 12248 33508 12300
rect 33560 12288 33566 12300
rect 33597 12291 33655 12297
rect 33597 12288 33609 12291
rect 33560 12260 33609 12288
rect 33560 12248 33566 12260
rect 33597 12257 33609 12260
rect 33643 12257 33655 12291
rect 33597 12251 33655 12257
rect 34606 12248 34612 12300
rect 34664 12288 34670 12300
rect 34664 12260 35020 12288
rect 34664 12248 34670 12260
rect 31205 12223 31263 12229
rect 31205 12189 31217 12223
rect 31251 12189 31263 12223
rect 31665 12223 31723 12229
rect 31665 12220 31677 12223
rect 31205 12183 31263 12189
rect 31312 12192 31677 12220
rect 29638 12152 29644 12164
rect 28828 12124 29644 12152
rect 29638 12112 29644 12124
rect 29696 12112 29702 12164
rect 29730 12112 29736 12164
rect 29788 12112 29794 12164
rect 30466 12112 30472 12164
rect 30524 12152 30530 12164
rect 30944 12152 30972 12180
rect 30524 12124 30972 12152
rect 30524 12112 30530 12124
rect 21269 12087 21327 12093
rect 21269 12053 21281 12087
rect 21315 12053 21327 12087
rect 21269 12047 21327 12053
rect 21726 12044 21732 12096
rect 21784 12044 21790 12096
rect 23014 12044 23020 12096
rect 23072 12044 23078 12096
rect 24946 12044 24952 12096
rect 25004 12044 25010 12096
rect 25314 12044 25320 12096
rect 25372 12044 25378 12096
rect 25774 12044 25780 12096
rect 25832 12084 25838 12096
rect 31312 12084 31340 12192
rect 31665 12189 31677 12192
rect 31711 12189 31723 12223
rect 31665 12183 31723 12189
rect 31849 12223 31907 12229
rect 31849 12189 31861 12223
rect 31895 12220 31907 12223
rect 31938 12220 31944 12232
rect 31895 12192 31944 12220
rect 31895 12189 31907 12192
rect 31849 12183 31907 12189
rect 31938 12180 31944 12192
rect 31996 12180 32002 12232
rect 32401 12223 32459 12229
rect 32401 12189 32413 12223
rect 32447 12189 32459 12223
rect 32401 12183 32459 12189
rect 31386 12112 31392 12164
rect 31444 12152 31450 12164
rect 32416 12152 32444 12183
rect 33318 12180 33324 12232
rect 33376 12180 33382 12232
rect 33873 12223 33931 12229
rect 33873 12189 33885 12223
rect 33919 12220 33931 12223
rect 34790 12220 34796 12232
rect 33919 12192 34796 12220
rect 33919 12189 33931 12192
rect 33873 12183 33931 12189
rect 34790 12180 34796 12192
rect 34848 12180 34854 12232
rect 34885 12223 34943 12229
rect 34885 12189 34897 12223
rect 34931 12189 34943 12223
rect 34992 12220 35020 12260
rect 35141 12223 35199 12229
rect 35141 12220 35153 12223
rect 34992 12192 35153 12220
rect 34885 12183 34943 12189
rect 35141 12189 35153 12192
rect 35187 12189 35199 12223
rect 35141 12183 35199 12189
rect 31444 12124 32444 12152
rect 31444 12112 31450 12124
rect 33042 12112 33048 12164
rect 33100 12152 33106 12164
rect 34900 12152 34928 12183
rect 33100 12124 34928 12152
rect 33100 12112 33106 12124
rect 25832 12056 31340 12084
rect 25832 12044 25838 12056
rect 31754 12044 31760 12096
rect 31812 12044 31818 12096
rect 32306 12044 32312 12096
rect 32364 12084 32370 12096
rect 34514 12084 34520 12096
rect 32364 12056 34520 12084
rect 32364 12044 32370 12056
rect 34514 12044 34520 12056
rect 34572 12044 34578 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 20898 11840 20904 11892
rect 20956 11880 20962 11892
rect 20993 11883 21051 11889
rect 20993 11880 21005 11883
rect 20956 11852 21005 11880
rect 20956 11840 20962 11852
rect 20993 11849 21005 11852
rect 21039 11849 21051 11883
rect 20993 11843 21051 11849
rect 21085 11883 21143 11889
rect 21085 11849 21097 11883
rect 21131 11880 21143 11883
rect 21726 11880 21732 11892
rect 21131 11852 21732 11880
rect 21131 11849 21143 11852
rect 21085 11843 21143 11849
rect 21726 11840 21732 11852
rect 21784 11880 21790 11892
rect 21784 11852 22508 11880
rect 21784 11840 21790 11852
rect 22480 11821 22508 11852
rect 22646 11840 22652 11892
rect 22704 11880 22710 11892
rect 24302 11880 24308 11892
rect 22704 11852 24308 11880
rect 22704 11840 22710 11852
rect 24302 11840 24308 11852
rect 24360 11840 24366 11892
rect 25314 11840 25320 11892
rect 25372 11880 25378 11892
rect 25685 11883 25743 11889
rect 25685 11880 25697 11883
rect 25372 11852 25697 11880
rect 25372 11840 25378 11852
rect 25685 11849 25697 11852
rect 25731 11880 25743 11883
rect 25731 11852 26280 11880
rect 25731 11849 25743 11852
rect 25685 11843 25743 11849
rect 22465 11815 22523 11821
rect 22465 11781 22477 11815
rect 22511 11812 22523 11815
rect 23750 11812 23756 11824
rect 22511 11784 23756 11812
rect 22511 11781 22523 11784
rect 22465 11775 22523 11781
rect 23750 11772 23756 11784
rect 23808 11772 23814 11824
rect 24572 11815 24630 11821
rect 24572 11781 24584 11815
rect 24618 11812 24630 11815
rect 24946 11812 24952 11824
rect 24618 11784 24952 11812
rect 24618 11781 24630 11784
rect 24572 11775 24630 11781
rect 24946 11772 24952 11784
rect 25004 11772 25010 11824
rect 26050 11772 26056 11824
rect 26108 11812 26114 11824
rect 26145 11815 26203 11821
rect 26145 11812 26157 11815
rect 26108 11784 26157 11812
rect 26108 11772 26114 11784
rect 26145 11781 26157 11784
rect 26191 11781 26203 11815
rect 26252 11812 26280 11852
rect 26510 11840 26516 11892
rect 26568 11840 26574 11892
rect 26602 11840 26608 11892
rect 26660 11880 26666 11892
rect 27157 11883 27215 11889
rect 27157 11880 27169 11883
rect 26660 11852 27169 11880
rect 26660 11840 26666 11852
rect 27157 11849 27169 11852
rect 27203 11849 27215 11883
rect 27157 11843 27215 11849
rect 27246 11840 27252 11892
rect 27304 11880 27310 11892
rect 28353 11883 28411 11889
rect 28353 11880 28365 11883
rect 27304 11852 28365 11880
rect 27304 11840 27310 11852
rect 28353 11849 28365 11852
rect 28399 11849 28411 11883
rect 28353 11843 28411 11849
rect 28534 11840 28540 11892
rect 28592 11880 28598 11892
rect 28592 11852 28948 11880
rect 28592 11840 28598 11852
rect 27525 11815 27583 11821
rect 27525 11812 27537 11815
rect 26252 11784 27537 11812
rect 26145 11775 26203 11781
rect 27525 11781 27537 11784
rect 27571 11781 27583 11815
rect 28626 11812 28632 11824
rect 27525 11775 27583 11781
rect 27632 11784 28632 11812
rect 22370 11704 22376 11756
rect 22428 11704 22434 11756
rect 23198 11704 23204 11756
rect 23256 11704 23262 11756
rect 24854 11744 24860 11756
rect 23400 11716 24860 11744
rect 21269 11679 21327 11685
rect 21269 11645 21281 11679
rect 21315 11676 21327 11679
rect 22649 11679 22707 11685
rect 21315 11648 22140 11676
rect 21315 11645 21327 11648
rect 21269 11639 21327 11645
rect 20622 11500 20628 11552
rect 20680 11500 20686 11552
rect 22002 11500 22008 11552
rect 22060 11500 22066 11552
rect 22112 11540 22140 11648
rect 22649 11645 22661 11679
rect 22695 11676 22707 11679
rect 22738 11676 22744 11688
rect 22695 11648 22744 11676
rect 22695 11645 22707 11648
rect 22649 11639 22707 11645
rect 22738 11636 22744 11648
rect 22796 11636 22802 11688
rect 23400 11685 23428 11716
rect 24854 11704 24860 11716
rect 24912 11744 24918 11756
rect 24912 11716 25360 11744
rect 24912 11704 24918 11716
rect 23385 11679 23443 11685
rect 23385 11645 23397 11679
rect 23431 11645 23443 11679
rect 23385 11639 23443 11645
rect 22186 11568 22192 11620
rect 22244 11608 22250 11620
rect 23400 11608 23428 11639
rect 24302 11636 24308 11688
rect 24360 11636 24366 11688
rect 25332 11676 25360 11716
rect 25682 11704 25688 11756
rect 25740 11744 25746 11756
rect 26329 11747 26387 11753
rect 26329 11744 26341 11747
rect 25740 11716 26341 11744
rect 25740 11704 25746 11716
rect 26329 11713 26341 11716
rect 26375 11713 26387 11747
rect 27632 11744 27660 11784
rect 26329 11707 26387 11713
rect 26712 11716 27660 11744
rect 26712 11676 26740 11716
rect 25332 11648 26740 11676
rect 26786 11636 26792 11688
rect 26844 11676 26850 11688
rect 27816 11685 27844 11784
rect 28626 11772 28632 11784
rect 28684 11812 28690 11824
rect 28920 11812 28948 11852
rect 30006 11840 30012 11892
rect 30064 11880 30070 11892
rect 31754 11880 31760 11892
rect 30064 11852 31760 11880
rect 30064 11840 30070 11852
rect 31754 11840 31760 11852
rect 31812 11840 31818 11892
rect 31846 11840 31852 11892
rect 31904 11880 31910 11892
rect 33689 11883 33747 11889
rect 33689 11880 33701 11883
rect 31904 11852 33701 11880
rect 31904 11840 31910 11852
rect 33689 11849 33701 11852
rect 33735 11849 33747 11883
rect 33689 11843 33747 11849
rect 34790 11840 34796 11892
rect 34848 11880 34854 11892
rect 35342 11880 35348 11892
rect 34848 11852 35348 11880
rect 34848 11840 34854 11852
rect 35342 11840 35348 11852
rect 35400 11880 35406 11892
rect 35621 11883 35679 11889
rect 35621 11880 35633 11883
rect 35400 11852 35633 11880
rect 35400 11840 35406 11852
rect 35621 11849 35633 11852
rect 35667 11849 35679 11883
rect 35621 11843 35679 11849
rect 32490 11812 32496 11824
rect 28684 11784 28856 11812
rect 28920 11784 32496 11812
rect 28684 11772 28690 11784
rect 28718 11704 28724 11756
rect 28776 11704 28782 11756
rect 28828 11744 28856 11784
rect 29917 11747 29975 11753
rect 28828 11716 28948 11744
rect 28920 11685 28948 11716
rect 29917 11713 29929 11747
rect 29963 11744 29975 11747
rect 30374 11744 30380 11756
rect 29963 11716 30380 11744
rect 29963 11713 29975 11716
rect 29917 11707 29975 11713
rect 30374 11704 30380 11716
rect 30432 11704 30438 11756
rect 31018 11704 31024 11756
rect 31076 11744 31082 11756
rect 31113 11747 31171 11753
rect 31113 11744 31125 11747
rect 31076 11716 31125 11744
rect 31076 11704 31082 11716
rect 31113 11713 31125 11716
rect 31159 11713 31171 11747
rect 32306 11744 32312 11756
rect 31113 11707 31171 11713
rect 31220 11716 32312 11744
rect 27617 11679 27675 11685
rect 27617 11676 27629 11679
rect 26844 11648 27629 11676
rect 26844 11636 26850 11648
rect 27617 11645 27629 11648
rect 27663 11645 27675 11679
rect 27617 11639 27675 11645
rect 27801 11679 27859 11685
rect 27801 11645 27813 11679
rect 27847 11645 27859 11679
rect 27801 11639 27859 11645
rect 28813 11679 28871 11685
rect 28813 11645 28825 11679
rect 28859 11645 28871 11679
rect 28813 11639 28871 11645
rect 28905 11679 28963 11685
rect 28905 11645 28917 11679
rect 28951 11645 28963 11679
rect 30009 11679 30067 11685
rect 30009 11676 30021 11679
rect 28905 11639 28963 11645
rect 29472 11648 30021 11676
rect 22244 11580 23428 11608
rect 22244 11568 22250 11580
rect 27522 11568 27528 11620
rect 27580 11608 27586 11620
rect 28828 11608 28856 11639
rect 27580 11580 28856 11608
rect 27580 11568 27586 11580
rect 27062 11540 27068 11552
rect 22112 11512 27068 11540
rect 27062 11500 27068 11512
rect 27120 11500 27126 11552
rect 28166 11500 28172 11552
rect 28224 11540 28230 11552
rect 29472 11540 29500 11648
rect 30009 11645 30021 11648
rect 30055 11645 30067 11679
rect 30009 11639 30067 11645
rect 30024 11608 30052 11639
rect 30190 11636 30196 11688
rect 30248 11636 30254 11688
rect 31220 11685 31248 11716
rect 32306 11704 32312 11716
rect 32364 11704 32370 11756
rect 31205 11679 31263 11685
rect 31205 11645 31217 11679
rect 31251 11645 31263 11679
rect 31205 11639 31263 11645
rect 31220 11608 31248 11639
rect 31294 11636 31300 11688
rect 31352 11636 31358 11688
rect 30024 11580 31248 11608
rect 32416 11608 32444 11784
rect 32490 11772 32496 11784
rect 32548 11772 32554 11824
rect 32769 11747 32827 11753
rect 32769 11713 32781 11747
rect 32815 11744 32827 11747
rect 33134 11744 33140 11756
rect 32815 11716 33140 11744
rect 32815 11713 32827 11716
rect 32769 11707 32827 11713
rect 33134 11704 33140 11716
rect 33192 11704 33198 11756
rect 33594 11704 33600 11756
rect 33652 11704 33658 11756
rect 33778 11704 33784 11756
rect 33836 11704 33842 11756
rect 34508 11747 34566 11753
rect 34508 11713 34520 11747
rect 34554 11744 34566 11747
rect 34790 11744 34796 11756
rect 34554 11716 34796 11744
rect 34554 11713 34566 11716
rect 34508 11707 34566 11713
rect 34790 11704 34796 11716
rect 34848 11704 34854 11756
rect 32858 11636 32864 11688
rect 32916 11636 32922 11688
rect 32953 11679 33011 11685
rect 32953 11645 32965 11679
rect 32999 11645 33011 11679
rect 32953 11639 33011 11645
rect 34241 11679 34299 11685
rect 34241 11645 34253 11679
rect 34287 11645 34299 11679
rect 34241 11639 34299 11645
rect 32968 11608 32996 11639
rect 32416 11580 32996 11608
rect 28224 11512 29500 11540
rect 28224 11500 28230 11512
rect 29546 11500 29552 11552
rect 29604 11500 29610 11552
rect 30650 11500 30656 11552
rect 30708 11540 30714 11552
rect 30745 11543 30803 11549
rect 30745 11540 30757 11543
rect 30708 11512 30757 11540
rect 30708 11500 30714 11512
rect 30745 11509 30757 11512
rect 30791 11509 30803 11543
rect 30745 11503 30803 11509
rect 30834 11500 30840 11552
rect 30892 11540 30898 11552
rect 31386 11540 31392 11552
rect 30892 11512 31392 11540
rect 30892 11500 30898 11512
rect 31386 11500 31392 11512
rect 31444 11500 31450 11552
rect 32398 11500 32404 11552
rect 32456 11500 32462 11552
rect 32490 11500 32496 11552
rect 32548 11540 32554 11552
rect 33042 11540 33048 11552
rect 32548 11512 33048 11540
rect 32548 11500 32554 11512
rect 33042 11500 33048 11512
rect 33100 11540 33106 11552
rect 34256 11540 34284 11639
rect 33100 11512 34284 11540
rect 33100 11500 33106 11512
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 22370 11296 22376 11348
rect 22428 11296 22434 11348
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 25961 11339 26019 11345
rect 23256 11308 25912 11336
rect 23256 11296 23262 11308
rect 25884 11268 25912 11308
rect 25961 11305 25973 11339
rect 26007 11336 26019 11339
rect 26786 11336 26792 11348
rect 26007 11308 26792 11336
rect 26007 11305 26019 11308
rect 25961 11299 26019 11305
rect 26786 11296 26792 11308
rect 26844 11296 26850 11348
rect 27062 11296 27068 11348
rect 27120 11336 27126 11348
rect 29181 11339 29239 11345
rect 27120 11308 28764 11336
rect 27120 11296 27126 11308
rect 28736 11268 28764 11308
rect 29181 11305 29193 11339
rect 29227 11336 29239 11339
rect 30374 11336 30380 11348
rect 29227 11308 30380 11336
rect 29227 11305 29239 11308
rect 29181 11299 29239 11305
rect 30374 11296 30380 11308
rect 30432 11296 30438 11348
rect 31018 11296 31024 11348
rect 31076 11336 31082 11348
rect 31757 11339 31815 11345
rect 31757 11336 31769 11339
rect 31076 11308 31769 11336
rect 31076 11296 31082 11308
rect 31757 11305 31769 11308
rect 31803 11305 31815 11339
rect 32490 11336 32496 11348
rect 31757 11299 31815 11305
rect 32232 11308 32496 11336
rect 25884 11240 27752 11268
rect 28736 11240 29684 11268
rect 19426 11160 19432 11212
rect 19484 11200 19490 11212
rect 20993 11203 21051 11209
rect 20993 11200 21005 11203
rect 19484 11172 21005 11200
rect 19484 11160 19490 11172
rect 20993 11169 21005 11172
rect 21039 11169 21051 11203
rect 20993 11163 21051 11169
rect 23750 11160 23756 11212
rect 23808 11160 23814 11212
rect 23937 11203 23995 11209
rect 23937 11169 23949 11203
rect 23983 11200 23995 11203
rect 24210 11200 24216 11212
rect 23983 11172 24216 11200
rect 23983 11169 23995 11172
rect 23937 11163 23995 11169
rect 24210 11160 24216 11172
rect 24268 11160 24274 11212
rect 24302 11160 24308 11212
rect 24360 11200 24366 11212
rect 24581 11203 24639 11209
rect 24581 11200 24593 11203
rect 24360 11172 24593 11200
rect 24360 11160 24366 11172
rect 24581 11169 24593 11172
rect 24627 11169 24639 11203
rect 24581 11163 24639 11169
rect 26418 11160 26424 11212
rect 26476 11200 26482 11212
rect 26881 11203 26939 11209
rect 26881 11200 26893 11203
rect 26476 11172 26893 11200
rect 26476 11160 26482 11172
rect 26881 11169 26893 11172
rect 26927 11169 26939 11203
rect 26881 11163 26939 11169
rect 21260 11135 21318 11141
rect 21260 11101 21272 11135
rect 21306 11132 21318 11135
rect 22002 11132 22008 11144
rect 21306 11104 22008 11132
rect 21306 11101 21318 11104
rect 21260 11095 21318 11101
rect 22002 11092 22008 11104
rect 22060 11092 22066 11144
rect 24848 11135 24906 11141
rect 24848 11101 24860 11135
rect 24894 11132 24906 11135
rect 24894 11104 26372 11132
rect 24894 11101 24906 11104
rect 24848 11095 24906 11101
rect 23290 10956 23296 11008
rect 23348 10956 23354 11008
rect 23474 10956 23480 11008
rect 23532 10996 23538 11008
rect 23661 10999 23719 11005
rect 23661 10996 23673 10999
rect 23532 10968 23673 10996
rect 23532 10956 23538 10968
rect 23661 10965 23673 10968
rect 23707 10965 23719 10999
rect 26344 10996 26372 11104
rect 26786 11092 26792 11144
rect 26844 11092 26850 11144
rect 26896 11132 26924 11163
rect 27062 11160 27068 11212
rect 27120 11160 27126 11212
rect 27154 11132 27160 11144
rect 26896 11104 27160 11132
rect 27154 11092 27160 11104
rect 27212 11092 27218 11144
rect 27724 11064 27752 11240
rect 27798 11160 27804 11212
rect 27856 11160 27862 11212
rect 28068 11135 28126 11141
rect 28068 11101 28080 11135
rect 28114 11132 28126 11135
rect 29546 11132 29552 11144
rect 28114 11104 29552 11132
rect 28114 11101 28126 11104
rect 28068 11095 28126 11101
rect 29546 11092 29552 11104
rect 29604 11092 29610 11144
rect 29656 11132 29684 11240
rect 29822 11160 29828 11212
rect 29880 11200 29886 11212
rect 30377 11203 30435 11209
rect 30377 11200 30389 11203
rect 29880 11172 30389 11200
rect 29880 11160 29886 11172
rect 30377 11169 30389 11172
rect 30423 11169 30435 11203
rect 30377 11163 30435 11169
rect 32232 11141 32260 11308
rect 32490 11296 32496 11308
rect 32548 11296 32554 11348
rect 33134 11296 33140 11348
rect 33192 11336 33198 11348
rect 33597 11339 33655 11345
rect 33597 11336 33609 11339
rect 33192 11308 33609 11336
rect 33192 11296 33198 11308
rect 33597 11305 33609 11308
rect 33643 11305 33655 11339
rect 33597 11299 33655 11305
rect 34790 11296 34796 11348
rect 34848 11336 34854 11348
rect 34885 11339 34943 11345
rect 34885 11336 34897 11339
rect 34848 11308 34897 11336
rect 34848 11296 34854 11308
rect 34885 11305 34897 11308
rect 34931 11305 34943 11339
rect 34885 11299 34943 11305
rect 35434 11200 35440 11212
rect 33520 11172 35440 11200
rect 32217 11135 32275 11141
rect 29656 11104 31754 11132
rect 30466 11064 30472 11076
rect 27724 11036 30472 11064
rect 30466 11024 30472 11036
rect 30524 11024 30530 11076
rect 30650 11073 30656 11076
rect 30633 11067 30656 11073
rect 30633 11033 30645 11067
rect 30633 11027 30656 11033
rect 30650 11024 30656 11027
rect 30708 11024 30714 11076
rect 26421 10999 26479 11005
rect 26421 10996 26433 10999
rect 26344 10968 26433 10996
rect 23661 10959 23719 10965
rect 26421 10965 26433 10968
rect 26467 10965 26479 10999
rect 31726 10996 31754 11104
rect 32217 11101 32229 11135
rect 32263 11101 32275 11135
rect 32217 11095 32275 11101
rect 32484 11135 32542 11141
rect 32484 11101 32496 11135
rect 32530 11101 32542 11135
rect 32484 11095 32542 11101
rect 32398 11024 32404 11076
rect 32456 11064 32462 11076
rect 32508 11064 32536 11095
rect 32456 11036 32536 11064
rect 32456 11024 32462 11036
rect 32950 11024 32956 11076
rect 33008 11064 33014 11076
rect 33520 11064 33548 11172
rect 35434 11160 35440 11172
rect 35492 11160 35498 11212
rect 35253 11135 35311 11141
rect 35253 11101 35265 11135
rect 35299 11132 35311 11135
rect 35342 11132 35348 11144
rect 35299 11104 35348 11132
rect 35299 11101 35311 11104
rect 35253 11095 35311 11101
rect 35342 11092 35348 11104
rect 35400 11092 35406 11144
rect 37829 11135 37887 11141
rect 37829 11101 37841 11135
rect 37875 11132 37887 11135
rect 39206 11132 39212 11144
rect 37875 11104 39212 11132
rect 37875 11101 37887 11104
rect 37829 11095 37887 11101
rect 39206 11092 39212 11104
rect 39264 11092 39270 11144
rect 33008 11036 33548 11064
rect 33008 11024 33014 11036
rect 34514 11024 34520 11076
rect 34572 11064 34578 11076
rect 34572 11036 35388 11064
rect 34572 11024 34578 11036
rect 32968 10996 32996 11024
rect 35360 11005 35388 11036
rect 38102 11024 38108 11076
rect 38160 11024 38166 11076
rect 31726 10968 32996 10996
rect 35345 10999 35403 11005
rect 26421 10959 26479 10965
rect 35345 10965 35357 10999
rect 35391 10965 35403 10999
rect 35345 10959 35403 10965
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 20898 10752 20904 10804
rect 20956 10792 20962 10804
rect 21085 10795 21143 10801
rect 21085 10792 21097 10795
rect 20956 10764 21097 10792
rect 20956 10752 20962 10764
rect 21085 10761 21097 10764
rect 21131 10761 21143 10795
rect 21085 10755 21143 10761
rect 22281 10795 22339 10801
rect 22281 10761 22293 10795
rect 22327 10792 22339 10795
rect 23014 10792 23020 10804
rect 22327 10764 23020 10792
rect 22327 10761 22339 10764
rect 22281 10755 22339 10761
rect 23014 10752 23020 10764
rect 23072 10752 23078 10804
rect 26605 10795 26663 10801
rect 26605 10761 26617 10795
rect 26651 10792 26663 10795
rect 28718 10792 28724 10804
rect 26651 10764 28724 10792
rect 26651 10761 26663 10764
rect 26605 10755 26663 10761
rect 28718 10752 28724 10764
rect 28776 10752 28782 10804
rect 29638 10752 29644 10804
rect 29696 10792 29702 10804
rect 30282 10792 30288 10804
rect 29696 10764 30288 10792
rect 29696 10752 29702 10764
rect 30282 10752 30288 10764
rect 30340 10792 30346 10804
rect 31297 10795 31355 10801
rect 31297 10792 31309 10795
rect 30340 10764 31309 10792
rect 30340 10752 30346 10764
rect 31297 10761 31309 10764
rect 31343 10761 31355 10795
rect 31297 10755 31355 10761
rect 33686 10752 33692 10804
rect 33744 10752 33750 10804
rect 19972 10727 20030 10733
rect 19972 10693 19984 10727
rect 20018 10724 20030 10727
rect 20622 10724 20628 10736
rect 20018 10696 20628 10724
rect 20018 10693 20030 10696
rect 19972 10687 20030 10693
rect 20622 10684 20628 10696
rect 20680 10684 20686 10736
rect 25240 10696 27844 10724
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19705 10659 19763 10665
rect 19705 10656 19717 10659
rect 19484 10628 19717 10656
rect 19484 10616 19490 10628
rect 19705 10625 19717 10628
rect 19751 10625 19763 10659
rect 19705 10619 19763 10625
rect 20530 10616 20536 10668
rect 20588 10656 20594 10668
rect 22005 10659 22063 10665
rect 20588 10628 21956 10656
rect 20588 10616 20594 10628
rect 21928 10588 21956 10628
rect 22005 10625 22017 10659
rect 22051 10656 22063 10659
rect 22370 10656 22376 10668
rect 22051 10628 22376 10656
rect 22051 10625 22063 10628
rect 22005 10619 22063 10625
rect 22370 10616 22376 10628
rect 22428 10616 22434 10668
rect 22646 10616 22652 10668
rect 22704 10656 22710 10668
rect 22741 10659 22799 10665
rect 22741 10656 22753 10659
rect 22704 10628 22753 10656
rect 22704 10616 22710 10628
rect 22741 10625 22753 10628
rect 22787 10625 22799 10659
rect 22741 10619 22799 10625
rect 23008 10659 23066 10665
rect 23008 10625 23020 10659
rect 23054 10656 23066 10659
rect 23290 10656 23296 10668
rect 23054 10628 23296 10656
rect 23054 10625 23066 10628
rect 23008 10619 23066 10625
rect 23290 10616 23296 10628
rect 23348 10616 23354 10668
rect 25240 10665 25268 10696
rect 27816 10668 27844 10696
rect 29932 10696 31754 10724
rect 25225 10659 25283 10665
rect 25225 10625 25237 10659
rect 25271 10625 25283 10659
rect 25225 10619 25283 10625
rect 25492 10659 25550 10665
rect 25492 10625 25504 10659
rect 25538 10656 25550 10659
rect 27706 10656 27712 10668
rect 25538 10628 27712 10656
rect 25538 10625 25550 10628
rect 25492 10619 25550 10625
rect 27706 10616 27712 10628
rect 27764 10616 27770 10668
rect 27798 10616 27804 10668
rect 27856 10656 27862 10668
rect 28350 10665 28356 10668
rect 28077 10659 28135 10665
rect 28077 10656 28089 10659
rect 27856 10628 28089 10656
rect 27856 10616 27862 10628
rect 28077 10625 28089 10628
rect 28123 10625 28135 10659
rect 28077 10619 28135 10625
rect 28344 10619 28356 10665
rect 28350 10616 28356 10619
rect 28408 10616 28414 10668
rect 29822 10616 29828 10668
rect 29880 10656 29886 10668
rect 29932 10665 29960 10696
rect 30190 10665 30196 10668
rect 29917 10659 29975 10665
rect 29917 10656 29929 10659
rect 29880 10628 29929 10656
rect 29880 10616 29886 10628
rect 29917 10625 29929 10628
rect 29963 10625 29975 10659
rect 29917 10619 29975 10625
rect 30184 10619 30196 10665
rect 30190 10616 30196 10619
rect 30248 10616 30254 10668
rect 31726 10656 31754 10696
rect 32309 10659 32367 10665
rect 32309 10656 32321 10659
rect 31726 10628 32321 10656
rect 32309 10625 32321 10628
rect 32355 10625 32367 10659
rect 32309 10619 32367 10625
rect 32398 10616 32404 10668
rect 32456 10656 32462 10668
rect 32565 10659 32623 10665
rect 32565 10656 32577 10659
rect 32456 10628 32577 10656
rect 32456 10616 32462 10628
rect 32565 10625 32577 10628
rect 32611 10625 32623 10659
rect 32565 10619 32623 10625
rect 22097 10591 22155 10597
rect 22097 10588 22109 10591
rect 21928 10560 22109 10588
rect 22097 10557 22109 10560
rect 22143 10588 22155 10591
rect 22186 10588 22192 10600
rect 22143 10560 22192 10588
rect 22143 10557 22155 10560
rect 22097 10551 22155 10557
rect 22186 10548 22192 10560
rect 22244 10548 22250 10600
rect 22278 10548 22284 10600
rect 22336 10548 22342 10600
rect 23474 10412 23480 10464
rect 23532 10452 23538 10464
rect 24121 10455 24179 10461
rect 24121 10452 24133 10455
rect 23532 10424 24133 10452
rect 23532 10412 23538 10424
rect 24121 10421 24133 10424
rect 24167 10421 24179 10455
rect 24121 10415 24179 10421
rect 29454 10412 29460 10464
rect 29512 10412 29518 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 22094 10208 22100 10260
rect 22152 10208 22158 10260
rect 22278 10208 22284 10260
rect 22336 10248 22342 10260
rect 23109 10251 23167 10257
rect 23109 10248 23121 10251
rect 22336 10220 23121 10248
rect 22336 10208 22342 10220
rect 23109 10217 23121 10220
rect 23155 10217 23167 10251
rect 23109 10211 23167 10217
rect 27522 10208 27528 10260
rect 27580 10208 27586 10260
rect 27706 10208 27712 10260
rect 27764 10248 27770 10260
rect 27985 10251 28043 10257
rect 27985 10248 27997 10251
rect 27764 10220 27997 10248
rect 27764 10208 27770 10220
rect 27985 10217 27997 10220
rect 28031 10217 28043 10251
rect 27985 10211 28043 10217
rect 30190 10208 30196 10260
rect 30248 10208 30254 10260
rect 30374 10208 30380 10260
rect 30432 10248 30438 10260
rect 30432 10220 31616 10248
rect 30432 10208 30438 10220
rect 30282 10140 30288 10192
rect 30340 10180 30346 10192
rect 30340 10152 30604 10180
rect 30340 10140 30346 10152
rect 22020 10084 23612 10112
rect 22020 10053 22048 10084
rect 22005 10047 22063 10053
rect 22005 10013 22017 10047
rect 22051 10013 22063 10047
rect 22005 10007 22063 10013
rect 22189 10047 22247 10053
rect 22189 10013 22201 10047
rect 22235 10044 22247 10047
rect 23106 10044 23112 10056
rect 22235 10016 23112 10044
rect 22235 10013 22247 10016
rect 22189 10007 22247 10013
rect 23106 10004 23112 10016
rect 23164 10004 23170 10056
rect 23293 10047 23351 10053
rect 23293 10013 23305 10047
rect 23339 10044 23351 10047
rect 23474 10044 23480 10056
rect 23339 10016 23480 10044
rect 23339 10013 23351 10016
rect 23293 10007 23351 10013
rect 23474 10004 23480 10016
rect 23532 10004 23538 10056
rect 23584 10053 23612 10084
rect 27246 10072 27252 10124
rect 27304 10112 27310 10124
rect 28445 10115 28503 10121
rect 28445 10112 28457 10115
rect 27304 10084 28457 10112
rect 27304 10072 27310 10084
rect 28445 10081 28457 10084
rect 28491 10081 28503 10115
rect 28445 10075 28503 10081
rect 28629 10115 28687 10121
rect 28629 10081 28641 10115
rect 28675 10112 28687 10115
rect 30466 10112 30472 10124
rect 28675 10084 30472 10112
rect 28675 10081 28687 10084
rect 28629 10075 28687 10081
rect 30466 10072 30472 10084
rect 30524 10072 30530 10124
rect 23569 10047 23627 10053
rect 23569 10013 23581 10047
rect 23615 10044 23627 10047
rect 23842 10044 23848 10056
rect 23615 10016 23848 10044
rect 23615 10013 23627 10016
rect 23569 10007 23627 10013
rect 23842 10004 23848 10016
rect 23900 10004 23906 10056
rect 26145 10047 26203 10053
rect 26145 10013 26157 10047
rect 26191 10044 26203 10047
rect 27798 10044 27804 10056
rect 26191 10016 27804 10044
rect 26191 10013 26203 10016
rect 26145 10007 26203 10013
rect 27798 10004 27804 10016
rect 27856 10004 27862 10056
rect 28353 10047 28411 10053
rect 28353 10013 28365 10047
rect 28399 10044 28411 10047
rect 28718 10044 28724 10056
rect 28399 10016 28724 10044
rect 28399 10013 28411 10016
rect 28353 10007 28411 10013
rect 28718 10004 28724 10016
rect 28776 10004 28782 10056
rect 30576 10053 30604 10152
rect 30650 10072 30656 10124
rect 30708 10112 30714 10124
rect 30745 10115 30803 10121
rect 30745 10112 30757 10115
rect 30708 10084 30757 10112
rect 30708 10072 30714 10084
rect 30745 10081 30757 10084
rect 30791 10112 30803 10115
rect 31294 10112 31300 10124
rect 30791 10084 31300 10112
rect 30791 10081 30803 10084
rect 30745 10075 30803 10081
rect 31294 10072 31300 10084
rect 31352 10072 31358 10124
rect 31588 10053 31616 10220
rect 32398 10208 32404 10260
rect 32456 10208 32462 10260
rect 32858 10112 32864 10124
rect 31726 10084 32864 10112
rect 30561 10047 30619 10053
rect 30561 10013 30573 10047
rect 30607 10013 30619 10047
rect 30561 10007 30619 10013
rect 31573 10047 31631 10053
rect 31573 10013 31585 10047
rect 31619 10013 31631 10047
rect 31573 10007 31631 10013
rect 23124 9908 23152 10004
rect 26412 9979 26470 9985
rect 26412 9945 26424 9979
rect 26458 9976 26470 9979
rect 27154 9976 27160 9988
rect 26458 9948 27160 9976
rect 26458 9945 26470 9948
rect 26412 9939 26470 9945
rect 27154 9936 27160 9948
rect 27212 9936 27218 9988
rect 31389 9979 31447 9985
rect 31389 9976 31401 9979
rect 30576 9948 31401 9976
rect 23477 9911 23535 9917
rect 23477 9908 23489 9911
rect 23124 9880 23489 9908
rect 23477 9877 23489 9880
rect 23523 9877 23535 9911
rect 23477 9871 23535 9877
rect 29730 9868 29736 9920
rect 29788 9908 29794 9920
rect 30576 9908 30604 9948
rect 31389 9945 31401 9948
rect 31435 9945 31447 9979
rect 31726 9976 31754 10084
rect 32858 10072 32864 10084
rect 32916 10072 32922 10124
rect 32950 10072 32956 10124
rect 33008 10072 33014 10124
rect 32769 10047 32827 10053
rect 32769 10013 32781 10047
rect 32815 10044 32827 10047
rect 33686 10044 33692 10056
rect 32815 10016 33692 10044
rect 32815 10013 32827 10016
rect 32769 10007 32827 10013
rect 33686 10004 33692 10016
rect 33744 10004 33750 10056
rect 34330 10004 34336 10056
rect 34388 10044 34394 10056
rect 37829 10047 37887 10053
rect 37829 10044 37841 10047
rect 34388 10016 37841 10044
rect 34388 10004 34394 10016
rect 37829 10013 37841 10016
rect 37875 10013 37887 10047
rect 37829 10007 37887 10013
rect 31389 9939 31447 9945
rect 31496 9948 31754 9976
rect 29788 9880 30604 9908
rect 29788 9868 29794 9880
rect 30650 9868 30656 9920
rect 30708 9908 30714 9920
rect 31496 9908 31524 9948
rect 38102 9936 38108 9988
rect 38160 9936 38166 9988
rect 30708 9880 31524 9908
rect 30708 9868 30714 9880
rect 31754 9868 31760 9920
rect 31812 9868 31818 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 27154 9664 27160 9716
rect 27212 9664 27218 9716
rect 27522 9664 27528 9716
rect 27580 9664 27586 9716
rect 27617 9707 27675 9713
rect 27617 9673 27629 9707
rect 27663 9673 27675 9707
rect 27617 9667 27675 9673
rect 27246 9596 27252 9648
rect 27304 9636 27310 9648
rect 27632 9636 27660 9667
rect 28350 9664 28356 9716
rect 28408 9704 28414 9716
rect 28537 9707 28595 9713
rect 28537 9704 28549 9707
rect 28408 9676 28549 9704
rect 28408 9664 28414 9676
rect 28537 9673 28549 9676
rect 28583 9673 28595 9707
rect 28537 9667 28595 9673
rect 28810 9664 28816 9716
rect 28868 9704 28874 9716
rect 28997 9707 29055 9713
rect 28997 9704 29009 9707
rect 28868 9676 29009 9704
rect 28868 9664 28874 9676
rect 28997 9673 29009 9676
rect 29043 9704 29055 9707
rect 30650 9704 30656 9716
rect 29043 9676 30656 9704
rect 29043 9673 29055 9676
rect 28997 9667 29055 9673
rect 30650 9664 30656 9676
rect 30708 9664 30714 9716
rect 27304 9608 27660 9636
rect 28905 9639 28963 9645
rect 27304 9596 27310 9608
rect 28905 9605 28917 9639
rect 28951 9636 28963 9639
rect 29454 9636 29460 9648
rect 28951 9608 29460 9636
rect 28951 9605 28963 9608
rect 28905 9599 28963 9605
rect 29454 9596 29460 9608
rect 29512 9636 29518 9648
rect 29917 9639 29975 9645
rect 29917 9636 29929 9639
rect 29512 9608 29929 9636
rect 29512 9596 29518 9608
rect 29917 9605 29929 9608
rect 29963 9605 29975 9639
rect 29917 9599 29975 9605
rect 30745 9639 30803 9645
rect 30745 9605 30757 9639
rect 30791 9636 30803 9639
rect 30834 9636 30840 9648
rect 30791 9608 30840 9636
rect 30791 9605 30803 9608
rect 30745 9599 30803 9605
rect 30834 9596 30840 9608
rect 30892 9596 30898 9648
rect 27430 9528 27436 9580
rect 27488 9568 27494 9580
rect 27488 9540 29132 9568
rect 27488 9528 27494 9540
rect 27724 9509 27752 9540
rect 29104 9509 29132 9540
rect 29730 9528 29736 9580
rect 29788 9528 29794 9580
rect 31018 9528 31024 9580
rect 31076 9528 31082 9580
rect 31113 9571 31171 9577
rect 31113 9537 31125 9571
rect 31159 9537 31171 9571
rect 31113 9531 31171 9537
rect 31205 9571 31263 9577
rect 31205 9537 31217 9571
rect 31251 9537 31263 9571
rect 31205 9531 31263 9537
rect 31389 9571 31447 9577
rect 31389 9537 31401 9571
rect 31435 9568 31447 9571
rect 31754 9568 31760 9580
rect 31435 9540 31760 9568
rect 31435 9537 31447 9540
rect 31389 9531 31447 9537
rect 27709 9503 27767 9509
rect 27709 9469 27721 9503
rect 27755 9469 27767 9503
rect 27709 9463 27767 9469
rect 29089 9503 29147 9509
rect 29089 9469 29101 9503
rect 29135 9469 29147 9503
rect 29089 9463 29147 9469
rect 29178 9460 29184 9512
rect 29236 9500 29242 9512
rect 30101 9503 30159 9509
rect 30101 9500 30113 9503
rect 29236 9472 30113 9500
rect 29236 9460 29242 9472
rect 30101 9469 30113 9472
rect 30147 9469 30159 9503
rect 30101 9463 30159 9469
rect 30742 9460 30748 9512
rect 30800 9500 30806 9512
rect 31128 9500 31156 9531
rect 30800 9472 31156 9500
rect 30800 9460 30806 9472
rect 28994 9324 29000 9376
rect 29052 9364 29058 9376
rect 31220 9364 31248 9531
rect 31754 9528 31760 9540
rect 31812 9528 31818 9580
rect 29052 9336 31248 9364
rect 29052 9324 29058 9336
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 32582 8984 32588 9036
rect 32640 9024 32646 9036
rect 37274 9024 37280 9036
rect 32640 8996 37280 9024
rect 32640 8984 32646 8996
rect 37274 8984 37280 8996
rect 37332 8984 37338 9036
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 37829 8483 37887 8489
rect 37829 8449 37841 8483
rect 37875 8480 37887 8483
rect 38194 8480 38200 8492
rect 37875 8452 38200 8480
rect 37875 8449 37887 8452
rect 37829 8443 37887 8449
rect 38194 8440 38200 8452
rect 38252 8440 38258 8492
rect 38102 8372 38108 8424
rect 38160 8372 38166 8424
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 37826 7352 37832 7404
rect 37884 7352 37890 7404
rect 38102 7284 38108 7336
rect 38160 7284 38166 7336
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 37274 5652 37280 5704
rect 37332 5692 37338 5704
rect 37829 5695 37887 5701
rect 37829 5692 37841 5695
rect 37332 5664 37841 5692
rect 37332 5652 37338 5664
rect 37829 5661 37841 5664
rect 37875 5661 37887 5695
rect 37829 5655 37887 5661
rect 38102 5584 38108 5636
rect 38160 5584 38166 5636
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 37826 4564 37832 4616
rect 37884 4564 37890 4616
rect 38102 4496 38108 4548
rect 38160 4496 38166 4548
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 37366 3000 37372 3052
rect 37424 3040 37430 3052
rect 37829 3043 37887 3049
rect 37829 3040 37841 3043
rect 37424 3012 37841 3040
rect 37424 3000 37430 3012
rect 37829 3009 37841 3012
rect 37875 3009 37887 3043
rect 37829 3003 37887 3009
rect 38102 2932 38108 2984
rect 38160 2932 38166 2984
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 37826 2388 37832 2440
rect 37884 2388 37890 2440
rect 38102 2320 38108 2372
rect 38160 2320 38166 2372
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4988 39244 5040 39296
rect 5908 39176 5960 39228
rect 10508 39108 10560 39160
rect 11704 39108 11756 39160
rect 21640 39108 21692 39160
rect 22100 39108 22152 39160
rect 28264 39108 28316 39160
rect 31576 39108 31628 39160
rect 3976 38972 4028 39024
rect 23296 38972 23348 39024
rect 5264 38904 5316 38956
rect 18604 38904 18656 38956
rect 3332 38836 3384 38888
rect 23388 38836 23440 38888
rect 5540 38768 5592 38820
rect 16948 38768 17000 38820
rect 18144 38768 18196 38820
rect 20168 38768 20220 38820
rect 26884 38768 26936 38820
rect 6644 38700 6696 38752
rect 22284 38700 22336 38752
rect 23204 38700 23256 38752
rect 34244 38700 34296 38752
rect 13728 38632 13780 38684
rect 26792 38632 26844 38684
rect 6184 38564 6236 38616
rect 31944 38564 31996 38616
rect 3056 38496 3108 38548
rect 23664 38496 23716 38548
rect 6276 38428 6328 38480
rect 17960 38428 18012 38480
rect 18236 38428 18288 38480
rect 32496 38428 32548 38480
rect 7748 38360 7800 38412
rect 25964 38360 26016 38412
rect 7012 38292 7064 38344
rect 18144 38292 18196 38344
rect 26148 38292 26200 38344
rect 31760 38292 31812 38344
rect 6000 38224 6052 38276
rect 35716 38224 35768 38276
rect 5816 38156 5868 38208
rect 33692 38156 33744 38208
rect 6368 38088 6420 38140
rect 16488 38088 16540 38140
rect 20904 38088 20956 38140
rect 35348 38088 35400 38140
rect 4068 38020 4120 38072
rect 23020 38020 23072 38072
rect 25504 38020 25556 38072
rect 30564 38020 30616 38072
rect 30656 38020 30708 38072
rect 32772 38020 32824 38072
rect 2596 37952 2648 38004
rect 13728 37952 13780 38004
rect 21272 37952 21324 38004
rect 35440 37952 35492 38004
rect 7288 37884 7340 37936
rect 27528 37884 27580 37936
rect 4804 37816 4856 37868
rect 26332 37816 26384 37868
rect 26976 37816 27028 37868
rect 33324 37816 33376 37868
rect 6736 37748 6788 37800
rect 31392 37748 31444 37800
rect 6920 37680 6972 37732
rect 30656 37680 30708 37732
rect 3700 37612 3752 37664
rect 20720 37612 20772 37664
rect 21916 37612 21968 37664
rect 25504 37612 25556 37664
rect 26240 37612 26292 37664
rect 34152 37612 34204 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 1768 37204 1820 37256
rect 3424 37247 3476 37256
rect 3424 37213 3433 37247
rect 3433 37213 3467 37247
rect 3467 37213 3476 37247
rect 3424 37204 3476 37213
rect 4528 37247 4580 37256
rect 4528 37213 4537 37247
rect 4537 37213 4571 37247
rect 4571 37213 4580 37247
rect 4528 37204 4580 37213
rect 4620 37204 4672 37256
rect 5080 37204 5132 37256
rect 7012 37315 7064 37324
rect 7012 37281 7021 37315
rect 7021 37281 7055 37315
rect 7055 37281 7064 37315
rect 7012 37272 7064 37281
rect 5724 37136 5776 37188
rect 6552 37136 6604 37188
rect 7196 37247 7248 37256
rect 7196 37213 7205 37247
rect 7205 37213 7239 37247
rect 7239 37213 7248 37247
rect 11060 37408 11112 37460
rect 15200 37408 15252 37460
rect 8576 37340 8628 37392
rect 16488 37340 16540 37392
rect 9496 37272 9548 37324
rect 10968 37272 11020 37324
rect 14832 37272 14884 37324
rect 20076 37272 20128 37324
rect 20996 37408 21048 37460
rect 22560 37408 22612 37460
rect 25780 37408 25832 37460
rect 27620 37408 27672 37460
rect 24308 37340 24360 37392
rect 28448 37340 28500 37392
rect 32956 37408 33008 37460
rect 38476 37408 38528 37460
rect 34520 37340 34572 37392
rect 7196 37204 7248 37213
rect 8208 37204 8260 37256
rect 10508 37247 10560 37256
rect 10508 37213 10517 37247
rect 10517 37213 10551 37247
rect 10551 37213 10560 37247
rect 10508 37204 10560 37213
rect 3516 37068 3568 37120
rect 3792 37068 3844 37120
rect 4620 37068 4672 37120
rect 4712 37111 4764 37120
rect 4712 37077 4721 37111
rect 4721 37077 4755 37111
rect 4755 37077 4764 37111
rect 4712 37068 4764 37077
rect 7288 37068 7340 37120
rect 8484 37179 8536 37188
rect 8484 37145 8493 37179
rect 8493 37145 8527 37179
rect 8527 37145 8536 37179
rect 8484 37136 8536 37145
rect 9128 37111 9180 37120
rect 9128 37077 9137 37111
rect 9137 37077 9171 37111
rect 9171 37077 9180 37111
rect 9128 37068 9180 37077
rect 9680 37136 9732 37188
rect 9772 37136 9824 37188
rect 12440 37136 12492 37188
rect 14372 37247 14424 37256
rect 14372 37213 14381 37247
rect 14381 37213 14415 37247
rect 14415 37213 14424 37247
rect 14372 37204 14424 37213
rect 14648 37204 14700 37256
rect 15016 37204 15068 37256
rect 17040 37247 17092 37256
rect 17040 37213 17049 37247
rect 17049 37213 17083 37247
rect 17083 37213 17092 37247
rect 17040 37204 17092 37213
rect 18328 37204 18380 37256
rect 19248 37204 19300 37256
rect 22100 37247 22152 37256
rect 22100 37213 22109 37247
rect 22109 37213 22143 37247
rect 22143 37213 22152 37247
rect 22100 37204 22152 37213
rect 26976 37272 27028 37324
rect 28080 37272 28132 37324
rect 23572 37247 23624 37256
rect 23572 37213 23581 37247
rect 23581 37213 23615 37247
rect 23615 37213 23624 37247
rect 23572 37204 23624 37213
rect 24952 37204 25004 37256
rect 15752 37136 15804 37188
rect 15936 37179 15988 37188
rect 15936 37145 15945 37179
rect 15945 37145 15979 37179
rect 15979 37145 15988 37179
rect 15936 37136 15988 37145
rect 17316 37179 17368 37188
rect 17316 37145 17325 37179
rect 17325 37145 17359 37179
rect 17359 37145 17368 37179
rect 17316 37136 17368 37145
rect 18788 37179 18840 37188
rect 18788 37145 18797 37179
rect 18797 37145 18831 37179
rect 18831 37145 18840 37179
rect 18788 37136 18840 37145
rect 20720 37136 20772 37188
rect 9588 37111 9640 37120
rect 9588 37077 9597 37111
rect 9597 37077 9631 37111
rect 9631 37077 9640 37111
rect 9588 37068 9640 37077
rect 11796 37111 11848 37120
rect 11796 37077 11805 37111
rect 11805 37077 11839 37111
rect 11839 37077 11848 37111
rect 11796 37068 11848 37077
rect 12716 37068 12768 37120
rect 13084 37068 13136 37120
rect 13360 37111 13412 37120
rect 13360 37077 13369 37111
rect 13369 37077 13403 37111
rect 13403 37077 13412 37111
rect 13360 37068 13412 37077
rect 14280 37068 14332 37120
rect 14556 37111 14608 37120
rect 14556 37077 14565 37111
rect 14565 37077 14599 37111
rect 14599 37077 14608 37111
rect 14556 37068 14608 37077
rect 15016 37068 15068 37120
rect 22468 37136 22520 37188
rect 22652 37179 22704 37188
rect 22652 37145 22661 37179
rect 22661 37145 22695 37179
rect 22695 37145 22704 37179
rect 22652 37136 22704 37145
rect 23480 37068 23532 37120
rect 23848 37179 23900 37188
rect 23848 37145 23857 37179
rect 23857 37145 23891 37179
rect 23891 37145 23900 37179
rect 23848 37136 23900 37145
rect 24124 37136 24176 37188
rect 26608 37204 26660 37256
rect 27252 37204 27304 37256
rect 32404 37315 32456 37324
rect 32404 37281 32413 37315
rect 32413 37281 32447 37315
rect 32447 37281 32456 37315
rect 32404 37272 32456 37281
rect 33692 37315 33744 37324
rect 33692 37281 33701 37315
rect 33701 37281 33735 37315
rect 33735 37281 33744 37315
rect 33692 37272 33744 37281
rect 28264 37204 28316 37256
rect 29184 37247 29236 37256
rect 29184 37213 29193 37247
rect 29193 37213 29227 37247
rect 29227 37213 29236 37247
rect 29184 37204 29236 37213
rect 30288 37247 30340 37256
rect 30288 37213 30297 37247
rect 30297 37213 30331 37247
rect 30331 37213 30340 37247
rect 30288 37204 30340 37213
rect 32036 37204 32088 37256
rect 32312 37247 32364 37256
rect 32312 37213 32328 37247
rect 32328 37213 32362 37247
rect 32362 37213 32364 37247
rect 32312 37204 32364 37213
rect 32588 37247 32640 37256
rect 32588 37213 32597 37247
rect 32597 37213 32631 37247
rect 32631 37213 32640 37247
rect 32588 37204 32640 37213
rect 33140 37204 33192 37256
rect 25320 37136 25372 37188
rect 29460 37136 29512 37188
rect 31116 37136 31168 37188
rect 33784 37204 33836 37256
rect 34244 37247 34296 37256
rect 34244 37213 34253 37247
rect 34253 37213 34287 37247
rect 34287 37213 34296 37247
rect 34244 37204 34296 37213
rect 35164 37204 35216 37256
rect 35532 37204 35584 37256
rect 38108 37204 38160 37256
rect 26240 37068 26292 37120
rect 26516 37068 26568 37120
rect 26884 37068 26936 37120
rect 28356 37068 28408 37120
rect 29092 37111 29144 37120
rect 29092 37077 29101 37111
rect 29101 37077 29135 37111
rect 29135 37077 29144 37111
rect 29092 37068 29144 37077
rect 32220 37068 32272 37120
rect 37556 37136 37608 37188
rect 38016 37179 38068 37188
rect 38016 37145 38025 37179
rect 38025 37145 38059 37179
rect 38059 37145 38068 37179
rect 38016 37136 38068 37145
rect 35808 37068 35860 37120
rect 37372 37068 37424 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 3056 36907 3108 36916
rect 3056 36873 3065 36907
rect 3065 36873 3099 36907
rect 3099 36873 3108 36907
rect 3056 36864 3108 36873
rect 3700 36907 3752 36916
rect 3700 36873 3709 36907
rect 3709 36873 3743 36907
rect 3743 36873 3752 36907
rect 3700 36864 3752 36873
rect 4804 36864 4856 36916
rect 5448 36864 5500 36916
rect 6000 36907 6052 36916
rect 6000 36873 6009 36907
rect 6009 36873 6043 36907
rect 6043 36873 6052 36907
rect 6000 36864 6052 36873
rect 9588 36864 9640 36916
rect 1676 36771 1728 36780
rect 1676 36737 1685 36771
rect 1685 36737 1719 36771
rect 1719 36737 1728 36771
rect 1676 36728 1728 36737
rect 4988 36839 5040 36848
rect 4988 36805 4997 36839
rect 4997 36805 5031 36839
rect 5031 36805 5040 36839
rect 4988 36796 5040 36805
rect 5356 36796 5408 36848
rect 1768 36567 1820 36576
rect 1768 36533 1777 36567
rect 1777 36533 1811 36567
rect 1811 36533 1820 36567
rect 1768 36524 1820 36533
rect 2412 36567 2464 36576
rect 2412 36533 2421 36567
rect 2421 36533 2455 36567
rect 2455 36533 2464 36567
rect 2412 36524 2464 36533
rect 3240 36524 3292 36576
rect 5632 36728 5684 36780
rect 5724 36771 5776 36780
rect 5724 36737 5733 36771
rect 5733 36737 5767 36771
rect 5767 36737 5776 36771
rect 5724 36728 5776 36737
rect 7012 36728 7064 36780
rect 4528 36592 4580 36644
rect 4988 36592 5040 36644
rect 7656 36660 7708 36712
rect 9128 36728 9180 36780
rect 11704 36796 11756 36848
rect 10508 36728 10560 36780
rect 12440 36864 12492 36916
rect 13544 36864 13596 36916
rect 14280 36864 14332 36916
rect 15752 36864 15804 36916
rect 23848 36864 23900 36916
rect 12716 36796 12768 36848
rect 11704 36660 11756 36712
rect 13084 36728 13136 36780
rect 18512 36796 18564 36848
rect 18604 36796 18656 36848
rect 22560 36839 22612 36848
rect 22560 36805 22569 36839
rect 22569 36805 22603 36839
rect 22603 36805 22612 36839
rect 22560 36796 22612 36805
rect 24308 36839 24360 36848
rect 24308 36805 24317 36839
rect 24317 36805 24351 36839
rect 24351 36805 24360 36839
rect 24308 36796 24360 36805
rect 14924 36728 14976 36780
rect 17132 36771 17184 36780
rect 17132 36737 17141 36771
rect 17141 36737 17175 36771
rect 17175 36737 17184 36771
rect 17132 36728 17184 36737
rect 18420 36728 18472 36780
rect 18880 36728 18932 36780
rect 19156 36771 19208 36780
rect 19156 36737 19165 36771
rect 19165 36737 19199 36771
rect 19199 36737 19208 36771
rect 19156 36728 19208 36737
rect 12440 36703 12492 36712
rect 12440 36669 12449 36703
rect 12449 36669 12483 36703
rect 12483 36669 12492 36703
rect 12440 36660 12492 36669
rect 7840 36592 7892 36644
rect 9220 36592 9272 36644
rect 9772 36592 9824 36644
rect 5448 36524 5500 36576
rect 7472 36524 7524 36576
rect 11152 36567 11204 36576
rect 11152 36533 11161 36567
rect 11161 36533 11195 36567
rect 11195 36533 11204 36567
rect 11152 36524 11204 36533
rect 11980 36524 12032 36576
rect 15844 36592 15896 36644
rect 23664 36728 23716 36780
rect 15016 36524 15068 36576
rect 15200 36524 15252 36576
rect 17408 36524 17460 36576
rect 17776 36524 17828 36576
rect 18604 36524 18656 36576
rect 18972 36567 19024 36576
rect 18972 36533 18981 36567
rect 18981 36533 19015 36567
rect 19015 36533 19024 36567
rect 18972 36524 19024 36533
rect 19248 36524 19300 36576
rect 19984 36703 20036 36712
rect 19984 36669 19993 36703
rect 19993 36669 20027 36703
rect 20027 36669 20036 36703
rect 19984 36660 20036 36669
rect 21548 36660 21600 36712
rect 22560 36660 22612 36712
rect 25504 36796 25556 36848
rect 27712 36839 27764 36848
rect 27712 36805 27721 36839
rect 27721 36805 27755 36839
rect 27755 36805 27764 36839
rect 27712 36796 27764 36805
rect 24400 36660 24452 36712
rect 26240 36660 26292 36712
rect 28080 36728 28132 36780
rect 31852 36864 31904 36916
rect 28724 36839 28776 36848
rect 28724 36805 28733 36839
rect 28733 36805 28767 36839
rect 28767 36805 28776 36839
rect 28724 36796 28776 36805
rect 29000 36796 29052 36848
rect 32220 36728 32272 36780
rect 27620 36660 27672 36712
rect 31300 36660 31352 36712
rect 26148 36592 26200 36644
rect 26608 36592 26660 36644
rect 31668 36660 31720 36712
rect 35716 36839 35768 36848
rect 35716 36805 35750 36839
rect 35750 36805 35768 36839
rect 35716 36796 35768 36805
rect 35808 36796 35860 36848
rect 33048 36728 33100 36780
rect 34520 36771 34572 36780
rect 34520 36737 34529 36771
rect 34529 36737 34563 36771
rect 34563 36737 34572 36771
rect 34520 36728 34572 36737
rect 36084 36728 36136 36780
rect 34612 36703 34664 36712
rect 34612 36669 34621 36703
rect 34621 36669 34655 36703
rect 34655 36669 34664 36703
rect 34612 36660 34664 36669
rect 21456 36567 21508 36576
rect 21456 36533 21465 36567
rect 21465 36533 21499 36567
rect 21499 36533 21508 36567
rect 21456 36524 21508 36533
rect 23664 36524 23716 36576
rect 29092 36524 29144 36576
rect 29368 36524 29420 36576
rect 34152 36592 34204 36644
rect 38016 36660 38068 36712
rect 29920 36524 29972 36576
rect 32588 36524 32640 36576
rect 33232 36524 33284 36576
rect 36176 36524 36228 36576
rect 36452 36524 36504 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2596 36363 2648 36372
rect 2596 36329 2605 36363
rect 2605 36329 2639 36363
rect 2639 36329 2648 36363
rect 2596 36320 2648 36329
rect 3332 36363 3384 36372
rect 3332 36329 3341 36363
rect 3341 36329 3375 36363
rect 3375 36329 3384 36363
rect 3332 36320 3384 36329
rect 5264 36363 5316 36372
rect 5264 36329 5273 36363
rect 5273 36329 5307 36363
rect 5307 36329 5316 36363
rect 5264 36320 5316 36329
rect 6736 36363 6788 36372
rect 6736 36329 6745 36363
rect 6745 36329 6779 36363
rect 6779 36329 6788 36363
rect 6736 36320 6788 36329
rect 7748 36363 7800 36372
rect 7748 36329 7757 36363
rect 7757 36329 7791 36363
rect 7791 36329 7800 36363
rect 7748 36320 7800 36329
rect 7840 36320 7892 36372
rect 9864 36320 9916 36372
rect 10508 36363 10560 36372
rect 10508 36329 10517 36363
rect 10517 36329 10551 36363
rect 10551 36329 10560 36363
rect 10508 36320 10560 36329
rect 7196 36252 7248 36304
rect 8576 36295 8628 36304
rect 8576 36261 8585 36295
rect 8585 36261 8619 36295
rect 8619 36261 8628 36295
rect 8576 36252 8628 36261
rect 10416 36252 10468 36304
rect 3240 36159 3292 36168
rect 3240 36125 3249 36159
rect 3249 36125 3283 36159
rect 3283 36125 3292 36159
rect 3240 36116 3292 36125
rect 5080 36116 5132 36168
rect 5448 36116 5500 36168
rect 5908 36159 5960 36168
rect 5908 36125 5917 36159
rect 5917 36125 5951 36159
rect 5951 36125 5960 36159
rect 5908 36116 5960 36125
rect 5816 36048 5868 36100
rect 6092 36091 6144 36100
rect 6092 36057 6101 36091
rect 6101 36057 6135 36091
rect 6135 36057 6144 36091
rect 6092 36048 6144 36057
rect 7196 36048 7248 36100
rect 7472 36159 7524 36168
rect 7472 36125 7481 36159
rect 7481 36125 7515 36159
rect 7515 36125 7524 36159
rect 7472 36116 7524 36125
rect 9220 36184 9272 36236
rect 9588 36184 9640 36236
rect 9864 36227 9916 36236
rect 9864 36193 9873 36227
rect 9873 36193 9907 36227
rect 9907 36193 9916 36227
rect 9864 36184 9916 36193
rect 12716 36252 12768 36304
rect 14924 36252 14976 36304
rect 10968 36184 11020 36236
rect 11704 36227 11756 36236
rect 11704 36193 11713 36227
rect 11713 36193 11747 36227
rect 11747 36193 11756 36227
rect 11704 36184 11756 36193
rect 15844 36252 15896 36304
rect 18420 36252 18472 36304
rect 11796 36116 11848 36168
rect 15200 36227 15252 36236
rect 15200 36193 15209 36227
rect 15209 36193 15243 36227
rect 15243 36193 15252 36227
rect 15200 36184 15252 36193
rect 8116 36048 8168 36100
rect 8300 36048 8352 36100
rect 8484 36048 8536 36100
rect 11704 36048 11756 36100
rect 14832 36116 14884 36168
rect 17132 36116 17184 36168
rect 18604 36184 18656 36236
rect 20444 36252 20496 36304
rect 23572 36320 23624 36372
rect 26240 36320 26292 36372
rect 27712 36320 27764 36372
rect 29276 36320 29328 36372
rect 29828 36320 29880 36372
rect 32036 36320 32088 36372
rect 21548 36227 21600 36236
rect 3516 35980 3568 36032
rect 7012 35980 7064 36032
rect 7564 35980 7616 36032
rect 9680 36023 9732 36032
rect 9680 35989 9689 36023
rect 9689 35989 9723 36023
rect 9723 35989 9732 36023
rect 9680 35980 9732 35989
rect 11152 35980 11204 36032
rect 12072 35980 12124 36032
rect 13636 36023 13688 36032
rect 13636 35989 13645 36023
rect 13645 35989 13679 36023
rect 13679 35989 13688 36023
rect 13636 35980 13688 35989
rect 15752 35980 15804 36032
rect 16396 36048 16448 36100
rect 17316 36023 17368 36032
rect 17316 35989 17325 36023
rect 17325 35989 17359 36023
rect 17359 35989 17368 36023
rect 17316 35980 17368 35989
rect 18052 35980 18104 36032
rect 18420 36159 18472 36168
rect 18420 36125 18429 36159
rect 18429 36125 18463 36159
rect 18463 36125 18472 36159
rect 18420 36116 18472 36125
rect 18512 36116 18564 36168
rect 19248 36116 19300 36168
rect 21548 36193 21557 36227
rect 21557 36193 21591 36227
rect 21591 36193 21600 36227
rect 21548 36184 21600 36193
rect 22652 36184 22704 36236
rect 24676 36184 24728 36236
rect 20168 36116 20220 36168
rect 20904 36159 20956 36168
rect 20904 36125 20913 36159
rect 20913 36125 20947 36159
rect 20947 36125 20956 36159
rect 20904 36116 20956 36125
rect 23848 36159 23900 36168
rect 23848 36125 23857 36159
rect 23857 36125 23891 36159
rect 23891 36125 23900 36159
rect 23848 36116 23900 36125
rect 24216 36116 24268 36168
rect 24584 36159 24636 36168
rect 24584 36125 24593 36159
rect 24593 36125 24627 36159
rect 24627 36125 24636 36159
rect 24584 36116 24636 36125
rect 25412 36227 25464 36236
rect 25412 36193 25421 36227
rect 25421 36193 25455 36227
rect 25455 36193 25464 36227
rect 25412 36184 25464 36193
rect 25504 36184 25556 36236
rect 29460 36252 29512 36304
rect 29920 36252 29972 36304
rect 32864 36252 32916 36304
rect 34428 36320 34480 36372
rect 36084 36252 36136 36304
rect 38108 36295 38160 36304
rect 38108 36261 38117 36295
rect 38117 36261 38151 36295
rect 38151 36261 38160 36295
rect 38108 36252 38160 36261
rect 18604 36048 18656 36100
rect 18972 36048 19024 36100
rect 21180 36048 21232 36100
rect 22284 36048 22336 36100
rect 24676 36048 24728 36100
rect 26056 36116 26108 36168
rect 26608 36116 26660 36168
rect 26884 36159 26936 36168
rect 26884 36125 26893 36159
rect 26893 36125 26927 36159
rect 26927 36125 26936 36159
rect 26884 36116 26936 36125
rect 27620 36184 27672 36236
rect 28540 36184 28592 36236
rect 27804 36116 27856 36168
rect 30104 36184 30156 36236
rect 30380 36184 30432 36236
rect 31852 36227 31904 36236
rect 31852 36193 31861 36227
rect 31861 36193 31895 36227
rect 31895 36193 31904 36227
rect 31852 36184 31904 36193
rect 32956 36184 33008 36236
rect 25044 36048 25096 36100
rect 23112 35980 23164 36032
rect 23572 35980 23624 36032
rect 24860 36023 24912 36032
rect 24860 35989 24869 36023
rect 24869 35989 24903 36023
rect 24903 35989 24912 36023
rect 24860 35980 24912 35989
rect 25136 35980 25188 36032
rect 26056 36023 26108 36032
rect 26056 35989 26065 36023
rect 26065 35989 26099 36023
rect 26099 35989 26108 36023
rect 26056 35980 26108 35989
rect 26240 36048 26292 36100
rect 27620 36091 27672 36100
rect 27620 36057 27629 36091
rect 27629 36057 27663 36091
rect 27663 36057 27672 36091
rect 27620 36048 27672 36057
rect 26976 35980 27028 36032
rect 28080 35980 28132 36032
rect 28172 35980 28224 36032
rect 28816 36159 28868 36168
rect 28816 36125 28825 36159
rect 28825 36125 28859 36159
rect 28859 36125 28868 36159
rect 28816 36116 28868 36125
rect 28908 36116 28960 36168
rect 29092 36116 29144 36168
rect 30840 36116 30892 36168
rect 30104 36048 30156 36100
rect 31944 36048 31996 36100
rect 36084 36159 36136 36168
rect 36084 36125 36093 36159
rect 36093 36125 36127 36159
rect 36127 36125 36136 36159
rect 36084 36116 36136 36125
rect 36176 36116 36228 36168
rect 33324 35980 33376 36032
rect 33416 35980 33468 36032
rect 36544 36048 36596 36100
rect 37188 35980 37240 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4804 35776 4856 35828
rect 6184 35776 6236 35828
rect 6644 35819 6696 35828
rect 6644 35785 6653 35819
rect 6653 35785 6687 35819
rect 6687 35785 6696 35819
rect 6644 35776 6696 35785
rect 9588 35776 9640 35828
rect 15936 35776 15988 35828
rect 17316 35776 17368 35828
rect 3424 35708 3476 35760
rect 5356 35708 5408 35760
rect 5448 35708 5500 35760
rect 4344 35683 4396 35692
rect 4344 35649 4353 35683
rect 4353 35649 4387 35683
rect 4387 35649 4396 35683
rect 4344 35640 4396 35649
rect 4528 35683 4580 35692
rect 4528 35649 4537 35683
rect 4537 35649 4571 35683
rect 4571 35649 4580 35683
rect 4528 35640 4580 35649
rect 4804 35683 4856 35692
rect 4804 35649 4813 35683
rect 4813 35649 4847 35683
rect 4847 35649 4856 35683
rect 4804 35640 4856 35649
rect 4988 35683 5040 35692
rect 4988 35649 4997 35683
rect 4997 35649 5031 35683
rect 5031 35649 5040 35683
rect 4988 35640 5040 35649
rect 5264 35640 5316 35692
rect 5816 35640 5868 35692
rect 6920 35708 6972 35760
rect 7104 35640 7156 35692
rect 9772 35708 9824 35760
rect 10232 35751 10284 35760
rect 10232 35717 10241 35751
rect 10241 35717 10275 35751
rect 10275 35717 10284 35751
rect 10232 35708 10284 35717
rect 19156 35776 19208 35828
rect 19248 35776 19300 35828
rect 7380 35683 7432 35692
rect 7380 35649 7389 35683
rect 7389 35649 7423 35683
rect 7423 35649 7432 35683
rect 7380 35640 7432 35649
rect 6828 35572 6880 35624
rect 8116 35640 8168 35692
rect 9128 35640 9180 35692
rect 11704 35640 11756 35692
rect 12072 35683 12124 35692
rect 12072 35649 12081 35683
rect 12081 35649 12115 35683
rect 12115 35649 12124 35683
rect 12072 35640 12124 35649
rect 7656 35572 7708 35624
rect 9864 35572 9916 35624
rect 12440 35640 12492 35692
rect 13084 35640 13136 35692
rect 7932 35504 7984 35556
rect 12716 35615 12768 35624
rect 12716 35581 12725 35615
rect 12725 35581 12759 35615
rect 12759 35581 12768 35615
rect 12716 35572 12768 35581
rect 15200 35640 15252 35692
rect 15752 35640 15804 35692
rect 3700 35479 3752 35488
rect 3700 35445 3709 35479
rect 3709 35445 3743 35479
rect 3743 35445 3752 35479
rect 3700 35436 3752 35445
rect 4528 35436 4580 35488
rect 5448 35436 5500 35488
rect 5908 35436 5960 35488
rect 14096 35479 14148 35488
rect 14096 35445 14105 35479
rect 14105 35445 14139 35479
rect 14139 35445 14148 35479
rect 14096 35436 14148 35445
rect 14280 35504 14332 35556
rect 15476 35572 15528 35624
rect 18328 35640 18380 35692
rect 21456 35776 21508 35828
rect 21272 35751 21324 35760
rect 21272 35717 21281 35751
rect 21281 35717 21315 35751
rect 21315 35717 21324 35751
rect 21272 35708 21324 35717
rect 22376 35708 22428 35760
rect 23296 35776 23348 35828
rect 23940 35708 23992 35760
rect 16304 35615 16356 35624
rect 16304 35581 16313 35615
rect 16313 35581 16347 35615
rect 16347 35581 16356 35615
rect 16304 35572 16356 35581
rect 17960 35572 18012 35624
rect 17040 35504 17092 35556
rect 18512 35615 18564 35624
rect 18512 35581 18521 35615
rect 18521 35581 18555 35615
rect 18555 35581 18564 35615
rect 18512 35572 18564 35581
rect 22008 35683 22060 35692
rect 22008 35649 22017 35683
rect 22017 35649 22051 35683
rect 22051 35649 22060 35683
rect 22008 35640 22060 35649
rect 23756 35640 23808 35692
rect 24032 35640 24084 35692
rect 25964 35708 26016 35760
rect 19616 35504 19668 35556
rect 20536 35504 20588 35556
rect 21456 35572 21508 35624
rect 22928 35572 22980 35624
rect 25136 35640 25188 35692
rect 25504 35683 25556 35692
rect 25504 35649 25513 35683
rect 25513 35649 25547 35683
rect 25547 35649 25556 35683
rect 25504 35640 25556 35649
rect 27344 35776 27396 35828
rect 27804 35776 27856 35828
rect 28816 35776 28868 35828
rect 32312 35776 32364 35828
rect 32772 35776 32824 35828
rect 32956 35776 33008 35828
rect 33324 35776 33376 35828
rect 37556 35819 37608 35828
rect 37556 35785 37565 35819
rect 37565 35785 37599 35819
rect 37599 35785 37608 35819
rect 37556 35776 37608 35785
rect 24768 35572 24820 35624
rect 25228 35572 25280 35624
rect 25596 35572 25648 35624
rect 25504 35504 25556 35556
rect 26240 35504 26292 35556
rect 15292 35436 15344 35488
rect 18420 35436 18472 35488
rect 20352 35436 20404 35488
rect 23756 35436 23808 35488
rect 25964 35479 26016 35488
rect 25964 35445 25973 35479
rect 25973 35445 26007 35479
rect 26007 35445 26016 35479
rect 25964 35436 26016 35445
rect 26608 35615 26660 35624
rect 26608 35581 26617 35615
rect 26617 35581 26651 35615
rect 26651 35581 26660 35615
rect 26608 35572 26660 35581
rect 31760 35708 31812 35760
rect 28632 35640 28684 35692
rect 29828 35683 29880 35692
rect 29828 35649 29837 35683
rect 29837 35649 29871 35683
rect 29871 35649 29880 35683
rect 29828 35640 29880 35649
rect 29920 35683 29972 35692
rect 29920 35649 29929 35683
rect 29929 35649 29963 35683
rect 29963 35649 29972 35683
rect 29920 35640 29972 35649
rect 31208 35683 31260 35692
rect 31208 35649 31217 35683
rect 31217 35649 31251 35683
rect 31251 35649 31260 35683
rect 31208 35640 31260 35649
rect 32588 35708 32640 35760
rect 33968 35708 34020 35760
rect 36544 35708 36596 35760
rect 36912 35708 36964 35760
rect 33048 35640 33100 35692
rect 33324 35683 33376 35692
rect 33324 35649 33333 35683
rect 33333 35649 33367 35683
rect 33367 35649 33376 35683
rect 33324 35640 33376 35649
rect 33784 35640 33836 35692
rect 37004 35640 37056 35692
rect 37372 35640 37424 35692
rect 26792 35572 26844 35624
rect 27804 35615 27856 35624
rect 27804 35581 27813 35615
rect 27813 35581 27847 35615
rect 27847 35581 27856 35615
rect 27804 35572 27856 35581
rect 28080 35572 28132 35624
rect 29000 35572 29052 35624
rect 30380 35615 30432 35624
rect 30380 35581 30389 35615
rect 30389 35581 30423 35615
rect 30423 35581 30432 35615
rect 30380 35572 30432 35581
rect 30656 35572 30708 35624
rect 32128 35572 32180 35624
rect 32680 35572 32732 35624
rect 33232 35572 33284 35624
rect 34152 35615 34204 35624
rect 34152 35581 34161 35615
rect 34161 35581 34195 35615
rect 34195 35581 34204 35615
rect 34152 35572 34204 35581
rect 36360 35572 36412 35624
rect 38108 35615 38160 35624
rect 38108 35581 38117 35615
rect 38117 35581 38151 35615
rect 38151 35581 38160 35615
rect 38108 35572 38160 35581
rect 26700 35504 26752 35556
rect 26884 35436 26936 35488
rect 28264 35479 28316 35488
rect 28264 35445 28273 35479
rect 28273 35445 28307 35479
rect 28307 35445 28316 35479
rect 28264 35436 28316 35445
rect 28908 35436 28960 35488
rect 29460 35436 29512 35488
rect 30288 35479 30340 35488
rect 30288 35445 30297 35479
rect 30297 35445 30331 35479
rect 30331 35445 30340 35479
rect 30288 35436 30340 35445
rect 30472 35479 30524 35488
rect 30472 35445 30481 35479
rect 30481 35445 30515 35479
rect 30515 35445 30524 35479
rect 30472 35436 30524 35445
rect 32680 35479 32732 35488
rect 32680 35445 32689 35479
rect 32689 35445 32723 35479
rect 32723 35445 32732 35479
rect 32680 35436 32732 35445
rect 33600 35436 33652 35488
rect 36728 35504 36780 35556
rect 35348 35436 35400 35488
rect 36636 35436 36688 35488
rect 38936 35436 38988 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4344 35232 4396 35284
rect 4988 35232 5040 35284
rect 5264 35232 5316 35284
rect 8668 35232 8720 35284
rect 9128 35275 9180 35284
rect 9128 35241 9137 35275
rect 9137 35241 9171 35275
rect 9171 35241 9180 35275
rect 9128 35232 9180 35241
rect 5540 35164 5592 35216
rect 8024 35164 8076 35216
rect 13636 35232 13688 35284
rect 16396 35232 16448 35284
rect 18144 35232 18196 35284
rect 6920 35096 6972 35148
rect 7380 35096 7432 35148
rect 4344 35028 4396 35080
rect 4620 34892 4672 34944
rect 4804 34892 4856 34944
rect 5080 34935 5132 34944
rect 5080 34901 5105 34935
rect 5105 34901 5132 34935
rect 5080 34892 5132 34901
rect 5356 34892 5408 34944
rect 5540 35028 5592 35080
rect 5908 35071 5960 35080
rect 5908 35037 5917 35071
rect 5917 35037 5951 35071
rect 5951 35037 5960 35071
rect 5908 35028 5960 35037
rect 6736 35028 6788 35080
rect 6828 35071 6880 35080
rect 6828 35037 6837 35071
rect 6837 35037 6871 35071
rect 6871 35037 6880 35071
rect 6828 35028 6880 35037
rect 7472 35071 7524 35080
rect 7472 35037 7481 35071
rect 7481 35037 7515 35071
rect 7515 35037 7524 35071
rect 7472 35028 7524 35037
rect 7840 35028 7892 35080
rect 7288 34960 7340 35012
rect 7748 35003 7800 35012
rect 7748 34969 7757 35003
rect 7757 34969 7791 35003
rect 7791 34969 7800 35003
rect 7748 34960 7800 34969
rect 8208 35071 8260 35080
rect 8208 35037 8217 35071
rect 8217 35037 8251 35071
rect 8251 35037 8260 35071
rect 8208 35028 8260 35037
rect 8392 35071 8444 35080
rect 8392 35037 8401 35071
rect 8401 35037 8435 35071
rect 8435 35037 8444 35071
rect 8392 35028 8444 35037
rect 9588 35139 9640 35148
rect 9588 35105 9597 35139
rect 9597 35105 9631 35139
rect 9631 35105 9640 35139
rect 9588 35096 9640 35105
rect 9496 35028 9548 35080
rect 10048 35096 10100 35148
rect 11152 35096 11204 35148
rect 13084 35164 13136 35216
rect 9772 35028 9824 35080
rect 10324 35071 10376 35080
rect 10324 35037 10333 35071
rect 10333 35037 10367 35071
rect 10367 35037 10376 35071
rect 10324 35028 10376 35037
rect 10416 35071 10468 35080
rect 10416 35037 10425 35071
rect 10425 35037 10459 35071
rect 10459 35037 10468 35071
rect 10416 35028 10468 35037
rect 12716 35096 12768 35148
rect 14648 35164 14700 35216
rect 20352 35232 20404 35284
rect 20536 35232 20588 35284
rect 25872 35232 25924 35284
rect 26792 35275 26844 35284
rect 26792 35241 26801 35275
rect 26801 35241 26835 35275
rect 26835 35241 26844 35275
rect 26792 35232 26844 35241
rect 27160 35232 27212 35284
rect 28448 35275 28500 35284
rect 28448 35241 28457 35275
rect 28457 35241 28491 35275
rect 28491 35241 28500 35275
rect 28448 35232 28500 35241
rect 32128 35232 32180 35284
rect 32956 35232 33008 35284
rect 19984 35164 20036 35216
rect 20904 35164 20956 35216
rect 21456 35164 21508 35216
rect 23848 35164 23900 35216
rect 25136 35207 25188 35216
rect 25136 35173 25145 35207
rect 25145 35173 25179 35207
rect 25179 35173 25188 35207
rect 25136 35164 25188 35173
rect 12164 35028 12216 35080
rect 13268 35071 13320 35080
rect 13268 35037 13277 35071
rect 13277 35037 13311 35071
rect 13311 35037 13320 35071
rect 13268 35028 13320 35037
rect 14556 35028 14608 35080
rect 14832 35096 14884 35148
rect 17132 35139 17184 35148
rect 17132 35105 17141 35139
rect 17141 35105 17175 35139
rect 17175 35105 17184 35139
rect 17132 35096 17184 35105
rect 17408 35096 17460 35148
rect 18696 35096 18748 35148
rect 6000 34892 6052 34944
rect 6092 34935 6144 34944
rect 6092 34901 6101 34935
rect 6101 34901 6135 34935
rect 6135 34901 6144 34935
rect 6092 34892 6144 34901
rect 6552 34892 6604 34944
rect 7196 34892 7248 34944
rect 9680 34960 9732 35012
rect 9404 34892 9456 34944
rect 9588 34892 9640 34944
rect 12624 34960 12676 35012
rect 15568 35028 15620 35080
rect 16120 35028 16172 35080
rect 17316 35028 17368 35080
rect 18328 35028 18380 35080
rect 21272 35096 21324 35148
rect 23388 35096 23440 35148
rect 11612 34892 11664 34944
rect 14096 34892 14148 34944
rect 16856 34960 16908 35012
rect 17960 34960 18012 35012
rect 19616 35071 19668 35080
rect 19616 35037 19625 35071
rect 19625 35037 19659 35071
rect 19659 35037 19668 35071
rect 19616 35028 19668 35037
rect 19984 35071 20036 35080
rect 19984 35037 19993 35071
rect 19993 35037 20027 35071
rect 20027 35037 20036 35071
rect 19984 35028 20036 35037
rect 20444 35028 20496 35080
rect 20628 35071 20680 35080
rect 20628 35037 20637 35071
rect 20637 35037 20671 35071
rect 20671 35037 20680 35071
rect 20628 35028 20680 35037
rect 20720 35071 20772 35080
rect 20720 35037 20729 35071
rect 20729 35037 20763 35071
rect 20763 35037 20772 35071
rect 20720 35028 20772 35037
rect 20812 35071 20864 35080
rect 20812 35037 20821 35071
rect 20821 35037 20855 35071
rect 20855 35037 20864 35071
rect 20812 35028 20864 35037
rect 21640 35071 21692 35080
rect 21640 35037 21649 35071
rect 21649 35037 21683 35071
rect 21683 35037 21692 35071
rect 21640 35028 21692 35037
rect 22560 35071 22612 35080
rect 22560 35037 22569 35071
rect 22569 35037 22603 35071
rect 22603 35037 22612 35071
rect 22560 35028 22612 35037
rect 23480 35071 23532 35080
rect 23480 35037 23489 35071
rect 23489 35037 23523 35071
rect 23523 35037 23532 35071
rect 23480 35028 23532 35037
rect 23756 35028 23808 35080
rect 25044 35028 25096 35080
rect 25228 35139 25280 35148
rect 25228 35105 25237 35139
rect 25237 35105 25271 35139
rect 25271 35105 25280 35139
rect 25228 35096 25280 35105
rect 25504 35096 25556 35148
rect 28264 35164 28316 35216
rect 29000 35164 29052 35216
rect 34520 35232 34572 35284
rect 34796 35232 34848 35284
rect 37280 35232 37332 35284
rect 34060 35164 34112 35216
rect 36636 35164 36688 35216
rect 37740 35164 37792 35216
rect 27252 35096 27304 35148
rect 28632 35139 28684 35148
rect 28632 35105 28641 35139
rect 28641 35105 28675 35139
rect 28675 35105 28684 35139
rect 28632 35096 28684 35105
rect 26332 35071 26384 35080
rect 26332 35037 26341 35071
rect 26341 35037 26375 35071
rect 26375 35037 26384 35071
rect 26332 35028 26384 35037
rect 26884 35028 26936 35080
rect 27068 35071 27120 35080
rect 27068 35037 27077 35071
rect 27077 35037 27111 35071
rect 27111 35037 27120 35071
rect 27068 35028 27120 35037
rect 29184 35096 29236 35148
rect 29920 35096 29972 35148
rect 31852 35139 31904 35148
rect 31852 35105 31861 35139
rect 31861 35105 31895 35139
rect 31895 35105 31904 35139
rect 31852 35096 31904 35105
rect 32404 35096 32456 35148
rect 33876 35139 33928 35148
rect 33876 35105 33885 35139
rect 33885 35105 33919 35139
rect 33919 35105 33928 35139
rect 33876 35096 33928 35105
rect 19340 34960 19392 35012
rect 19432 35003 19484 35012
rect 19432 34969 19441 35003
rect 19441 34969 19475 35003
rect 19475 34969 19484 35003
rect 19432 34960 19484 34969
rect 15660 34892 15712 34944
rect 21088 34960 21140 35012
rect 20444 34935 20496 34944
rect 20444 34901 20453 34935
rect 20453 34901 20487 34935
rect 20487 34901 20496 34935
rect 20444 34892 20496 34901
rect 20720 34892 20772 34944
rect 21732 34892 21784 34944
rect 22468 34960 22520 35012
rect 24032 34960 24084 35012
rect 24676 34960 24728 35012
rect 25412 34960 25464 35012
rect 25872 34960 25924 35012
rect 29276 35028 29328 35080
rect 31484 35071 31536 35080
rect 31484 35037 31493 35071
rect 31493 35037 31527 35071
rect 31527 35037 31536 35071
rect 31484 35028 31536 35037
rect 32772 35028 32824 35080
rect 22560 34892 22612 34944
rect 25136 34892 25188 34944
rect 25688 34892 25740 34944
rect 27252 34960 27304 35012
rect 26332 34892 26384 34944
rect 27804 34892 27856 34944
rect 28816 34892 28868 34944
rect 29184 34960 29236 35012
rect 30104 35003 30156 35012
rect 30104 34969 30113 35003
rect 30113 34969 30147 35003
rect 30147 34969 30156 35003
rect 30104 34960 30156 34969
rect 30748 34935 30800 34944
rect 30748 34901 30757 34935
rect 30757 34901 30791 34935
rect 30791 34901 30800 34935
rect 30748 34892 30800 34901
rect 31300 35003 31352 35012
rect 31300 34969 31309 35003
rect 31309 34969 31343 35003
rect 31343 34969 31352 35003
rect 31300 34960 31352 34969
rect 32680 34960 32732 35012
rect 34704 35096 34756 35148
rect 34428 35028 34480 35080
rect 36544 35096 36596 35148
rect 38384 35096 38436 35148
rect 35256 35028 35308 35080
rect 35440 35028 35492 35080
rect 36084 35028 36136 35080
rect 36176 35028 36228 35080
rect 37372 35028 37424 35080
rect 37464 35071 37516 35080
rect 37464 35037 37473 35071
rect 37473 35037 37507 35071
rect 37507 35037 37516 35071
rect 37464 35028 37516 35037
rect 33048 34935 33100 34944
rect 33048 34901 33057 34935
rect 33057 34901 33091 34935
rect 33091 34901 33100 34935
rect 33048 34892 33100 34901
rect 36728 34960 36780 35012
rect 37924 35028 37976 35080
rect 37648 35003 37700 35012
rect 37648 34969 37657 35003
rect 37657 34969 37691 35003
rect 37691 34969 37700 35003
rect 37648 34960 37700 34969
rect 34980 34892 35032 34944
rect 35072 34935 35124 34944
rect 35072 34901 35081 34935
rect 35081 34901 35115 34935
rect 35115 34901 35124 34935
rect 35072 34892 35124 34901
rect 36820 34892 36872 34944
rect 37372 34892 37424 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 3608 34731 3660 34740
rect 3608 34697 3617 34731
rect 3617 34697 3651 34731
rect 3651 34697 3660 34731
rect 3608 34688 3660 34697
rect 4896 34688 4948 34740
rect 5172 34688 5224 34740
rect 6552 34688 6604 34740
rect 3516 34595 3568 34604
rect 3516 34561 3525 34595
rect 3525 34561 3559 34595
rect 3559 34561 3568 34595
rect 3516 34552 3568 34561
rect 4160 34595 4212 34604
rect 4160 34561 4169 34595
rect 4169 34561 4203 34595
rect 4203 34561 4212 34595
rect 4160 34552 4212 34561
rect 5908 34620 5960 34672
rect 5540 34552 5592 34604
rect 5724 34595 5776 34604
rect 5724 34561 5733 34595
rect 5733 34561 5767 34595
rect 5767 34561 5776 34595
rect 5724 34552 5776 34561
rect 11980 34688 12032 34740
rect 7196 34620 7248 34672
rect 5908 34527 5960 34536
rect 5908 34493 5917 34527
rect 5917 34493 5951 34527
rect 5951 34493 5960 34527
rect 5908 34484 5960 34493
rect 6920 34552 6972 34604
rect 7012 34552 7064 34604
rect 7196 34484 7248 34536
rect 7840 34552 7892 34604
rect 8024 34552 8076 34604
rect 9036 34552 9088 34604
rect 9404 34552 9456 34604
rect 5540 34416 5592 34468
rect 7380 34416 7432 34468
rect 7564 34416 7616 34468
rect 8576 34459 8628 34468
rect 8576 34425 8585 34459
rect 8585 34425 8619 34459
rect 8619 34425 8628 34459
rect 8576 34416 8628 34425
rect 9772 34484 9824 34536
rect 10048 34595 10100 34604
rect 10048 34561 10057 34595
rect 10057 34561 10091 34595
rect 10091 34561 10100 34595
rect 10048 34552 10100 34561
rect 14280 34620 14332 34672
rect 15200 34688 15252 34740
rect 15476 34731 15528 34740
rect 15476 34697 15485 34731
rect 15485 34697 15519 34731
rect 15519 34697 15528 34731
rect 15476 34688 15528 34697
rect 17132 34688 17184 34740
rect 19892 34688 19944 34740
rect 20076 34688 20128 34740
rect 20904 34688 20956 34740
rect 21180 34688 21232 34740
rect 22652 34731 22704 34740
rect 22652 34697 22661 34731
rect 22661 34697 22695 34731
rect 22695 34697 22704 34731
rect 22652 34688 22704 34697
rect 23848 34688 23900 34740
rect 20444 34663 20496 34672
rect 10324 34552 10376 34604
rect 11980 34552 12032 34604
rect 12164 34595 12216 34604
rect 12164 34561 12173 34595
rect 12173 34561 12207 34595
rect 12207 34561 12216 34595
rect 12164 34552 12216 34561
rect 14004 34552 14056 34604
rect 12440 34484 12492 34536
rect 14188 34595 14240 34604
rect 14188 34561 14197 34595
rect 14197 34561 14231 34595
rect 14231 34561 14240 34595
rect 14188 34552 14240 34561
rect 14372 34595 14424 34604
rect 14372 34561 14381 34595
rect 14381 34561 14415 34595
rect 14415 34561 14424 34595
rect 14372 34552 14424 34561
rect 14648 34552 14700 34604
rect 15016 34552 15068 34604
rect 15108 34484 15160 34536
rect 16856 34552 16908 34604
rect 17500 34595 17552 34604
rect 17500 34561 17509 34595
rect 17509 34561 17543 34595
rect 17543 34561 17552 34595
rect 17500 34552 17552 34561
rect 17684 34552 17736 34604
rect 17960 34552 18012 34604
rect 19616 34595 19668 34604
rect 19616 34561 19625 34595
rect 19625 34561 19659 34595
rect 19659 34561 19668 34595
rect 19616 34552 19668 34561
rect 19708 34595 19760 34604
rect 19708 34561 19717 34595
rect 19717 34561 19751 34595
rect 19751 34561 19760 34595
rect 19708 34552 19760 34561
rect 20444 34629 20453 34663
rect 20453 34629 20487 34663
rect 20487 34629 20496 34663
rect 20444 34620 20496 34629
rect 23388 34620 23440 34672
rect 20996 34552 21048 34604
rect 17776 34484 17828 34536
rect 21364 34484 21416 34536
rect 21456 34484 21508 34536
rect 23020 34552 23072 34604
rect 23296 34595 23348 34604
rect 23296 34561 23305 34595
rect 23305 34561 23339 34595
rect 23339 34561 23348 34595
rect 23296 34552 23348 34561
rect 25596 34620 25648 34672
rect 24216 34595 24268 34604
rect 24216 34561 24225 34595
rect 24225 34561 24259 34595
rect 24259 34561 24268 34595
rect 24216 34552 24268 34561
rect 26608 34620 26660 34672
rect 27160 34620 27212 34672
rect 26424 34552 26476 34604
rect 26792 34552 26844 34604
rect 27804 34620 27856 34672
rect 27896 34663 27948 34672
rect 27896 34629 27905 34663
rect 27905 34629 27939 34663
rect 27939 34629 27948 34663
rect 27896 34620 27948 34629
rect 27528 34595 27580 34604
rect 27528 34561 27537 34595
rect 27537 34561 27571 34595
rect 27571 34561 27580 34595
rect 27528 34552 27580 34561
rect 28264 34552 28316 34604
rect 31852 34688 31904 34740
rect 33876 34688 33928 34740
rect 34612 34688 34664 34740
rect 36912 34731 36964 34740
rect 36912 34697 36921 34731
rect 36921 34697 36955 34731
rect 36955 34697 36964 34731
rect 36912 34688 36964 34697
rect 37096 34688 37148 34740
rect 29000 34620 29052 34672
rect 27804 34527 27856 34536
rect 27804 34493 27813 34527
rect 27813 34493 27847 34527
rect 27847 34493 27856 34527
rect 30104 34552 30156 34604
rect 30380 34552 30432 34604
rect 30656 34552 30708 34604
rect 30748 34595 30800 34604
rect 30748 34561 30757 34595
rect 30757 34561 30791 34595
rect 30791 34561 30800 34595
rect 30748 34552 30800 34561
rect 27804 34484 27856 34493
rect 29552 34527 29604 34536
rect 29552 34493 29561 34527
rect 29561 34493 29595 34527
rect 29595 34493 29604 34527
rect 29552 34484 29604 34493
rect 31024 34527 31076 34536
rect 31024 34493 31033 34527
rect 31033 34493 31067 34527
rect 31067 34493 31076 34527
rect 31024 34484 31076 34493
rect 31300 34484 31352 34536
rect 32864 34552 32916 34604
rect 32680 34527 32732 34536
rect 32680 34493 32689 34527
rect 32689 34493 32723 34527
rect 32723 34493 32732 34527
rect 32680 34484 32732 34493
rect 33692 34620 33744 34672
rect 34336 34620 34388 34672
rect 33508 34595 33560 34604
rect 33508 34561 33517 34595
rect 33517 34561 33551 34595
rect 33551 34561 33560 34595
rect 33508 34552 33560 34561
rect 33600 34595 33652 34604
rect 33600 34561 33610 34595
rect 33610 34561 33644 34595
rect 33644 34561 33652 34595
rect 33600 34552 33652 34561
rect 33416 34484 33468 34536
rect 34152 34552 34204 34604
rect 35072 34595 35124 34604
rect 35072 34561 35081 34595
rect 35081 34561 35115 34595
rect 35115 34561 35124 34595
rect 35072 34552 35124 34561
rect 35164 34595 35216 34604
rect 35164 34561 35178 34595
rect 35178 34561 35212 34595
rect 35212 34561 35216 34595
rect 35164 34552 35216 34561
rect 35624 34552 35676 34604
rect 35440 34484 35492 34536
rect 36176 34484 36228 34536
rect 36544 34595 36596 34604
rect 36544 34561 36553 34595
rect 36553 34561 36587 34595
rect 36587 34561 36596 34595
rect 36544 34552 36596 34561
rect 37188 34620 37240 34672
rect 9496 34416 9548 34468
rect 10876 34416 10928 34468
rect 12808 34416 12860 34468
rect 12900 34416 12952 34468
rect 4160 34348 4212 34400
rect 7104 34348 7156 34400
rect 9588 34348 9640 34400
rect 10140 34348 10192 34400
rect 13268 34391 13320 34400
rect 13268 34357 13277 34391
rect 13277 34357 13311 34391
rect 13311 34357 13320 34391
rect 13268 34348 13320 34357
rect 13544 34416 13596 34468
rect 16028 34416 16080 34468
rect 13636 34391 13688 34400
rect 13636 34357 13645 34391
rect 13645 34357 13679 34391
rect 13679 34357 13688 34391
rect 13636 34348 13688 34357
rect 13820 34348 13872 34400
rect 14464 34348 14516 34400
rect 14648 34348 14700 34400
rect 17960 34348 18012 34400
rect 18328 34416 18380 34468
rect 19340 34416 19392 34468
rect 25228 34416 25280 34468
rect 25596 34416 25648 34468
rect 25872 34416 25924 34468
rect 32404 34416 32456 34468
rect 32864 34416 32916 34468
rect 33140 34416 33192 34468
rect 34428 34416 34480 34468
rect 34704 34416 34756 34468
rect 35164 34416 35216 34468
rect 36728 34595 36780 34604
rect 36728 34561 36742 34595
rect 36742 34561 36776 34595
rect 36776 34561 36780 34595
rect 36728 34552 36780 34561
rect 37832 34595 37884 34604
rect 37832 34561 37841 34595
rect 37841 34561 37875 34595
rect 37875 34561 37884 34595
rect 37832 34552 37884 34561
rect 38108 34527 38160 34536
rect 38108 34493 38117 34527
rect 38117 34493 38151 34527
rect 38151 34493 38160 34527
rect 38108 34484 38160 34493
rect 36728 34416 36780 34468
rect 36820 34416 36872 34468
rect 37188 34416 37240 34468
rect 20720 34348 20772 34400
rect 20812 34391 20864 34400
rect 20812 34357 20821 34391
rect 20821 34357 20855 34391
rect 20855 34357 20864 34391
rect 20812 34348 20864 34357
rect 21088 34348 21140 34400
rect 21824 34348 21876 34400
rect 22100 34391 22152 34400
rect 22100 34357 22109 34391
rect 22109 34357 22143 34391
rect 22143 34357 22152 34391
rect 22100 34348 22152 34357
rect 22652 34348 22704 34400
rect 24216 34348 24268 34400
rect 25504 34391 25556 34400
rect 25504 34357 25513 34391
rect 25513 34357 25547 34391
rect 25547 34357 25556 34391
rect 25504 34348 25556 34357
rect 27252 34391 27304 34400
rect 27252 34357 27261 34391
rect 27261 34357 27295 34391
rect 27295 34357 27304 34391
rect 27252 34348 27304 34357
rect 27896 34348 27948 34400
rect 28816 34348 28868 34400
rect 30840 34391 30892 34400
rect 30840 34357 30849 34391
rect 30849 34357 30883 34391
rect 30883 34357 30892 34391
rect 30840 34348 30892 34357
rect 32496 34348 32548 34400
rect 33876 34348 33928 34400
rect 37464 34348 37516 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 4988 34144 5040 34196
rect 6828 34144 6880 34196
rect 7564 34187 7616 34196
rect 7564 34153 7573 34187
rect 7573 34153 7607 34187
rect 7607 34153 7616 34187
rect 7564 34144 7616 34153
rect 8208 34144 8260 34196
rect 8576 34144 8628 34196
rect 9680 34144 9732 34196
rect 7932 34076 7984 34128
rect 8024 34076 8076 34128
rect 13084 34144 13136 34196
rect 4068 33983 4120 33992
rect 4068 33949 4077 33983
rect 4077 33949 4111 33983
rect 4111 33949 4120 33983
rect 4068 33940 4120 33949
rect 5172 34008 5224 34060
rect 4988 33983 5040 33992
rect 4988 33949 4997 33983
rect 4997 33949 5031 33983
rect 5031 33949 5040 33983
rect 4988 33940 5040 33949
rect 4896 33872 4948 33924
rect 5540 34008 5592 34060
rect 6092 34008 6144 34060
rect 6552 34008 6604 34060
rect 6184 33940 6236 33992
rect 6644 33940 6696 33992
rect 7288 33940 7340 33992
rect 7472 33983 7524 33992
rect 7472 33949 7481 33983
rect 7481 33949 7515 33983
rect 7515 33949 7524 33983
rect 7472 33940 7524 33949
rect 7840 33940 7892 33992
rect 8944 34008 8996 34060
rect 8392 33983 8444 33992
rect 8392 33949 8401 33983
rect 8401 33949 8435 33983
rect 8435 33949 8444 33983
rect 8392 33940 8444 33949
rect 6552 33915 6604 33924
rect 6552 33881 6561 33915
rect 6561 33881 6595 33915
rect 6595 33881 6604 33915
rect 6552 33872 6604 33881
rect 6736 33915 6788 33924
rect 6736 33881 6745 33915
rect 6745 33881 6779 33915
rect 6779 33881 6788 33915
rect 6736 33872 6788 33881
rect 6920 33915 6972 33924
rect 6920 33881 6929 33915
rect 6929 33881 6963 33915
rect 6963 33881 6972 33915
rect 6920 33872 6972 33881
rect 7104 33872 7156 33924
rect 9036 33872 9088 33924
rect 13176 34076 13228 34128
rect 9680 34008 9732 34060
rect 13360 34144 13412 34196
rect 14556 34187 14608 34196
rect 14556 34153 14565 34187
rect 14565 34153 14599 34187
rect 14599 34153 14608 34187
rect 14556 34144 14608 34153
rect 14740 34187 14792 34196
rect 14740 34153 14749 34187
rect 14749 34153 14783 34187
rect 14783 34153 14792 34187
rect 14740 34144 14792 34153
rect 15844 34144 15896 34196
rect 14372 34051 14424 34060
rect 14372 34017 14381 34051
rect 14381 34017 14415 34051
rect 14415 34017 14424 34051
rect 14372 34008 14424 34017
rect 17500 34076 17552 34128
rect 18880 34076 18932 34128
rect 15568 34008 15620 34060
rect 15752 34051 15804 34060
rect 15752 34017 15761 34051
rect 15761 34017 15795 34051
rect 15795 34017 15804 34051
rect 15752 34008 15804 34017
rect 15844 34051 15896 34060
rect 15844 34017 15853 34051
rect 15853 34017 15887 34051
rect 15887 34017 15896 34051
rect 15844 34008 15896 34017
rect 9772 33940 9824 33992
rect 10324 33983 10376 33992
rect 10324 33949 10333 33983
rect 10333 33949 10367 33983
rect 10367 33949 10376 33983
rect 10324 33940 10376 33949
rect 10876 33940 10928 33992
rect 11152 33940 11204 33992
rect 11520 33940 11572 33992
rect 12440 33940 12492 33992
rect 12532 33983 12584 33992
rect 12532 33949 12541 33983
rect 12541 33949 12575 33983
rect 12575 33949 12584 33983
rect 12532 33940 12584 33949
rect 13176 33915 13228 33924
rect 13176 33881 13185 33915
rect 13185 33881 13219 33915
rect 13219 33881 13228 33915
rect 13176 33872 13228 33881
rect 13636 33983 13688 33992
rect 13636 33949 13645 33983
rect 13645 33949 13679 33983
rect 13679 33949 13688 33983
rect 13636 33940 13688 33949
rect 13820 33940 13872 33992
rect 14648 33940 14700 33992
rect 14832 33940 14884 33992
rect 14924 33940 14976 33992
rect 15108 33940 15160 33992
rect 15660 33983 15712 33992
rect 15660 33949 15669 33983
rect 15669 33949 15703 33983
rect 15703 33949 15712 33983
rect 15660 33940 15712 33949
rect 16028 33983 16080 33992
rect 16028 33949 16037 33983
rect 16037 33949 16071 33983
rect 16071 33949 16080 33983
rect 16028 33940 16080 33949
rect 16672 33983 16724 33992
rect 16672 33949 16681 33983
rect 16681 33949 16715 33983
rect 16715 33949 16724 33983
rect 16672 33940 16724 33949
rect 18236 34008 18288 34060
rect 19708 34076 19760 34128
rect 20628 34144 20680 34196
rect 21640 34144 21692 34196
rect 21824 34144 21876 34196
rect 22100 34144 22152 34196
rect 21364 34076 21416 34128
rect 19524 34008 19576 34060
rect 17960 33940 18012 33992
rect 4068 33804 4120 33856
rect 6092 33847 6144 33856
rect 6092 33813 6101 33847
rect 6101 33813 6135 33847
rect 6135 33813 6144 33847
rect 6092 33804 6144 33813
rect 6184 33804 6236 33856
rect 7472 33804 7524 33856
rect 7748 33847 7800 33856
rect 7748 33813 7757 33847
rect 7757 33813 7791 33847
rect 7791 33813 7800 33847
rect 7748 33804 7800 33813
rect 7932 33804 7984 33856
rect 12348 33804 12400 33856
rect 12992 33804 13044 33856
rect 13452 33804 13504 33856
rect 14004 33804 14056 33856
rect 14188 33872 14240 33924
rect 17592 33915 17644 33924
rect 17592 33881 17601 33915
rect 17601 33881 17635 33915
rect 17635 33881 17644 33915
rect 17592 33872 17644 33881
rect 18880 33940 18932 33992
rect 20352 34008 20404 34060
rect 20628 33940 20680 33992
rect 21272 33983 21324 33992
rect 21272 33949 21281 33983
rect 21281 33949 21315 33983
rect 21315 33949 21324 33983
rect 21272 33940 21324 33949
rect 21548 33940 21600 33992
rect 22100 34051 22152 34060
rect 22100 34017 22109 34051
rect 22109 34017 22143 34051
rect 22143 34017 22152 34051
rect 23020 34144 23072 34196
rect 23940 34144 23992 34196
rect 24400 34144 24452 34196
rect 24860 34187 24912 34196
rect 24860 34153 24869 34187
rect 24869 34153 24903 34187
rect 24903 34153 24912 34187
rect 24860 34144 24912 34153
rect 24952 34144 25004 34196
rect 25780 34144 25832 34196
rect 27712 34144 27764 34196
rect 31576 34144 31628 34196
rect 31852 34144 31904 34196
rect 33140 34144 33192 34196
rect 34152 34144 34204 34196
rect 34244 34144 34296 34196
rect 34428 34144 34480 34196
rect 34612 34144 34664 34196
rect 34704 34144 34756 34196
rect 22100 34008 22152 34017
rect 20720 33872 20772 33924
rect 25320 34076 25372 34128
rect 27436 34076 27488 34128
rect 22928 34051 22980 34060
rect 22928 34017 22937 34051
rect 22937 34017 22971 34051
rect 22971 34017 22980 34051
rect 22928 34008 22980 34017
rect 23112 34051 23164 34060
rect 23112 34017 23121 34051
rect 23121 34017 23155 34051
rect 23155 34017 23164 34051
rect 23112 34008 23164 34017
rect 23756 34051 23808 34060
rect 23756 34017 23765 34051
rect 23765 34017 23799 34051
rect 23799 34017 23808 34051
rect 23756 34008 23808 34017
rect 23940 34008 23992 34060
rect 28080 34076 28132 34128
rect 31024 34076 31076 34128
rect 31208 34076 31260 34128
rect 22652 33940 22704 33992
rect 23020 33940 23072 33992
rect 24952 33983 25004 33992
rect 24952 33949 24961 33983
rect 24961 33949 24995 33983
rect 24995 33949 25004 33983
rect 24952 33940 25004 33949
rect 25320 33940 25372 33992
rect 15476 33804 15528 33856
rect 16856 33847 16908 33856
rect 16856 33813 16865 33847
rect 16865 33813 16899 33847
rect 16899 33813 16908 33847
rect 16856 33804 16908 33813
rect 16948 33804 17000 33856
rect 18788 33804 18840 33856
rect 18880 33847 18932 33856
rect 18880 33813 18889 33847
rect 18889 33813 18923 33847
rect 18923 33813 18932 33847
rect 18880 33804 18932 33813
rect 20904 33804 20956 33856
rect 22744 33872 22796 33924
rect 24124 33872 24176 33924
rect 24400 33872 24452 33924
rect 24584 33915 24636 33924
rect 24584 33881 24593 33915
rect 24593 33881 24627 33915
rect 24627 33881 24636 33915
rect 24584 33872 24636 33881
rect 25412 33872 25464 33924
rect 26148 33983 26200 33992
rect 26148 33949 26157 33983
rect 26157 33949 26191 33983
rect 26191 33949 26200 33983
rect 26148 33940 26200 33949
rect 26240 33983 26292 33992
rect 26240 33949 26249 33983
rect 26249 33949 26283 33983
rect 26283 33949 26292 33983
rect 26240 33940 26292 33949
rect 26424 33940 26476 33992
rect 27160 33940 27212 33992
rect 27528 33940 27580 33992
rect 27620 33940 27672 33992
rect 31852 34008 31904 34060
rect 32128 34076 32180 34128
rect 32496 34008 32548 34060
rect 26516 33872 26568 33924
rect 27804 33872 27856 33924
rect 27896 33872 27948 33924
rect 28172 33983 28224 33992
rect 28172 33949 28181 33983
rect 28181 33949 28215 33983
rect 28215 33949 28224 33983
rect 28172 33940 28224 33949
rect 28816 33940 28868 33992
rect 29092 33940 29144 33992
rect 29276 33940 29328 33992
rect 28356 33872 28408 33924
rect 28632 33872 28684 33924
rect 30288 33983 30340 33992
rect 30288 33949 30297 33983
rect 30297 33949 30331 33983
rect 30331 33949 30340 33983
rect 30288 33940 30340 33949
rect 30012 33915 30064 33924
rect 30012 33881 30021 33915
rect 30021 33881 30055 33915
rect 30055 33881 30064 33915
rect 30012 33872 30064 33881
rect 22376 33847 22428 33856
rect 22376 33813 22385 33847
rect 22385 33813 22419 33847
rect 22419 33813 22428 33847
rect 22376 33804 22428 33813
rect 22560 33804 22612 33856
rect 23020 33804 23072 33856
rect 25596 33804 25648 33856
rect 25688 33804 25740 33856
rect 27160 33804 27212 33856
rect 28172 33804 28224 33856
rect 28724 33804 28776 33856
rect 29092 33847 29144 33856
rect 29092 33813 29101 33847
rect 29101 33813 29135 33847
rect 29135 33813 29144 33847
rect 29092 33804 29144 33813
rect 29460 33804 29512 33856
rect 31208 33940 31260 33992
rect 31392 33983 31444 33992
rect 31392 33949 31401 33983
rect 31401 33949 31435 33983
rect 31435 33949 31444 33983
rect 31392 33940 31444 33949
rect 32864 33940 32916 33992
rect 33232 33940 33284 33992
rect 33416 33983 33468 33992
rect 33416 33949 33425 33983
rect 33425 33949 33459 33983
rect 33459 33949 33468 33983
rect 33416 33940 33468 33949
rect 33692 34008 33744 34060
rect 35716 34144 35768 34196
rect 38292 34144 38344 34196
rect 34888 34076 34940 34128
rect 30748 33872 30800 33924
rect 34060 33940 34112 33992
rect 35256 34008 35308 34060
rect 34520 33940 34572 33992
rect 35716 34008 35768 34060
rect 36084 34008 36136 34060
rect 36820 34051 36872 34060
rect 36820 34017 36829 34051
rect 36829 34017 36863 34051
rect 36863 34017 36872 34051
rect 36820 34008 36872 34017
rect 33692 33872 33744 33924
rect 35992 33983 36044 33992
rect 35992 33949 36001 33983
rect 36001 33949 36035 33983
rect 36035 33949 36044 33983
rect 35992 33940 36044 33949
rect 37096 33983 37148 33992
rect 37096 33949 37130 33983
rect 37130 33949 37148 33983
rect 35716 33872 35768 33924
rect 37096 33940 37148 33949
rect 36268 33872 36320 33924
rect 37832 33872 37884 33924
rect 30472 33804 30524 33856
rect 33600 33804 33652 33856
rect 34336 33804 34388 33856
rect 34612 33804 34664 33856
rect 35808 33804 35860 33856
rect 36176 33804 36228 33856
rect 36452 33804 36504 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4804 33600 4856 33652
rect 4988 33600 5040 33652
rect 8576 33600 8628 33652
rect 3976 33532 4028 33584
rect 7748 33532 7800 33584
rect 9956 33643 10008 33652
rect 9956 33609 9965 33643
rect 9965 33609 9999 33643
rect 9999 33609 10008 33643
rect 9956 33600 10008 33609
rect 8944 33532 8996 33584
rect 4804 33464 4856 33516
rect 5356 33507 5408 33516
rect 5356 33473 5365 33507
rect 5365 33473 5399 33507
rect 5399 33473 5408 33507
rect 5356 33464 5408 33473
rect 5816 33507 5868 33516
rect 5816 33473 5825 33507
rect 5825 33473 5859 33507
rect 5859 33473 5868 33507
rect 5816 33464 5868 33473
rect 4896 33396 4948 33448
rect 5632 33396 5684 33448
rect 6552 33396 6604 33448
rect 7104 33464 7156 33516
rect 8760 33464 8812 33516
rect 9496 33464 9548 33516
rect 11060 33532 11112 33584
rect 13452 33600 13504 33652
rect 13544 33643 13596 33652
rect 13544 33609 13553 33643
rect 13553 33609 13587 33643
rect 13587 33609 13596 33643
rect 13544 33600 13596 33609
rect 14924 33600 14976 33652
rect 15108 33643 15160 33652
rect 15108 33609 15117 33643
rect 15117 33609 15151 33643
rect 15151 33609 15160 33643
rect 15108 33600 15160 33609
rect 12348 33532 12400 33584
rect 13268 33532 13320 33584
rect 10968 33507 11020 33516
rect 7656 33439 7708 33448
rect 7656 33405 7665 33439
rect 7665 33405 7699 33439
rect 7699 33405 7708 33439
rect 7656 33396 7708 33405
rect 8668 33396 8720 33448
rect 9864 33396 9916 33448
rect 10048 33439 10100 33448
rect 10048 33405 10057 33439
rect 10057 33405 10091 33439
rect 10091 33405 10100 33439
rect 10048 33396 10100 33405
rect 10968 33473 10977 33507
rect 10977 33473 11011 33507
rect 11011 33473 11020 33507
rect 10968 33464 11020 33473
rect 11704 33507 11756 33516
rect 11704 33473 11713 33507
rect 11713 33473 11747 33507
rect 11747 33473 11756 33507
rect 11704 33464 11756 33473
rect 11888 33464 11940 33516
rect 12624 33507 12676 33516
rect 12624 33473 12633 33507
rect 12633 33473 12667 33507
rect 12667 33473 12676 33507
rect 12624 33464 12676 33473
rect 10692 33396 10744 33448
rect 13636 33464 13688 33516
rect 14648 33532 14700 33584
rect 15752 33600 15804 33652
rect 16948 33643 17000 33652
rect 16948 33609 16957 33643
rect 16957 33609 16991 33643
rect 16991 33609 17000 33643
rect 16948 33600 17000 33609
rect 17408 33643 17460 33652
rect 17408 33609 17417 33643
rect 17417 33609 17451 33643
rect 17451 33609 17460 33643
rect 17408 33600 17460 33609
rect 17592 33600 17644 33652
rect 17868 33600 17920 33652
rect 18880 33600 18932 33652
rect 21272 33600 21324 33652
rect 21456 33643 21508 33652
rect 21456 33609 21465 33643
rect 21465 33609 21499 33643
rect 21499 33609 21508 33643
rect 21456 33600 21508 33609
rect 22192 33600 22244 33652
rect 24124 33600 24176 33652
rect 14004 33507 14056 33516
rect 14004 33473 14013 33507
rect 14013 33473 14047 33507
rect 14047 33473 14056 33507
rect 14004 33464 14056 33473
rect 14556 33464 14608 33516
rect 15108 33464 15160 33516
rect 13176 33396 13228 33448
rect 13544 33396 13596 33448
rect 13820 33439 13872 33448
rect 13820 33405 13829 33439
rect 13829 33405 13863 33439
rect 13863 33405 13872 33439
rect 13820 33396 13872 33405
rect 7288 33328 7340 33380
rect 7380 33328 7432 33380
rect 9956 33328 10008 33380
rect 12072 33328 12124 33380
rect 14280 33328 14332 33380
rect 15568 33575 15620 33584
rect 15568 33541 15577 33575
rect 15577 33541 15611 33575
rect 15611 33541 15620 33575
rect 15568 33532 15620 33541
rect 15660 33532 15712 33584
rect 15752 33507 15804 33516
rect 15752 33473 15761 33507
rect 15761 33473 15795 33507
rect 15795 33473 15804 33507
rect 15752 33464 15804 33473
rect 15936 33464 15988 33516
rect 16488 33464 16540 33516
rect 17592 33464 17644 33516
rect 16948 33396 17000 33448
rect 17684 33439 17736 33448
rect 17684 33405 17693 33439
rect 17693 33405 17727 33439
rect 17727 33405 17736 33439
rect 17684 33396 17736 33405
rect 18420 33464 18472 33516
rect 3884 33303 3936 33312
rect 3884 33269 3893 33303
rect 3893 33269 3927 33303
rect 3927 33269 3936 33303
rect 3884 33260 3936 33269
rect 4804 33303 4856 33312
rect 4804 33269 4813 33303
rect 4813 33269 4847 33303
rect 4847 33269 4856 33303
rect 4804 33260 4856 33269
rect 4896 33260 4948 33312
rect 5816 33303 5868 33312
rect 5816 33269 5825 33303
rect 5825 33269 5859 33303
rect 5859 33269 5868 33303
rect 5816 33260 5868 33269
rect 6552 33260 6604 33312
rect 6828 33260 6880 33312
rect 8576 33260 8628 33312
rect 10140 33260 10192 33312
rect 11704 33303 11756 33312
rect 11704 33269 11713 33303
rect 11713 33269 11747 33303
rect 11747 33269 11756 33303
rect 11704 33260 11756 33269
rect 12808 33260 12860 33312
rect 13728 33260 13780 33312
rect 13820 33260 13872 33312
rect 15016 33260 15068 33312
rect 17408 33328 17460 33380
rect 20076 33532 20128 33584
rect 24860 33532 24912 33584
rect 27252 33600 27304 33652
rect 27344 33600 27396 33652
rect 30196 33643 30248 33652
rect 30196 33609 30205 33643
rect 30205 33609 30239 33643
rect 30239 33609 30248 33643
rect 30196 33600 30248 33609
rect 30564 33643 30616 33652
rect 30564 33609 30573 33643
rect 30573 33609 30607 33643
rect 30607 33609 30616 33643
rect 30564 33600 30616 33609
rect 32864 33600 32916 33652
rect 20444 33464 20496 33516
rect 19432 33396 19484 33448
rect 17776 33260 17828 33312
rect 17960 33260 18012 33312
rect 20260 33328 20312 33380
rect 21456 33464 21508 33516
rect 21916 33464 21968 33516
rect 21088 33439 21140 33448
rect 21088 33405 21097 33439
rect 21097 33405 21131 33439
rect 21131 33405 21140 33439
rect 21088 33396 21140 33405
rect 22284 33507 22336 33516
rect 22284 33473 22293 33507
rect 22293 33473 22327 33507
rect 22327 33473 22336 33507
rect 22284 33464 22336 33473
rect 22560 33507 22612 33516
rect 22560 33473 22569 33507
rect 22569 33473 22603 33507
rect 22603 33473 22612 33507
rect 22560 33464 22612 33473
rect 22744 33464 22796 33516
rect 23296 33464 23348 33516
rect 24032 33464 24084 33516
rect 24584 33507 24636 33516
rect 24584 33473 24593 33507
rect 24593 33473 24627 33507
rect 24627 33473 24636 33507
rect 24584 33464 24636 33473
rect 25688 33575 25740 33584
rect 25688 33541 25697 33575
rect 25697 33541 25731 33575
rect 25731 33541 25740 33575
rect 25688 33532 25740 33541
rect 28908 33532 28960 33584
rect 25044 33507 25096 33516
rect 25044 33473 25053 33507
rect 25053 33473 25087 33507
rect 25087 33473 25096 33507
rect 25044 33464 25096 33473
rect 25596 33464 25648 33516
rect 23204 33396 23256 33448
rect 23572 33396 23624 33448
rect 23848 33396 23900 33448
rect 24124 33396 24176 33448
rect 25688 33396 25740 33448
rect 25872 33396 25924 33448
rect 26148 33507 26200 33516
rect 26148 33473 26157 33507
rect 26157 33473 26191 33507
rect 26191 33473 26200 33507
rect 26148 33464 26200 33473
rect 26792 33464 26844 33516
rect 27436 33507 27488 33516
rect 27436 33473 27445 33507
rect 27445 33473 27479 33507
rect 27479 33473 27488 33507
rect 27436 33464 27488 33473
rect 27528 33464 27580 33516
rect 29644 33532 29696 33584
rect 29828 33532 29880 33584
rect 30012 33464 30064 33516
rect 22008 33328 22060 33380
rect 22284 33328 22336 33380
rect 22468 33328 22520 33380
rect 23480 33328 23532 33380
rect 27896 33396 27948 33448
rect 30380 33464 30432 33516
rect 32496 33532 32548 33584
rect 33140 33575 33192 33584
rect 33140 33541 33149 33575
rect 33149 33541 33183 33575
rect 33183 33541 33192 33575
rect 33140 33532 33192 33541
rect 31024 33507 31076 33516
rect 31024 33473 31033 33507
rect 31033 33473 31067 33507
rect 31067 33473 31076 33507
rect 31024 33464 31076 33473
rect 30196 33396 30248 33448
rect 32864 33507 32916 33516
rect 32864 33473 32873 33507
rect 32873 33473 32907 33507
rect 32907 33473 32916 33507
rect 32864 33464 32916 33473
rect 33692 33532 33744 33584
rect 33876 33464 33928 33516
rect 32588 33328 32640 33380
rect 18880 33303 18932 33312
rect 18880 33269 18889 33303
rect 18889 33269 18923 33303
rect 18923 33269 18932 33303
rect 18880 33260 18932 33269
rect 21180 33303 21232 33312
rect 21180 33269 21189 33303
rect 21189 33269 21223 33303
rect 21223 33269 21232 33303
rect 21180 33260 21232 33269
rect 21272 33260 21324 33312
rect 22100 33260 22152 33312
rect 22928 33260 22980 33312
rect 24032 33260 24084 33312
rect 24400 33260 24452 33312
rect 25136 33260 25188 33312
rect 25228 33303 25280 33312
rect 25228 33269 25237 33303
rect 25237 33269 25271 33303
rect 25271 33269 25280 33303
rect 25228 33260 25280 33269
rect 25688 33260 25740 33312
rect 26056 33260 26108 33312
rect 26332 33303 26384 33312
rect 26332 33269 26341 33303
rect 26341 33269 26375 33303
rect 26375 33269 26384 33303
rect 26332 33260 26384 33269
rect 27160 33303 27212 33312
rect 27160 33269 27169 33303
rect 27169 33269 27203 33303
rect 27203 33269 27212 33303
rect 27160 33260 27212 33269
rect 27344 33260 27396 33312
rect 27896 33260 27948 33312
rect 28172 33303 28224 33312
rect 28172 33269 28181 33303
rect 28181 33269 28215 33303
rect 28215 33269 28224 33303
rect 28172 33260 28224 33269
rect 28632 33260 28684 33312
rect 29276 33260 29328 33312
rect 29644 33303 29696 33312
rect 29644 33269 29653 33303
rect 29653 33269 29687 33303
rect 29687 33269 29696 33303
rect 29644 33260 29696 33269
rect 30656 33260 30708 33312
rect 32772 33260 32824 33312
rect 33692 33396 33744 33448
rect 34244 33507 34296 33516
rect 34244 33473 34253 33507
rect 34253 33473 34287 33507
rect 34287 33473 34296 33507
rect 34244 33464 34296 33473
rect 34336 33507 34388 33516
rect 34336 33473 34345 33507
rect 34345 33473 34379 33507
rect 34379 33473 34388 33507
rect 34336 33464 34388 33473
rect 34796 33532 34848 33584
rect 35624 33643 35676 33652
rect 35624 33609 35633 33643
rect 35633 33609 35667 33643
rect 35667 33609 35676 33643
rect 35624 33600 35676 33609
rect 35808 33532 35860 33584
rect 34888 33396 34940 33448
rect 34428 33328 34480 33380
rect 35072 33507 35124 33516
rect 35072 33473 35081 33507
rect 35081 33473 35115 33507
rect 35115 33473 35124 33507
rect 35072 33464 35124 33473
rect 35256 33507 35308 33516
rect 35256 33473 35265 33507
rect 35265 33473 35299 33507
rect 35299 33473 35308 33507
rect 35256 33464 35308 33473
rect 37372 33532 37424 33584
rect 36268 33507 36320 33516
rect 36268 33473 36275 33507
rect 36275 33473 36320 33507
rect 36268 33464 36320 33473
rect 35716 33396 35768 33448
rect 35900 33396 35952 33448
rect 36452 33507 36504 33516
rect 36452 33473 36461 33507
rect 36461 33473 36495 33507
rect 36495 33473 36504 33507
rect 36452 33464 36504 33473
rect 36636 33464 36688 33516
rect 36912 33396 36964 33448
rect 37648 33507 37700 33516
rect 37648 33473 37657 33507
rect 37657 33473 37691 33507
rect 37691 33473 37700 33507
rect 37648 33464 37700 33473
rect 38292 33600 38344 33652
rect 37924 33464 37976 33516
rect 39396 33396 39448 33448
rect 36176 33328 36228 33380
rect 36268 33328 36320 33380
rect 36544 33328 36596 33380
rect 33600 33260 33652 33312
rect 34060 33260 34112 33312
rect 36728 33303 36780 33312
rect 36728 33269 36737 33303
rect 36737 33269 36771 33303
rect 36771 33269 36780 33303
rect 36728 33260 36780 33269
rect 37372 33260 37424 33312
rect 38016 33303 38068 33312
rect 38016 33269 38025 33303
rect 38025 33269 38059 33303
rect 38059 33269 38068 33303
rect 38016 33260 38068 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 7840 33056 7892 33108
rect 10048 33056 10100 33108
rect 10968 33056 11020 33108
rect 11888 33056 11940 33108
rect 12624 33099 12676 33108
rect 12624 33065 12633 33099
rect 12633 33065 12667 33099
rect 12667 33065 12676 33099
rect 12624 33056 12676 33065
rect 12900 33056 12952 33108
rect 13268 33099 13320 33108
rect 13268 33065 13277 33099
rect 13277 33065 13311 33099
rect 13311 33065 13320 33099
rect 13268 33056 13320 33065
rect 13544 33056 13596 33108
rect 14004 33056 14056 33108
rect 4620 32988 4672 33040
rect 6184 32988 6236 33040
rect 6460 32988 6512 33040
rect 8024 32988 8076 33040
rect 8484 32988 8536 33040
rect 12164 32988 12216 33040
rect 13360 32988 13412 33040
rect 15292 33099 15344 33108
rect 15292 33065 15301 33099
rect 15301 33065 15335 33099
rect 15335 33065 15344 33099
rect 15292 33056 15344 33065
rect 15660 33056 15712 33108
rect 15844 33056 15896 33108
rect 16120 33056 16172 33108
rect 16488 33099 16540 33108
rect 16488 33065 16497 33099
rect 16497 33065 16531 33099
rect 16531 33065 16540 33099
rect 16488 33056 16540 33065
rect 17224 33056 17276 33108
rect 17868 33056 17920 33108
rect 18972 33056 19024 33108
rect 19984 33056 20036 33108
rect 20352 33099 20404 33108
rect 20352 33065 20361 33099
rect 20361 33065 20395 33099
rect 20395 33065 20404 33099
rect 20352 33056 20404 33065
rect 20628 33056 20680 33108
rect 8208 32920 8260 32972
rect 8576 32963 8628 32972
rect 8576 32929 8585 32963
rect 8585 32929 8619 32963
rect 8619 32929 8628 32963
rect 8576 32920 8628 32929
rect 8668 32920 8720 32972
rect 9220 32920 9272 32972
rect 9680 32920 9732 32972
rect 4988 32852 5040 32904
rect 5172 32716 5224 32768
rect 5632 32852 5684 32904
rect 5724 32852 5776 32904
rect 6368 32852 6420 32904
rect 6460 32852 6512 32904
rect 6736 32852 6788 32904
rect 7196 32852 7248 32904
rect 7840 32852 7892 32904
rect 8484 32895 8536 32904
rect 8484 32861 8493 32895
rect 8493 32861 8527 32895
rect 8527 32861 8536 32895
rect 8484 32852 8536 32861
rect 6920 32784 6972 32836
rect 7932 32784 7984 32836
rect 8852 32852 8904 32904
rect 9496 32895 9548 32904
rect 9496 32861 9505 32895
rect 9505 32861 9539 32895
rect 9539 32861 9548 32895
rect 9496 32852 9548 32861
rect 9588 32895 9640 32904
rect 9588 32861 9597 32895
rect 9597 32861 9631 32895
rect 9631 32861 9640 32895
rect 9588 32852 9640 32861
rect 10416 32895 10468 32904
rect 10416 32861 10425 32895
rect 10425 32861 10459 32895
rect 10459 32861 10468 32895
rect 10416 32852 10468 32861
rect 10692 32895 10744 32904
rect 10692 32861 10701 32895
rect 10701 32861 10735 32895
rect 10735 32861 10744 32895
rect 10692 32852 10744 32861
rect 11428 32852 11480 32904
rect 11612 32895 11664 32904
rect 11612 32861 11621 32895
rect 11621 32861 11655 32895
rect 11655 32861 11664 32895
rect 11612 32852 11664 32861
rect 11796 32895 11848 32904
rect 11796 32861 11805 32895
rect 11805 32861 11839 32895
rect 11839 32861 11848 32895
rect 11796 32852 11848 32861
rect 12072 32920 12124 32972
rect 14096 32920 14148 32972
rect 14648 32920 14700 32972
rect 15016 32920 15068 32972
rect 12348 32827 12400 32836
rect 5448 32716 5500 32768
rect 12348 32793 12357 32827
rect 12357 32793 12391 32827
rect 12391 32793 12400 32827
rect 12348 32784 12400 32793
rect 12440 32784 12492 32836
rect 12716 32852 12768 32904
rect 13544 32852 13596 32904
rect 14188 32852 14240 32904
rect 15752 32920 15804 32972
rect 15384 32895 15436 32904
rect 15384 32861 15393 32895
rect 15393 32861 15427 32895
rect 15427 32861 15436 32895
rect 15384 32852 15436 32861
rect 15476 32852 15528 32904
rect 17316 32988 17368 33040
rect 17684 32988 17736 33040
rect 18420 32988 18472 33040
rect 21824 32988 21876 33040
rect 18880 32920 18932 32972
rect 22100 32988 22152 33040
rect 22376 33099 22428 33108
rect 22376 33065 22385 33099
rect 22385 33065 22419 33099
rect 22419 33065 22428 33099
rect 22376 33056 22428 33065
rect 23756 33056 23808 33108
rect 24492 33056 24544 33108
rect 25044 33056 25096 33108
rect 26700 33056 26752 33108
rect 25228 32988 25280 33040
rect 25320 32988 25372 33040
rect 25872 32988 25924 33040
rect 26792 32988 26844 33040
rect 27896 32988 27948 33040
rect 16856 32852 16908 32904
rect 9128 32759 9180 32768
rect 9128 32725 9137 32759
rect 9137 32725 9171 32759
rect 9171 32725 9180 32759
rect 9128 32716 9180 32725
rect 9312 32716 9364 32768
rect 10416 32716 10468 32768
rect 11796 32716 11848 32768
rect 11888 32716 11940 32768
rect 12900 32716 12952 32768
rect 14188 32716 14240 32768
rect 14280 32716 14332 32768
rect 19432 32852 19484 32904
rect 20628 32852 20680 32904
rect 21088 32852 21140 32904
rect 21180 32852 21232 32904
rect 18328 32827 18380 32836
rect 18328 32793 18337 32827
rect 18337 32793 18371 32827
rect 18371 32793 18380 32827
rect 18328 32784 18380 32793
rect 18420 32784 18472 32836
rect 21272 32784 21324 32836
rect 22744 32963 22796 32972
rect 22744 32929 22753 32963
rect 22753 32929 22787 32963
rect 22787 32929 22796 32963
rect 22744 32920 22796 32929
rect 23756 32963 23808 32972
rect 23756 32929 23765 32963
rect 23765 32929 23799 32963
rect 23799 32929 23808 32963
rect 23756 32920 23808 32929
rect 26884 32920 26936 32972
rect 28356 33056 28408 33108
rect 30472 33056 30524 33108
rect 30656 33056 30708 33108
rect 30932 33056 30984 33108
rect 32496 33056 32548 33108
rect 33324 33056 33376 33108
rect 28448 32988 28500 33040
rect 31760 32988 31812 33040
rect 32128 32988 32180 33040
rect 29368 32920 29420 32972
rect 29552 32920 29604 32972
rect 29736 32920 29788 32972
rect 30380 32963 30432 32972
rect 30380 32929 30389 32963
rect 30389 32929 30423 32963
rect 30423 32929 30432 32963
rect 30380 32920 30432 32929
rect 31024 32920 31076 32972
rect 31484 32920 31536 32972
rect 23296 32852 23348 32904
rect 23664 32852 23716 32904
rect 23848 32895 23900 32904
rect 23848 32861 23857 32895
rect 23857 32861 23891 32895
rect 23891 32861 23900 32895
rect 23848 32852 23900 32861
rect 24400 32852 24452 32904
rect 24768 32852 24820 32904
rect 24952 32895 25004 32904
rect 24952 32861 24961 32895
rect 24961 32861 24995 32895
rect 24995 32861 25004 32895
rect 24952 32852 25004 32861
rect 25044 32895 25096 32904
rect 25044 32861 25053 32895
rect 25053 32861 25087 32895
rect 25087 32861 25096 32895
rect 25044 32852 25096 32861
rect 25228 32895 25280 32904
rect 25228 32861 25237 32895
rect 25237 32861 25271 32895
rect 25271 32861 25280 32895
rect 25228 32852 25280 32861
rect 26056 32852 26108 32904
rect 27436 32895 27488 32904
rect 27436 32861 27445 32895
rect 27445 32861 27479 32895
rect 27479 32861 27488 32895
rect 27436 32852 27488 32861
rect 27528 32895 27580 32904
rect 27528 32861 27537 32895
rect 27537 32861 27571 32895
rect 27571 32861 27580 32895
rect 27528 32852 27580 32861
rect 28172 32852 28224 32904
rect 28356 32895 28408 32904
rect 28356 32861 28365 32895
rect 28365 32861 28399 32895
rect 28399 32861 28408 32895
rect 28356 32852 28408 32861
rect 28816 32895 28868 32904
rect 28816 32861 28825 32895
rect 28825 32861 28859 32895
rect 28859 32861 28868 32895
rect 28816 32852 28868 32861
rect 22928 32784 22980 32836
rect 23480 32784 23532 32836
rect 24676 32784 24728 32836
rect 25320 32784 25372 32836
rect 29276 32784 29328 32836
rect 29736 32784 29788 32836
rect 30196 32895 30248 32904
rect 30196 32861 30205 32895
rect 30205 32861 30239 32895
rect 30239 32861 30248 32895
rect 30196 32852 30248 32861
rect 19064 32716 19116 32768
rect 19156 32716 19208 32768
rect 20812 32716 20864 32768
rect 20904 32759 20956 32768
rect 20904 32725 20913 32759
rect 20913 32725 20947 32759
rect 20947 32725 20956 32759
rect 20904 32716 20956 32725
rect 21456 32716 21508 32768
rect 22100 32716 22152 32768
rect 22560 32716 22612 32768
rect 23204 32716 23256 32768
rect 26148 32716 26200 32768
rect 28908 32716 28960 32768
rect 32128 32852 32180 32904
rect 32312 32895 32364 32904
rect 32312 32861 32321 32895
rect 32321 32861 32355 32895
rect 32355 32861 32364 32895
rect 32312 32852 32364 32861
rect 32588 32852 32640 32904
rect 32680 32852 32732 32904
rect 32864 32852 32916 32904
rect 34520 33056 34572 33108
rect 34152 32988 34204 33040
rect 33140 32852 33192 32904
rect 33324 32895 33376 32904
rect 33324 32861 33333 32895
rect 33333 32861 33367 32895
rect 33367 32861 33376 32895
rect 33324 32852 33376 32861
rect 33416 32895 33468 32904
rect 34336 32963 34388 32972
rect 34336 32929 34345 32963
rect 34345 32929 34379 32963
rect 34379 32929 34388 32963
rect 34336 32920 34388 32929
rect 33416 32861 33430 32895
rect 33430 32861 33464 32895
rect 33464 32861 33468 32895
rect 33416 32852 33468 32861
rect 34520 32852 34572 32904
rect 35072 32895 35124 32904
rect 35072 32861 35081 32895
rect 35081 32861 35115 32895
rect 35115 32861 35124 32895
rect 35072 32852 35124 32861
rect 38016 33056 38068 33108
rect 35716 32920 35768 32972
rect 36728 32920 36780 32972
rect 36636 32852 36688 32904
rect 31760 32716 31812 32768
rect 35808 32827 35860 32836
rect 35808 32793 35817 32827
rect 35817 32793 35851 32827
rect 35851 32793 35860 32827
rect 35808 32784 35860 32793
rect 34704 32716 34756 32768
rect 35348 32716 35400 32768
rect 35716 32716 35768 32768
rect 36544 32784 36596 32836
rect 37464 32784 37516 32836
rect 36176 32759 36228 32768
rect 36176 32725 36185 32759
rect 36185 32725 36219 32759
rect 36219 32725 36228 32759
rect 36176 32716 36228 32725
rect 37832 32716 37884 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 8484 32512 8536 32564
rect 7104 32444 7156 32496
rect 9128 32444 9180 32496
rect 4528 32376 4580 32428
rect 2688 32308 2740 32360
rect 5816 32419 5868 32428
rect 5816 32385 5825 32419
rect 5825 32385 5859 32419
rect 5859 32385 5868 32419
rect 5816 32376 5868 32385
rect 6000 32419 6052 32428
rect 6000 32385 6009 32419
rect 6009 32385 6043 32419
rect 6043 32385 6052 32419
rect 6000 32376 6052 32385
rect 6736 32419 6788 32428
rect 6736 32385 6745 32419
rect 6745 32385 6779 32419
rect 6779 32385 6788 32419
rect 6736 32376 6788 32385
rect 6920 32419 6972 32428
rect 6920 32385 6929 32419
rect 6929 32385 6963 32419
rect 6963 32385 6972 32419
rect 6920 32376 6972 32385
rect 8300 32376 8352 32428
rect 9036 32376 9088 32428
rect 6368 32308 6420 32360
rect 7012 32308 7064 32360
rect 7380 32308 7432 32360
rect 8760 32308 8812 32360
rect 9404 32308 9456 32360
rect 9956 32419 10008 32428
rect 9956 32385 9965 32419
rect 9965 32385 9999 32419
rect 9999 32385 10008 32419
rect 9956 32376 10008 32385
rect 10140 32419 10192 32428
rect 10140 32385 10149 32419
rect 10149 32385 10183 32419
rect 10183 32385 10192 32419
rect 10140 32376 10192 32385
rect 13820 32512 13872 32564
rect 14004 32512 14056 32564
rect 15844 32512 15896 32564
rect 16120 32512 16172 32564
rect 19156 32512 19208 32564
rect 19432 32512 19484 32564
rect 22100 32512 22152 32564
rect 22192 32512 22244 32564
rect 11796 32487 11848 32496
rect 11796 32453 11805 32487
rect 11805 32453 11839 32487
rect 11839 32453 11848 32487
rect 11796 32444 11848 32453
rect 11244 32376 11296 32428
rect 11336 32376 11388 32428
rect 10508 32308 10560 32360
rect 11796 32308 11848 32360
rect 12532 32308 12584 32360
rect 12992 32444 13044 32496
rect 14832 32444 14884 32496
rect 15200 32487 15252 32496
rect 15200 32453 15209 32487
rect 15209 32453 15243 32487
rect 15243 32453 15252 32487
rect 15200 32444 15252 32453
rect 17960 32487 18012 32496
rect 17960 32453 17969 32487
rect 17969 32453 18003 32487
rect 18003 32453 18012 32487
rect 17960 32444 18012 32453
rect 18328 32444 18380 32496
rect 12808 32376 12860 32428
rect 14096 32376 14148 32428
rect 15476 32419 15528 32428
rect 15476 32385 15485 32419
rect 15485 32385 15519 32419
rect 15519 32385 15528 32419
rect 15476 32376 15528 32385
rect 16948 32419 17000 32428
rect 16948 32385 16957 32419
rect 16957 32385 16991 32419
rect 16991 32385 17000 32419
rect 16948 32376 17000 32385
rect 17132 32419 17184 32428
rect 17132 32385 17141 32419
rect 17141 32385 17175 32419
rect 17175 32385 17184 32419
rect 17132 32376 17184 32385
rect 17500 32376 17552 32428
rect 17776 32419 17828 32428
rect 17776 32385 17785 32419
rect 17785 32385 17819 32419
rect 17819 32385 17828 32419
rect 17776 32376 17828 32385
rect 18236 32376 18288 32428
rect 20720 32444 20772 32496
rect 20812 32487 20864 32496
rect 20812 32453 20821 32487
rect 20821 32453 20855 32487
rect 20855 32453 20864 32487
rect 20812 32444 20864 32453
rect 23756 32512 23808 32564
rect 24768 32512 24820 32564
rect 25412 32512 25464 32564
rect 25504 32555 25556 32564
rect 25504 32521 25513 32555
rect 25513 32521 25547 32555
rect 25547 32521 25556 32555
rect 25504 32512 25556 32521
rect 19984 32376 20036 32428
rect 12992 32308 13044 32360
rect 13084 32351 13136 32360
rect 13084 32317 13093 32351
rect 13093 32317 13127 32351
rect 13127 32317 13136 32351
rect 13084 32308 13136 32317
rect 5172 32240 5224 32292
rect 5632 32240 5684 32292
rect 7104 32283 7156 32292
rect 7104 32249 7113 32283
rect 7113 32249 7147 32283
rect 7147 32249 7156 32283
rect 7104 32240 7156 32249
rect 4068 32172 4120 32224
rect 4620 32172 4672 32224
rect 4712 32215 4764 32224
rect 4712 32181 4721 32215
rect 4721 32181 4755 32215
rect 4755 32181 4764 32215
rect 4712 32172 4764 32181
rect 5816 32172 5868 32224
rect 9680 32240 9732 32292
rect 11244 32240 11296 32292
rect 15016 32308 15068 32360
rect 13268 32240 13320 32292
rect 15384 32240 15436 32292
rect 19340 32308 19392 32360
rect 20352 32419 20404 32428
rect 20352 32385 20361 32419
rect 20361 32385 20395 32419
rect 20395 32385 20404 32419
rect 20352 32376 20404 32385
rect 21640 32376 21692 32428
rect 22192 32376 22244 32428
rect 22468 32419 22520 32428
rect 22468 32385 22477 32419
rect 22477 32385 22511 32419
rect 22511 32385 22520 32419
rect 22468 32376 22520 32385
rect 23480 32444 23532 32496
rect 22836 32376 22888 32428
rect 8576 32172 8628 32224
rect 8760 32172 8812 32224
rect 8944 32215 8996 32224
rect 8944 32181 8953 32215
rect 8953 32181 8987 32215
rect 8987 32181 8996 32215
rect 8944 32172 8996 32181
rect 9036 32172 9088 32224
rect 9772 32172 9824 32224
rect 9864 32172 9916 32224
rect 11060 32215 11112 32224
rect 11060 32181 11069 32215
rect 11069 32181 11103 32215
rect 11103 32181 11112 32215
rect 11060 32172 11112 32181
rect 11612 32172 11664 32224
rect 15108 32172 15160 32224
rect 15660 32215 15712 32224
rect 15660 32181 15669 32215
rect 15669 32181 15703 32215
rect 15703 32181 15712 32215
rect 15660 32172 15712 32181
rect 18052 32240 18104 32292
rect 18880 32240 18932 32292
rect 17868 32172 17920 32224
rect 18236 32172 18288 32224
rect 18788 32172 18840 32224
rect 19248 32215 19300 32224
rect 19248 32181 19257 32215
rect 19257 32181 19291 32215
rect 19291 32181 19300 32215
rect 19248 32172 19300 32181
rect 19340 32172 19392 32224
rect 20536 32172 20588 32224
rect 20996 32215 21048 32224
rect 20996 32181 21005 32215
rect 21005 32181 21039 32215
rect 21039 32181 21048 32215
rect 20996 32172 21048 32181
rect 21732 32240 21784 32292
rect 22468 32240 22520 32292
rect 22744 32351 22796 32360
rect 22744 32317 22753 32351
rect 22753 32317 22787 32351
rect 22787 32317 22796 32351
rect 27344 32444 27396 32496
rect 24032 32376 24084 32428
rect 25136 32376 25188 32428
rect 25320 32419 25372 32428
rect 25320 32385 25329 32419
rect 25329 32385 25363 32419
rect 25363 32385 25372 32419
rect 25320 32376 25372 32385
rect 27528 32376 27580 32428
rect 36176 32512 36228 32564
rect 37464 32555 37516 32564
rect 37464 32521 37473 32555
rect 37473 32521 37507 32555
rect 37507 32521 37516 32555
rect 37464 32512 37516 32521
rect 37832 32555 37884 32564
rect 37832 32521 37841 32555
rect 37841 32521 37875 32555
rect 37875 32521 37884 32555
rect 37832 32512 37884 32521
rect 27804 32376 27856 32428
rect 22744 32308 22796 32317
rect 24124 32351 24176 32360
rect 24124 32317 24133 32351
rect 24133 32317 24167 32351
rect 24167 32317 24176 32351
rect 24124 32308 24176 32317
rect 24768 32308 24820 32360
rect 25412 32308 25464 32360
rect 25780 32308 25832 32360
rect 28264 32376 28316 32428
rect 28724 32419 28776 32428
rect 28724 32385 28730 32419
rect 28730 32385 28776 32419
rect 28724 32376 28776 32385
rect 28908 32351 28960 32360
rect 22836 32240 22888 32292
rect 23848 32240 23900 32292
rect 24584 32240 24636 32292
rect 24676 32240 24728 32292
rect 25044 32240 25096 32292
rect 25412 32172 25464 32224
rect 26516 32172 26568 32224
rect 28908 32317 28917 32351
rect 28917 32317 28951 32351
rect 28951 32317 28960 32351
rect 28908 32308 28960 32317
rect 29000 32351 29052 32360
rect 29000 32317 29009 32351
rect 29009 32317 29043 32351
rect 29043 32317 29052 32351
rect 29000 32308 29052 32317
rect 28172 32240 28224 32292
rect 29828 32444 29880 32496
rect 30288 32444 30340 32496
rect 31208 32444 31260 32496
rect 29460 32376 29512 32428
rect 30104 32376 30156 32428
rect 30656 32419 30708 32428
rect 30656 32385 30665 32419
rect 30665 32385 30699 32419
rect 30699 32385 30708 32419
rect 30656 32376 30708 32385
rect 31024 32419 31076 32428
rect 31024 32385 31033 32419
rect 31033 32385 31067 32419
rect 31067 32385 31076 32419
rect 31024 32376 31076 32385
rect 31576 32419 31628 32428
rect 31576 32385 31585 32419
rect 31585 32385 31619 32419
rect 31619 32385 31628 32419
rect 31576 32376 31628 32385
rect 31944 32376 31996 32428
rect 32312 32419 32364 32428
rect 32312 32385 32321 32419
rect 32321 32385 32355 32419
rect 32355 32385 32364 32419
rect 32312 32376 32364 32385
rect 33232 32444 33284 32496
rect 34428 32444 34480 32496
rect 32588 32376 32640 32428
rect 29276 32308 29328 32360
rect 30932 32308 30984 32360
rect 33048 32419 33100 32428
rect 33048 32385 33057 32419
rect 33057 32385 33091 32419
rect 33091 32385 33100 32419
rect 33048 32376 33100 32385
rect 33324 32376 33376 32428
rect 34612 32376 34664 32428
rect 34888 32376 34940 32428
rect 34796 32308 34848 32360
rect 35624 32308 35676 32360
rect 35808 32308 35860 32360
rect 36176 32419 36228 32428
rect 36176 32385 36185 32419
rect 36185 32385 36219 32419
rect 36219 32385 36228 32419
rect 36176 32376 36228 32385
rect 29276 32172 29328 32224
rect 29828 32172 29880 32224
rect 32404 32215 32456 32224
rect 32404 32181 32413 32215
rect 32413 32181 32447 32215
rect 32447 32181 32456 32215
rect 32404 32172 32456 32181
rect 32956 32172 33008 32224
rect 33876 32240 33928 32292
rect 36084 32240 36136 32292
rect 38016 32351 38068 32360
rect 38016 32317 38025 32351
rect 38025 32317 38059 32351
rect 38059 32317 38068 32351
rect 38016 32308 38068 32317
rect 36728 32240 36780 32292
rect 37924 32240 37976 32292
rect 34980 32172 35032 32224
rect 35348 32172 35400 32224
rect 35900 32172 35952 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 6368 31968 6420 32020
rect 7012 31968 7064 32020
rect 8484 31968 8536 32020
rect 4436 31875 4488 31884
rect 4436 31841 4445 31875
rect 4445 31841 4479 31875
rect 4479 31841 4488 31875
rect 4436 31832 4488 31841
rect 5816 31900 5868 31952
rect 9404 31968 9456 32020
rect 10140 31968 10192 32020
rect 12256 31968 12308 32020
rect 9588 31900 9640 31952
rect 9772 31900 9824 31952
rect 13084 31968 13136 32020
rect 5448 31832 5500 31884
rect 4988 31764 5040 31816
rect 5356 31807 5408 31816
rect 5356 31773 5365 31807
rect 5365 31773 5399 31807
rect 5399 31773 5408 31807
rect 5356 31764 5408 31773
rect 5816 31807 5868 31816
rect 5816 31773 5825 31807
rect 5825 31773 5859 31807
rect 5859 31773 5868 31807
rect 5816 31764 5868 31773
rect 6000 31807 6052 31816
rect 6000 31773 6009 31807
rect 6009 31773 6043 31807
rect 6043 31773 6052 31807
rect 6000 31764 6052 31773
rect 6368 31764 6420 31816
rect 6184 31696 6236 31748
rect 4620 31628 4672 31680
rect 4896 31628 4948 31680
rect 5540 31628 5592 31680
rect 6552 31807 6604 31816
rect 6552 31773 6561 31807
rect 6561 31773 6595 31807
rect 6595 31773 6604 31807
rect 6552 31764 6604 31773
rect 6644 31807 6696 31816
rect 6644 31773 6653 31807
rect 6653 31773 6687 31807
rect 6687 31773 6696 31807
rect 6644 31764 6696 31773
rect 7932 31832 7984 31884
rect 9404 31875 9456 31884
rect 9404 31841 9413 31875
rect 9413 31841 9447 31875
rect 9447 31841 9456 31875
rect 9404 31832 9456 31841
rect 9496 31875 9548 31884
rect 9496 31841 9505 31875
rect 9505 31841 9539 31875
rect 9539 31841 9548 31875
rect 9496 31832 9548 31841
rect 10140 31832 10192 31884
rect 8024 31764 8076 31816
rect 8300 31764 8352 31816
rect 7564 31696 7616 31748
rect 7656 31696 7708 31748
rect 8576 31764 8628 31816
rect 9220 31764 9272 31816
rect 8668 31696 8720 31748
rect 9772 31764 9824 31816
rect 10416 31807 10468 31816
rect 10416 31773 10425 31807
rect 10425 31773 10459 31807
rect 10459 31773 10468 31807
rect 10416 31764 10468 31773
rect 10508 31764 10560 31816
rect 11336 31832 11388 31884
rect 10784 31807 10836 31816
rect 10784 31773 10793 31807
rect 10793 31773 10827 31807
rect 10827 31773 10836 31807
rect 10784 31764 10836 31773
rect 11520 31807 11572 31816
rect 11520 31773 11529 31807
rect 11529 31773 11563 31807
rect 11563 31773 11572 31807
rect 11520 31764 11572 31773
rect 12992 31900 13044 31952
rect 13912 31968 13964 32020
rect 14464 31968 14516 32020
rect 14924 32011 14976 32020
rect 14924 31977 14933 32011
rect 14933 31977 14967 32011
rect 14967 31977 14976 32011
rect 14924 31968 14976 31977
rect 16212 32011 16264 32020
rect 16212 31977 16221 32011
rect 16221 31977 16255 32011
rect 16255 31977 16264 32011
rect 16212 31968 16264 31977
rect 16856 31968 16908 32020
rect 17500 31968 17552 32020
rect 13452 31943 13504 31952
rect 13452 31909 13461 31943
rect 13461 31909 13495 31943
rect 13495 31909 13504 31943
rect 13452 31900 13504 31909
rect 15292 31900 15344 31952
rect 12532 31832 12584 31884
rect 12992 31764 13044 31816
rect 13176 31764 13228 31816
rect 14188 31832 14240 31884
rect 15016 31875 15068 31884
rect 15016 31841 15025 31875
rect 15025 31841 15059 31875
rect 15059 31841 15068 31875
rect 15016 31832 15068 31841
rect 16580 31900 16632 31952
rect 17960 31900 18012 31952
rect 17500 31832 17552 31884
rect 18788 31968 18840 32020
rect 19892 31968 19944 32020
rect 18420 31900 18472 31952
rect 18880 31900 18932 31952
rect 20996 31968 21048 32020
rect 22376 31968 22428 32020
rect 22468 31968 22520 32020
rect 22652 31968 22704 32020
rect 24768 32011 24820 32020
rect 24768 31977 24777 32011
rect 24777 31977 24811 32011
rect 24811 31977 24820 32011
rect 24768 31968 24820 31977
rect 20628 31900 20680 31952
rect 21272 31900 21324 31952
rect 21364 31943 21416 31952
rect 21364 31909 21373 31943
rect 21373 31909 21407 31943
rect 21407 31909 21416 31943
rect 21364 31900 21416 31909
rect 26516 31968 26568 32020
rect 26884 31968 26936 32020
rect 27620 31968 27672 32020
rect 28356 31968 28408 32020
rect 13360 31764 13412 31816
rect 13636 31764 13688 31816
rect 14280 31807 14332 31816
rect 14280 31773 14289 31807
rect 14289 31773 14323 31807
rect 14323 31773 14332 31807
rect 14280 31764 14332 31773
rect 14464 31807 14516 31816
rect 14464 31773 14473 31807
rect 14473 31773 14507 31807
rect 14507 31773 14516 31807
rect 14464 31764 14516 31773
rect 15476 31764 15528 31816
rect 16120 31807 16172 31816
rect 16120 31773 16129 31807
rect 16129 31773 16163 31807
rect 16163 31773 16172 31807
rect 16120 31764 16172 31773
rect 16304 31807 16356 31816
rect 16304 31773 16313 31807
rect 16313 31773 16347 31807
rect 16347 31773 16356 31807
rect 16304 31764 16356 31773
rect 6644 31628 6696 31680
rect 6736 31628 6788 31680
rect 7932 31628 7984 31680
rect 8208 31628 8260 31680
rect 9036 31628 9088 31680
rect 10692 31628 10744 31680
rect 12348 31628 12400 31680
rect 13452 31628 13504 31680
rect 14372 31671 14424 31680
rect 14372 31637 14381 31671
rect 14381 31637 14415 31671
rect 14415 31637 14424 31671
rect 14372 31628 14424 31637
rect 14832 31696 14884 31748
rect 15292 31696 15344 31748
rect 17776 31764 17828 31816
rect 17408 31696 17460 31748
rect 18604 31764 18656 31816
rect 20812 31832 20864 31884
rect 19892 31764 19944 31816
rect 21732 31832 21784 31884
rect 23020 31832 23072 31884
rect 24952 31875 25004 31884
rect 24952 31841 24961 31875
rect 24961 31841 24995 31875
rect 24995 31841 25004 31875
rect 24952 31832 25004 31841
rect 25044 31875 25096 31884
rect 25044 31841 25053 31875
rect 25053 31841 25087 31875
rect 25087 31841 25096 31875
rect 25044 31832 25096 31841
rect 25320 31900 25372 31952
rect 25688 31900 25740 31952
rect 26976 31900 27028 31952
rect 27528 31900 27580 31952
rect 31760 31968 31812 32020
rect 31944 31968 31996 32020
rect 29000 31943 29052 31952
rect 29000 31909 29009 31943
rect 29009 31909 29043 31943
rect 29043 31909 29052 31943
rect 29000 31900 29052 31909
rect 25412 31832 25464 31884
rect 20996 31807 21048 31816
rect 20996 31773 21005 31807
rect 21005 31773 21039 31807
rect 21039 31773 21048 31807
rect 20996 31764 21048 31773
rect 17040 31628 17092 31680
rect 17132 31671 17184 31680
rect 17132 31637 17157 31671
rect 17157 31637 17184 31671
rect 17132 31628 17184 31637
rect 17776 31628 17828 31680
rect 18052 31628 18104 31680
rect 20076 31696 20128 31748
rect 20536 31696 20588 31748
rect 21916 31807 21968 31816
rect 21916 31773 21925 31807
rect 21925 31773 21959 31807
rect 21959 31773 21968 31807
rect 21916 31764 21968 31773
rect 22100 31807 22152 31816
rect 22100 31773 22109 31807
rect 22109 31773 22143 31807
rect 22143 31773 22152 31807
rect 22100 31764 22152 31773
rect 22560 31764 22612 31816
rect 23388 31764 23440 31816
rect 25780 31875 25832 31884
rect 25780 31841 25789 31875
rect 25789 31841 25823 31875
rect 25823 31841 25832 31875
rect 25780 31832 25832 31841
rect 26056 31832 26108 31884
rect 26424 31832 26476 31884
rect 26516 31832 26568 31884
rect 28448 31764 28500 31816
rect 28632 31807 28684 31816
rect 28632 31773 28641 31807
rect 28641 31773 28675 31807
rect 28675 31773 28684 31807
rect 28632 31764 28684 31773
rect 21456 31696 21508 31748
rect 18880 31628 18932 31680
rect 24032 31696 24084 31748
rect 24584 31696 24636 31748
rect 25044 31696 25096 31748
rect 23388 31628 23440 31680
rect 23940 31671 23992 31680
rect 23940 31637 23949 31671
rect 23949 31637 23983 31671
rect 23983 31637 23992 31671
rect 23940 31628 23992 31637
rect 24492 31628 24544 31680
rect 26056 31628 26108 31680
rect 27712 31739 27764 31748
rect 27712 31705 27721 31739
rect 27721 31705 27755 31739
rect 27755 31705 27764 31739
rect 27712 31696 27764 31705
rect 27896 31696 27948 31748
rect 28540 31696 28592 31748
rect 29552 31764 29604 31816
rect 30012 31900 30064 31952
rect 32496 31900 32548 31952
rect 32864 31900 32916 31952
rect 33508 31968 33560 32020
rect 34612 31968 34664 32020
rect 34060 31943 34112 31952
rect 34060 31909 34069 31943
rect 34069 31909 34103 31943
rect 34103 31909 34112 31943
rect 34060 31900 34112 31909
rect 29828 31875 29880 31884
rect 29828 31841 29837 31875
rect 29837 31841 29871 31875
rect 29871 31841 29880 31875
rect 29828 31832 29880 31841
rect 30104 31832 30156 31884
rect 30288 31832 30340 31884
rect 30472 31832 30524 31884
rect 30932 31832 30984 31884
rect 31208 31832 31260 31884
rect 31852 31832 31904 31884
rect 35532 31968 35584 32020
rect 36544 31968 36596 32020
rect 37004 31968 37056 32020
rect 30012 31807 30064 31816
rect 30012 31773 30021 31807
rect 30021 31773 30055 31807
rect 30055 31773 30064 31807
rect 30012 31764 30064 31773
rect 30196 31764 30248 31816
rect 31484 31807 31536 31816
rect 31484 31773 31493 31807
rect 31493 31773 31527 31807
rect 31527 31773 31536 31807
rect 31484 31764 31536 31773
rect 32956 31807 33008 31816
rect 32956 31773 32965 31807
rect 32965 31773 32999 31807
rect 32999 31773 33008 31807
rect 32956 31764 33008 31773
rect 27252 31628 27304 31680
rect 28264 31628 28316 31680
rect 32220 31696 32272 31748
rect 33416 31807 33468 31816
rect 33416 31773 33430 31807
rect 33430 31773 33464 31807
rect 33464 31773 33468 31807
rect 33416 31764 33468 31773
rect 33600 31764 33652 31816
rect 33232 31739 33284 31748
rect 33232 31705 33241 31739
rect 33241 31705 33275 31739
rect 33275 31705 33284 31739
rect 33232 31696 33284 31705
rect 33324 31739 33376 31748
rect 33324 31705 33333 31739
rect 33333 31705 33367 31739
rect 33367 31705 33376 31739
rect 33324 31696 33376 31705
rect 33968 31764 34020 31816
rect 36452 31900 36504 31952
rect 34520 31696 34572 31748
rect 34704 31696 34756 31748
rect 34888 31696 34940 31748
rect 35164 31807 35216 31816
rect 35164 31773 35198 31807
rect 35198 31773 35216 31807
rect 35164 31764 35216 31773
rect 36820 31875 36872 31884
rect 36820 31841 36829 31875
rect 36829 31841 36863 31875
rect 36863 31841 36872 31875
rect 36820 31832 36872 31841
rect 37464 31764 37516 31816
rect 29552 31628 29604 31680
rect 30196 31628 30248 31680
rect 31576 31628 31628 31680
rect 32956 31628 33008 31680
rect 38016 31696 38068 31748
rect 33508 31628 33560 31680
rect 34428 31628 34480 31680
rect 34612 31628 34664 31680
rect 35256 31628 35308 31680
rect 35808 31628 35860 31680
rect 36360 31628 36412 31680
rect 36820 31628 36872 31680
rect 37188 31628 37240 31680
rect 37832 31628 37884 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 5172 31331 5224 31340
rect 5172 31297 5181 31331
rect 5181 31297 5215 31331
rect 5215 31297 5224 31331
rect 5172 31288 5224 31297
rect 5080 31220 5132 31272
rect 5724 31288 5776 31340
rect 6736 31288 6788 31340
rect 10876 31424 10928 31476
rect 10968 31424 11020 31476
rect 12716 31424 12768 31476
rect 13636 31424 13688 31476
rect 14372 31424 14424 31476
rect 20996 31424 21048 31476
rect 21180 31424 21232 31476
rect 22192 31424 22244 31476
rect 23112 31424 23164 31476
rect 7840 31356 7892 31408
rect 7196 31288 7248 31340
rect 7656 31288 7708 31340
rect 7932 31331 7984 31340
rect 7932 31297 7941 31331
rect 7941 31297 7975 31331
rect 7975 31297 7984 31331
rect 7932 31288 7984 31297
rect 8024 31331 8076 31340
rect 8024 31297 8033 31331
rect 8033 31297 8067 31331
rect 8067 31297 8076 31331
rect 8024 31288 8076 31297
rect 8944 31356 8996 31408
rect 9220 31356 9272 31408
rect 9496 31356 9548 31408
rect 5908 31263 5960 31272
rect 5908 31229 5917 31263
rect 5917 31229 5951 31263
rect 5951 31229 5960 31263
rect 5908 31220 5960 31229
rect 7748 31220 7800 31272
rect 8760 31220 8812 31272
rect 7656 31152 7708 31204
rect 7840 31152 7892 31204
rect 9404 31288 9456 31340
rect 10692 31356 10744 31408
rect 11336 31356 11388 31408
rect 9312 31220 9364 31272
rect 10876 31331 10928 31340
rect 10876 31297 10885 31331
rect 10885 31297 10919 31331
rect 10919 31297 10928 31331
rect 10876 31288 10928 31297
rect 11060 31331 11112 31340
rect 11060 31297 11069 31331
rect 11069 31297 11103 31331
rect 11103 31297 11112 31331
rect 11060 31288 11112 31297
rect 12348 31331 12400 31340
rect 12348 31297 12357 31331
rect 12357 31297 12391 31331
rect 12391 31297 12400 31331
rect 12348 31288 12400 31297
rect 12440 31288 12492 31340
rect 13728 31356 13780 31408
rect 13084 31288 13136 31340
rect 9864 31263 9916 31272
rect 9864 31229 9873 31263
rect 9873 31229 9907 31263
rect 9907 31229 9916 31263
rect 9864 31220 9916 31229
rect 8944 31152 8996 31204
rect 5448 31084 5500 31136
rect 8300 31084 8352 31136
rect 9036 31084 9088 31136
rect 9128 31084 9180 31136
rect 9772 31195 9824 31204
rect 9772 31161 9781 31195
rect 9781 31161 9815 31195
rect 9815 31161 9824 31195
rect 9772 31152 9824 31161
rect 10416 31152 10468 31204
rect 11060 31152 11112 31204
rect 11520 31220 11572 31272
rect 12624 31220 12676 31272
rect 13268 31220 13320 31272
rect 13544 31288 13596 31340
rect 13820 31288 13872 31340
rect 13912 31331 13964 31340
rect 13912 31297 13921 31331
rect 13921 31297 13955 31331
rect 13955 31297 13964 31331
rect 13912 31288 13964 31297
rect 15200 31356 15252 31408
rect 15936 31356 15988 31408
rect 17592 31356 17644 31408
rect 18236 31356 18288 31408
rect 20444 31356 20496 31408
rect 13728 31220 13780 31272
rect 14372 31220 14424 31272
rect 11980 31152 12032 31204
rect 12808 31152 12860 31204
rect 14924 31288 14976 31340
rect 16856 31331 16908 31340
rect 16856 31297 16865 31331
rect 16865 31297 16899 31331
rect 16899 31297 16908 31331
rect 16856 31288 16908 31297
rect 15016 31220 15068 31272
rect 17132 31288 17184 31340
rect 17408 31288 17460 31340
rect 19432 31288 19484 31340
rect 20260 31331 20312 31340
rect 20260 31297 20294 31331
rect 20294 31297 20312 31331
rect 20260 31288 20312 31297
rect 22468 31331 22520 31340
rect 22468 31297 22477 31331
rect 22477 31297 22511 31331
rect 22511 31297 22520 31331
rect 22468 31288 22520 31297
rect 9956 31084 10008 31136
rect 10876 31084 10928 31136
rect 12256 31084 12308 31136
rect 12624 31084 12676 31136
rect 12716 31084 12768 31136
rect 15200 31152 15252 31204
rect 16580 31152 16632 31204
rect 16856 31152 16908 31204
rect 19340 31220 19392 31272
rect 22652 31331 22704 31340
rect 22652 31297 22661 31331
rect 22661 31297 22695 31331
rect 22695 31297 22704 31331
rect 22652 31288 22704 31297
rect 23204 31288 23256 31340
rect 23664 31356 23716 31408
rect 23388 31288 23440 31340
rect 25504 31331 25556 31340
rect 25504 31297 25513 31331
rect 25513 31297 25547 31331
rect 25547 31297 25556 31331
rect 25504 31288 25556 31297
rect 25596 31331 25648 31340
rect 25596 31297 25605 31331
rect 25605 31297 25639 31331
rect 25639 31297 25648 31331
rect 25596 31288 25648 31297
rect 23112 31220 23164 31272
rect 32036 31424 32088 31476
rect 32496 31424 32548 31476
rect 27620 31356 27672 31408
rect 29092 31356 29144 31408
rect 26976 31288 27028 31340
rect 21272 31152 21324 31204
rect 24952 31152 25004 31204
rect 16120 31084 16172 31136
rect 17224 31084 17276 31136
rect 18144 31084 18196 31136
rect 18512 31084 18564 31136
rect 19064 31084 19116 31136
rect 19984 31084 20036 31136
rect 20628 31084 20680 31136
rect 21824 31084 21876 31136
rect 21916 31084 21968 31136
rect 22560 31084 22612 31136
rect 22744 31127 22796 31136
rect 22744 31093 22753 31127
rect 22753 31093 22787 31127
rect 22787 31093 22796 31127
rect 22744 31084 22796 31093
rect 27160 31152 27212 31204
rect 26148 31127 26200 31136
rect 26148 31093 26157 31127
rect 26157 31093 26191 31127
rect 26191 31093 26200 31127
rect 26148 31084 26200 31093
rect 27528 31263 27580 31272
rect 27528 31229 27537 31263
rect 27537 31229 27571 31263
rect 27571 31229 27580 31263
rect 27528 31220 27580 31229
rect 28632 31288 28684 31340
rect 29276 31288 29328 31340
rect 29736 31356 29788 31408
rect 30196 31356 30248 31408
rect 33324 31424 33376 31476
rect 34060 31424 34112 31476
rect 34520 31424 34572 31476
rect 37464 31467 37516 31476
rect 37464 31433 37473 31467
rect 37473 31433 37507 31467
rect 37507 31433 37516 31467
rect 37464 31424 37516 31433
rect 30656 31288 30708 31340
rect 31392 31288 31444 31340
rect 28540 31263 28592 31272
rect 28540 31229 28549 31263
rect 28549 31229 28583 31263
rect 28583 31229 28592 31263
rect 28540 31220 28592 31229
rect 30840 31152 30892 31204
rect 31208 31220 31260 31272
rect 32312 31288 32364 31340
rect 32496 31288 32548 31340
rect 32864 31331 32916 31340
rect 32864 31297 32873 31331
rect 32873 31297 32907 31331
rect 32907 31297 32916 31331
rect 32864 31288 32916 31297
rect 33508 31356 33560 31408
rect 34244 31399 34296 31408
rect 34244 31365 34253 31399
rect 34253 31365 34287 31399
rect 34287 31365 34296 31399
rect 34244 31356 34296 31365
rect 34704 31356 34756 31408
rect 37832 31399 37884 31408
rect 37832 31365 37841 31399
rect 37841 31365 37875 31399
rect 37875 31365 37884 31399
rect 37832 31356 37884 31365
rect 31760 31220 31812 31272
rect 33140 31220 33192 31272
rect 33232 31220 33284 31272
rect 33416 31220 33468 31272
rect 32128 31152 32180 31204
rect 34428 31331 34480 31340
rect 34428 31297 34442 31331
rect 34442 31297 34476 31331
rect 34476 31297 34480 31331
rect 34428 31288 34480 31297
rect 34796 31288 34848 31340
rect 35256 31331 35308 31340
rect 35256 31297 35265 31331
rect 35265 31297 35299 31331
rect 35299 31297 35308 31331
rect 35256 31288 35308 31297
rect 35440 31331 35492 31340
rect 35440 31297 35449 31331
rect 35449 31297 35483 31331
rect 35483 31297 35492 31331
rect 35440 31288 35492 31297
rect 36084 31288 36136 31340
rect 36360 31331 36412 31340
rect 36360 31297 36367 31331
rect 36367 31297 36412 31331
rect 36360 31288 36412 31297
rect 35808 31220 35860 31272
rect 36636 31331 36688 31340
rect 36636 31297 36650 31331
rect 36650 31297 36684 31331
rect 36684 31297 36688 31331
rect 36636 31288 36688 31297
rect 36820 31288 36872 31340
rect 29276 31084 29328 31136
rect 29736 31084 29788 31136
rect 30196 31084 30248 31136
rect 30472 31127 30524 31136
rect 30472 31093 30481 31127
rect 30481 31093 30515 31127
rect 30515 31093 30524 31127
rect 30472 31084 30524 31093
rect 31208 31084 31260 31136
rect 34152 31084 34204 31136
rect 34428 31084 34480 31136
rect 34980 31084 35032 31136
rect 35716 31084 35768 31136
rect 36176 31152 36228 31204
rect 36636 31152 36688 31204
rect 36268 31084 36320 31136
rect 36820 31127 36872 31136
rect 36820 31093 36829 31127
rect 36829 31093 36863 31127
rect 36863 31093 36872 31127
rect 38108 31263 38160 31272
rect 38108 31229 38117 31263
rect 38117 31229 38151 31263
rect 38151 31229 38160 31263
rect 38108 31220 38160 31229
rect 36820 31084 36872 31093
rect 37372 31084 37424 31136
rect 37924 31084 37976 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 6000 30880 6052 30932
rect 8208 30880 8260 30932
rect 11060 30880 11112 30932
rect 12164 30880 12216 30932
rect 9036 30812 9088 30864
rect 12256 30812 12308 30864
rect 5356 30719 5408 30728
rect 5356 30685 5365 30719
rect 5365 30685 5399 30719
rect 5399 30685 5408 30719
rect 5356 30676 5408 30685
rect 7104 30744 7156 30796
rect 8484 30744 8536 30796
rect 8944 30744 8996 30796
rect 6644 30676 6696 30728
rect 6920 30676 6972 30728
rect 7288 30676 7340 30728
rect 9680 30744 9732 30796
rect 10140 30744 10192 30796
rect 11428 30744 11480 30796
rect 14464 30880 14516 30932
rect 14832 30880 14884 30932
rect 5080 30540 5132 30592
rect 7472 30540 7524 30592
rect 8484 30608 8536 30660
rect 8760 30608 8812 30660
rect 9496 30676 9548 30728
rect 10232 30719 10284 30728
rect 10232 30685 10241 30719
rect 10241 30685 10275 30719
rect 10275 30685 10284 30719
rect 10232 30676 10284 30685
rect 12624 30744 12676 30796
rect 14464 30744 14516 30796
rect 15752 30744 15804 30796
rect 17592 30880 17644 30932
rect 20260 30880 20312 30932
rect 21088 30880 21140 30932
rect 21732 30880 21784 30932
rect 18052 30812 18104 30864
rect 23756 30880 23808 30932
rect 23940 30880 23992 30932
rect 22284 30812 22336 30864
rect 22652 30812 22704 30864
rect 8392 30540 8444 30592
rect 9588 30608 9640 30660
rect 11336 30651 11388 30660
rect 11336 30617 11345 30651
rect 11345 30617 11379 30651
rect 11379 30617 11388 30651
rect 11336 30608 11388 30617
rect 11520 30651 11572 30660
rect 11520 30617 11545 30651
rect 11545 30617 11572 30651
rect 11520 30608 11572 30617
rect 12072 30608 12124 30660
rect 12992 30676 13044 30728
rect 13176 30719 13228 30728
rect 13176 30685 13185 30719
rect 13185 30685 13219 30719
rect 13219 30685 13228 30719
rect 13176 30676 13228 30685
rect 13360 30719 13412 30728
rect 13360 30685 13369 30719
rect 13369 30685 13403 30719
rect 13403 30685 13412 30719
rect 13360 30676 13412 30685
rect 13452 30719 13504 30728
rect 13452 30685 13487 30719
rect 13487 30685 13504 30719
rect 13452 30676 13504 30685
rect 12900 30608 12952 30660
rect 13820 30676 13872 30728
rect 15292 30719 15344 30728
rect 15292 30685 15301 30719
rect 15301 30685 15335 30719
rect 15335 30685 15344 30719
rect 15292 30676 15344 30685
rect 15384 30676 15436 30728
rect 18144 30676 18196 30728
rect 20536 30719 20588 30728
rect 20536 30685 20545 30719
rect 20545 30685 20579 30719
rect 20579 30685 20588 30719
rect 20536 30676 20588 30685
rect 22836 30744 22888 30796
rect 9496 30540 9548 30592
rect 10232 30540 10284 30592
rect 11796 30540 11848 30592
rect 13728 30608 13780 30660
rect 13452 30540 13504 30592
rect 15016 30608 15068 30660
rect 16488 30608 16540 30660
rect 16948 30608 17000 30660
rect 14832 30583 14884 30592
rect 14832 30549 14841 30583
rect 14841 30549 14875 30583
rect 14875 30549 14884 30583
rect 14832 30540 14884 30549
rect 17592 30540 17644 30592
rect 17960 30651 18012 30660
rect 17960 30617 17969 30651
rect 17969 30617 18003 30651
rect 18003 30617 18012 30651
rect 17960 30608 18012 30617
rect 18328 30608 18380 30660
rect 18512 30608 18564 30660
rect 20628 30608 20680 30660
rect 22008 30719 22060 30728
rect 22008 30685 22017 30719
rect 22017 30685 22051 30719
rect 22051 30685 22060 30719
rect 22008 30676 22060 30685
rect 22100 30719 22152 30728
rect 22100 30685 22109 30719
rect 22109 30685 22143 30719
rect 22143 30685 22152 30719
rect 22100 30676 22152 30685
rect 22376 30676 22428 30728
rect 22652 30719 22704 30728
rect 22652 30685 22661 30719
rect 22661 30685 22695 30719
rect 22695 30685 22704 30719
rect 22652 30676 22704 30685
rect 23480 30744 23532 30796
rect 24308 30744 24360 30796
rect 24768 30787 24820 30796
rect 24768 30753 24777 30787
rect 24777 30753 24811 30787
rect 24811 30753 24820 30787
rect 24768 30744 24820 30753
rect 26056 30812 26108 30864
rect 25780 30744 25832 30796
rect 20904 30540 20956 30592
rect 22468 30608 22520 30660
rect 22560 30608 22612 30660
rect 22192 30540 22244 30592
rect 24768 30608 24820 30660
rect 25504 30676 25556 30728
rect 26608 30676 26660 30728
rect 27344 30812 27396 30864
rect 27068 30744 27120 30796
rect 27528 30880 27580 30932
rect 28632 30880 28684 30932
rect 29276 30880 29328 30932
rect 30840 30880 30892 30932
rect 31208 30923 31260 30932
rect 31208 30889 31217 30923
rect 31217 30889 31251 30923
rect 31251 30889 31260 30923
rect 31208 30880 31260 30889
rect 31760 30880 31812 30932
rect 32128 30880 32180 30932
rect 32496 30880 32548 30932
rect 36084 30880 36136 30932
rect 37556 30880 37608 30932
rect 38200 30880 38252 30932
rect 28172 30812 28224 30864
rect 28356 30812 28408 30864
rect 28816 30812 28868 30864
rect 29000 30812 29052 30864
rect 27436 30719 27488 30728
rect 27436 30685 27445 30719
rect 27445 30685 27479 30719
rect 27479 30685 27488 30719
rect 27436 30676 27488 30685
rect 26424 30608 26476 30660
rect 28172 30608 28224 30660
rect 28632 30676 28684 30728
rect 29552 30744 29604 30796
rect 30012 30744 30064 30796
rect 30104 30744 30156 30796
rect 30380 30744 30432 30796
rect 31484 30812 31536 30864
rect 31668 30744 31720 30796
rect 28816 30676 28868 30728
rect 29828 30676 29880 30728
rect 31760 30719 31812 30728
rect 31760 30685 31769 30719
rect 31769 30685 31803 30719
rect 31803 30685 31812 30719
rect 31760 30676 31812 30685
rect 31852 30719 31904 30728
rect 31852 30685 31861 30719
rect 31861 30685 31895 30719
rect 31895 30685 31904 30719
rect 31852 30676 31904 30685
rect 32312 30812 32364 30864
rect 32312 30676 32364 30728
rect 32864 30812 32916 30864
rect 33140 30812 33192 30864
rect 36820 30812 36872 30864
rect 32956 30744 33008 30796
rect 30380 30608 30432 30660
rect 24032 30540 24084 30592
rect 25780 30540 25832 30592
rect 26332 30540 26384 30592
rect 26884 30583 26936 30592
rect 26884 30549 26893 30583
rect 26893 30549 26927 30583
rect 26927 30549 26936 30583
rect 26884 30540 26936 30549
rect 27620 30540 27672 30592
rect 27712 30540 27764 30592
rect 28540 30540 28592 30592
rect 28724 30540 28776 30592
rect 28908 30583 28960 30592
rect 28908 30549 28917 30583
rect 28917 30549 28951 30583
rect 28951 30549 28960 30583
rect 28908 30540 28960 30549
rect 29828 30540 29880 30592
rect 31392 30540 31444 30592
rect 32588 30540 32640 30592
rect 33232 30719 33284 30728
rect 33232 30685 33246 30719
rect 33246 30685 33280 30719
rect 33280 30685 33284 30719
rect 33968 30744 34020 30796
rect 37096 30787 37148 30796
rect 37096 30753 37105 30787
rect 37105 30753 37139 30787
rect 37139 30753 37148 30787
rect 37096 30744 37148 30753
rect 37372 30744 37424 30796
rect 38292 30787 38344 30796
rect 38292 30753 38301 30787
rect 38301 30753 38335 30787
rect 38335 30753 38344 30787
rect 38292 30744 38344 30753
rect 33232 30676 33284 30685
rect 33140 30651 33192 30660
rect 33140 30617 33149 30651
rect 33149 30617 33183 30651
rect 33183 30617 33192 30651
rect 33140 30608 33192 30617
rect 33784 30608 33836 30660
rect 34888 30719 34940 30728
rect 34888 30685 34897 30719
rect 34897 30685 34931 30719
rect 34931 30685 34940 30719
rect 34888 30676 34940 30685
rect 35440 30676 35492 30728
rect 35900 30719 35952 30728
rect 35900 30685 35909 30719
rect 35909 30685 35943 30719
rect 35943 30685 35952 30719
rect 35900 30676 35952 30685
rect 36084 30719 36136 30728
rect 36084 30685 36091 30719
rect 36091 30685 36136 30719
rect 36084 30676 36136 30685
rect 36544 30676 36596 30728
rect 36636 30676 36688 30728
rect 36820 30676 36872 30728
rect 37188 30719 37240 30728
rect 37188 30685 37197 30719
rect 37197 30685 37231 30719
rect 37231 30685 37240 30719
rect 37188 30676 37240 30685
rect 38384 30676 38436 30728
rect 33324 30540 33376 30592
rect 33508 30540 33560 30592
rect 33600 30540 33652 30592
rect 34060 30540 34112 30592
rect 36176 30651 36228 30660
rect 36176 30617 36185 30651
rect 36185 30617 36219 30651
rect 36219 30617 36228 30651
rect 36176 30608 36228 30617
rect 36268 30651 36320 30660
rect 36268 30617 36277 30651
rect 36277 30617 36311 30651
rect 36311 30617 36320 30651
rect 36268 30608 36320 30617
rect 37648 30540 37700 30592
rect 38016 30540 38068 30592
rect 38292 30583 38344 30592
rect 38292 30549 38301 30583
rect 38301 30549 38335 30583
rect 38335 30549 38344 30583
rect 38292 30540 38344 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 6000 30336 6052 30388
rect 11336 30336 11388 30388
rect 8024 30268 8076 30320
rect 8484 30268 8536 30320
rect 9128 30268 9180 30320
rect 9220 30268 9272 30320
rect 6644 29996 6696 30048
rect 8116 30200 8168 30252
rect 8944 30200 8996 30252
rect 9772 30243 9824 30252
rect 9772 30209 9781 30243
rect 9781 30209 9815 30243
rect 9815 30209 9824 30243
rect 9772 30200 9824 30209
rect 11152 30268 11204 30320
rect 11244 30268 11296 30320
rect 13176 30336 13228 30388
rect 12900 30268 12952 30320
rect 7380 30175 7432 30184
rect 7380 30141 7389 30175
rect 7389 30141 7423 30175
rect 7423 30141 7432 30175
rect 7380 30132 7432 30141
rect 8576 30132 8628 30184
rect 7748 29996 7800 30048
rect 8024 29996 8076 30048
rect 8760 30039 8812 30048
rect 8760 30005 8769 30039
rect 8769 30005 8803 30039
rect 8803 30005 8812 30039
rect 8760 29996 8812 30005
rect 9128 29996 9180 30048
rect 9496 29996 9548 30048
rect 9680 29996 9732 30048
rect 11520 30200 11572 30252
rect 11704 30243 11756 30252
rect 11704 30209 11713 30243
rect 11713 30209 11747 30243
rect 11747 30209 11756 30243
rect 11704 30200 11756 30209
rect 12440 30200 12492 30252
rect 15108 30336 15160 30388
rect 20168 30336 20220 30388
rect 21180 30336 21232 30388
rect 13636 30243 13688 30252
rect 13636 30209 13645 30243
rect 13645 30209 13679 30243
rect 13679 30209 13688 30243
rect 13636 30200 13688 30209
rect 14832 30200 14884 30252
rect 15016 30200 15068 30252
rect 16212 30200 16264 30252
rect 16396 30200 16448 30252
rect 11796 30132 11848 30184
rect 10508 30064 10560 30116
rect 12624 30175 12676 30184
rect 12624 30141 12633 30175
rect 12633 30141 12667 30175
rect 12667 30141 12676 30175
rect 12624 30132 12676 30141
rect 12716 30175 12768 30184
rect 12716 30141 12725 30175
rect 12725 30141 12759 30175
rect 12759 30141 12768 30175
rect 12716 30132 12768 30141
rect 12808 30175 12860 30184
rect 12808 30141 12817 30175
rect 12817 30141 12851 30175
rect 12851 30141 12860 30175
rect 12808 30132 12860 30141
rect 13728 30132 13780 30184
rect 17592 30268 17644 30320
rect 20628 30268 20680 30320
rect 17040 30243 17092 30252
rect 17040 30209 17049 30243
rect 17049 30209 17083 30243
rect 17083 30209 17092 30243
rect 17040 30200 17092 30209
rect 17224 30243 17276 30252
rect 17224 30209 17233 30243
rect 17233 30209 17267 30243
rect 17267 30209 17276 30243
rect 17224 30200 17276 30209
rect 17316 30200 17368 30252
rect 19340 30200 19392 30252
rect 18328 30132 18380 30184
rect 18420 30175 18472 30184
rect 18420 30141 18429 30175
rect 18429 30141 18463 30175
rect 18463 30141 18472 30175
rect 18420 30132 18472 30141
rect 20904 30243 20956 30252
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 20904 30200 20956 30209
rect 21088 30200 21140 30252
rect 21272 30243 21324 30252
rect 21272 30209 21281 30243
rect 21281 30209 21315 30243
rect 21315 30209 21324 30243
rect 21272 30200 21324 30209
rect 21456 30268 21508 30320
rect 23756 30336 23808 30388
rect 26240 30336 26292 30388
rect 22192 30268 22244 30320
rect 22560 30268 22612 30320
rect 23112 30268 23164 30320
rect 21180 30132 21232 30184
rect 22008 30200 22060 30252
rect 22284 30243 22336 30252
rect 22284 30209 22293 30243
rect 22293 30209 22327 30243
rect 22327 30209 22336 30243
rect 22284 30200 22336 30209
rect 22468 30243 22520 30252
rect 22468 30209 22477 30243
rect 22477 30209 22511 30243
rect 22511 30209 22520 30243
rect 22468 30200 22520 30209
rect 24584 30311 24636 30320
rect 24584 30277 24593 30311
rect 24593 30277 24627 30311
rect 24627 30277 24636 30311
rect 24584 30268 24636 30277
rect 25044 30268 25096 30320
rect 25596 30268 25648 30320
rect 26056 30268 26108 30320
rect 26792 30268 26844 30320
rect 23480 30200 23532 30252
rect 24492 30200 24544 30252
rect 24860 30200 24912 30252
rect 27344 30336 27396 30388
rect 29828 30336 29880 30388
rect 30104 30336 30156 30388
rect 30196 30336 30248 30388
rect 34612 30336 34664 30388
rect 36084 30336 36136 30388
rect 38200 30336 38252 30388
rect 27068 30268 27120 30320
rect 27712 30268 27764 30320
rect 16488 30064 16540 30116
rect 10876 29996 10928 30048
rect 10968 30039 11020 30048
rect 10968 30005 10977 30039
rect 10977 30005 11011 30039
rect 11011 30005 11020 30039
rect 10968 29996 11020 30005
rect 11244 29996 11296 30048
rect 12348 30039 12400 30048
rect 12348 30005 12357 30039
rect 12357 30005 12391 30039
rect 12391 30005 12400 30039
rect 12348 29996 12400 30005
rect 13084 29996 13136 30048
rect 13820 30039 13872 30048
rect 13820 30005 13829 30039
rect 13829 30005 13863 30039
rect 13863 30005 13872 30039
rect 13820 29996 13872 30005
rect 15936 29996 15988 30048
rect 22008 30064 22060 30116
rect 23572 30132 23624 30184
rect 25596 30175 25648 30184
rect 25596 30141 25605 30175
rect 25605 30141 25639 30175
rect 25639 30141 25648 30175
rect 25596 30132 25648 30141
rect 28448 30200 28500 30252
rect 27344 30175 27396 30184
rect 22560 30064 22612 30116
rect 23112 30064 23164 30116
rect 25228 30064 25280 30116
rect 25320 30064 25372 30116
rect 25872 30107 25924 30116
rect 25872 30073 25881 30107
rect 25881 30073 25915 30107
rect 25915 30073 25924 30107
rect 25872 30064 25924 30073
rect 19708 30039 19760 30048
rect 19708 30005 19717 30039
rect 19717 30005 19751 30039
rect 19751 30005 19760 30039
rect 19708 29996 19760 30005
rect 21088 29996 21140 30048
rect 21456 29996 21508 30048
rect 22468 29996 22520 30048
rect 24584 29996 24636 30048
rect 25412 29996 25464 30048
rect 27344 30141 27353 30175
rect 27353 30141 27387 30175
rect 27387 30141 27396 30175
rect 27344 30132 27396 30141
rect 27712 30132 27764 30184
rect 28080 30132 28132 30184
rect 28172 30175 28224 30184
rect 28172 30141 28181 30175
rect 28181 30141 28215 30175
rect 28215 30141 28224 30175
rect 28172 30132 28224 30141
rect 26332 30064 26384 30116
rect 27804 30064 27856 30116
rect 30288 30200 30340 30252
rect 28632 30107 28684 30116
rect 28632 30073 28641 30107
rect 28641 30073 28675 30107
rect 28675 30073 28684 30107
rect 28632 30064 28684 30073
rect 27160 30039 27212 30048
rect 27160 30005 27169 30039
rect 27169 30005 27203 30039
rect 27203 30005 27212 30039
rect 27160 29996 27212 30005
rect 27344 29996 27396 30048
rect 27436 29996 27488 30048
rect 29092 30175 29144 30184
rect 29092 30141 29101 30175
rect 29101 30141 29135 30175
rect 29135 30141 29144 30175
rect 29092 30132 29144 30141
rect 29552 30132 29604 30184
rect 29828 30132 29880 30184
rect 30104 30107 30156 30116
rect 30104 30073 30113 30107
rect 30113 30073 30147 30107
rect 30147 30073 30156 30107
rect 30104 30064 30156 30073
rect 31668 30268 31720 30320
rect 34244 30268 34296 30320
rect 33232 30200 33284 30252
rect 33508 30243 33560 30252
rect 33508 30209 33517 30243
rect 33517 30209 33551 30243
rect 33551 30209 33560 30243
rect 33508 30200 33560 30209
rect 31760 30132 31812 30184
rect 31944 30132 31996 30184
rect 32956 30132 33008 30184
rect 33876 30243 33928 30252
rect 33876 30209 33885 30243
rect 33885 30209 33919 30243
rect 33919 30209 33928 30243
rect 33876 30200 33928 30209
rect 34152 30200 34204 30252
rect 34428 30200 34480 30252
rect 36728 30268 36780 30320
rect 37556 30268 37608 30320
rect 35348 30243 35400 30252
rect 35348 30209 35382 30243
rect 35382 30209 35400 30243
rect 35348 30200 35400 30209
rect 32312 30064 32364 30116
rect 33508 30064 33560 30116
rect 33692 30064 33744 30116
rect 38108 30175 38160 30184
rect 38108 30141 38117 30175
rect 38117 30141 38151 30175
rect 38151 30141 38160 30175
rect 38108 30132 38160 30141
rect 30196 29996 30248 30048
rect 30656 29996 30708 30048
rect 31208 30039 31260 30048
rect 31208 30005 31217 30039
rect 31217 30005 31251 30039
rect 31251 30005 31260 30039
rect 31208 29996 31260 30005
rect 31668 30039 31720 30048
rect 31668 30005 31677 30039
rect 31677 30005 31711 30039
rect 31711 30005 31720 30039
rect 31668 29996 31720 30005
rect 32128 29996 32180 30048
rect 32864 29996 32916 30048
rect 33140 29996 33192 30048
rect 34888 29996 34940 30048
rect 35808 29996 35860 30048
rect 36360 29996 36412 30048
rect 37464 30039 37516 30048
rect 37464 30005 37473 30039
rect 37473 30005 37507 30039
rect 37507 30005 37516 30039
rect 37464 29996 37516 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3976 29792 4028 29844
rect 4528 29792 4580 29844
rect 8116 29835 8168 29844
rect 8116 29801 8125 29835
rect 8125 29801 8159 29835
rect 8159 29801 8168 29835
rect 8116 29792 8168 29801
rect 8208 29792 8260 29844
rect 10416 29792 10468 29844
rect 9404 29724 9456 29776
rect 9496 29724 9548 29776
rect 11152 29724 11204 29776
rect 12716 29792 12768 29844
rect 13268 29792 13320 29844
rect 7196 29656 7248 29708
rect 7012 29631 7064 29640
rect 7012 29597 7021 29631
rect 7021 29597 7055 29631
rect 7055 29597 7064 29631
rect 7012 29588 7064 29597
rect 7104 29588 7156 29640
rect 7564 29656 7616 29708
rect 8760 29656 8812 29708
rect 9128 29699 9180 29708
rect 9128 29665 9137 29699
rect 9137 29665 9171 29699
rect 9171 29665 9180 29699
rect 9128 29656 9180 29665
rect 9588 29699 9640 29708
rect 9588 29665 9597 29699
rect 9597 29665 9631 29699
rect 9631 29665 9640 29699
rect 10508 29699 10560 29708
rect 9588 29656 9640 29665
rect 10508 29665 10517 29699
rect 10517 29665 10551 29699
rect 10551 29665 10560 29699
rect 10508 29656 10560 29665
rect 11980 29724 12032 29776
rect 12440 29724 12492 29776
rect 16028 29792 16080 29844
rect 16212 29835 16264 29844
rect 16212 29801 16221 29835
rect 16221 29801 16255 29835
rect 16255 29801 16264 29835
rect 16212 29792 16264 29801
rect 16488 29792 16540 29844
rect 15384 29724 15436 29776
rect 17040 29724 17092 29776
rect 18604 29724 18656 29776
rect 19708 29724 19760 29776
rect 20904 29724 20956 29776
rect 13636 29656 13688 29708
rect 8300 29631 8352 29640
rect 8300 29597 8309 29631
rect 8309 29597 8343 29631
rect 8343 29597 8352 29631
rect 8300 29588 8352 29597
rect 8484 29631 8536 29640
rect 8484 29597 8493 29631
rect 8493 29597 8527 29631
rect 8527 29597 8536 29631
rect 8484 29588 8536 29597
rect 9312 29588 9364 29640
rect 10140 29588 10192 29640
rect 10232 29631 10284 29640
rect 10232 29597 10241 29631
rect 10241 29597 10275 29631
rect 10275 29597 10284 29631
rect 10232 29588 10284 29597
rect 10692 29631 10744 29640
rect 10692 29597 10701 29631
rect 10701 29597 10735 29631
rect 10735 29597 10744 29631
rect 10692 29588 10744 29597
rect 12992 29588 13044 29640
rect 13728 29588 13780 29640
rect 14740 29588 14792 29640
rect 15936 29631 15988 29640
rect 15936 29597 15945 29631
rect 15945 29597 15979 29631
rect 15979 29597 15988 29631
rect 15936 29588 15988 29597
rect 16028 29631 16080 29640
rect 16028 29597 16037 29631
rect 16037 29597 16071 29631
rect 16071 29597 16080 29631
rect 16028 29588 16080 29597
rect 10876 29520 10928 29572
rect 11244 29520 11296 29572
rect 12256 29520 12308 29572
rect 12440 29563 12492 29572
rect 12440 29529 12449 29563
rect 12449 29529 12483 29563
rect 12483 29529 12492 29563
rect 12440 29520 12492 29529
rect 12624 29563 12676 29572
rect 12624 29529 12633 29563
rect 12633 29529 12667 29563
rect 12667 29529 12676 29563
rect 12624 29520 12676 29529
rect 13084 29520 13136 29572
rect 14280 29563 14332 29572
rect 14280 29529 14289 29563
rect 14289 29529 14323 29563
rect 14323 29529 14332 29563
rect 14280 29520 14332 29529
rect 15016 29563 15068 29572
rect 15016 29529 15025 29563
rect 15025 29529 15059 29563
rect 15059 29529 15068 29563
rect 15016 29520 15068 29529
rect 15476 29520 15528 29572
rect 16396 29520 16448 29572
rect 16948 29588 17000 29640
rect 17316 29588 17368 29640
rect 17960 29588 18012 29640
rect 19156 29588 19208 29640
rect 17592 29520 17644 29572
rect 8208 29452 8260 29504
rect 8668 29452 8720 29504
rect 9772 29495 9824 29504
rect 9772 29461 9781 29495
rect 9781 29461 9815 29495
rect 9815 29461 9824 29495
rect 9772 29452 9824 29461
rect 12716 29452 12768 29504
rect 13452 29452 13504 29504
rect 13728 29452 13780 29504
rect 16856 29452 16908 29504
rect 18972 29452 19024 29504
rect 19340 29520 19392 29572
rect 20260 29563 20312 29572
rect 20260 29529 20269 29563
rect 20269 29529 20303 29563
rect 20303 29529 20312 29563
rect 20260 29520 20312 29529
rect 21548 29724 21600 29776
rect 22652 29724 22704 29776
rect 24492 29792 24544 29844
rect 27068 29792 27120 29844
rect 27344 29835 27396 29844
rect 27344 29801 27353 29835
rect 27353 29801 27387 29835
rect 27387 29801 27396 29835
rect 27344 29792 27396 29801
rect 28172 29792 28224 29844
rect 29828 29792 29880 29844
rect 30288 29835 30340 29844
rect 30288 29801 30297 29835
rect 30297 29801 30331 29835
rect 30331 29801 30340 29835
rect 30288 29792 30340 29801
rect 30472 29792 30524 29844
rect 34520 29792 34572 29844
rect 34980 29835 35032 29844
rect 34980 29801 34989 29835
rect 34989 29801 35023 29835
rect 35023 29801 35032 29835
rect 34980 29792 35032 29801
rect 36084 29792 36136 29844
rect 36452 29792 36504 29844
rect 21916 29699 21968 29708
rect 21916 29665 21925 29699
rect 21925 29665 21959 29699
rect 21959 29665 21968 29699
rect 21916 29656 21968 29665
rect 22008 29656 22060 29708
rect 25780 29724 25832 29776
rect 30564 29724 30616 29776
rect 21456 29588 21508 29640
rect 22192 29631 22244 29640
rect 22192 29597 22201 29631
rect 22201 29597 22235 29631
rect 22235 29597 22244 29631
rect 22192 29588 22244 29597
rect 23480 29631 23532 29640
rect 21640 29520 21692 29572
rect 23480 29597 23489 29631
rect 23489 29597 23523 29631
rect 23523 29597 23532 29631
rect 23480 29588 23532 29597
rect 23664 29631 23716 29640
rect 23664 29597 23673 29631
rect 23673 29597 23707 29631
rect 23707 29597 23716 29631
rect 23664 29588 23716 29597
rect 23756 29631 23808 29640
rect 23756 29597 23765 29631
rect 23765 29597 23799 29631
rect 23799 29597 23808 29631
rect 23756 29588 23808 29597
rect 23940 29631 23992 29640
rect 23940 29597 23949 29631
rect 23949 29597 23983 29631
rect 23983 29597 23992 29631
rect 23940 29588 23992 29597
rect 24768 29656 24820 29708
rect 25136 29656 25188 29708
rect 25228 29656 25280 29708
rect 25964 29656 26016 29708
rect 24860 29588 24912 29640
rect 25596 29588 25648 29640
rect 26976 29588 27028 29640
rect 26608 29563 26660 29572
rect 26608 29529 26617 29563
rect 26617 29529 26651 29563
rect 26651 29529 26660 29563
rect 26608 29520 26660 29529
rect 27252 29588 27304 29640
rect 30196 29656 30248 29708
rect 30380 29699 30432 29708
rect 30380 29665 30389 29699
rect 30389 29665 30423 29699
rect 30423 29665 30432 29699
rect 30380 29656 30432 29665
rect 33140 29724 33192 29776
rect 33324 29724 33376 29776
rect 32588 29656 32640 29708
rect 28172 29588 28224 29640
rect 28448 29588 28500 29640
rect 28724 29631 28776 29640
rect 28724 29597 28733 29631
rect 28733 29597 28767 29631
rect 28767 29597 28776 29631
rect 28724 29588 28776 29597
rect 28908 29588 28960 29640
rect 27160 29520 27212 29572
rect 27436 29520 27488 29572
rect 23296 29495 23348 29504
rect 23296 29461 23305 29495
rect 23305 29461 23339 29495
rect 23339 29461 23348 29495
rect 23296 29452 23348 29461
rect 23572 29452 23624 29504
rect 27712 29452 27764 29504
rect 27804 29495 27856 29504
rect 27804 29461 27813 29495
rect 27813 29461 27847 29495
rect 27847 29461 27856 29495
rect 27804 29452 27856 29461
rect 28632 29520 28684 29572
rect 29368 29588 29420 29640
rect 30564 29631 30616 29640
rect 30564 29597 30573 29631
rect 30573 29597 30607 29631
rect 30607 29597 30616 29631
rect 30564 29588 30616 29597
rect 31300 29631 31352 29640
rect 31300 29597 31309 29631
rect 31309 29597 31343 29631
rect 31343 29597 31352 29631
rect 31300 29588 31352 29597
rect 31392 29588 31444 29640
rect 32312 29588 32364 29640
rect 33692 29656 33744 29708
rect 34612 29724 34664 29776
rect 38200 29835 38252 29844
rect 38200 29801 38209 29835
rect 38209 29801 38243 29835
rect 38243 29801 38252 29835
rect 38200 29792 38252 29801
rect 34796 29656 34848 29708
rect 38292 29724 38344 29776
rect 35532 29656 35584 29708
rect 29184 29520 29236 29572
rect 29828 29520 29880 29572
rect 30104 29563 30156 29572
rect 30104 29529 30113 29563
rect 30113 29529 30147 29563
rect 30147 29529 30156 29563
rect 30104 29520 30156 29529
rect 30656 29520 30708 29572
rect 30748 29520 30800 29572
rect 33876 29588 33928 29640
rect 34428 29588 34480 29640
rect 35716 29631 35768 29640
rect 35716 29597 35725 29631
rect 35725 29597 35759 29631
rect 35759 29597 35768 29631
rect 35716 29588 35768 29597
rect 36360 29656 36412 29708
rect 36544 29588 36596 29640
rect 36636 29588 36688 29640
rect 36912 29588 36964 29640
rect 37464 29588 37516 29640
rect 29736 29495 29788 29504
rect 29736 29461 29745 29495
rect 29745 29461 29779 29495
rect 29779 29461 29788 29495
rect 29736 29452 29788 29461
rect 30472 29452 30524 29504
rect 31484 29452 31536 29504
rect 33232 29452 33284 29504
rect 34704 29520 34756 29572
rect 33692 29495 33744 29504
rect 33692 29461 33701 29495
rect 33701 29461 33735 29495
rect 33735 29461 33744 29495
rect 33692 29452 33744 29461
rect 34612 29452 34664 29504
rect 36176 29452 36228 29504
rect 36360 29495 36412 29504
rect 36360 29461 36369 29495
rect 36369 29461 36403 29495
rect 36403 29461 36412 29495
rect 36360 29452 36412 29461
rect 37556 29520 37608 29572
rect 36544 29452 36596 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 7472 29291 7524 29300
rect 7472 29257 7481 29291
rect 7481 29257 7515 29291
rect 7515 29257 7524 29291
rect 7472 29248 7524 29257
rect 8116 29291 8168 29300
rect 8116 29257 8125 29291
rect 8125 29257 8159 29291
rect 8159 29257 8168 29291
rect 8116 29248 8168 29257
rect 8392 29248 8444 29300
rect 9588 29248 9640 29300
rect 9680 29248 9732 29300
rect 12716 29248 12768 29300
rect 7380 29180 7432 29232
rect 13912 29248 13964 29300
rect 14832 29248 14884 29300
rect 7564 29112 7616 29164
rect 7932 29155 7984 29164
rect 7932 29121 7941 29155
rect 7941 29121 7975 29155
rect 7975 29121 7984 29155
rect 7932 29112 7984 29121
rect 8208 29112 8260 29164
rect 8392 29044 8444 29096
rect 4620 28976 4672 29028
rect 7012 28976 7064 29028
rect 4528 28908 4580 28960
rect 7196 28908 7248 28960
rect 7840 28908 7892 28960
rect 8760 29155 8812 29164
rect 8760 29121 8769 29155
rect 8769 29121 8803 29155
rect 8803 29121 8812 29155
rect 8760 29112 8812 29121
rect 8852 29112 8904 29164
rect 9772 29112 9824 29164
rect 10416 29155 10468 29164
rect 10416 29121 10425 29155
rect 10425 29121 10459 29155
rect 10459 29121 10468 29155
rect 10416 29112 10468 29121
rect 10600 29112 10652 29164
rect 10784 29112 10836 29164
rect 11704 29112 11756 29164
rect 9220 29087 9272 29096
rect 9220 29053 9229 29087
rect 9229 29053 9263 29087
rect 9263 29053 9272 29087
rect 9220 29044 9272 29053
rect 9404 29087 9456 29096
rect 9404 29053 9413 29087
rect 9413 29053 9447 29087
rect 9447 29053 9456 29087
rect 9404 29044 9456 29053
rect 9588 29087 9640 29096
rect 8668 29019 8720 29028
rect 8668 28985 8677 29019
rect 8677 28985 8711 29019
rect 8711 28985 8720 29019
rect 8668 28976 8720 28985
rect 8852 28976 8904 29028
rect 8944 28976 8996 29028
rect 9588 29053 9597 29087
rect 9597 29053 9631 29087
rect 9631 29053 9640 29087
rect 9588 29044 9640 29053
rect 11520 29044 11572 29096
rect 12624 29044 12676 29096
rect 13268 29112 13320 29164
rect 15016 29180 15068 29232
rect 17776 29248 17828 29300
rect 17040 29180 17092 29232
rect 14740 29112 14792 29164
rect 15568 29112 15620 29164
rect 16028 29112 16080 29164
rect 16856 29155 16908 29164
rect 16856 29121 16865 29155
rect 16865 29121 16899 29155
rect 16899 29121 16908 29155
rect 16856 29112 16908 29121
rect 17132 29112 17184 29164
rect 18512 29112 18564 29164
rect 20260 29180 20312 29232
rect 19248 29112 19300 29164
rect 20720 29248 20772 29300
rect 21272 29248 21324 29300
rect 22468 29291 22520 29300
rect 22468 29257 22477 29291
rect 22477 29257 22511 29291
rect 22511 29257 22520 29291
rect 22468 29248 22520 29257
rect 22928 29248 22980 29300
rect 24584 29248 24636 29300
rect 24768 29248 24820 29300
rect 24952 29248 25004 29300
rect 26424 29248 26476 29300
rect 26608 29248 26660 29300
rect 21272 29112 21324 29164
rect 22100 29112 22152 29164
rect 22376 29155 22428 29164
rect 22376 29121 22385 29155
rect 22385 29121 22419 29155
rect 22419 29121 22428 29155
rect 22376 29112 22428 29121
rect 9680 28976 9732 29028
rect 10508 28976 10560 29028
rect 11980 28976 12032 29028
rect 13084 28976 13136 29028
rect 17224 29044 17276 29096
rect 20996 29044 21048 29096
rect 23480 29044 23532 29096
rect 9864 28908 9916 28960
rect 10416 28908 10468 28960
rect 10968 28908 11020 28960
rect 15016 28951 15068 28960
rect 15016 28917 15025 28951
rect 15025 28917 15059 28951
rect 15059 28917 15068 28951
rect 15016 28908 15068 28917
rect 15200 28908 15252 28960
rect 15936 28908 15988 28960
rect 18604 29019 18656 29028
rect 18604 28985 18613 29019
rect 18613 28985 18647 29019
rect 18647 28985 18656 29019
rect 18604 28976 18656 28985
rect 23756 28976 23808 29028
rect 24216 29155 24268 29164
rect 24216 29121 24225 29155
rect 24225 29121 24259 29155
rect 24259 29121 24268 29155
rect 24216 29112 24268 29121
rect 24860 29155 24912 29164
rect 24860 29121 24869 29155
rect 24869 29121 24903 29155
rect 24903 29121 24912 29155
rect 24860 29112 24912 29121
rect 25688 29223 25740 29232
rect 25688 29189 25697 29223
rect 25697 29189 25731 29223
rect 25731 29189 25740 29223
rect 25688 29180 25740 29189
rect 25044 29155 25096 29164
rect 25044 29121 25053 29155
rect 25053 29121 25087 29155
rect 25087 29121 25096 29155
rect 25044 29112 25096 29121
rect 25504 29112 25556 29164
rect 27896 29180 27948 29232
rect 26884 29112 26936 29164
rect 27068 29112 27120 29164
rect 27344 29155 27396 29164
rect 27344 29121 27353 29155
rect 27353 29121 27387 29155
rect 27387 29121 27396 29155
rect 27344 29112 27396 29121
rect 28172 29155 28224 29164
rect 28172 29121 28181 29155
rect 28181 29121 28215 29155
rect 28215 29121 28224 29155
rect 28172 29112 28224 29121
rect 28264 29112 28316 29164
rect 26240 29087 26292 29096
rect 26240 29053 26249 29087
rect 26249 29053 26283 29087
rect 26283 29053 26292 29087
rect 29276 29248 29328 29300
rect 29184 29180 29236 29232
rect 29368 29155 29420 29164
rect 29368 29121 29377 29155
rect 29377 29121 29411 29155
rect 29411 29121 29420 29155
rect 29368 29112 29420 29121
rect 31944 29248 31996 29300
rect 32680 29248 32732 29300
rect 33232 29248 33284 29300
rect 29828 29180 29880 29232
rect 30472 29155 30524 29164
rect 30472 29121 30481 29155
rect 30481 29121 30515 29155
rect 30515 29121 30524 29155
rect 30472 29112 30524 29121
rect 30564 29155 30616 29164
rect 30564 29121 30573 29155
rect 30573 29121 30607 29155
rect 30607 29121 30616 29155
rect 30564 29112 30616 29121
rect 30656 29155 30708 29164
rect 30656 29121 30665 29155
rect 30665 29121 30699 29155
rect 30699 29121 30708 29155
rect 30656 29112 30708 29121
rect 30932 29180 30984 29232
rect 33048 29223 33100 29232
rect 33048 29189 33057 29223
rect 33057 29189 33091 29223
rect 33091 29189 33100 29223
rect 33048 29180 33100 29189
rect 31300 29155 31352 29164
rect 31300 29121 31309 29155
rect 31309 29121 31343 29155
rect 31343 29121 31352 29155
rect 31300 29112 31352 29121
rect 32772 29112 32824 29164
rect 26240 29044 26292 29053
rect 16396 28908 16448 28960
rect 16672 28908 16724 28960
rect 17684 28908 17736 28960
rect 20076 28908 20128 28960
rect 22008 28951 22060 28960
rect 22008 28917 22017 28951
rect 22017 28917 22051 28951
rect 22051 28917 22060 28951
rect 22008 28908 22060 28917
rect 22284 28908 22336 28960
rect 23664 28908 23716 28960
rect 25688 28976 25740 29028
rect 31024 29044 31076 29096
rect 31484 29044 31536 29096
rect 33876 29248 33928 29300
rect 33508 29180 33560 29232
rect 34244 29248 34296 29300
rect 34060 29223 34112 29232
rect 34060 29189 34069 29223
rect 34069 29189 34103 29223
rect 34103 29189 34112 29223
rect 34060 29180 34112 29189
rect 33692 29155 33744 29164
rect 33692 29121 33701 29155
rect 33701 29121 33735 29155
rect 33735 29121 33744 29155
rect 33692 29112 33744 29121
rect 34152 29155 34204 29164
rect 34152 29121 34166 29155
rect 34166 29121 34200 29155
rect 34200 29121 34204 29155
rect 34152 29112 34204 29121
rect 34244 29044 34296 29096
rect 35532 29248 35584 29300
rect 36360 29248 36412 29300
rect 35072 29155 35124 29164
rect 35072 29121 35081 29155
rect 35081 29121 35115 29155
rect 35115 29121 35124 29155
rect 35072 29112 35124 29121
rect 36452 29180 36504 29232
rect 37188 29180 37240 29232
rect 38200 29180 38252 29232
rect 34520 29044 34572 29096
rect 34888 29044 34940 29096
rect 35716 29112 35768 29164
rect 35992 29155 36044 29164
rect 35992 29121 36001 29155
rect 36001 29121 36035 29155
rect 36035 29121 36044 29155
rect 35992 29112 36044 29121
rect 35900 29044 35952 29096
rect 37924 29044 37976 29096
rect 38108 29087 38160 29096
rect 38108 29053 38117 29087
rect 38117 29053 38151 29087
rect 38151 29053 38160 29087
rect 38108 29044 38160 29053
rect 30564 28976 30616 29028
rect 33692 28976 33744 29028
rect 35440 28976 35492 29028
rect 26516 28908 26568 28960
rect 27068 28908 27120 28960
rect 27344 28908 27396 28960
rect 27896 28908 27948 28960
rect 29276 28908 29328 28960
rect 29368 28908 29420 28960
rect 30472 28908 30524 28960
rect 31208 28908 31260 28960
rect 32772 28908 32824 28960
rect 35716 28908 35768 28960
rect 35992 28908 36044 28960
rect 37464 28951 37516 28960
rect 37464 28917 37473 28951
rect 37473 28917 37507 28951
rect 37507 28917 37516 28951
rect 37464 28908 37516 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 5816 28704 5868 28756
rect 7104 28500 7156 28552
rect 9312 28543 9364 28552
rect 9312 28509 9321 28543
rect 9321 28509 9355 28543
rect 9355 28509 9364 28543
rect 9312 28500 9364 28509
rect 10600 28636 10652 28688
rect 10692 28679 10744 28688
rect 10692 28645 10701 28679
rect 10701 28645 10735 28679
rect 10735 28645 10744 28679
rect 10692 28636 10744 28645
rect 9772 28568 9824 28620
rect 9864 28500 9916 28552
rect 8024 28432 8076 28484
rect 9772 28432 9824 28484
rect 12532 28568 12584 28620
rect 14372 28704 14424 28756
rect 15016 28704 15068 28756
rect 18880 28704 18932 28756
rect 24216 28704 24268 28756
rect 24308 28704 24360 28756
rect 26056 28704 26108 28756
rect 10048 28500 10100 28552
rect 8392 28364 8444 28416
rect 9128 28407 9180 28416
rect 9128 28373 9137 28407
rect 9137 28373 9171 28407
rect 9171 28373 9180 28407
rect 9128 28364 9180 28373
rect 10784 28543 10836 28552
rect 10784 28509 10793 28543
rect 10793 28509 10827 28543
rect 10827 28509 10836 28543
rect 10784 28500 10836 28509
rect 10968 28500 11020 28552
rect 10692 28432 10744 28484
rect 11520 28500 11572 28552
rect 12256 28500 12308 28552
rect 12348 28500 12400 28552
rect 12716 28543 12768 28552
rect 12716 28509 12725 28543
rect 12725 28509 12759 28543
rect 12759 28509 12768 28543
rect 12716 28500 12768 28509
rect 15200 28636 15252 28688
rect 17040 28679 17092 28688
rect 17040 28645 17049 28679
rect 17049 28645 17083 28679
rect 17083 28645 17092 28679
rect 17040 28636 17092 28645
rect 17684 28636 17736 28688
rect 21732 28636 21784 28688
rect 24584 28636 24636 28688
rect 26976 28747 27028 28756
rect 26976 28713 26985 28747
rect 26985 28713 27019 28747
rect 27019 28713 27028 28747
rect 26976 28704 27028 28713
rect 27068 28747 27120 28756
rect 27068 28713 27077 28747
rect 27077 28713 27111 28747
rect 27111 28713 27120 28747
rect 27068 28704 27120 28713
rect 27804 28636 27856 28688
rect 14188 28500 14240 28552
rect 14280 28543 14332 28552
rect 14280 28509 14289 28543
rect 14289 28509 14323 28543
rect 14323 28509 14332 28543
rect 14280 28500 14332 28509
rect 18144 28611 18196 28620
rect 18144 28577 18153 28611
rect 18153 28577 18187 28611
rect 18187 28577 18196 28611
rect 18144 28568 18196 28577
rect 19984 28568 20036 28620
rect 21824 28568 21876 28620
rect 15936 28543 15988 28552
rect 15936 28509 15970 28543
rect 15970 28509 15988 28543
rect 15936 28500 15988 28509
rect 17868 28500 17920 28552
rect 18236 28500 18288 28552
rect 18880 28500 18932 28552
rect 21088 28500 21140 28552
rect 11428 28432 11480 28484
rect 12808 28432 12860 28484
rect 13728 28475 13780 28484
rect 13728 28441 13737 28475
rect 13737 28441 13771 28475
rect 13771 28441 13780 28475
rect 13728 28432 13780 28441
rect 15292 28432 15344 28484
rect 16120 28432 16172 28484
rect 21732 28500 21784 28552
rect 24032 28568 24084 28620
rect 22192 28543 22244 28552
rect 22192 28509 22201 28543
rect 22201 28509 22235 28543
rect 22235 28509 22244 28543
rect 22192 28500 22244 28509
rect 22652 28543 22704 28552
rect 22652 28509 22661 28543
rect 22661 28509 22695 28543
rect 22695 28509 22704 28543
rect 22652 28500 22704 28509
rect 22928 28543 22980 28552
rect 22928 28509 22937 28543
rect 22937 28509 22971 28543
rect 22971 28509 22980 28543
rect 22928 28500 22980 28509
rect 23848 28543 23900 28552
rect 23848 28509 23857 28543
rect 23857 28509 23891 28543
rect 23891 28509 23900 28543
rect 23848 28500 23900 28509
rect 24584 28543 24636 28552
rect 24584 28509 24593 28543
rect 24593 28509 24627 28543
rect 24627 28509 24636 28543
rect 24584 28500 24636 28509
rect 25412 28500 25464 28552
rect 26240 28568 26292 28620
rect 26424 28568 26476 28620
rect 28264 28568 28316 28620
rect 11060 28364 11112 28416
rect 11704 28364 11756 28416
rect 12348 28364 12400 28416
rect 13452 28407 13504 28416
rect 13452 28373 13461 28407
rect 13461 28373 13495 28407
rect 13495 28373 13504 28407
rect 13452 28364 13504 28373
rect 13544 28364 13596 28416
rect 16580 28364 16632 28416
rect 17500 28407 17552 28416
rect 17500 28373 17509 28407
rect 17509 28373 17543 28407
rect 17543 28373 17552 28407
rect 17500 28364 17552 28373
rect 17592 28364 17644 28416
rect 20536 28364 20588 28416
rect 20812 28407 20864 28416
rect 20812 28373 20821 28407
rect 20821 28373 20855 28407
rect 20855 28373 20864 28407
rect 20812 28364 20864 28373
rect 21456 28364 21508 28416
rect 22560 28432 22612 28484
rect 23388 28475 23440 28484
rect 23388 28441 23397 28475
rect 23397 28441 23431 28475
rect 23431 28441 23440 28475
rect 23388 28432 23440 28441
rect 23480 28432 23532 28484
rect 24768 28432 24820 28484
rect 25688 28432 25740 28484
rect 25872 28475 25924 28484
rect 25872 28441 25881 28475
rect 25881 28441 25915 28475
rect 25915 28441 25924 28475
rect 25872 28432 25924 28441
rect 26148 28543 26200 28552
rect 26148 28509 26157 28543
rect 26157 28509 26191 28543
rect 26191 28509 26200 28543
rect 26148 28500 26200 28509
rect 27160 28543 27212 28552
rect 27160 28509 27169 28543
rect 27169 28509 27203 28543
rect 27203 28509 27212 28543
rect 27160 28500 27212 28509
rect 27528 28500 27580 28552
rect 30380 28704 30432 28756
rect 31024 28704 31076 28756
rect 31484 28704 31536 28756
rect 33048 28704 33100 28756
rect 33508 28747 33560 28756
rect 33508 28713 33517 28747
rect 33517 28713 33551 28747
rect 33551 28713 33560 28747
rect 33508 28704 33560 28713
rect 33876 28704 33928 28756
rect 32956 28636 33008 28688
rect 33692 28636 33744 28688
rect 36084 28704 36136 28756
rect 38200 28747 38252 28756
rect 38200 28713 38209 28747
rect 38209 28713 38243 28747
rect 38243 28713 38252 28747
rect 38200 28704 38252 28713
rect 29184 28611 29236 28620
rect 29184 28577 29193 28611
rect 29193 28577 29227 28611
rect 29227 28577 29236 28611
rect 29184 28568 29236 28577
rect 29276 28568 29328 28620
rect 31300 28568 31352 28620
rect 27804 28432 27856 28484
rect 21640 28364 21692 28416
rect 23572 28364 23624 28416
rect 25412 28364 25464 28416
rect 25964 28364 26016 28416
rect 30380 28500 30432 28552
rect 30656 28543 30708 28552
rect 30656 28509 30665 28543
rect 30665 28509 30699 28543
rect 30699 28509 30708 28543
rect 34888 28611 34940 28620
rect 34888 28577 34897 28611
rect 34897 28577 34931 28611
rect 34931 28577 34940 28611
rect 34888 28568 34940 28577
rect 30656 28500 30708 28509
rect 28908 28432 28960 28484
rect 31668 28500 31720 28552
rect 33692 28500 33744 28552
rect 37464 28500 37516 28552
rect 32680 28432 32732 28484
rect 28816 28364 28868 28416
rect 31024 28364 31076 28416
rect 33692 28364 33744 28416
rect 34244 28364 34296 28416
rect 38384 28432 38436 28484
rect 35716 28364 35768 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 8024 28203 8076 28212
rect 8024 28169 8033 28203
rect 8033 28169 8067 28203
rect 8067 28169 8076 28203
rect 8024 28160 8076 28169
rect 9128 28160 9180 28212
rect 10140 28160 10192 28212
rect 10784 28160 10836 28212
rect 12716 28160 12768 28212
rect 8300 28092 8352 28144
rect 8392 28067 8444 28076
rect 8392 28033 8401 28067
rect 8401 28033 8435 28067
rect 8435 28033 8444 28067
rect 8392 28024 8444 28033
rect 8484 27956 8536 28008
rect 10508 28092 10560 28144
rect 10048 28067 10100 28076
rect 10048 28033 10057 28067
rect 10057 28033 10091 28067
rect 10091 28033 10100 28067
rect 10048 28024 10100 28033
rect 10876 28067 10928 28076
rect 10876 28033 10885 28067
rect 10885 28033 10919 28067
rect 10919 28033 10928 28067
rect 10876 28024 10928 28033
rect 14188 28092 14240 28144
rect 12072 28067 12124 28076
rect 12072 28033 12095 28067
rect 12095 28033 12124 28067
rect 10140 27956 10192 28008
rect 10692 27956 10744 28008
rect 12072 28024 12124 28033
rect 12164 28067 12216 28076
rect 12164 28033 12173 28067
rect 12173 28033 12207 28067
rect 12207 28033 12216 28067
rect 12164 28024 12216 28033
rect 12256 28067 12308 28076
rect 12256 28033 12265 28067
rect 12265 28033 12299 28067
rect 12299 28033 12308 28067
rect 12256 28024 12308 28033
rect 12440 28067 12492 28076
rect 12440 28033 12449 28067
rect 12449 28033 12483 28067
rect 12483 28033 12492 28067
rect 12440 28024 12492 28033
rect 13176 28067 13228 28076
rect 13176 28033 13210 28067
rect 13210 28033 13228 28067
rect 13176 28024 13228 28033
rect 13636 28024 13688 28076
rect 15568 28135 15620 28144
rect 12900 27999 12952 28008
rect 12900 27965 12909 27999
rect 12909 27965 12943 27999
rect 12943 27965 12952 27999
rect 12900 27956 12952 27965
rect 15568 28101 15577 28135
rect 15577 28101 15611 28135
rect 15611 28101 15620 28135
rect 15568 28092 15620 28101
rect 17132 28092 17184 28144
rect 20720 28160 20772 28212
rect 21088 28160 21140 28212
rect 21548 28160 21600 28212
rect 22008 28160 22060 28212
rect 23204 28160 23256 28212
rect 15016 28024 15068 28076
rect 15384 28067 15436 28076
rect 15384 28033 15393 28067
rect 15393 28033 15427 28067
rect 15427 28033 15436 28067
rect 15384 28024 15436 28033
rect 16028 28024 16080 28076
rect 16856 28067 16908 28076
rect 16856 28033 16865 28067
rect 16865 28033 16899 28067
rect 16899 28033 16908 28067
rect 16856 28024 16908 28033
rect 17316 28024 17368 28076
rect 18328 28024 18380 28076
rect 17684 27956 17736 28008
rect 18880 27956 18932 28008
rect 19156 27999 19208 28008
rect 19156 27965 19165 27999
rect 19165 27965 19199 27999
rect 19199 27965 19208 27999
rect 19156 27956 19208 27965
rect 20076 28024 20128 28076
rect 21088 28067 21140 28076
rect 19524 27956 19576 28008
rect 21088 28033 21097 28067
rect 21097 28033 21131 28067
rect 21131 28033 21140 28067
rect 21088 28024 21140 28033
rect 21364 28024 21416 28076
rect 22928 28024 22980 28076
rect 22100 27956 22152 28008
rect 7564 27888 7616 27940
rect 9772 27888 9824 27940
rect 10048 27888 10100 27940
rect 12532 27888 12584 27940
rect 14096 27888 14148 27940
rect 16856 27888 16908 27940
rect 19892 27888 19944 27940
rect 21364 27931 21416 27940
rect 21364 27897 21373 27931
rect 21373 27897 21407 27931
rect 21407 27897 21416 27931
rect 21364 27888 21416 27897
rect 22744 27956 22796 28008
rect 23296 28092 23348 28144
rect 23480 28024 23532 28076
rect 23572 28067 23624 28076
rect 23572 28033 23581 28067
rect 23581 28033 23615 28067
rect 23615 28033 23624 28067
rect 23572 28024 23624 28033
rect 24124 28160 24176 28212
rect 25596 28160 25648 28212
rect 23848 28092 23900 28144
rect 24860 28024 24912 28076
rect 25320 28024 25372 28076
rect 25412 28067 25464 28076
rect 25412 28033 25421 28067
rect 25421 28033 25455 28067
rect 25455 28033 25464 28067
rect 25412 28024 25464 28033
rect 26056 28092 26108 28144
rect 27528 28160 27580 28212
rect 28632 28160 28684 28212
rect 30564 28160 30616 28212
rect 25504 27956 25556 28008
rect 27160 28024 27212 28076
rect 28724 28092 28776 28144
rect 31668 28092 31720 28144
rect 31852 28092 31904 28144
rect 28172 28024 28224 28076
rect 28540 28024 28592 28076
rect 29000 28067 29052 28076
rect 29000 28033 29009 28067
rect 29009 28033 29043 28067
rect 29043 28033 29052 28067
rect 29000 28024 29052 28033
rect 29092 28024 29144 28076
rect 9588 27863 9640 27872
rect 9588 27829 9597 27863
rect 9597 27829 9631 27863
rect 9631 27829 9640 27863
rect 9588 27820 9640 27829
rect 10140 27820 10192 27872
rect 12716 27820 12768 27872
rect 15108 27820 15160 27872
rect 15936 27863 15988 27872
rect 15936 27829 15945 27863
rect 15945 27829 15979 27863
rect 15979 27829 15988 27863
rect 15936 27820 15988 27829
rect 18328 27820 18380 27872
rect 18420 27820 18472 27872
rect 18696 27820 18748 27872
rect 23020 27888 23072 27940
rect 22008 27863 22060 27872
rect 22008 27829 22017 27863
rect 22017 27829 22051 27863
rect 22051 27829 22060 27863
rect 22008 27820 22060 27829
rect 23204 27863 23256 27872
rect 23204 27829 23213 27863
rect 23213 27829 23247 27863
rect 23247 27829 23256 27863
rect 23204 27820 23256 27829
rect 23480 27931 23532 27940
rect 23480 27897 23489 27931
rect 23489 27897 23523 27931
rect 23523 27897 23532 27931
rect 23480 27888 23532 27897
rect 25596 27888 25648 27940
rect 26056 27956 26108 28008
rect 26148 27956 26200 28008
rect 27712 27956 27764 28008
rect 28264 27956 28316 28008
rect 30656 28067 30708 28076
rect 30656 28033 30665 28067
rect 30665 28033 30699 28067
rect 30699 28033 30708 28067
rect 30656 28024 30708 28033
rect 31576 28067 31628 28076
rect 31576 28033 31585 28067
rect 31585 28033 31619 28067
rect 31619 28033 31628 28067
rect 31576 28024 31628 28033
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 34796 28092 34848 28144
rect 30472 27956 30524 28008
rect 30840 27956 30892 28008
rect 32772 27956 32824 28008
rect 33876 28024 33928 28076
rect 34060 28067 34112 28076
rect 34060 28033 34069 28067
rect 34069 28033 34103 28067
rect 34103 28033 34112 28067
rect 34060 28024 34112 28033
rect 34152 28024 34204 28076
rect 34428 28024 34480 28076
rect 35348 28160 35400 28212
rect 37372 28092 37424 28144
rect 24492 27863 24544 27872
rect 24492 27829 24501 27863
rect 24501 27829 24535 27863
rect 24535 27829 24544 27863
rect 24492 27820 24544 27829
rect 24676 27820 24728 27872
rect 33324 27888 33376 27940
rect 35164 28024 35216 28076
rect 37464 28024 37516 28076
rect 38016 27999 38068 28008
rect 38016 27965 38025 27999
rect 38025 27965 38059 27999
rect 38059 27965 38068 27999
rect 38016 27956 38068 27965
rect 26148 27863 26200 27872
rect 26148 27829 26157 27863
rect 26157 27829 26191 27863
rect 26191 27829 26200 27863
rect 26148 27820 26200 27829
rect 26332 27820 26384 27872
rect 29644 27820 29696 27872
rect 29736 27820 29788 27872
rect 33508 27820 33560 27872
rect 34060 27820 34112 27872
rect 34428 27820 34480 27872
rect 34612 27820 34664 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4712 27616 4764 27668
rect 6920 27616 6972 27668
rect 9312 27616 9364 27668
rect 10048 27659 10100 27668
rect 10048 27625 10057 27659
rect 10057 27625 10091 27659
rect 10091 27625 10100 27659
rect 10048 27616 10100 27625
rect 3516 27548 3568 27600
rect 5356 27548 5408 27600
rect 7104 27523 7156 27532
rect 7104 27489 7113 27523
rect 7113 27489 7147 27523
rect 7147 27489 7156 27523
rect 7104 27480 7156 27489
rect 10692 27480 10744 27532
rect 8208 27412 8260 27464
rect 8576 27412 8628 27464
rect 9680 27412 9732 27464
rect 8024 27344 8076 27396
rect 10876 27412 10928 27464
rect 11060 27455 11112 27464
rect 11060 27421 11069 27455
rect 11069 27421 11103 27455
rect 11103 27421 11112 27455
rect 12256 27616 12308 27668
rect 12072 27548 12124 27600
rect 11704 27480 11756 27532
rect 11060 27412 11112 27421
rect 12348 27480 12400 27532
rect 12716 27616 12768 27668
rect 13084 27616 13136 27668
rect 13176 27616 13228 27668
rect 17868 27659 17920 27668
rect 17868 27625 17877 27659
rect 17877 27625 17911 27659
rect 17911 27625 17920 27659
rect 17868 27616 17920 27625
rect 19892 27616 19944 27668
rect 22192 27616 22244 27668
rect 23112 27659 23164 27668
rect 23112 27625 23121 27659
rect 23121 27625 23155 27659
rect 23155 27625 23164 27659
rect 23112 27616 23164 27625
rect 23296 27616 23348 27668
rect 23480 27616 23532 27668
rect 24492 27616 24544 27668
rect 26056 27616 26108 27668
rect 13360 27548 13412 27600
rect 14556 27548 14608 27600
rect 17132 27548 17184 27600
rect 12440 27412 12492 27464
rect 12716 27455 12768 27464
rect 12716 27421 12725 27455
rect 12725 27421 12759 27455
rect 12759 27421 12768 27455
rect 12716 27412 12768 27421
rect 12808 27412 12860 27464
rect 13084 27455 13136 27464
rect 13084 27421 13093 27455
rect 13093 27421 13127 27455
rect 13127 27421 13136 27455
rect 13084 27412 13136 27421
rect 13452 27412 13504 27464
rect 15568 27480 15620 27532
rect 18328 27523 18380 27532
rect 18328 27489 18337 27523
rect 18337 27489 18371 27523
rect 18371 27489 18380 27523
rect 18328 27480 18380 27489
rect 18420 27523 18472 27532
rect 18420 27489 18429 27523
rect 18429 27489 18463 27523
rect 18463 27489 18472 27523
rect 18420 27480 18472 27489
rect 20168 27480 20220 27532
rect 14556 27455 14608 27464
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 15200 27412 15252 27464
rect 15292 27412 15344 27464
rect 15660 27455 15712 27464
rect 15660 27421 15669 27455
rect 15669 27421 15703 27455
rect 15703 27421 15712 27455
rect 15660 27412 15712 27421
rect 15936 27455 15988 27464
rect 15936 27421 15970 27455
rect 15970 27421 15988 27455
rect 15936 27412 15988 27421
rect 16488 27412 16540 27464
rect 17960 27412 18012 27464
rect 18236 27412 18288 27464
rect 14096 27344 14148 27396
rect 8576 27276 8628 27328
rect 10416 27276 10468 27328
rect 11888 27276 11940 27328
rect 11980 27276 12032 27328
rect 19248 27344 19300 27396
rect 14832 27319 14884 27328
rect 14832 27285 14841 27319
rect 14841 27285 14875 27319
rect 14875 27285 14884 27319
rect 14832 27276 14884 27285
rect 18052 27276 18104 27328
rect 18696 27276 18748 27328
rect 19064 27276 19116 27328
rect 21272 27548 21324 27600
rect 22376 27548 22428 27600
rect 22008 27480 22060 27532
rect 23204 27480 23256 27532
rect 25872 27548 25924 27600
rect 26792 27616 26844 27668
rect 28356 27616 28408 27668
rect 28540 27616 28592 27668
rect 30564 27616 30616 27668
rect 34796 27616 34848 27668
rect 20444 27344 20496 27396
rect 22100 27412 22152 27464
rect 23020 27455 23072 27464
rect 23020 27421 23029 27455
rect 23029 27421 23063 27455
rect 23063 27421 23072 27455
rect 23020 27412 23072 27421
rect 23112 27455 23164 27464
rect 23112 27421 23121 27455
rect 23121 27421 23155 27455
rect 23155 27421 23164 27455
rect 23112 27412 23164 27421
rect 21548 27344 21600 27396
rect 23572 27344 23624 27396
rect 24032 27455 24084 27464
rect 24032 27421 24041 27455
rect 24041 27421 24075 27455
rect 24075 27421 24084 27455
rect 24032 27412 24084 27421
rect 24492 27480 24544 27532
rect 24400 27344 24452 27396
rect 24584 27387 24636 27396
rect 24584 27353 24593 27387
rect 24593 27353 24627 27387
rect 24627 27353 24636 27387
rect 24584 27344 24636 27353
rect 25320 27412 25372 27464
rect 26056 27480 26108 27532
rect 27344 27480 27396 27532
rect 26608 27412 26660 27464
rect 26240 27344 26292 27396
rect 26332 27387 26384 27396
rect 26332 27353 26366 27387
rect 26366 27353 26384 27387
rect 27896 27548 27948 27600
rect 28080 27548 28132 27600
rect 30012 27548 30064 27600
rect 30656 27548 30708 27600
rect 35992 27591 36044 27600
rect 35992 27557 36001 27591
rect 36001 27557 36035 27591
rect 36035 27557 36044 27591
rect 35992 27548 36044 27557
rect 27804 27480 27856 27532
rect 28724 27480 28776 27532
rect 28080 27412 28132 27464
rect 29184 27480 29236 27532
rect 32220 27523 32272 27532
rect 32220 27489 32229 27523
rect 32229 27489 32263 27523
rect 32263 27489 32272 27523
rect 32220 27480 32272 27489
rect 28908 27455 28960 27464
rect 28908 27421 28917 27455
rect 28917 27421 28951 27455
rect 28951 27421 28960 27455
rect 28908 27412 28960 27421
rect 29276 27412 29328 27464
rect 30012 27412 30064 27464
rect 30380 27455 30432 27464
rect 30380 27421 30389 27455
rect 30389 27421 30423 27455
rect 30423 27421 30432 27455
rect 30380 27412 30432 27421
rect 30564 27455 30616 27464
rect 30564 27421 30573 27455
rect 30573 27421 30607 27455
rect 30607 27421 30616 27455
rect 30564 27412 30616 27421
rect 26332 27344 26384 27353
rect 20720 27276 20772 27328
rect 21824 27319 21876 27328
rect 21824 27285 21833 27319
rect 21833 27285 21867 27319
rect 21867 27285 21876 27319
rect 21824 27276 21876 27285
rect 23480 27276 23532 27328
rect 25228 27319 25280 27328
rect 25228 27285 25237 27319
rect 25237 27285 25271 27319
rect 25271 27285 25280 27319
rect 25228 27276 25280 27285
rect 27252 27276 27304 27328
rect 28632 27319 28684 27328
rect 28632 27285 28641 27319
rect 28641 27285 28675 27319
rect 28675 27285 28684 27319
rect 28632 27276 28684 27285
rect 31024 27344 31076 27396
rect 31300 27344 31352 27396
rect 33140 27344 33192 27396
rect 33416 27412 33468 27464
rect 33692 27412 33744 27464
rect 34888 27455 34940 27464
rect 34888 27421 34897 27455
rect 34897 27421 34931 27455
rect 34931 27421 34940 27455
rect 34888 27412 34940 27421
rect 34428 27344 34480 27396
rect 34796 27344 34848 27396
rect 35072 27412 35124 27464
rect 35164 27387 35216 27396
rect 35164 27353 35173 27387
rect 35173 27353 35207 27387
rect 35207 27353 35216 27387
rect 35164 27344 35216 27353
rect 32772 27276 32824 27328
rect 33324 27276 33376 27328
rect 34520 27276 34572 27328
rect 36084 27344 36136 27396
rect 36636 27412 36688 27464
rect 36728 27455 36780 27464
rect 36728 27421 36737 27455
rect 36737 27421 36771 27455
rect 36771 27421 36780 27455
rect 36728 27412 36780 27421
rect 37464 27344 37516 27396
rect 35808 27276 35860 27328
rect 36636 27276 36688 27328
rect 38108 27319 38160 27328
rect 38108 27285 38117 27319
rect 38117 27285 38151 27319
rect 38151 27285 38160 27319
rect 38108 27276 38160 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 8024 27115 8076 27124
rect 8024 27081 8033 27115
rect 8033 27081 8067 27115
rect 8067 27081 8076 27115
rect 8024 27072 8076 27081
rect 9312 27072 9364 27124
rect 8576 27004 8628 27056
rect 11060 27004 11112 27056
rect 9588 26979 9640 26988
rect 9588 26945 9597 26979
rect 9597 26945 9631 26979
rect 9631 26945 9640 26979
rect 9588 26936 9640 26945
rect 9864 26979 9916 26988
rect 9864 26945 9873 26979
rect 9873 26945 9907 26979
rect 9907 26945 9916 26979
rect 9864 26936 9916 26945
rect 9956 26800 10008 26852
rect 10140 26868 10192 26920
rect 10508 26868 10560 26920
rect 10968 26936 11020 26988
rect 10876 26868 10928 26920
rect 12808 27004 12860 27056
rect 12992 27072 13044 27124
rect 13452 27072 13504 27124
rect 18144 27072 18196 27124
rect 19248 27072 19300 27124
rect 14832 27004 14884 27056
rect 13360 26936 13412 26988
rect 13452 26979 13504 26988
rect 13452 26945 13461 26979
rect 13461 26945 13495 26979
rect 13495 26945 13504 26979
rect 13452 26936 13504 26945
rect 14464 26936 14516 26988
rect 19340 27004 19392 27056
rect 16948 26979 17000 26988
rect 16948 26945 16957 26979
rect 16957 26945 16991 26979
rect 16991 26945 17000 26979
rect 16948 26936 17000 26945
rect 17500 26936 17552 26988
rect 17592 26936 17644 26988
rect 13176 26868 13228 26920
rect 13912 26911 13964 26920
rect 13912 26877 13921 26911
rect 13921 26877 13955 26911
rect 13955 26877 13964 26911
rect 13912 26868 13964 26877
rect 15384 26868 15436 26920
rect 16028 26868 16080 26920
rect 10140 26775 10192 26784
rect 10140 26741 10149 26775
rect 10149 26741 10183 26775
rect 10183 26741 10192 26775
rect 10140 26732 10192 26741
rect 10600 26732 10652 26784
rect 12256 26775 12308 26784
rect 12256 26741 12265 26775
rect 12265 26741 12299 26775
rect 12299 26741 12308 26775
rect 12256 26732 12308 26741
rect 13268 26775 13320 26784
rect 13268 26741 13277 26775
rect 13277 26741 13311 26775
rect 13311 26741 13320 26775
rect 13268 26732 13320 26741
rect 15200 26800 15252 26852
rect 14924 26732 14976 26784
rect 15292 26775 15344 26784
rect 15292 26741 15301 26775
rect 15301 26741 15335 26775
rect 15335 26741 15344 26775
rect 15292 26732 15344 26741
rect 15568 26732 15620 26784
rect 16120 26775 16172 26784
rect 16120 26741 16129 26775
rect 16129 26741 16163 26775
rect 16163 26741 16172 26775
rect 16120 26732 16172 26741
rect 18236 26732 18288 26784
rect 18604 26936 18656 26988
rect 18880 26936 18932 26988
rect 19064 26979 19116 26988
rect 19064 26945 19073 26979
rect 19073 26945 19107 26979
rect 19107 26945 19116 26979
rect 19064 26936 19116 26945
rect 19248 26936 19300 26988
rect 20076 27072 20128 27124
rect 20628 27047 20680 27056
rect 20628 27013 20637 27047
rect 20637 27013 20671 27047
rect 20671 27013 20680 27047
rect 20628 27004 20680 27013
rect 21364 27072 21416 27124
rect 22008 27072 22060 27124
rect 25228 27072 25280 27124
rect 21824 27004 21876 27056
rect 22468 26936 22520 26988
rect 19892 26868 19944 26920
rect 20536 26868 20588 26920
rect 20904 26911 20956 26920
rect 18512 26800 18564 26852
rect 20904 26877 20913 26911
rect 20913 26877 20947 26911
rect 20947 26877 20956 26911
rect 20904 26868 20956 26877
rect 21364 26868 21416 26920
rect 23296 26936 23348 26988
rect 23848 27004 23900 27056
rect 24124 27004 24176 27056
rect 24492 27004 24544 27056
rect 26424 27072 26476 27124
rect 27988 27072 28040 27124
rect 28080 27072 28132 27124
rect 26056 27004 26108 27056
rect 27712 27047 27764 27056
rect 27712 27013 27721 27047
rect 27721 27013 27755 27047
rect 27755 27013 27764 27047
rect 27712 27004 27764 27013
rect 27896 27004 27948 27056
rect 23756 26868 23808 26920
rect 25228 26936 25280 26988
rect 25596 26979 25648 26988
rect 25596 26945 25605 26979
rect 25605 26945 25639 26979
rect 25639 26945 25648 26979
rect 25596 26936 25648 26945
rect 26700 26936 26752 26988
rect 27252 26979 27304 26988
rect 27252 26945 27261 26979
rect 27261 26945 27295 26979
rect 27295 26945 27304 26979
rect 27252 26936 27304 26945
rect 28172 26936 28224 26988
rect 29000 27004 29052 27056
rect 29092 26936 29144 26988
rect 31024 26979 31076 26988
rect 31024 26945 31033 26979
rect 31033 26945 31067 26979
rect 31067 26945 31076 26979
rect 31024 26936 31076 26945
rect 34888 27072 34940 27124
rect 37096 27072 37148 27124
rect 37464 27115 37516 27124
rect 37464 27081 37473 27115
rect 37473 27081 37507 27115
rect 37507 27081 37516 27115
rect 37464 27072 37516 27081
rect 37740 27072 37792 27124
rect 27436 26868 27488 26920
rect 29000 26868 29052 26920
rect 30748 26868 30800 26920
rect 31116 26868 31168 26920
rect 31852 26936 31904 26988
rect 32404 26936 32456 26988
rect 32496 26936 32548 26988
rect 18880 26732 18932 26784
rect 20628 26732 20680 26784
rect 20812 26732 20864 26784
rect 25872 26800 25924 26852
rect 26884 26800 26936 26852
rect 29736 26800 29788 26852
rect 30012 26800 30064 26852
rect 32220 26868 32272 26920
rect 33416 26936 33468 26988
rect 33784 26979 33836 26988
rect 33784 26945 33793 26979
rect 33793 26945 33827 26979
rect 33827 26945 33836 26979
rect 33784 26936 33836 26945
rect 34612 27004 34664 27056
rect 35716 27004 35768 27056
rect 35808 27004 35860 27056
rect 34060 26979 34112 26988
rect 34060 26945 34069 26979
rect 34069 26945 34103 26979
rect 34103 26945 34112 26979
rect 34060 26936 34112 26945
rect 34980 26979 35032 26988
rect 34980 26945 34989 26979
rect 34989 26945 35023 26979
rect 35023 26945 35032 26979
rect 34980 26936 35032 26945
rect 35440 26936 35492 26988
rect 35900 26936 35952 26988
rect 36360 27004 36412 27056
rect 35808 26868 35860 26920
rect 33876 26800 33928 26852
rect 36360 26868 36412 26920
rect 23756 26775 23808 26784
rect 23756 26741 23765 26775
rect 23765 26741 23799 26775
rect 23799 26741 23808 26775
rect 23756 26732 23808 26741
rect 24492 26732 24544 26784
rect 24860 26732 24912 26784
rect 27436 26732 27488 26784
rect 30380 26732 30432 26784
rect 31852 26732 31904 26784
rect 32496 26732 32548 26784
rect 36636 26800 36688 26852
rect 34152 26732 34204 26784
rect 34428 26732 34480 26784
rect 34704 26732 34756 26784
rect 35808 26732 35860 26784
rect 38108 26936 38160 26988
rect 38016 26911 38068 26920
rect 38016 26877 38025 26911
rect 38025 26877 38059 26911
rect 38059 26877 38068 26911
rect 38016 26868 38068 26877
rect 38476 26868 38528 26920
rect 39120 26868 39172 26920
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 11336 26571 11388 26580
rect 11336 26537 11345 26571
rect 11345 26537 11379 26571
rect 11379 26537 11388 26571
rect 18512 26571 18564 26580
rect 11336 26528 11388 26537
rect 18512 26537 18521 26571
rect 18521 26537 18555 26571
rect 18555 26537 18564 26571
rect 18512 26528 18564 26537
rect 20260 26528 20312 26580
rect 13176 26503 13228 26512
rect 13176 26469 13185 26503
rect 13185 26469 13219 26503
rect 13219 26469 13228 26503
rect 13176 26460 13228 26469
rect 15200 26460 15252 26512
rect 15568 26460 15620 26512
rect 16856 26460 16908 26512
rect 8208 26392 8260 26444
rect 15660 26392 15712 26444
rect 17408 26392 17460 26444
rect 11704 26324 11756 26376
rect 12900 26324 12952 26376
rect 13912 26324 13964 26376
rect 14740 26367 14792 26376
rect 14740 26333 14749 26367
rect 14749 26333 14783 26367
rect 14783 26333 14792 26367
rect 14740 26324 14792 26333
rect 14832 26324 14884 26376
rect 10968 26256 11020 26308
rect 12256 26256 12308 26308
rect 12440 26256 12492 26308
rect 14464 26256 14516 26308
rect 14924 26299 14976 26308
rect 14924 26265 14933 26299
rect 14933 26265 14967 26299
rect 14967 26265 14976 26299
rect 14924 26256 14976 26265
rect 15200 26324 15252 26376
rect 15568 26324 15620 26376
rect 17776 26367 17828 26376
rect 17776 26333 17785 26367
rect 17785 26333 17819 26367
rect 17819 26333 17828 26367
rect 17776 26324 17828 26333
rect 17868 26367 17920 26376
rect 17868 26333 17877 26367
rect 17877 26333 17911 26367
rect 17911 26333 17920 26367
rect 17868 26324 17920 26333
rect 18052 26435 18104 26444
rect 18052 26401 18061 26435
rect 18061 26401 18095 26435
rect 18095 26401 18104 26435
rect 18052 26392 18104 26401
rect 18696 26392 18748 26444
rect 19340 26460 19392 26512
rect 18236 26324 18288 26376
rect 19340 26324 19392 26376
rect 20076 26324 20128 26376
rect 20536 26324 20588 26376
rect 16580 26256 16632 26308
rect 19892 26256 19944 26308
rect 21732 26392 21784 26444
rect 22652 26528 22704 26580
rect 25964 26528 26016 26580
rect 28080 26528 28132 26580
rect 28264 26528 28316 26580
rect 30472 26528 30524 26580
rect 30748 26528 30800 26580
rect 23572 26460 23624 26512
rect 23848 26503 23900 26512
rect 23848 26469 23857 26503
rect 23857 26469 23891 26503
rect 23891 26469 23900 26503
rect 23848 26460 23900 26469
rect 24584 26460 24636 26512
rect 26148 26392 26200 26444
rect 21640 26367 21692 26376
rect 21640 26333 21649 26367
rect 21649 26333 21683 26367
rect 21683 26333 21692 26367
rect 21640 26324 21692 26333
rect 5264 26188 5316 26240
rect 11060 26188 11112 26240
rect 11980 26188 12032 26240
rect 12532 26188 12584 26240
rect 12992 26188 13044 26240
rect 16488 26188 16540 26240
rect 17224 26188 17276 26240
rect 17868 26188 17920 26240
rect 18512 26188 18564 26240
rect 21456 26188 21508 26240
rect 23756 26324 23808 26376
rect 24676 26367 24728 26376
rect 24676 26333 24685 26367
rect 24685 26333 24719 26367
rect 24719 26333 24728 26367
rect 24676 26324 24728 26333
rect 24860 26367 24912 26376
rect 24860 26333 24869 26367
rect 24869 26333 24903 26367
rect 24903 26333 24912 26367
rect 24860 26324 24912 26333
rect 28080 26392 28132 26444
rect 30656 26460 30708 26512
rect 31024 26460 31076 26512
rect 32956 26528 33008 26580
rect 35808 26528 35860 26580
rect 36452 26571 36504 26580
rect 36452 26537 36461 26571
rect 36461 26537 36495 26571
rect 36495 26537 36504 26571
rect 36452 26528 36504 26537
rect 28264 26435 28316 26444
rect 28264 26401 28273 26435
rect 28273 26401 28307 26435
rect 28307 26401 28316 26435
rect 28264 26392 28316 26401
rect 28540 26392 28592 26444
rect 28816 26392 28868 26444
rect 28448 26324 28500 26376
rect 29184 26367 29236 26376
rect 29184 26333 29193 26367
rect 29193 26333 29227 26367
rect 29227 26333 29236 26367
rect 29184 26324 29236 26333
rect 29276 26324 29328 26376
rect 22468 26256 22520 26308
rect 23572 26256 23624 26308
rect 25136 26256 25188 26308
rect 25228 26299 25280 26308
rect 25228 26265 25237 26299
rect 25237 26265 25271 26299
rect 25271 26265 25280 26299
rect 25228 26256 25280 26265
rect 25872 26256 25924 26308
rect 26240 26256 26292 26308
rect 26332 26299 26384 26308
rect 26332 26265 26341 26299
rect 26341 26265 26375 26299
rect 26375 26265 26384 26299
rect 26332 26256 26384 26265
rect 26516 26299 26568 26308
rect 26516 26265 26525 26299
rect 26525 26265 26559 26299
rect 26559 26265 26568 26299
rect 26516 26256 26568 26265
rect 26976 26256 27028 26308
rect 27068 26256 27120 26308
rect 29736 26299 29788 26308
rect 29736 26265 29745 26299
rect 29745 26265 29779 26299
rect 29779 26265 29788 26299
rect 29736 26256 29788 26265
rect 33600 26392 33652 26444
rect 33784 26392 33836 26444
rect 30748 26367 30800 26376
rect 30748 26333 30755 26367
rect 30755 26333 30800 26367
rect 30748 26324 30800 26333
rect 30932 26367 30984 26376
rect 30932 26333 30941 26367
rect 30941 26333 30975 26367
rect 30975 26333 30984 26367
rect 30932 26324 30984 26333
rect 31208 26324 31260 26376
rect 31392 26324 31444 26376
rect 32864 26324 32916 26376
rect 33508 26324 33560 26376
rect 33876 26367 33928 26376
rect 33876 26333 33885 26367
rect 33885 26333 33919 26367
rect 33919 26333 33928 26367
rect 33876 26324 33928 26333
rect 34888 26367 34940 26376
rect 34888 26333 34897 26367
rect 34897 26333 34931 26367
rect 34931 26333 34940 26367
rect 34888 26324 34940 26333
rect 35900 26460 35952 26512
rect 35808 26392 35860 26444
rect 31576 26256 31628 26308
rect 32404 26256 32456 26308
rect 33048 26256 33100 26308
rect 35072 26299 35124 26308
rect 35072 26265 35081 26299
rect 35081 26265 35115 26299
rect 35115 26265 35124 26299
rect 35072 26256 35124 26265
rect 35164 26299 35216 26308
rect 35164 26265 35173 26299
rect 35173 26265 35207 26299
rect 35207 26265 35216 26299
rect 35164 26256 35216 26265
rect 35348 26256 35400 26308
rect 35900 26367 35952 26376
rect 35900 26333 35909 26367
rect 35909 26333 35943 26367
rect 35943 26333 35952 26367
rect 35900 26324 35952 26333
rect 36544 26392 36596 26444
rect 36176 26367 36228 26376
rect 36176 26333 36185 26367
rect 36185 26333 36219 26367
rect 36219 26333 36228 26367
rect 36176 26324 36228 26333
rect 36268 26367 36320 26376
rect 36268 26333 36277 26367
rect 36277 26333 36311 26367
rect 36311 26333 36320 26367
rect 36268 26324 36320 26333
rect 36912 26367 36964 26376
rect 36912 26333 36921 26367
rect 36921 26333 36955 26367
rect 36955 26333 36964 26367
rect 36912 26324 36964 26333
rect 36820 26256 36872 26308
rect 37464 26256 37516 26308
rect 25504 26188 25556 26240
rect 27712 26188 27764 26240
rect 27896 26188 27948 26240
rect 28908 26188 28960 26240
rect 30472 26188 30524 26240
rect 30748 26188 30800 26240
rect 31208 26231 31260 26240
rect 31208 26197 31217 26231
rect 31217 26197 31251 26231
rect 31251 26197 31260 26231
rect 31208 26188 31260 26197
rect 32864 26188 32916 26240
rect 34796 26188 34848 26240
rect 35900 26188 35952 26240
rect 37740 26188 37792 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 2412 25984 2464 26036
rect 10140 25916 10192 25968
rect 10968 26027 11020 26036
rect 10968 25993 10977 26027
rect 10977 25993 11011 26027
rect 11011 25993 11020 26027
rect 10968 25984 11020 25993
rect 11060 25984 11112 26036
rect 12992 25984 13044 26036
rect 15844 25984 15896 26036
rect 16488 25984 16540 26036
rect 18512 25984 18564 26036
rect 18788 26027 18840 26036
rect 18788 25993 18797 26027
rect 18797 25993 18831 26027
rect 18831 25993 18840 26027
rect 18788 25984 18840 25993
rect 19064 25984 19116 26036
rect 8300 25848 8352 25900
rect 10416 25891 10468 25900
rect 10416 25857 10425 25891
rect 10425 25857 10459 25891
rect 10459 25857 10468 25891
rect 10416 25848 10468 25857
rect 10600 25891 10652 25900
rect 10600 25857 10609 25891
rect 10609 25857 10643 25891
rect 10643 25857 10652 25891
rect 10600 25848 10652 25857
rect 10876 25848 10928 25900
rect 11704 25891 11756 25900
rect 11704 25857 11713 25891
rect 11713 25857 11747 25891
rect 11747 25857 11756 25891
rect 11704 25848 11756 25857
rect 11980 25891 12032 25900
rect 11980 25857 12014 25891
rect 12014 25857 12032 25891
rect 11980 25848 12032 25857
rect 12716 25916 12768 25968
rect 14740 25916 14792 25968
rect 11336 25780 11388 25832
rect 13728 25848 13780 25900
rect 14096 25848 14148 25900
rect 14188 25891 14240 25900
rect 14188 25857 14197 25891
rect 14197 25857 14231 25891
rect 14231 25857 14240 25891
rect 14188 25848 14240 25857
rect 14464 25848 14516 25900
rect 15568 25848 15620 25900
rect 17040 25848 17092 25900
rect 13912 25780 13964 25832
rect 9864 25712 9916 25764
rect 11704 25644 11756 25696
rect 14096 25644 14148 25696
rect 17592 25712 17644 25764
rect 16212 25687 16264 25696
rect 16212 25653 16221 25687
rect 16221 25653 16255 25687
rect 16255 25653 16264 25687
rect 16212 25644 16264 25653
rect 17408 25687 17460 25696
rect 17408 25653 17417 25687
rect 17417 25653 17451 25687
rect 17451 25653 17460 25687
rect 17408 25644 17460 25653
rect 17960 25916 18012 25968
rect 20536 25916 20588 25968
rect 22008 25959 22060 25968
rect 22008 25925 22017 25959
rect 22017 25925 22051 25959
rect 22051 25925 22060 25959
rect 22008 25916 22060 25925
rect 22192 26027 22244 26036
rect 22192 25993 22201 26027
rect 22201 25993 22235 26027
rect 22235 25993 22244 26027
rect 22192 25984 22244 25993
rect 26700 25916 26752 25968
rect 17868 25891 17920 25900
rect 17868 25857 17877 25891
rect 17877 25857 17911 25891
rect 17911 25857 17920 25891
rect 17868 25848 17920 25857
rect 18604 25891 18656 25900
rect 18604 25857 18613 25891
rect 18613 25857 18647 25891
rect 18647 25857 18656 25891
rect 18604 25848 18656 25857
rect 19432 25891 19484 25900
rect 19432 25857 19441 25891
rect 19441 25857 19475 25891
rect 19475 25857 19484 25891
rect 19432 25848 19484 25857
rect 19616 25891 19668 25900
rect 19616 25857 19625 25891
rect 19625 25857 19659 25891
rect 19659 25857 19668 25891
rect 19616 25848 19668 25857
rect 20168 25891 20220 25900
rect 20168 25857 20177 25891
rect 20177 25857 20211 25891
rect 20211 25857 20220 25891
rect 20168 25848 20220 25857
rect 20352 25891 20404 25900
rect 20352 25857 20361 25891
rect 20361 25857 20395 25891
rect 20395 25857 20404 25891
rect 20352 25848 20404 25857
rect 20628 25848 20680 25900
rect 18420 25823 18472 25832
rect 18420 25789 18429 25823
rect 18429 25789 18463 25823
rect 18463 25789 18472 25823
rect 18420 25780 18472 25789
rect 19064 25780 19116 25832
rect 19340 25780 19392 25832
rect 19248 25712 19300 25764
rect 19892 25780 19944 25832
rect 20996 25823 21048 25832
rect 20996 25789 21005 25823
rect 21005 25789 21039 25823
rect 21039 25789 21048 25823
rect 20996 25780 21048 25789
rect 21732 25848 21784 25900
rect 25964 25848 26016 25900
rect 20352 25712 20404 25764
rect 20536 25712 20588 25764
rect 22100 25712 22152 25764
rect 22192 25712 22244 25764
rect 23204 25780 23256 25832
rect 24768 25780 24820 25832
rect 26700 25780 26752 25832
rect 27620 25891 27672 25900
rect 27620 25857 27629 25891
rect 27629 25857 27663 25891
rect 27663 25857 27672 25891
rect 27620 25848 27672 25857
rect 27988 25891 28040 25900
rect 27988 25857 27997 25891
rect 27997 25857 28031 25891
rect 28031 25857 28040 25891
rect 27988 25848 28040 25857
rect 32864 25984 32916 26036
rect 32956 25984 33008 26036
rect 35072 25984 35124 26036
rect 35164 25984 35216 26036
rect 36360 25984 36412 26036
rect 37464 26027 37516 26036
rect 37464 25993 37473 26027
rect 37473 25993 37507 26027
rect 37507 25993 37516 26027
rect 37464 25984 37516 25993
rect 29644 25916 29696 25968
rect 28908 25848 28960 25900
rect 29184 25891 29236 25900
rect 29184 25857 29193 25891
rect 29193 25857 29227 25891
rect 29227 25857 29236 25891
rect 29184 25848 29236 25857
rect 30196 25916 30248 25968
rect 31760 25916 31812 25968
rect 32220 25916 32272 25968
rect 32404 25959 32456 25968
rect 32404 25925 32413 25959
rect 32413 25925 32447 25959
rect 32447 25925 32456 25959
rect 32404 25916 32456 25925
rect 27712 25780 27764 25832
rect 27896 25780 27948 25832
rect 28172 25823 28224 25832
rect 28172 25789 28181 25823
rect 28181 25789 28215 25823
rect 28215 25789 28224 25823
rect 28172 25780 28224 25789
rect 28724 25780 28776 25832
rect 32496 25848 32548 25900
rect 30748 25823 30800 25832
rect 30748 25789 30757 25823
rect 30757 25789 30791 25823
rect 30791 25789 30800 25823
rect 30748 25780 30800 25789
rect 19984 25644 20036 25696
rect 20168 25644 20220 25696
rect 20904 25687 20956 25696
rect 20904 25653 20913 25687
rect 20913 25653 20947 25687
rect 20947 25653 20956 25687
rect 20904 25644 20956 25653
rect 20996 25644 21048 25696
rect 21272 25644 21324 25696
rect 23388 25712 23440 25764
rect 24124 25755 24176 25764
rect 24124 25721 24133 25755
rect 24133 25721 24167 25755
rect 24167 25721 24176 25755
rect 24124 25712 24176 25721
rect 26332 25712 26384 25764
rect 30196 25712 30248 25764
rect 30564 25712 30616 25764
rect 31392 25780 31444 25832
rect 33048 25916 33100 25968
rect 32772 25848 32824 25900
rect 33968 25848 34020 25900
rect 32404 25712 32456 25764
rect 33876 25755 33928 25764
rect 33876 25721 33885 25755
rect 33885 25721 33919 25755
rect 33919 25721 33928 25755
rect 33876 25712 33928 25721
rect 22744 25644 22796 25696
rect 26884 25644 26936 25696
rect 27988 25644 28040 25696
rect 28356 25644 28408 25696
rect 30380 25644 30432 25696
rect 30472 25644 30524 25696
rect 32220 25644 32272 25696
rect 33968 25644 34020 25696
rect 34428 25823 34480 25832
rect 34428 25789 34437 25823
rect 34437 25789 34471 25823
rect 34471 25789 34480 25823
rect 34428 25780 34480 25789
rect 35072 25780 35124 25832
rect 36912 25916 36964 25968
rect 37372 25916 37424 25968
rect 37740 25916 37792 25968
rect 38016 25823 38068 25832
rect 38016 25789 38025 25823
rect 38025 25789 38059 25823
rect 38059 25789 38068 25823
rect 38016 25780 38068 25789
rect 38568 25712 38620 25764
rect 36728 25644 36780 25696
rect 36820 25687 36872 25696
rect 36820 25653 36829 25687
rect 36829 25653 36863 25687
rect 36863 25653 36872 25687
rect 36820 25644 36872 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 15476 25440 15528 25492
rect 15568 25483 15620 25492
rect 15568 25449 15577 25483
rect 15577 25449 15611 25483
rect 15611 25449 15620 25483
rect 15568 25440 15620 25449
rect 16580 25483 16632 25492
rect 16580 25449 16589 25483
rect 16589 25449 16623 25483
rect 16623 25449 16632 25483
rect 16580 25440 16632 25449
rect 17040 25483 17092 25492
rect 17040 25449 17049 25483
rect 17049 25449 17083 25483
rect 17083 25449 17092 25483
rect 17040 25440 17092 25449
rect 20444 25440 20496 25492
rect 20628 25440 20680 25492
rect 23572 25440 23624 25492
rect 25688 25440 25740 25492
rect 25872 25483 25924 25492
rect 25872 25449 25881 25483
rect 25881 25449 25915 25483
rect 25915 25449 25924 25483
rect 25872 25440 25924 25449
rect 10140 25372 10192 25424
rect 9496 25304 9548 25356
rect 10508 25304 10560 25356
rect 8852 25236 8904 25288
rect 11428 25304 11480 25356
rect 13912 25372 13964 25424
rect 14740 25372 14792 25424
rect 15108 25372 15160 25424
rect 19800 25372 19852 25424
rect 19892 25372 19944 25424
rect 10876 25236 10928 25288
rect 11060 25168 11112 25220
rect 11612 25236 11664 25288
rect 13452 25279 13504 25288
rect 13452 25245 13461 25279
rect 13461 25245 13495 25279
rect 13495 25245 13504 25279
rect 13452 25236 13504 25245
rect 15200 25304 15252 25356
rect 14648 25236 14700 25288
rect 15016 25279 15068 25288
rect 15016 25245 15025 25279
rect 15025 25245 15059 25279
rect 15059 25245 15068 25279
rect 15016 25236 15068 25245
rect 16212 25304 16264 25356
rect 17592 25304 17644 25356
rect 18604 25304 18656 25356
rect 15384 25279 15436 25288
rect 15384 25245 15393 25279
rect 15393 25245 15427 25279
rect 15427 25245 15436 25279
rect 16580 25279 16632 25288
rect 15384 25236 15436 25245
rect 16580 25245 16589 25279
rect 16589 25245 16623 25279
rect 16623 25245 16632 25279
rect 16580 25236 16632 25245
rect 16856 25279 16908 25288
rect 16856 25245 16865 25279
rect 16865 25245 16899 25279
rect 16899 25245 16908 25279
rect 16856 25236 16908 25245
rect 16948 25236 17000 25288
rect 19064 25304 19116 25356
rect 18788 25236 18840 25288
rect 12072 25168 12124 25220
rect 14464 25211 14516 25220
rect 14464 25177 14473 25211
rect 14473 25177 14507 25211
rect 14507 25177 14516 25211
rect 14464 25168 14516 25177
rect 14924 25168 14976 25220
rect 9128 25143 9180 25152
rect 9128 25109 9137 25143
rect 9137 25109 9171 25143
rect 9171 25109 9180 25143
rect 9128 25100 9180 25109
rect 9496 25143 9548 25152
rect 9496 25109 9505 25143
rect 9505 25109 9539 25143
rect 9539 25109 9548 25143
rect 9496 25100 9548 25109
rect 10232 25100 10284 25152
rect 11704 25100 11756 25152
rect 15292 25100 15344 25152
rect 18512 25168 18564 25220
rect 17500 25143 17552 25152
rect 17500 25109 17509 25143
rect 17509 25109 17543 25143
rect 17543 25109 17552 25143
rect 17500 25100 17552 25109
rect 20352 25304 20404 25356
rect 21456 25347 21508 25356
rect 21456 25313 21465 25347
rect 21465 25313 21499 25347
rect 21499 25313 21508 25347
rect 21456 25304 21508 25313
rect 22652 25347 22704 25356
rect 22652 25313 22661 25347
rect 22661 25313 22695 25347
rect 22695 25313 22704 25347
rect 22652 25304 22704 25313
rect 20352 25168 20404 25220
rect 20628 25168 20680 25220
rect 22468 25279 22520 25288
rect 22468 25245 22477 25279
rect 22477 25245 22511 25279
rect 22511 25245 22520 25279
rect 22468 25236 22520 25245
rect 23664 25372 23716 25424
rect 24032 25372 24084 25424
rect 23572 25347 23624 25356
rect 23572 25313 23581 25347
rect 23581 25313 23615 25347
rect 23615 25313 23624 25347
rect 23572 25304 23624 25313
rect 24952 25372 25004 25424
rect 25044 25372 25096 25424
rect 26240 25372 26292 25424
rect 24584 25304 24636 25356
rect 24860 25304 24912 25356
rect 23112 25236 23164 25288
rect 25320 25236 25372 25288
rect 25872 25304 25924 25356
rect 27988 25372 28040 25424
rect 28908 25440 28960 25492
rect 29552 25440 29604 25492
rect 26516 25279 26568 25288
rect 26516 25245 26525 25279
rect 26525 25245 26559 25279
rect 26559 25245 26568 25279
rect 26516 25236 26568 25245
rect 26608 25279 26660 25288
rect 26608 25245 26617 25279
rect 26617 25245 26651 25279
rect 26651 25245 26660 25279
rect 26608 25236 26660 25245
rect 27620 25279 27672 25288
rect 27620 25245 27629 25279
rect 27629 25245 27663 25279
rect 27663 25245 27672 25279
rect 27620 25236 27672 25245
rect 28080 25236 28132 25288
rect 28908 25304 28960 25356
rect 22560 25168 22612 25220
rect 20076 25100 20128 25152
rect 20996 25143 21048 25152
rect 20996 25109 21005 25143
rect 21005 25109 21039 25143
rect 21039 25109 21048 25143
rect 20996 25100 21048 25109
rect 21364 25143 21416 25152
rect 21364 25109 21373 25143
rect 21373 25109 21407 25143
rect 21407 25109 21416 25143
rect 21364 25100 21416 25109
rect 21456 25100 21508 25152
rect 24860 25168 24912 25220
rect 25044 25100 25096 25152
rect 25136 25100 25188 25152
rect 27988 25168 28040 25220
rect 30288 25483 30340 25492
rect 30288 25449 30297 25483
rect 30297 25449 30331 25483
rect 30331 25449 30340 25483
rect 30288 25440 30340 25449
rect 30472 25440 30524 25492
rect 31392 25440 31444 25492
rect 33508 25440 33560 25492
rect 36084 25440 36136 25492
rect 36636 25440 36688 25492
rect 36728 25440 36780 25492
rect 39304 25440 39356 25492
rect 30932 25372 30984 25424
rect 33416 25372 33468 25424
rect 29920 25304 29972 25356
rect 31392 25304 31444 25356
rect 32956 25304 33008 25356
rect 35532 25372 35584 25424
rect 33784 25304 33836 25356
rect 28356 25211 28408 25220
rect 28356 25177 28365 25211
rect 28365 25177 28399 25211
rect 28399 25177 28408 25211
rect 28356 25168 28408 25177
rect 27252 25143 27304 25152
rect 27252 25109 27261 25143
rect 27261 25109 27295 25143
rect 27295 25109 27304 25143
rect 27252 25100 27304 25109
rect 27896 25100 27948 25152
rect 30196 25236 30248 25288
rect 30288 25236 30340 25288
rect 31484 25236 31536 25288
rect 32220 25279 32272 25288
rect 32220 25245 32229 25279
rect 32229 25245 32263 25279
rect 32263 25245 32272 25279
rect 32220 25236 32272 25245
rect 32404 25279 32456 25288
rect 29184 25168 29236 25220
rect 28908 25100 28960 25152
rect 29000 25100 29052 25152
rect 29552 25168 29604 25220
rect 30472 25168 30524 25220
rect 30564 25168 30616 25220
rect 31576 25168 31628 25220
rect 30196 25100 30248 25152
rect 31116 25100 31168 25152
rect 32404 25245 32413 25279
rect 32413 25245 32447 25279
rect 32447 25245 32456 25279
rect 32404 25236 32456 25245
rect 32864 25236 32916 25288
rect 33232 25236 33284 25288
rect 34428 25304 34480 25356
rect 35624 25304 35676 25356
rect 35256 25279 35308 25288
rect 35256 25245 35265 25279
rect 35265 25245 35299 25279
rect 35299 25245 35308 25279
rect 35256 25236 35308 25245
rect 36084 25279 36136 25288
rect 36084 25245 36093 25279
rect 36093 25245 36127 25279
rect 36127 25245 36136 25279
rect 36084 25236 36136 25245
rect 36176 25279 36228 25288
rect 36176 25245 36185 25279
rect 36185 25245 36219 25279
rect 36219 25245 36228 25279
rect 36176 25236 36228 25245
rect 36912 25347 36964 25356
rect 36912 25313 36921 25347
rect 36921 25313 36955 25347
rect 36955 25313 36964 25347
rect 36912 25304 36964 25313
rect 37648 25236 37700 25288
rect 33600 25168 33652 25220
rect 34980 25168 35032 25220
rect 33140 25100 33192 25152
rect 33876 25100 33928 25152
rect 34796 25100 34848 25152
rect 35808 25168 35860 25220
rect 37004 25168 37056 25220
rect 37188 25211 37240 25220
rect 37188 25177 37222 25211
rect 37222 25177 37240 25211
rect 37188 25168 37240 25177
rect 35348 25100 35400 25152
rect 35440 25143 35492 25152
rect 35440 25109 35449 25143
rect 35449 25109 35483 25143
rect 35483 25109 35492 25143
rect 35440 25100 35492 25109
rect 36820 25100 36872 25152
rect 37832 25100 37884 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9496 24896 9548 24948
rect 15108 24939 15160 24948
rect 9128 24828 9180 24880
rect 15108 24905 15117 24939
rect 15117 24905 15151 24939
rect 15151 24905 15160 24939
rect 15108 24896 15160 24905
rect 16304 24896 16356 24948
rect 17316 24896 17368 24948
rect 17500 24896 17552 24948
rect 19524 24896 19576 24948
rect 18788 24828 18840 24880
rect 5356 24760 5408 24812
rect 10140 24760 10192 24812
rect 10232 24803 10284 24812
rect 10232 24769 10241 24803
rect 10241 24769 10275 24803
rect 10275 24769 10284 24803
rect 10232 24760 10284 24769
rect 10324 24803 10376 24812
rect 10324 24769 10333 24803
rect 10333 24769 10367 24803
rect 10367 24769 10376 24803
rect 10324 24760 10376 24769
rect 10876 24760 10928 24812
rect 11704 24803 11756 24812
rect 11704 24769 11713 24803
rect 11713 24769 11747 24803
rect 11747 24769 11756 24803
rect 11704 24760 11756 24769
rect 11888 24803 11940 24812
rect 11888 24769 11897 24803
rect 11897 24769 11931 24803
rect 11931 24769 11940 24803
rect 11888 24760 11940 24769
rect 11980 24803 12032 24812
rect 11980 24769 11989 24803
rect 11989 24769 12023 24803
rect 12023 24769 12032 24803
rect 11980 24760 12032 24769
rect 12072 24803 12124 24812
rect 12072 24769 12081 24803
rect 12081 24769 12115 24803
rect 12115 24769 12124 24803
rect 12072 24760 12124 24769
rect 8208 24735 8260 24744
rect 8208 24701 8217 24735
rect 8217 24701 8251 24735
rect 8251 24701 8260 24735
rect 8208 24692 8260 24701
rect 11428 24692 11480 24744
rect 12900 24735 12952 24744
rect 12900 24701 12909 24735
rect 12909 24701 12943 24735
rect 12943 24701 12952 24735
rect 12900 24692 12952 24701
rect 10876 24624 10928 24676
rect 14372 24692 14424 24744
rect 10048 24599 10100 24608
rect 10048 24565 10057 24599
rect 10057 24565 10091 24599
rect 10091 24565 10100 24599
rect 10048 24556 10100 24565
rect 12256 24599 12308 24608
rect 12256 24565 12265 24599
rect 12265 24565 12299 24599
rect 12299 24565 12308 24599
rect 12256 24556 12308 24565
rect 15016 24624 15068 24676
rect 16212 24760 16264 24812
rect 16856 24760 16908 24812
rect 17316 24760 17368 24812
rect 17684 24803 17736 24812
rect 17684 24769 17693 24803
rect 17693 24769 17727 24803
rect 17727 24769 17736 24803
rect 17684 24760 17736 24769
rect 19800 24871 19852 24880
rect 19800 24837 19809 24871
rect 19809 24837 19843 24871
rect 19843 24837 19852 24871
rect 19800 24828 19852 24837
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 19616 24760 19668 24812
rect 20996 24939 21048 24948
rect 20996 24905 21005 24939
rect 21005 24905 21039 24939
rect 21039 24905 21048 24939
rect 20996 24896 21048 24905
rect 22652 24896 22704 24948
rect 26148 24896 26200 24948
rect 27620 24896 27672 24948
rect 28356 24896 28408 24948
rect 21364 24828 21416 24880
rect 20260 24760 20312 24812
rect 20904 24803 20956 24812
rect 18328 24692 18380 24744
rect 15844 24624 15896 24676
rect 19800 24692 19852 24744
rect 20904 24769 20913 24803
rect 20913 24769 20947 24803
rect 20947 24769 20956 24803
rect 20904 24760 20956 24769
rect 21824 24760 21876 24812
rect 23940 24803 23992 24812
rect 23940 24769 23949 24803
rect 23949 24769 23983 24803
rect 23983 24769 23992 24803
rect 23940 24760 23992 24769
rect 24676 24760 24728 24812
rect 25780 24828 25832 24880
rect 25964 24803 26016 24812
rect 20536 24692 20588 24744
rect 22008 24735 22060 24744
rect 22008 24701 22017 24735
rect 22017 24701 22051 24735
rect 22051 24701 22060 24735
rect 22008 24692 22060 24701
rect 25964 24769 25973 24803
rect 25973 24769 26007 24803
rect 26007 24769 26016 24803
rect 25964 24760 26016 24769
rect 26056 24760 26108 24812
rect 26240 24803 26292 24812
rect 26240 24769 26249 24803
rect 26249 24769 26283 24803
rect 26283 24769 26292 24803
rect 26240 24760 26292 24769
rect 27344 24828 27396 24880
rect 29184 24896 29236 24948
rect 31208 24896 31260 24948
rect 31484 24896 31536 24948
rect 29092 24828 29144 24880
rect 27620 24803 27672 24812
rect 27620 24769 27629 24803
rect 27629 24769 27663 24803
rect 27663 24769 27672 24803
rect 27620 24760 27672 24769
rect 26884 24692 26936 24744
rect 27896 24760 27948 24812
rect 29184 24760 29236 24812
rect 29460 24828 29512 24880
rect 30288 24828 30340 24880
rect 30472 24828 30524 24880
rect 31300 24828 31352 24880
rect 32864 24871 32916 24880
rect 32864 24837 32873 24871
rect 32873 24837 32907 24871
rect 32907 24837 32916 24871
rect 32864 24828 32916 24837
rect 33140 24828 33192 24880
rect 33508 24828 33560 24880
rect 29552 24803 29604 24812
rect 29552 24769 29561 24803
rect 29561 24769 29595 24803
rect 29595 24769 29604 24803
rect 29552 24760 29604 24769
rect 29644 24803 29696 24812
rect 29644 24769 29653 24803
rect 29653 24769 29687 24803
rect 29687 24769 29696 24803
rect 29644 24760 29696 24769
rect 30196 24760 30248 24812
rect 30380 24803 30432 24812
rect 30380 24769 30389 24803
rect 30389 24769 30423 24803
rect 30423 24769 30432 24803
rect 30380 24760 30432 24769
rect 30656 24803 30708 24812
rect 30656 24769 30665 24803
rect 30665 24769 30699 24803
rect 30699 24769 30708 24803
rect 30656 24760 30708 24769
rect 31392 24803 31444 24812
rect 31392 24769 31401 24803
rect 31401 24769 31435 24803
rect 31435 24769 31444 24803
rect 31392 24760 31444 24769
rect 27988 24692 28040 24744
rect 28540 24735 28592 24744
rect 28540 24701 28549 24735
rect 28549 24701 28583 24735
rect 28583 24701 28592 24735
rect 28540 24692 28592 24701
rect 31116 24692 31168 24744
rect 20168 24624 20220 24676
rect 25504 24624 25556 24676
rect 16764 24556 16816 24608
rect 17316 24599 17368 24608
rect 17316 24565 17325 24599
rect 17325 24565 17359 24599
rect 17359 24565 17368 24599
rect 17316 24556 17368 24565
rect 20536 24599 20588 24608
rect 20536 24565 20545 24599
rect 20545 24565 20579 24599
rect 20579 24565 20588 24599
rect 20536 24556 20588 24565
rect 20720 24556 20772 24608
rect 22652 24556 22704 24608
rect 23848 24556 23900 24608
rect 25320 24599 25372 24608
rect 25320 24565 25329 24599
rect 25329 24565 25363 24599
rect 25363 24565 25372 24599
rect 25320 24556 25372 24565
rect 25964 24556 26016 24608
rect 26424 24556 26476 24608
rect 27896 24556 27948 24608
rect 29000 24556 29052 24608
rect 29644 24556 29696 24608
rect 30288 24556 30340 24608
rect 30380 24599 30432 24608
rect 30380 24565 30389 24599
rect 30389 24565 30423 24599
rect 30423 24565 30432 24599
rect 30380 24556 30432 24565
rect 30472 24556 30524 24608
rect 30840 24556 30892 24608
rect 31208 24599 31260 24608
rect 31208 24565 31217 24599
rect 31217 24565 31251 24599
rect 31251 24565 31260 24599
rect 31208 24556 31260 24565
rect 31760 24624 31812 24676
rect 32220 24624 32272 24676
rect 34980 24896 35032 24948
rect 35624 24896 35676 24948
rect 35992 24896 36044 24948
rect 37556 24896 37608 24948
rect 37832 24939 37884 24948
rect 37832 24905 37841 24939
rect 37841 24905 37875 24939
rect 37875 24905 37884 24939
rect 37832 24896 37884 24905
rect 32404 24692 32456 24744
rect 33876 24760 33928 24812
rect 34612 24803 34664 24812
rect 34612 24769 34621 24803
rect 34621 24769 34655 24803
rect 34655 24769 34664 24803
rect 34612 24760 34664 24769
rect 34888 24803 34940 24812
rect 34888 24769 34897 24803
rect 34897 24769 34931 24803
rect 34931 24769 34940 24803
rect 34888 24760 34940 24769
rect 32956 24735 33008 24744
rect 32956 24701 32965 24735
rect 32965 24701 32999 24735
rect 32999 24701 33008 24735
rect 32956 24692 33008 24701
rect 33140 24692 33192 24744
rect 34060 24692 34112 24744
rect 35348 24760 35400 24812
rect 35532 24760 35584 24812
rect 35808 24803 35860 24812
rect 35808 24769 35818 24803
rect 35818 24769 35852 24803
rect 35852 24769 35860 24803
rect 35808 24760 35860 24769
rect 35992 24803 36044 24812
rect 35992 24769 36001 24803
rect 36001 24769 36035 24803
rect 36035 24769 36044 24803
rect 35992 24760 36044 24769
rect 36268 24760 36320 24812
rect 39580 24760 39632 24812
rect 36452 24692 36504 24744
rect 38016 24735 38068 24744
rect 38016 24701 38025 24735
rect 38025 24701 38059 24735
rect 38059 24701 38068 24735
rect 38016 24692 38068 24701
rect 35440 24624 35492 24676
rect 33416 24599 33468 24608
rect 33416 24565 33425 24599
rect 33425 24565 33459 24599
rect 33459 24565 33468 24599
rect 33416 24556 33468 24565
rect 33876 24556 33928 24608
rect 34244 24556 34296 24608
rect 35808 24556 35860 24608
rect 37188 24624 37240 24676
rect 37372 24556 37424 24608
rect 37648 24556 37700 24608
rect 37924 24556 37976 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2688 24352 2740 24404
rect 15292 24352 15344 24404
rect 16212 24352 16264 24404
rect 18696 24395 18748 24404
rect 18696 24361 18705 24395
rect 18705 24361 18739 24395
rect 18739 24361 18748 24395
rect 18696 24352 18748 24361
rect 18880 24352 18932 24404
rect 19616 24352 19668 24404
rect 11980 24216 12032 24268
rect 14740 24284 14792 24336
rect 12900 24216 12952 24268
rect 13452 24216 13504 24268
rect 8208 24148 8260 24200
rect 11428 24148 11480 24200
rect 12348 24148 12400 24200
rect 12256 24080 12308 24132
rect 13728 24191 13780 24200
rect 13728 24157 13737 24191
rect 13737 24157 13771 24191
rect 13771 24157 13780 24191
rect 13728 24148 13780 24157
rect 14832 24148 14884 24200
rect 15660 24148 15712 24200
rect 19340 24284 19392 24336
rect 17316 24259 17368 24268
rect 17316 24225 17325 24259
rect 17325 24225 17359 24259
rect 17359 24225 17368 24259
rect 17316 24216 17368 24225
rect 17408 24259 17460 24268
rect 17408 24225 17417 24259
rect 17417 24225 17451 24259
rect 17451 24225 17460 24259
rect 17408 24216 17460 24225
rect 16580 24148 16632 24200
rect 20904 24352 20956 24404
rect 21824 24352 21876 24404
rect 22468 24352 22520 24404
rect 30380 24352 30432 24404
rect 31760 24395 31812 24404
rect 31760 24361 31769 24395
rect 31769 24361 31803 24395
rect 31803 24361 31812 24395
rect 31760 24352 31812 24361
rect 32680 24395 32732 24404
rect 32680 24361 32689 24395
rect 32689 24361 32723 24395
rect 32723 24361 32732 24395
rect 32680 24352 32732 24361
rect 33232 24352 33284 24404
rect 20812 24284 20864 24336
rect 22468 24216 22520 24268
rect 22560 24259 22612 24268
rect 22560 24225 22569 24259
rect 22569 24225 22603 24259
rect 22603 24225 22612 24259
rect 22560 24216 22612 24225
rect 18420 24191 18472 24200
rect 18420 24157 18429 24191
rect 18429 24157 18463 24191
rect 18463 24157 18472 24191
rect 18420 24148 18472 24157
rect 14004 24080 14056 24132
rect 15016 24080 15068 24132
rect 15936 24080 15988 24132
rect 12992 24012 13044 24064
rect 13084 24055 13136 24064
rect 13084 24021 13093 24055
rect 13093 24021 13127 24055
rect 13127 24021 13136 24055
rect 13084 24012 13136 24021
rect 13360 24012 13412 24064
rect 16856 24055 16908 24064
rect 16856 24021 16865 24055
rect 16865 24021 16899 24055
rect 16899 24021 16908 24055
rect 16856 24012 16908 24021
rect 17132 24012 17184 24064
rect 18420 24012 18472 24064
rect 18604 24148 18656 24200
rect 19064 24148 19116 24200
rect 22008 24148 22060 24200
rect 23480 24191 23532 24200
rect 23480 24157 23489 24191
rect 23489 24157 23523 24191
rect 23523 24157 23532 24191
rect 23480 24148 23532 24157
rect 26700 24284 26752 24336
rect 28356 24284 28408 24336
rect 29644 24284 29696 24336
rect 24860 24216 24912 24268
rect 24952 24148 25004 24200
rect 25688 24216 25740 24268
rect 27160 24216 27212 24268
rect 27804 24216 27856 24268
rect 20536 24080 20588 24132
rect 20076 24012 20128 24064
rect 20260 24012 20312 24064
rect 23848 24080 23900 24132
rect 23940 24080 23992 24132
rect 25872 24148 25924 24200
rect 26240 24148 26292 24200
rect 25688 24080 25740 24132
rect 26608 24191 26660 24200
rect 26608 24157 26617 24191
rect 26617 24157 26651 24191
rect 26651 24157 26660 24191
rect 26608 24148 26660 24157
rect 27068 24148 27120 24200
rect 27896 24191 27948 24200
rect 27896 24157 27905 24191
rect 27905 24157 27939 24191
rect 27939 24157 27948 24191
rect 27896 24148 27948 24157
rect 27988 24191 28040 24200
rect 27988 24157 27997 24191
rect 27997 24157 28031 24191
rect 28031 24157 28040 24191
rect 27988 24148 28040 24157
rect 29276 24148 29328 24200
rect 29552 24148 29604 24200
rect 26700 24080 26752 24132
rect 30472 24284 30524 24336
rect 32128 24216 32180 24268
rect 30196 24148 30248 24200
rect 30288 24148 30340 24200
rect 23572 24055 23624 24064
rect 23572 24021 23581 24055
rect 23581 24021 23615 24055
rect 23615 24021 23624 24055
rect 23572 24012 23624 24021
rect 25872 24012 25924 24064
rect 26516 24012 26568 24064
rect 29092 24055 29144 24064
rect 29092 24021 29101 24055
rect 29101 24021 29135 24055
rect 29135 24021 29144 24055
rect 29092 24012 29144 24021
rect 30656 24080 30708 24132
rect 31852 24148 31904 24200
rect 33784 24352 33836 24404
rect 35348 24352 35400 24404
rect 36268 24352 36320 24404
rect 33600 24284 33652 24336
rect 34428 24284 34480 24336
rect 35624 24284 35676 24336
rect 35716 24284 35768 24336
rect 36728 24284 36780 24336
rect 33508 24148 33560 24200
rect 33784 24191 33836 24200
rect 33784 24157 33793 24191
rect 33793 24157 33827 24191
rect 33827 24157 33836 24191
rect 33784 24148 33836 24157
rect 32220 24080 32272 24132
rect 32496 24123 32548 24132
rect 32496 24089 32505 24123
rect 32505 24089 32539 24123
rect 32539 24089 32548 24123
rect 32496 24080 32548 24089
rect 32588 24080 32640 24132
rect 30840 24012 30892 24064
rect 31116 24012 31168 24064
rect 31668 24012 31720 24064
rect 32128 24012 32180 24064
rect 32864 24055 32916 24064
rect 32864 24021 32873 24055
rect 32873 24021 32907 24055
rect 32907 24021 32916 24055
rect 32864 24012 32916 24021
rect 33416 24080 33468 24132
rect 34888 24191 34940 24200
rect 34888 24157 34897 24191
rect 34897 24157 34931 24191
rect 34931 24157 34940 24191
rect 34888 24148 34940 24157
rect 35072 24148 35124 24200
rect 35808 24191 35860 24200
rect 35808 24157 35817 24191
rect 35817 24157 35851 24191
rect 35851 24157 35860 24191
rect 35808 24148 35860 24157
rect 36912 24259 36964 24268
rect 36912 24225 36921 24259
rect 36921 24225 36955 24259
rect 36955 24225 36964 24259
rect 36912 24216 36964 24225
rect 35992 24148 36044 24200
rect 36268 24148 36320 24200
rect 35256 24080 35308 24132
rect 36452 24080 36504 24132
rect 37464 24080 37516 24132
rect 36636 24012 36688 24064
rect 37832 24012 37884 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 10876 23851 10928 23860
rect 10876 23817 10885 23851
rect 10885 23817 10919 23851
rect 10919 23817 10928 23851
rect 10876 23808 10928 23817
rect 12348 23808 12400 23860
rect 10048 23740 10100 23792
rect 8208 23672 8260 23724
rect 12808 23672 12860 23724
rect 13084 23740 13136 23792
rect 13452 23715 13504 23724
rect 13452 23681 13461 23715
rect 13461 23681 13495 23715
rect 13495 23681 13504 23715
rect 13452 23672 13504 23681
rect 11060 23604 11112 23656
rect 12256 23604 12308 23656
rect 14004 23672 14056 23724
rect 15936 23851 15988 23860
rect 15936 23817 15945 23851
rect 15945 23817 15979 23851
rect 15979 23817 15988 23851
rect 15936 23808 15988 23817
rect 18880 23808 18932 23860
rect 19616 23808 19668 23860
rect 20260 23808 20312 23860
rect 20444 23851 20496 23860
rect 20444 23817 20453 23851
rect 20453 23817 20487 23851
rect 20487 23817 20496 23851
rect 20444 23808 20496 23817
rect 20536 23808 20588 23860
rect 20996 23808 21048 23860
rect 23296 23808 23348 23860
rect 26332 23808 26384 23860
rect 16120 23740 16172 23792
rect 15660 23715 15712 23724
rect 15660 23681 15669 23715
rect 15669 23681 15703 23715
rect 15703 23681 15712 23715
rect 15660 23672 15712 23681
rect 16396 23672 16448 23724
rect 17040 23672 17092 23724
rect 17316 23715 17368 23724
rect 17316 23681 17325 23715
rect 17325 23681 17359 23715
rect 17359 23681 17368 23715
rect 17316 23672 17368 23681
rect 19432 23672 19484 23724
rect 19708 23715 19760 23724
rect 19708 23681 19717 23715
rect 19717 23681 19751 23715
rect 19751 23681 19760 23715
rect 19708 23672 19760 23681
rect 20536 23672 20588 23724
rect 20628 23715 20680 23724
rect 20628 23681 20637 23715
rect 20637 23681 20671 23715
rect 20671 23681 20680 23715
rect 20628 23672 20680 23681
rect 20904 23715 20956 23724
rect 20904 23681 20913 23715
rect 20913 23681 20947 23715
rect 20947 23681 20956 23715
rect 20904 23672 20956 23681
rect 16672 23536 16724 23588
rect 18972 23604 19024 23656
rect 19892 23604 19944 23656
rect 20076 23604 20128 23656
rect 22376 23783 22428 23792
rect 22376 23749 22385 23783
rect 22385 23749 22419 23783
rect 22419 23749 22428 23783
rect 22376 23740 22428 23749
rect 24584 23740 24636 23792
rect 25136 23740 25188 23792
rect 25964 23740 26016 23792
rect 26608 23808 26660 23860
rect 27804 23808 27856 23860
rect 28908 23808 28960 23860
rect 29460 23808 29512 23860
rect 29552 23808 29604 23860
rect 21088 23672 21140 23724
rect 22284 23715 22336 23724
rect 22284 23681 22293 23715
rect 22293 23681 22327 23715
rect 22327 23681 22336 23715
rect 22284 23672 22336 23681
rect 22836 23715 22888 23724
rect 22836 23681 22845 23715
rect 22845 23681 22879 23715
rect 22879 23681 22888 23715
rect 22836 23672 22888 23681
rect 23296 23672 23348 23724
rect 25504 23715 25556 23724
rect 25504 23681 25513 23715
rect 25513 23681 25547 23715
rect 25547 23681 25556 23715
rect 25504 23672 25556 23681
rect 11980 23511 12032 23520
rect 11980 23477 11989 23511
rect 11989 23477 12023 23511
rect 12023 23477 12032 23511
rect 11980 23468 12032 23477
rect 13728 23468 13780 23520
rect 17224 23511 17276 23520
rect 17224 23477 17233 23511
rect 17233 23477 17267 23511
rect 17267 23477 17276 23511
rect 17224 23468 17276 23477
rect 17776 23511 17828 23520
rect 17776 23477 17785 23511
rect 17785 23477 17819 23511
rect 17819 23477 17828 23511
rect 17776 23468 17828 23477
rect 18604 23536 18656 23588
rect 19616 23536 19668 23588
rect 19708 23536 19760 23588
rect 22192 23536 22244 23588
rect 24308 23579 24360 23588
rect 24308 23545 24317 23579
rect 24317 23545 24351 23579
rect 24351 23545 24360 23579
rect 26148 23715 26200 23724
rect 26148 23681 26157 23715
rect 26157 23681 26191 23715
rect 26191 23681 26200 23715
rect 26148 23672 26200 23681
rect 29276 23740 29328 23792
rect 27436 23672 27488 23724
rect 26516 23604 26568 23656
rect 28448 23672 28500 23724
rect 28540 23715 28592 23724
rect 28540 23681 28549 23715
rect 28549 23681 28583 23715
rect 28583 23681 28592 23715
rect 28540 23672 28592 23681
rect 28264 23604 28316 23656
rect 29092 23672 29144 23724
rect 30104 23783 30156 23792
rect 30104 23749 30113 23783
rect 30113 23749 30147 23783
rect 30147 23749 30156 23783
rect 30104 23740 30156 23749
rect 33416 23808 33468 23860
rect 31392 23740 31444 23792
rect 32956 23740 33008 23792
rect 33600 23740 33652 23792
rect 34796 23808 34848 23860
rect 34888 23808 34940 23860
rect 37464 23851 37516 23860
rect 37464 23817 37473 23851
rect 37473 23817 37507 23851
rect 37507 23817 37516 23851
rect 37464 23808 37516 23817
rect 37832 23851 37884 23860
rect 37832 23817 37841 23851
rect 37841 23817 37875 23851
rect 37875 23817 37884 23851
rect 37832 23808 37884 23817
rect 29276 23647 29328 23656
rect 29276 23613 29285 23647
rect 29285 23613 29319 23647
rect 29319 23613 29328 23647
rect 29276 23604 29328 23613
rect 24308 23536 24360 23545
rect 20536 23468 20588 23520
rect 20628 23468 20680 23520
rect 21640 23468 21692 23520
rect 25136 23511 25188 23520
rect 25136 23477 25145 23511
rect 25145 23477 25179 23511
rect 25179 23477 25188 23511
rect 25136 23468 25188 23477
rect 29736 23536 29788 23588
rect 30196 23715 30248 23724
rect 30196 23681 30210 23715
rect 30210 23681 30244 23715
rect 30244 23681 30248 23715
rect 30196 23672 30248 23681
rect 30380 23672 30432 23724
rect 30932 23672 30984 23724
rect 31300 23672 31352 23724
rect 32128 23672 32180 23724
rect 32312 23672 32364 23724
rect 32588 23672 32640 23724
rect 32772 23672 32824 23724
rect 33784 23672 33836 23724
rect 33876 23715 33928 23724
rect 33876 23681 33885 23715
rect 33885 23681 33919 23715
rect 33919 23681 33928 23715
rect 33876 23672 33928 23681
rect 34244 23715 34296 23724
rect 34244 23681 34253 23715
rect 34253 23681 34287 23715
rect 34287 23681 34296 23715
rect 34244 23672 34296 23681
rect 34612 23672 34664 23724
rect 34796 23672 34848 23724
rect 35716 23740 35768 23792
rect 35256 23715 35308 23724
rect 35256 23681 35265 23715
rect 35265 23681 35299 23715
rect 35299 23681 35308 23715
rect 35256 23672 35308 23681
rect 32036 23604 32088 23656
rect 33508 23604 33560 23656
rect 33600 23604 33652 23656
rect 34152 23604 34204 23656
rect 35440 23715 35492 23724
rect 35440 23681 35454 23715
rect 35454 23681 35488 23715
rect 35488 23681 35492 23715
rect 35440 23672 35492 23681
rect 35900 23672 35952 23724
rect 36360 23715 36412 23724
rect 36360 23681 36369 23715
rect 36369 23681 36403 23715
rect 36403 23681 36412 23715
rect 36360 23672 36412 23681
rect 36636 23715 36688 23724
rect 36636 23681 36645 23715
rect 36645 23681 36679 23715
rect 36679 23681 36688 23715
rect 36636 23672 36688 23681
rect 37464 23672 37516 23724
rect 35992 23604 36044 23656
rect 38016 23647 38068 23656
rect 38016 23613 38025 23647
rect 38025 23613 38059 23647
rect 38059 23613 38068 23647
rect 38016 23604 38068 23613
rect 30656 23536 30708 23588
rect 32864 23536 32916 23588
rect 36268 23536 36320 23588
rect 36544 23579 36596 23588
rect 36544 23545 36553 23579
rect 36553 23545 36587 23579
rect 36587 23545 36596 23579
rect 36544 23536 36596 23545
rect 36728 23536 36780 23588
rect 25780 23468 25832 23520
rect 27344 23468 27396 23520
rect 27712 23468 27764 23520
rect 28816 23511 28868 23520
rect 28816 23477 28825 23511
rect 28825 23477 28859 23511
rect 28859 23477 28868 23511
rect 28816 23468 28868 23477
rect 29644 23468 29696 23520
rect 30380 23511 30432 23520
rect 30380 23477 30389 23511
rect 30389 23477 30423 23511
rect 30423 23477 30432 23511
rect 30380 23468 30432 23477
rect 31392 23511 31444 23520
rect 31392 23477 31401 23511
rect 31401 23477 31435 23511
rect 31435 23477 31444 23511
rect 31392 23468 31444 23477
rect 33232 23468 33284 23520
rect 34336 23468 34388 23520
rect 34520 23511 34572 23520
rect 34520 23477 34529 23511
rect 34529 23477 34563 23511
rect 34563 23477 34572 23511
rect 34520 23468 34572 23477
rect 35256 23468 35308 23520
rect 36084 23468 36136 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 7196 23264 7248 23316
rect 11244 23264 11296 23316
rect 12808 23307 12860 23316
rect 12808 23273 12817 23307
rect 12817 23273 12851 23307
rect 12851 23273 12860 23307
rect 12808 23264 12860 23273
rect 15016 23307 15068 23316
rect 15016 23273 15025 23307
rect 15025 23273 15059 23307
rect 15059 23273 15068 23307
rect 15016 23264 15068 23273
rect 17316 23264 17368 23316
rect 18880 23239 18932 23248
rect 18880 23205 18889 23239
rect 18889 23205 18923 23239
rect 18923 23205 18932 23239
rect 18880 23196 18932 23205
rect 19892 23196 19944 23248
rect 20628 23196 20680 23248
rect 11428 23171 11480 23180
rect 11428 23137 11437 23171
rect 11437 23137 11471 23171
rect 11471 23137 11480 23171
rect 11428 23128 11480 23137
rect 19340 23128 19392 23180
rect 20168 23128 20220 23180
rect 23572 23264 23624 23316
rect 23756 23264 23808 23316
rect 24768 23264 24820 23316
rect 27988 23264 28040 23316
rect 23664 23128 23716 23180
rect 11980 23060 12032 23112
rect 13820 23060 13872 23112
rect 15108 23103 15160 23112
rect 15108 23069 15117 23103
rect 15117 23069 15151 23103
rect 15151 23069 15160 23103
rect 15108 23060 15160 23069
rect 15476 23060 15528 23112
rect 19156 23060 19208 23112
rect 19616 23103 19668 23112
rect 19616 23069 19625 23103
rect 19625 23069 19659 23103
rect 19659 23069 19668 23103
rect 19616 23060 19668 23069
rect 19708 23060 19760 23112
rect 20352 23060 20404 23112
rect 20720 23103 20772 23112
rect 20720 23069 20729 23103
rect 20729 23069 20763 23103
rect 20763 23069 20772 23103
rect 20720 23060 20772 23069
rect 22008 23060 22060 23112
rect 22928 23060 22980 23112
rect 23756 23060 23808 23112
rect 24860 23128 24912 23180
rect 28448 23239 28500 23248
rect 28448 23205 28457 23239
rect 28457 23205 28491 23239
rect 28491 23205 28500 23239
rect 28448 23196 28500 23205
rect 28540 23196 28592 23248
rect 29276 23196 29328 23248
rect 25320 23128 25372 23180
rect 24216 23060 24268 23112
rect 24308 23060 24360 23112
rect 24768 23060 24820 23112
rect 25504 23060 25556 23112
rect 25688 23060 25740 23112
rect 16856 22992 16908 23044
rect 17767 23035 17819 23044
rect 17767 23001 17799 23035
rect 17799 23001 17819 23035
rect 17767 22992 17819 23001
rect 18604 22992 18656 23044
rect 23664 23035 23716 23044
rect 23664 23001 23673 23035
rect 23673 23001 23707 23035
rect 23707 23001 23716 23035
rect 23664 22992 23716 23001
rect 25228 22992 25280 23044
rect 13084 22924 13136 22976
rect 16672 22924 16724 22976
rect 17132 22924 17184 22976
rect 17868 22924 17920 22976
rect 17960 22924 18012 22976
rect 19708 22924 19760 22976
rect 20812 22924 20864 22976
rect 22744 22924 22796 22976
rect 23940 22924 23992 22976
rect 24308 22924 24360 22976
rect 24492 22924 24544 22976
rect 26148 22924 26200 22976
rect 26332 22967 26384 22976
rect 26332 22933 26341 22967
rect 26341 22933 26375 22967
rect 26375 22933 26384 22967
rect 26332 22924 26384 22933
rect 30380 23128 30432 23180
rect 26792 23060 26844 23112
rect 27344 23060 27396 23112
rect 29276 23060 29328 23112
rect 29736 23103 29788 23112
rect 29736 23069 29745 23103
rect 29745 23069 29779 23103
rect 29779 23069 29788 23103
rect 29736 23060 29788 23069
rect 27436 23035 27488 23044
rect 27436 23001 27445 23035
rect 27445 23001 27479 23035
rect 27479 23001 27488 23035
rect 27436 22992 27488 23001
rect 27988 22992 28040 23044
rect 28356 22992 28408 23044
rect 28724 22992 28776 23044
rect 30012 23103 30064 23112
rect 30012 23069 30021 23103
rect 30021 23069 30055 23103
rect 30055 23069 30064 23103
rect 30012 23060 30064 23069
rect 30196 23103 30248 23112
rect 30196 23069 30210 23103
rect 30210 23069 30244 23103
rect 30244 23069 30248 23103
rect 30196 23060 30248 23069
rect 30840 23307 30892 23316
rect 30840 23273 30849 23307
rect 30849 23273 30883 23307
rect 30883 23273 30892 23307
rect 30840 23264 30892 23273
rect 32772 23264 32824 23316
rect 33876 23264 33928 23316
rect 34428 23264 34480 23316
rect 35164 23264 35216 23316
rect 35900 23264 35952 23316
rect 31576 23196 31628 23248
rect 37464 23264 37516 23316
rect 31024 23060 31076 23112
rect 31576 23060 31628 23112
rect 31852 23103 31904 23112
rect 31852 23069 31861 23103
rect 31861 23069 31895 23103
rect 31895 23069 31904 23103
rect 31852 23060 31904 23069
rect 32220 23060 32272 23112
rect 32772 23103 32824 23112
rect 32772 23069 32781 23103
rect 32781 23069 32815 23103
rect 32815 23069 32824 23103
rect 32772 23060 32824 23069
rect 28632 22924 28684 22976
rect 30012 22924 30064 22976
rect 32404 22992 32456 23044
rect 33416 23060 33468 23112
rect 30288 22924 30340 22976
rect 30380 22967 30432 22976
rect 30380 22933 30389 22967
rect 30389 22933 30423 22967
rect 30423 22933 30432 22967
rect 30380 22924 30432 22933
rect 30564 22924 30616 22976
rect 32956 22924 33008 22976
rect 33140 23035 33192 23044
rect 33140 23001 33149 23035
rect 33149 23001 33183 23035
rect 33183 23001 33192 23035
rect 33140 22992 33192 23001
rect 34244 23103 34296 23112
rect 34244 23069 34253 23103
rect 34253 23069 34287 23103
rect 34287 23069 34296 23103
rect 34244 23060 34296 23069
rect 39304 23196 39356 23248
rect 34796 23060 34848 23112
rect 35532 23128 35584 23180
rect 33232 22924 33284 22976
rect 33508 22924 33560 22976
rect 34428 22992 34480 23044
rect 34612 22992 34664 23044
rect 35164 23103 35216 23112
rect 35164 23069 35173 23103
rect 35173 23069 35207 23103
rect 35207 23069 35216 23103
rect 35164 23060 35216 23069
rect 35348 23103 35400 23112
rect 35348 23069 35362 23103
rect 35362 23069 35396 23103
rect 35396 23069 35400 23103
rect 35348 23060 35400 23069
rect 35808 23060 35860 23112
rect 36912 23060 36964 23112
rect 37004 23060 37056 23112
rect 38292 23103 38344 23112
rect 38292 23069 38301 23103
rect 38301 23069 38335 23103
rect 38335 23069 38344 23103
rect 38292 23060 38344 23069
rect 35716 22992 35768 23044
rect 36728 22992 36780 23044
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 15108 22720 15160 22772
rect 13084 22695 13136 22704
rect 13084 22661 13118 22695
rect 13118 22661 13136 22695
rect 13084 22652 13136 22661
rect 14280 22652 14332 22704
rect 16764 22652 16816 22704
rect 18604 22763 18656 22772
rect 18604 22729 18613 22763
rect 18613 22729 18647 22763
rect 18647 22729 18656 22763
rect 18604 22720 18656 22729
rect 19340 22720 19392 22772
rect 20444 22763 20496 22772
rect 20444 22729 20453 22763
rect 20453 22729 20487 22763
rect 20487 22729 20496 22763
rect 20444 22720 20496 22729
rect 22560 22720 22612 22772
rect 20352 22652 20404 22704
rect 24492 22720 24544 22772
rect 12900 22584 12952 22636
rect 15292 22584 15344 22636
rect 16212 22584 16264 22636
rect 16488 22584 16540 22636
rect 16580 22584 16632 22636
rect 15568 22559 15620 22568
rect 15568 22525 15577 22559
rect 15577 22525 15611 22559
rect 15611 22525 15620 22559
rect 15568 22516 15620 22525
rect 15844 22516 15896 22568
rect 17500 22627 17552 22636
rect 17500 22593 17509 22627
rect 17509 22593 17543 22627
rect 17543 22593 17552 22627
rect 17500 22584 17552 22593
rect 17316 22516 17368 22568
rect 18696 22584 18748 22636
rect 19156 22584 19208 22636
rect 20720 22584 20772 22636
rect 24216 22652 24268 22704
rect 27068 22720 27120 22772
rect 27344 22763 27396 22772
rect 27344 22729 27353 22763
rect 27353 22729 27387 22763
rect 27387 22729 27396 22763
rect 27344 22720 27396 22729
rect 27528 22720 27580 22772
rect 28632 22763 28684 22772
rect 28632 22729 28641 22763
rect 28641 22729 28675 22763
rect 28675 22729 28684 22763
rect 28632 22720 28684 22729
rect 29092 22720 29144 22772
rect 30472 22720 30524 22772
rect 17868 22516 17920 22568
rect 18788 22516 18840 22568
rect 13452 22380 13504 22432
rect 17408 22448 17460 22500
rect 17960 22448 18012 22500
rect 22192 22627 22244 22636
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 22284 22584 22336 22636
rect 22744 22584 22796 22636
rect 24032 22584 24084 22636
rect 25228 22584 25280 22636
rect 30380 22652 30432 22704
rect 25964 22627 26016 22636
rect 25964 22593 25973 22627
rect 25973 22593 26007 22627
rect 26007 22593 26016 22627
rect 25964 22584 26016 22593
rect 26056 22584 26108 22636
rect 16672 22380 16724 22432
rect 19524 22380 19576 22432
rect 22284 22491 22336 22500
rect 22284 22457 22293 22491
rect 22293 22457 22327 22491
rect 22327 22457 22336 22491
rect 22284 22448 22336 22457
rect 22836 22559 22888 22568
rect 22836 22525 22845 22559
rect 22845 22525 22879 22559
rect 22879 22525 22888 22559
rect 22836 22516 22888 22525
rect 23296 22516 23348 22568
rect 25688 22516 25740 22568
rect 26608 22584 26660 22636
rect 27160 22584 27212 22636
rect 27620 22584 27672 22636
rect 28264 22627 28316 22636
rect 28264 22593 28273 22627
rect 28273 22593 28307 22627
rect 28307 22593 28316 22627
rect 28264 22584 28316 22593
rect 24676 22448 24728 22500
rect 25412 22491 25464 22500
rect 25412 22457 25421 22491
rect 25421 22457 25455 22491
rect 25455 22457 25464 22491
rect 25412 22448 25464 22457
rect 25596 22448 25648 22500
rect 26056 22448 26108 22500
rect 26884 22516 26936 22568
rect 27068 22516 27120 22568
rect 28724 22584 28776 22636
rect 23296 22380 23348 22432
rect 23664 22380 23716 22432
rect 24860 22380 24912 22432
rect 27068 22380 27120 22432
rect 28448 22448 28500 22500
rect 29460 22584 29512 22636
rect 29644 22584 29696 22636
rect 30840 22627 30892 22636
rect 30840 22593 30849 22627
rect 30849 22593 30883 22627
rect 30883 22593 30892 22627
rect 30840 22584 30892 22593
rect 31300 22652 31352 22704
rect 31576 22652 31628 22704
rect 32680 22652 32732 22704
rect 36360 22720 36412 22772
rect 34152 22652 34204 22704
rect 35164 22652 35216 22704
rect 35532 22652 35584 22704
rect 32772 22627 32824 22636
rect 32772 22593 32779 22627
rect 32779 22593 32813 22627
rect 32813 22593 32824 22627
rect 32772 22584 32824 22593
rect 33140 22584 33192 22636
rect 33876 22627 33928 22636
rect 33876 22593 33886 22627
rect 33886 22593 33920 22627
rect 33920 22593 33928 22627
rect 33876 22584 33928 22593
rect 33968 22627 34020 22636
rect 33968 22593 33978 22627
rect 33978 22593 34012 22627
rect 34012 22593 34020 22627
rect 33968 22584 34020 22593
rect 30932 22516 30984 22568
rect 31300 22559 31352 22568
rect 31300 22525 31309 22559
rect 31309 22525 31343 22559
rect 31343 22525 31352 22559
rect 31300 22516 31352 22525
rect 31392 22516 31444 22568
rect 33600 22516 33652 22568
rect 35348 22627 35400 22636
rect 35348 22593 35357 22627
rect 35357 22593 35391 22627
rect 35391 22593 35400 22627
rect 35348 22584 35400 22593
rect 34428 22516 34480 22568
rect 35716 22627 35768 22636
rect 35716 22593 35725 22627
rect 35725 22593 35759 22627
rect 35759 22593 35768 22627
rect 35716 22584 35768 22593
rect 37004 22584 37056 22636
rect 37464 22627 37516 22636
rect 37464 22593 37473 22627
rect 37473 22593 37507 22627
rect 37507 22593 37516 22627
rect 37464 22584 37516 22593
rect 35624 22516 35676 22568
rect 35900 22516 35952 22568
rect 36728 22559 36780 22568
rect 36728 22525 36737 22559
rect 36737 22525 36771 22559
rect 36771 22525 36780 22559
rect 36728 22516 36780 22525
rect 29552 22448 29604 22500
rect 29276 22380 29328 22432
rect 32220 22380 32272 22432
rect 34520 22448 34572 22500
rect 37924 22448 37976 22500
rect 33324 22380 33376 22432
rect 36176 22380 36228 22432
rect 36544 22380 36596 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 17316 22219 17368 22228
rect 17316 22185 17325 22219
rect 17325 22185 17359 22219
rect 17359 22185 17368 22219
rect 17316 22176 17368 22185
rect 18788 22219 18840 22228
rect 18788 22185 18797 22219
rect 18797 22185 18831 22219
rect 18831 22185 18840 22219
rect 18788 22176 18840 22185
rect 19432 22219 19484 22228
rect 19432 22185 19441 22219
rect 19441 22185 19475 22219
rect 19475 22185 19484 22219
rect 19432 22176 19484 22185
rect 17868 22108 17920 22160
rect 22468 22176 22520 22228
rect 22560 22176 22612 22228
rect 19800 22151 19852 22160
rect 19800 22117 19809 22151
rect 19809 22117 19843 22151
rect 19843 22117 19852 22151
rect 19800 22108 19852 22117
rect 12900 22040 12952 22092
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 15292 22083 15344 22092
rect 15292 22049 15301 22083
rect 15301 22049 15335 22083
rect 15335 22049 15344 22083
rect 15292 22040 15344 22049
rect 15384 22040 15436 22092
rect 17224 22040 17276 22092
rect 19340 22040 19392 22092
rect 11060 21972 11112 22024
rect 14280 21972 14332 22024
rect 14832 22015 14884 22024
rect 14832 21981 14841 22015
rect 14841 21981 14875 22015
rect 14875 21981 14884 22015
rect 14832 21972 14884 21981
rect 15200 21972 15252 22024
rect 15568 21972 15620 22024
rect 18236 21972 18288 22024
rect 19524 21972 19576 22024
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 20168 21972 20220 22024
rect 22284 22108 22336 22160
rect 23204 22108 23256 22160
rect 23848 22176 23900 22228
rect 27344 22176 27396 22228
rect 24768 22108 24820 22160
rect 24860 22151 24912 22160
rect 24860 22117 24869 22151
rect 24869 22117 24903 22151
rect 24903 22117 24912 22151
rect 24860 22108 24912 22117
rect 26516 22151 26568 22160
rect 26516 22117 26525 22151
rect 26525 22117 26559 22151
rect 26559 22117 26568 22151
rect 26516 22108 26568 22117
rect 22836 22040 22888 22092
rect 11796 21904 11848 21956
rect 16764 21904 16816 21956
rect 21088 21904 21140 21956
rect 22744 21972 22796 22024
rect 23388 21972 23440 22024
rect 22192 21904 22244 21956
rect 22284 21904 22336 21956
rect 23940 21972 23992 22024
rect 24768 21972 24820 22024
rect 27068 22040 27120 22092
rect 27896 22176 27948 22228
rect 27988 22176 28040 22228
rect 28632 22108 28684 22160
rect 30012 22176 30064 22228
rect 33140 22176 33192 22228
rect 34428 22176 34480 22228
rect 35624 22176 35676 22228
rect 30840 22108 30892 22160
rect 27804 22083 27856 22092
rect 27804 22049 27813 22083
rect 27813 22049 27847 22083
rect 27847 22049 27856 22083
rect 27804 22040 27856 22049
rect 28540 22083 28592 22092
rect 28540 22049 28563 22083
rect 28563 22049 28592 22083
rect 28540 22040 28592 22049
rect 29552 22040 29604 22092
rect 27528 22015 27580 22024
rect 27528 21981 27537 22015
rect 27537 21981 27571 22015
rect 27571 21981 27580 22015
rect 27528 21972 27580 21981
rect 28080 21972 28132 22024
rect 29000 22015 29052 22024
rect 29000 21981 29009 22015
rect 29009 21981 29043 22015
rect 29043 21981 29052 22015
rect 29000 21972 29052 21981
rect 25412 21904 25464 21956
rect 28448 21904 28500 21956
rect 28540 21904 28592 21956
rect 28908 21947 28960 21956
rect 28908 21913 28917 21947
rect 28917 21913 28951 21947
rect 28951 21913 28960 21947
rect 28908 21904 28960 21913
rect 30104 21972 30156 22024
rect 31024 22015 31076 22024
rect 31024 21981 31033 22015
rect 31033 21981 31067 22015
rect 31067 21981 31076 22015
rect 31024 21972 31076 21981
rect 31116 22015 31168 22024
rect 31116 21981 31126 22015
rect 31126 21981 31160 22015
rect 31160 21981 31168 22015
rect 31116 21972 31168 21981
rect 32496 22108 32548 22160
rect 32956 22108 33008 22160
rect 33416 22108 33468 22160
rect 34888 22108 34940 22160
rect 38844 22176 38896 22228
rect 31484 22015 31536 22024
rect 31484 21981 31498 22015
rect 31498 21981 31532 22015
rect 31532 21981 31536 22015
rect 31484 21972 31536 21981
rect 32312 22015 32364 22024
rect 32312 21981 32319 22015
rect 32319 21981 32364 22015
rect 32312 21972 32364 21981
rect 33784 22083 33836 22092
rect 33784 22049 33793 22083
rect 33793 22049 33827 22083
rect 33827 22049 33836 22083
rect 33784 22040 33836 22049
rect 33876 22083 33928 22092
rect 33876 22049 33885 22083
rect 33885 22049 33919 22083
rect 33919 22049 33928 22083
rect 33876 22040 33928 22049
rect 34152 22040 34204 22092
rect 32680 21972 32732 22024
rect 32772 21972 32824 22024
rect 33232 21972 33284 22024
rect 33416 22015 33468 22024
rect 33416 21981 33425 22015
rect 33425 21981 33459 22015
rect 33459 21981 33468 22015
rect 33416 21972 33468 21981
rect 33692 21972 33744 22024
rect 33968 21972 34020 22024
rect 34796 21972 34848 22024
rect 35072 22015 35124 22024
rect 35072 21981 35079 22015
rect 35079 21981 35124 22015
rect 35072 21972 35124 21981
rect 35532 22040 35584 22092
rect 36912 22083 36964 22092
rect 36912 22049 36921 22083
rect 36921 22049 36955 22083
rect 36955 22049 36964 22083
rect 36912 22040 36964 22049
rect 35808 21972 35860 22024
rect 35992 22015 36044 22024
rect 35992 21981 36001 22015
rect 36001 21981 36035 22015
rect 36035 21981 36044 22015
rect 35992 21972 36044 21981
rect 30380 21904 30432 21956
rect 30564 21904 30616 21956
rect 12348 21879 12400 21888
rect 12348 21845 12357 21879
rect 12357 21845 12391 21879
rect 12391 21845 12400 21879
rect 12348 21836 12400 21845
rect 13084 21836 13136 21888
rect 18144 21836 18196 21888
rect 18604 21836 18656 21888
rect 22376 21836 22428 21888
rect 23204 21836 23256 21888
rect 24124 21836 24176 21888
rect 24216 21836 24268 21888
rect 26424 21836 26476 21888
rect 28264 21836 28316 21888
rect 28356 21879 28408 21888
rect 28356 21845 28365 21879
rect 28365 21845 28399 21879
rect 28399 21845 28408 21879
rect 28356 21836 28408 21845
rect 29000 21836 29052 21888
rect 31576 21836 31628 21888
rect 32036 21836 32088 21888
rect 32128 21836 32180 21888
rect 32772 21879 32824 21888
rect 32772 21845 32781 21879
rect 32781 21845 32815 21879
rect 32815 21845 32824 21879
rect 32772 21836 32824 21845
rect 35256 21947 35308 21956
rect 35256 21913 35265 21947
rect 35265 21913 35299 21947
rect 35299 21913 35308 21947
rect 35256 21904 35308 21913
rect 37188 21947 37240 21956
rect 37188 21913 37222 21947
rect 37222 21913 37240 21947
rect 37188 21904 37240 21913
rect 37556 21972 37608 22024
rect 38292 21972 38344 22024
rect 38200 21836 38252 21888
rect 38292 21879 38344 21888
rect 38292 21845 38301 21879
rect 38301 21845 38335 21879
rect 38335 21845 38344 21879
rect 38292 21836 38344 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 11796 21675 11848 21684
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 12164 21632 12216 21684
rect 15844 21632 15896 21684
rect 18236 21675 18288 21684
rect 18236 21641 18245 21675
rect 18245 21641 18279 21675
rect 18279 21641 18288 21675
rect 18236 21632 18288 21641
rect 12348 21564 12400 21616
rect 13820 21564 13872 21616
rect 14280 21564 14332 21616
rect 17960 21564 18012 21616
rect 19248 21632 19300 21684
rect 20260 21675 20312 21684
rect 20260 21641 20269 21675
rect 20269 21641 20303 21675
rect 20303 21641 20312 21675
rect 20260 21632 20312 21641
rect 20628 21632 20680 21684
rect 22192 21632 22244 21684
rect 23388 21632 23440 21684
rect 23848 21675 23900 21684
rect 23848 21641 23857 21675
rect 23857 21641 23891 21675
rect 23891 21641 23900 21675
rect 23848 21632 23900 21641
rect 23940 21675 23992 21684
rect 23940 21641 23949 21675
rect 23949 21641 23983 21675
rect 23983 21641 23992 21675
rect 23940 21632 23992 21641
rect 24400 21632 24452 21684
rect 26608 21632 26660 21684
rect 27160 21632 27212 21684
rect 28080 21675 28132 21684
rect 28080 21641 28089 21675
rect 28089 21641 28123 21675
rect 28123 21641 28132 21675
rect 28080 21632 28132 21641
rect 19156 21564 19208 21616
rect 12256 21428 12308 21480
rect 5172 21360 5224 21412
rect 13084 21360 13136 21412
rect 6920 21292 6972 21344
rect 11060 21292 11112 21344
rect 13636 21496 13688 21548
rect 14832 21496 14884 21548
rect 13452 21471 13504 21480
rect 13452 21437 13461 21471
rect 13461 21437 13495 21471
rect 13495 21437 13504 21471
rect 13452 21428 13504 21437
rect 15568 21539 15620 21548
rect 15568 21505 15577 21539
rect 15577 21505 15611 21539
rect 15611 21505 15620 21539
rect 15568 21496 15620 21505
rect 20996 21564 21048 21616
rect 15660 21428 15712 21480
rect 16764 21428 16816 21480
rect 20076 21496 20128 21548
rect 22744 21564 22796 21616
rect 24124 21607 24176 21616
rect 24124 21573 24133 21607
rect 24133 21573 24167 21607
rect 24167 21573 24176 21607
rect 24124 21564 24176 21573
rect 25596 21564 25648 21616
rect 26148 21607 26200 21616
rect 26148 21573 26157 21607
rect 26157 21573 26191 21607
rect 26191 21573 26200 21607
rect 26148 21564 26200 21573
rect 29000 21632 29052 21684
rect 29828 21632 29880 21684
rect 30012 21632 30064 21684
rect 31024 21632 31076 21684
rect 18512 21428 18564 21480
rect 19156 21428 19208 21480
rect 21456 21539 21508 21548
rect 21456 21505 21465 21539
rect 21465 21505 21499 21539
rect 21499 21505 21508 21539
rect 21456 21496 21508 21505
rect 22284 21539 22336 21548
rect 22284 21505 22293 21539
rect 22293 21505 22327 21539
rect 22327 21505 22336 21539
rect 22284 21496 22336 21505
rect 22376 21539 22428 21548
rect 22376 21505 22385 21539
rect 22385 21505 22419 21539
rect 22419 21505 22428 21539
rect 22376 21496 22428 21505
rect 22560 21496 22612 21548
rect 18696 21360 18748 21412
rect 20444 21360 20496 21412
rect 21088 21428 21140 21480
rect 23572 21496 23624 21548
rect 23756 21539 23808 21548
rect 23756 21505 23765 21539
rect 23765 21505 23799 21539
rect 23799 21505 23808 21539
rect 23756 21496 23808 21505
rect 24492 21496 24544 21548
rect 25044 21496 25096 21548
rect 25412 21496 25464 21548
rect 24308 21428 24360 21480
rect 25596 21428 25648 21480
rect 25872 21428 25924 21480
rect 26884 21496 26936 21548
rect 27068 21496 27120 21548
rect 28632 21564 28684 21616
rect 28448 21539 28500 21548
rect 28448 21505 28457 21539
rect 28457 21505 28491 21539
rect 28491 21505 28500 21539
rect 28448 21496 28500 21505
rect 28540 21539 28592 21548
rect 28540 21505 28549 21539
rect 28549 21505 28583 21539
rect 28583 21505 28592 21539
rect 28540 21496 28592 21505
rect 26056 21428 26108 21480
rect 21640 21360 21692 21412
rect 22744 21360 22796 21412
rect 22836 21360 22888 21412
rect 27160 21428 27212 21480
rect 27804 21428 27856 21480
rect 28264 21471 28316 21480
rect 28264 21437 28273 21471
rect 28273 21437 28307 21471
rect 28307 21437 28316 21471
rect 29276 21564 29328 21616
rect 30196 21564 30248 21616
rect 30288 21607 30340 21616
rect 30288 21573 30297 21607
rect 30297 21573 30331 21607
rect 30331 21573 30340 21607
rect 30288 21564 30340 21573
rect 29000 21496 29052 21548
rect 29184 21496 29236 21548
rect 28264 21428 28316 21437
rect 28816 21428 28868 21480
rect 15568 21292 15620 21344
rect 17776 21292 17828 21344
rect 19984 21292 20036 21344
rect 20076 21335 20128 21344
rect 20076 21301 20085 21335
rect 20085 21301 20119 21335
rect 20119 21301 20128 21335
rect 20076 21292 20128 21301
rect 20168 21292 20220 21344
rect 20536 21292 20588 21344
rect 20628 21335 20680 21344
rect 20628 21301 20637 21335
rect 20637 21301 20671 21335
rect 20671 21301 20680 21335
rect 20628 21292 20680 21301
rect 22008 21335 22060 21344
rect 22008 21301 22017 21335
rect 22017 21301 22051 21335
rect 22051 21301 22060 21335
rect 22008 21292 22060 21301
rect 22468 21292 22520 21344
rect 24584 21335 24636 21344
rect 24584 21301 24593 21335
rect 24593 21301 24627 21335
rect 24627 21301 24636 21335
rect 24584 21292 24636 21301
rect 26516 21335 26568 21344
rect 26516 21301 26525 21335
rect 26525 21301 26559 21335
rect 26559 21301 26568 21335
rect 26516 21292 26568 21301
rect 29000 21360 29052 21412
rect 29460 21428 29512 21480
rect 30656 21496 30708 21548
rect 32128 21564 32180 21616
rect 31116 21539 31168 21548
rect 31116 21505 31125 21539
rect 31125 21505 31159 21539
rect 31159 21505 31168 21539
rect 31116 21496 31168 21505
rect 31392 21496 31444 21548
rect 32496 21607 32548 21616
rect 32496 21573 32505 21607
rect 32505 21573 32539 21607
rect 32539 21573 32548 21607
rect 32496 21564 32548 21573
rect 33324 21632 33376 21684
rect 34612 21632 34664 21684
rect 37188 21632 37240 21684
rect 38292 21632 38344 21684
rect 32312 21539 32364 21548
rect 32312 21505 32321 21539
rect 32321 21505 32355 21539
rect 32355 21505 32364 21539
rect 32312 21496 32364 21505
rect 32680 21539 32732 21548
rect 32680 21505 32689 21539
rect 32689 21505 32723 21539
rect 32723 21505 32732 21539
rect 32680 21496 32732 21505
rect 32772 21496 32824 21548
rect 33600 21496 33652 21548
rect 34520 21539 34572 21548
rect 34520 21505 34529 21539
rect 34529 21505 34563 21539
rect 34563 21505 34572 21539
rect 34520 21496 34572 21505
rect 35256 21564 35308 21616
rect 35440 21564 35492 21616
rect 26976 21292 27028 21344
rect 27528 21292 27580 21344
rect 28448 21292 28500 21344
rect 29552 21292 29604 21344
rect 30472 21360 30524 21412
rect 30748 21360 30800 21412
rect 34428 21428 34480 21480
rect 34704 21428 34756 21480
rect 34888 21539 34940 21548
rect 34888 21505 34897 21539
rect 34897 21505 34931 21539
rect 34931 21505 34940 21539
rect 34888 21496 34940 21505
rect 35348 21496 35400 21548
rect 36084 21564 36136 21616
rect 36452 21539 36504 21548
rect 36452 21505 36461 21539
rect 36461 21505 36495 21539
rect 36495 21505 36504 21539
rect 36452 21496 36504 21505
rect 37648 21496 37700 21548
rect 38936 21496 38988 21548
rect 37924 21471 37976 21480
rect 37924 21437 37933 21471
rect 37933 21437 37967 21471
rect 37967 21437 37976 21471
rect 37924 21428 37976 21437
rect 38108 21471 38160 21480
rect 38108 21437 38117 21471
rect 38117 21437 38151 21471
rect 38151 21437 38160 21471
rect 38108 21428 38160 21437
rect 32588 21360 32640 21412
rect 30196 21292 30248 21344
rect 31208 21292 31260 21344
rect 31576 21292 31628 21344
rect 32312 21292 32364 21344
rect 33508 21335 33560 21344
rect 33508 21301 33517 21335
rect 33517 21301 33551 21335
rect 33551 21301 33560 21335
rect 33508 21292 33560 21301
rect 33968 21292 34020 21344
rect 34060 21292 34112 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 13636 21131 13688 21140
rect 13636 21097 13645 21131
rect 13645 21097 13679 21131
rect 13679 21097 13688 21131
rect 13636 21088 13688 21097
rect 16764 21020 16816 21072
rect 11244 20927 11296 20936
rect 11244 20893 11253 20927
rect 11253 20893 11287 20927
rect 11287 20893 11296 20927
rect 11244 20884 11296 20893
rect 12624 20884 12676 20936
rect 15292 20952 15344 21004
rect 15476 20995 15528 21004
rect 15476 20961 15485 20995
rect 15485 20961 15519 20995
rect 15519 20961 15528 20995
rect 15476 20952 15528 20961
rect 15016 20927 15068 20936
rect 15016 20893 15025 20927
rect 15025 20893 15059 20927
rect 15059 20893 15068 20927
rect 15016 20884 15068 20893
rect 15200 20884 15252 20936
rect 22008 21088 22060 21140
rect 22560 21131 22612 21140
rect 22560 21097 22569 21131
rect 22569 21097 22603 21131
rect 22603 21097 22612 21131
rect 22560 21088 22612 21097
rect 23756 21088 23808 21140
rect 25688 21088 25740 21140
rect 25872 21088 25924 21140
rect 26056 21088 26108 21140
rect 26976 21088 27028 21140
rect 30564 21088 30616 21140
rect 19156 21020 19208 21072
rect 19248 21020 19300 21072
rect 19984 21020 20036 21072
rect 15568 20816 15620 20868
rect 17132 20859 17184 20868
rect 17132 20825 17141 20859
rect 17141 20825 17175 20859
rect 17175 20825 17184 20859
rect 17132 20816 17184 20825
rect 19248 20884 19300 20936
rect 19340 20884 19392 20936
rect 20168 20884 20220 20936
rect 20628 21020 20680 21072
rect 23296 21020 23348 21072
rect 20444 20952 20496 21004
rect 22100 20952 22152 21004
rect 22192 20952 22244 21004
rect 22928 20952 22980 21004
rect 21088 20884 21140 20936
rect 21456 20884 21508 20936
rect 24216 20952 24268 21004
rect 25228 20995 25280 21004
rect 25228 20961 25237 20995
rect 25237 20961 25271 20995
rect 25271 20961 25280 20995
rect 25228 20952 25280 20961
rect 27620 21020 27672 21072
rect 29276 21020 29328 21072
rect 26240 20952 26292 21004
rect 22100 20816 22152 20868
rect 22652 20816 22704 20868
rect 23388 20927 23440 20936
rect 23388 20893 23397 20927
rect 23397 20893 23431 20927
rect 23431 20893 23440 20927
rect 23388 20884 23440 20893
rect 23480 20927 23532 20936
rect 23480 20893 23489 20927
rect 23489 20893 23523 20927
rect 23523 20893 23532 20927
rect 23480 20884 23532 20893
rect 26700 20884 26752 20936
rect 27804 20952 27856 21004
rect 29552 20952 29604 21004
rect 30012 20952 30064 21004
rect 24676 20816 24728 20868
rect 25872 20816 25924 20868
rect 17776 20791 17828 20800
rect 17776 20757 17785 20791
rect 17785 20757 17819 20791
rect 17819 20757 17828 20791
rect 17776 20748 17828 20757
rect 18512 20791 18564 20800
rect 18512 20757 18521 20791
rect 18521 20757 18555 20791
rect 18555 20757 18564 20791
rect 18512 20748 18564 20757
rect 22928 20748 22980 20800
rect 24860 20748 24912 20800
rect 24952 20791 25004 20800
rect 24952 20757 24961 20791
rect 24961 20757 24995 20791
rect 24995 20757 25004 20791
rect 24952 20748 25004 20757
rect 25044 20791 25096 20800
rect 25044 20757 25053 20791
rect 25053 20757 25087 20791
rect 25087 20757 25096 20791
rect 25044 20748 25096 20757
rect 25320 20748 25372 20800
rect 25964 20791 26016 20800
rect 25964 20757 25989 20791
rect 25989 20757 26016 20791
rect 25964 20748 26016 20757
rect 26700 20748 26752 20800
rect 28816 20884 28868 20936
rect 29460 20884 29512 20936
rect 27344 20816 27396 20868
rect 30380 20952 30432 21004
rect 31484 20952 31536 21004
rect 30564 20884 30616 20936
rect 31300 20884 31352 20936
rect 32036 20952 32088 21004
rect 32220 20927 32272 20936
rect 32220 20893 32229 20927
rect 32229 20893 32263 20927
rect 32263 20893 32272 20927
rect 32220 20884 32272 20893
rect 32312 20927 32364 20936
rect 32312 20893 32321 20927
rect 32321 20893 32355 20927
rect 32355 20893 32364 20927
rect 32312 20884 32364 20893
rect 32588 20884 32640 20936
rect 30748 20816 30800 20868
rect 31116 20859 31168 20868
rect 31116 20825 31125 20859
rect 31125 20825 31159 20859
rect 31159 20825 31168 20859
rect 31116 20816 31168 20825
rect 26976 20791 27028 20800
rect 26976 20757 26985 20791
rect 26985 20757 27019 20791
rect 27019 20757 27028 20791
rect 26976 20748 27028 20757
rect 27712 20791 27764 20800
rect 27712 20757 27721 20791
rect 27721 20757 27755 20791
rect 27755 20757 27764 20791
rect 27712 20748 27764 20757
rect 28816 20748 28868 20800
rect 32680 20816 32732 20868
rect 33324 21020 33376 21072
rect 33232 20927 33284 20936
rect 33232 20893 33241 20927
rect 33241 20893 33275 20927
rect 33275 20893 33284 20927
rect 33232 20884 33284 20893
rect 33324 20927 33376 20936
rect 33324 20893 33333 20927
rect 33333 20893 33367 20927
rect 33367 20893 33376 20927
rect 33324 20884 33376 20893
rect 37280 21088 37332 21140
rect 34428 20952 34480 21004
rect 34612 20952 34664 21004
rect 35532 20995 35584 21004
rect 35532 20961 35541 20995
rect 35541 20961 35575 20995
rect 35575 20961 35584 20995
rect 35532 20952 35584 20961
rect 34060 20927 34112 20936
rect 34060 20893 34069 20927
rect 34069 20893 34103 20927
rect 34103 20893 34112 20927
rect 34060 20884 34112 20893
rect 34152 20884 34204 20936
rect 35256 20884 35308 20936
rect 31300 20791 31352 20800
rect 31300 20757 31309 20791
rect 31309 20757 31343 20791
rect 31343 20757 31352 20791
rect 31300 20748 31352 20757
rect 31944 20791 31996 20800
rect 31944 20757 31953 20791
rect 31953 20757 31987 20791
rect 31987 20757 31996 20791
rect 31944 20748 31996 20757
rect 32956 20748 33008 20800
rect 35716 20816 35768 20868
rect 36360 20884 36412 20936
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 12440 20544 12492 20596
rect 15016 20544 15068 20596
rect 15108 20544 15160 20596
rect 16212 20587 16264 20596
rect 16212 20553 16221 20587
rect 16221 20553 16255 20587
rect 16255 20553 16264 20587
rect 16212 20544 16264 20553
rect 16948 20544 17000 20596
rect 17040 20544 17092 20596
rect 15752 20476 15804 20528
rect 15292 20408 15344 20460
rect 13268 20383 13320 20392
rect 13268 20349 13277 20383
rect 13277 20349 13311 20383
rect 13311 20349 13320 20383
rect 13268 20340 13320 20349
rect 13452 20340 13504 20392
rect 15016 20340 15068 20392
rect 15476 20383 15528 20392
rect 15476 20349 15485 20383
rect 15485 20349 15519 20383
rect 15519 20349 15528 20383
rect 15476 20340 15528 20349
rect 15568 20340 15620 20392
rect 16580 20408 16632 20460
rect 16948 20408 17000 20460
rect 17500 20408 17552 20460
rect 17776 20451 17828 20460
rect 17776 20417 17785 20451
rect 17785 20417 17819 20451
rect 17819 20417 17828 20451
rect 17776 20408 17828 20417
rect 20536 20544 20588 20596
rect 20720 20544 20772 20596
rect 22284 20544 22336 20596
rect 23848 20544 23900 20596
rect 25228 20544 25280 20596
rect 18512 20476 18564 20528
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 20260 20408 20312 20460
rect 21272 20451 21324 20460
rect 21272 20417 21281 20451
rect 21281 20417 21315 20451
rect 21315 20417 21324 20451
rect 21272 20408 21324 20417
rect 21456 20451 21508 20460
rect 21456 20417 21465 20451
rect 21465 20417 21499 20451
rect 21499 20417 21508 20451
rect 21456 20408 21508 20417
rect 22192 20408 22244 20460
rect 22468 20451 22520 20460
rect 22468 20417 22477 20451
rect 22477 20417 22511 20451
rect 22511 20417 22520 20451
rect 22468 20408 22520 20417
rect 22744 20451 22796 20460
rect 22744 20417 22753 20451
rect 22753 20417 22787 20451
rect 22787 20417 22796 20451
rect 22744 20408 22796 20417
rect 22836 20451 22888 20460
rect 22836 20417 22845 20451
rect 22845 20417 22879 20451
rect 22879 20417 22888 20451
rect 22836 20408 22888 20417
rect 23112 20451 23164 20460
rect 23112 20417 23121 20451
rect 23121 20417 23155 20451
rect 23155 20417 23164 20451
rect 23112 20408 23164 20417
rect 23296 20451 23348 20460
rect 23296 20417 23305 20451
rect 23305 20417 23339 20451
rect 23339 20417 23348 20451
rect 23296 20408 23348 20417
rect 23664 20408 23716 20460
rect 20076 20340 20128 20392
rect 12348 20272 12400 20324
rect 14004 20272 14056 20324
rect 19432 20315 19484 20324
rect 19432 20281 19441 20315
rect 19441 20281 19475 20315
rect 19475 20281 19484 20315
rect 19432 20272 19484 20281
rect 20168 20315 20220 20324
rect 20168 20281 20177 20315
rect 20177 20281 20211 20315
rect 20211 20281 20220 20315
rect 20168 20272 20220 20281
rect 20904 20340 20956 20392
rect 20996 20340 21048 20392
rect 25412 20476 25464 20528
rect 25964 20476 26016 20528
rect 25688 20408 25740 20460
rect 26240 20476 26292 20528
rect 28356 20519 28408 20528
rect 28356 20485 28365 20519
rect 28365 20485 28399 20519
rect 28399 20485 28408 20519
rect 28356 20476 28408 20485
rect 28540 20587 28592 20596
rect 28540 20553 28549 20587
rect 28549 20553 28583 20587
rect 28583 20553 28592 20587
rect 28540 20544 28592 20553
rect 30748 20544 30800 20596
rect 33324 20544 33376 20596
rect 33784 20544 33836 20596
rect 35808 20544 35860 20596
rect 36268 20544 36320 20596
rect 28908 20476 28960 20528
rect 27068 20408 27120 20460
rect 14648 20204 14700 20256
rect 15108 20204 15160 20256
rect 15292 20247 15344 20256
rect 15292 20213 15301 20247
rect 15301 20213 15335 20247
rect 15335 20213 15344 20247
rect 15292 20204 15344 20213
rect 16028 20247 16080 20256
rect 16028 20213 16037 20247
rect 16037 20213 16071 20247
rect 16071 20213 16080 20247
rect 16028 20204 16080 20213
rect 17224 20247 17276 20256
rect 17224 20213 17233 20247
rect 17233 20213 17267 20247
rect 17267 20213 17276 20247
rect 17224 20204 17276 20213
rect 17500 20204 17552 20256
rect 19340 20204 19392 20256
rect 20076 20204 20128 20256
rect 22100 20315 22152 20324
rect 22100 20281 22109 20315
rect 22109 20281 22143 20315
rect 22143 20281 22152 20315
rect 22100 20272 22152 20281
rect 25228 20340 25280 20392
rect 26332 20340 26384 20392
rect 26608 20340 26660 20392
rect 27436 20340 27488 20392
rect 27988 20340 28040 20392
rect 28724 20408 28776 20460
rect 29276 20451 29328 20460
rect 29276 20417 29285 20451
rect 29285 20417 29319 20451
rect 29319 20417 29328 20451
rect 29276 20408 29328 20417
rect 30380 20476 30432 20528
rect 28540 20340 28592 20392
rect 29368 20383 29420 20392
rect 29368 20349 29377 20383
rect 29377 20349 29411 20383
rect 29411 20349 29420 20383
rect 29368 20340 29420 20349
rect 29736 20340 29788 20392
rect 30656 20451 30708 20460
rect 30656 20417 30665 20451
rect 30665 20417 30699 20451
rect 30699 20417 30708 20451
rect 30656 20408 30708 20417
rect 30748 20340 30800 20392
rect 26516 20272 26568 20324
rect 27896 20272 27948 20324
rect 28356 20315 28408 20324
rect 28356 20281 28365 20315
rect 28365 20281 28399 20315
rect 28399 20281 28408 20315
rect 28356 20272 28408 20281
rect 31392 20340 31444 20392
rect 31852 20340 31904 20392
rect 21272 20204 21324 20256
rect 22192 20204 22244 20256
rect 22468 20204 22520 20256
rect 27528 20204 27580 20256
rect 31484 20272 31536 20324
rect 29644 20247 29696 20256
rect 29644 20213 29653 20247
rect 29653 20213 29687 20247
rect 29687 20213 29696 20247
rect 29644 20204 29696 20213
rect 30840 20204 30892 20256
rect 32404 20272 32456 20324
rect 31852 20204 31904 20256
rect 32680 20451 32732 20460
rect 32680 20417 32689 20451
rect 32689 20417 32723 20451
rect 32723 20417 32732 20451
rect 32680 20408 32732 20417
rect 33140 20408 33192 20460
rect 33324 20408 33376 20460
rect 33784 20408 33836 20460
rect 34060 20408 34112 20460
rect 34152 20451 34204 20460
rect 34152 20417 34161 20451
rect 34161 20417 34195 20451
rect 34195 20417 34204 20451
rect 34152 20408 34204 20417
rect 32956 20340 33008 20392
rect 33232 20340 33284 20392
rect 34428 20408 34480 20460
rect 34980 20451 35032 20460
rect 34980 20417 34989 20451
rect 34989 20417 35023 20451
rect 35023 20417 35032 20451
rect 34980 20408 35032 20417
rect 35624 20408 35676 20460
rect 35256 20340 35308 20392
rect 35716 20340 35768 20392
rect 32864 20272 32916 20324
rect 35992 20408 36044 20460
rect 36452 20408 36504 20460
rect 37372 20476 37424 20528
rect 37832 20451 37884 20460
rect 37832 20417 37841 20451
rect 37841 20417 37875 20451
rect 37875 20417 37884 20451
rect 37832 20408 37884 20417
rect 36084 20383 36136 20392
rect 36084 20349 36093 20383
rect 36093 20349 36127 20383
rect 36127 20349 36136 20383
rect 36084 20340 36136 20349
rect 38016 20476 38068 20528
rect 38108 20383 38160 20392
rect 38108 20349 38117 20383
rect 38117 20349 38151 20383
rect 38151 20349 38160 20383
rect 38108 20340 38160 20349
rect 32956 20247 33008 20256
rect 32956 20213 32965 20247
rect 32965 20213 32999 20247
rect 32999 20213 33008 20247
rect 32956 20204 33008 20213
rect 33140 20204 33192 20256
rect 33416 20204 33468 20256
rect 34428 20204 34480 20256
rect 36176 20204 36228 20256
rect 37464 20247 37516 20256
rect 37464 20213 37473 20247
rect 37473 20213 37507 20247
rect 37507 20213 37516 20247
rect 37464 20204 37516 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 12624 20043 12676 20052
rect 12624 20009 12633 20043
rect 12633 20009 12667 20043
rect 12667 20009 12676 20043
rect 12624 20000 12676 20009
rect 13268 20043 13320 20052
rect 13268 20009 13277 20043
rect 13277 20009 13311 20043
rect 13311 20009 13320 20043
rect 13268 20000 13320 20009
rect 14740 20000 14792 20052
rect 15476 20000 15528 20052
rect 16580 20043 16632 20052
rect 16580 20009 16589 20043
rect 16589 20009 16623 20043
rect 16623 20009 16632 20043
rect 16580 20000 16632 20009
rect 20444 20043 20496 20052
rect 20444 20009 20453 20043
rect 20453 20009 20487 20043
rect 20487 20009 20496 20043
rect 20444 20000 20496 20009
rect 23296 20000 23348 20052
rect 23480 20000 23532 20052
rect 24032 20000 24084 20052
rect 26608 20000 26660 20052
rect 11244 19839 11296 19848
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 12348 19796 12400 19848
rect 16028 19932 16080 19984
rect 15292 19864 15344 19916
rect 14740 19839 14792 19848
rect 14740 19805 14749 19839
rect 14749 19805 14783 19839
rect 14783 19805 14792 19839
rect 14740 19796 14792 19805
rect 14924 19796 14976 19848
rect 14464 19728 14516 19780
rect 15108 19839 15160 19848
rect 15108 19805 15117 19839
rect 15117 19805 15151 19839
rect 15151 19805 15160 19839
rect 18052 19864 18104 19916
rect 19984 19975 20036 19984
rect 19984 19941 19993 19975
rect 19993 19941 20027 19975
rect 20027 19941 20036 19975
rect 19984 19932 20036 19941
rect 20260 19932 20312 19984
rect 20812 19932 20864 19984
rect 20904 19932 20956 19984
rect 21640 19932 21692 19984
rect 21732 19864 21784 19916
rect 15108 19796 15160 19805
rect 15660 19796 15712 19848
rect 16672 19796 16724 19848
rect 17960 19839 18012 19848
rect 17960 19805 17969 19839
rect 17969 19805 18003 19839
rect 18003 19805 18012 19839
rect 17960 19796 18012 19805
rect 20536 19796 20588 19848
rect 20720 19839 20772 19848
rect 20720 19805 20729 19839
rect 20729 19805 20763 19839
rect 20763 19805 20772 19839
rect 20720 19796 20772 19805
rect 20812 19839 20864 19848
rect 20812 19805 20821 19839
rect 20821 19805 20855 19839
rect 20855 19805 20864 19839
rect 20812 19796 20864 19805
rect 20904 19839 20956 19848
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 22744 19932 22796 19984
rect 22008 19864 22060 19916
rect 15752 19728 15804 19780
rect 15936 19660 15988 19712
rect 16488 19660 16540 19712
rect 18052 19660 18104 19712
rect 18696 19771 18748 19780
rect 18696 19737 18705 19771
rect 18705 19737 18739 19771
rect 18739 19737 18748 19771
rect 18696 19728 18748 19737
rect 18880 19728 18932 19780
rect 22192 19839 22244 19848
rect 22192 19805 22201 19839
rect 22201 19805 22235 19839
rect 22235 19805 22244 19839
rect 22192 19796 22244 19805
rect 22376 19839 22428 19848
rect 22376 19805 22385 19839
rect 22385 19805 22419 19839
rect 22419 19805 22428 19839
rect 22376 19796 22428 19805
rect 22284 19728 22336 19780
rect 23020 19796 23072 19848
rect 23572 19864 23624 19916
rect 24860 19932 24912 19984
rect 23664 19796 23716 19848
rect 20352 19660 20404 19712
rect 23020 19660 23072 19712
rect 23480 19728 23532 19780
rect 24216 19796 24268 19848
rect 25412 19796 25464 19848
rect 26056 19796 26108 19848
rect 26332 19796 26384 19848
rect 31300 20000 31352 20052
rect 32036 20000 32088 20052
rect 33232 20000 33284 20052
rect 34152 20000 34204 20052
rect 34704 20000 34756 20052
rect 34980 20000 35032 20052
rect 35256 20000 35308 20052
rect 35532 20000 35584 20052
rect 27344 19932 27396 19984
rect 28724 19932 28776 19984
rect 29000 19932 29052 19984
rect 31024 19932 31076 19984
rect 26884 19864 26936 19916
rect 27252 19864 27304 19916
rect 23388 19660 23440 19712
rect 24768 19660 24820 19712
rect 26516 19728 26568 19780
rect 27436 19796 27488 19848
rect 28908 19796 28960 19848
rect 33048 19864 33100 19916
rect 26792 19728 26844 19780
rect 27252 19728 27304 19780
rect 26056 19660 26108 19712
rect 26240 19660 26292 19712
rect 29460 19728 29512 19780
rect 29644 19728 29696 19780
rect 30472 19728 30524 19780
rect 33692 19864 33744 19916
rect 35624 19975 35676 19984
rect 35624 19941 35633 19975
rect 35633 19941 35667 19975
rect 35667 19941 35676 19975
rect 35624 19932 35676 19941
rect 36360 19864 36412 19916
rect 33232 19796 33284 19848
rect 33876 19796 33928 19848
rect 34796 19796 34848 19848
rect 35072 19839 35124 19848
rect 35072 19805 35082 19839
rect 35082 19805 35116 19839
rect 35116 19805 35124 19839
rect 35072 19796 35124 19805
rect 35256 19839 35308 19848
rect 35256 19805 35265 19839
rect 35265 19805 35299 19839
rect 35299 19805 35308 19839
rect 35256 19796 35308 19805
rect 35532 19796 35584 19848
rect 35808 19796 35860 19848
rect 35992 19796 36044 19848
rect 36176 19796 36228 19848
rect 36544 19796 36596 19848
rect 37464 19796 37516 19848
rect 32036 19728 32088 19780
rect 33508 19728 33560 19780
rect 33600 19771 33652 19780
rect 33600 19737 33609 19771
rect 33609 19737 33643 19771
rect 33643 19737 33652 19771
rect 33600 19728 33652 19737
rect 28264 19703 28316 19712
rect 28264 19669 28273 19703
rect 28273 19669 28307 19703
rect 28307 19669 28316 19703
rect 28264 19660 28316 19669
rect 31300 19660 31352 19712
rect 31668 19660 31720 19712
rect 32404 19660 32456 19712
rect 34888 19660 34940 19712
rect 37832 19728 37884 19780
rect 36636 19660 36688 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 13820 19499 13872 19508
rect 13820 19465 13829 19499
rect 13829 19465 13863 19499
rect 13863 19465 13872 19499
rect 13820 19456 13872 19465
rect 14740 19456 14792 19508
rect 20260 19456 20312 19508
rect 20812 19456 20864 19508
rect 21272 19456 21324 19508
rect 23204 19456 23256 19508
rect 24676 19456 24728 19508
rect 25044 19456 25096 19508
rect 26424 19456 26476 19508
rect 27160 19456 27212 19508
rect 27344 19456 27396 19508
rect 16672 19388 16724 19440
rect 19616 19388 19668 19440
rect 20536 19388 20588 19440
rect 22100 19388 22152 19440
rect 24400 19388 24452 19440
rect 12348 19320 12400 19372
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 16580 19320 16632 19372
rect 17132 19363 17184 19372
rect 17132 19329 17141 19363
rect 17141 19329 17175 19363
rect 17175 19329 17184 19363
rect 17132 19320 17184 19329
rect 17684 19320 17736 19372
rect 17776 19320 17828 19372
rect 18052 19320 18104 19372
rect 20628 19320 20680 19372
rect 21456 19320 21508 19372
rect 23480 19320 23532 19372
rect 23756 19320 23808 19372
rect 24308 19363 24360 19372
rect 24308 19329 24317 19363
rect 24317 19329 24351 19363
rect 24351 19329 24360 19363
rect 24308 19320 24360 19329
rect 24492 19363 24544 19372
rect 24492 19329 24501 19363
rect 24501 19329 24535 19363
rect 24535 19329 24544 19363
rect 24492 19320 24544 19329
rect 14372 19252 14424 19304
rect 14464 19252 14516 19304
rect 15200 19295 15252 19304
rect 15200 19261 15209 19295
rect 15209 19261 15243 19295
rect 15243 19261 15252 19295
rect 15200 19252 15252 19261
rect 15384 19252 15436 19304
rect 13544 19184 13596 19236
rect 14464 19116 14516 19168
rect 15936 19116 15988 19168
rect 16764 19184 16816 19236
rect 17040 19184 17092 19236
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 18512 19252 18564 19304
rect 19340 19252 19392 19304
rect 20996 19252 21048 19304
rect 21088 19184 21140 19236
rect 18512 19116 18564 19168
rect 18972 19159 19024 19168
rect 18972 19125 18981 19159
rect 18981 19125 19015 19159
rect 19015 19125 19024 19159
rect 18972 19116 19024 19125
rect 21732 19252 21784 19304
rect 22008 19252 22060 19304
rect 21916 19184 21968 19236
rect 23940 19252 23992 19304
rect 24216 19252 24268 19304
rect 24676 19363 24728 19372
rect 24676 19329 24685 19363
rect 24685 19329 24719 19363
rect 24719 19329 24728 19363
rect 24676 19320 24728 19329
rect 24768 19320 24820 19372
rect 25964 19363 26016 19372
rect 25964 19329 25973 19363
rect 25973 19329 26007 19363
rect 26007 19329 26016 19363
rect 25964 19320 26016 19329
rect 26148 19363 26200 19372
rect 26148 19329 26157 19363
rect 26157 19329 26191 19363
rect 26191 19329 26200 19363
rect 26148 19320 26200 19329
rect 26240 19363 26292 19372
rect 26240 19329 26249 19363
rect 26249 19329 26283 19363
rect 26283 19329 26292 19363
rect 26240 19320 26292 19329
rect 26884 19320 26936 19372
rect 27252 19320 27304 19372
rect 30012 19456 30064 19508
rect 28724 19388 28776 19440
rect 29000 19431 29052 19440
rect 29000 19397 29009 19431
rect 29009 19397 29043 19431
rect 29043 19397 29052 19431
rect 29000 19388 29052 19397
rect 29460 19388 29512 19440
rect 31024 19456 31076 19508
rect 31116 19456 31168 19508
rect 32864 19499 32916 19508
rect 32864 19465 32873 19499
rect 32873 19465 32907 19499
rect 32907 19465 32916 19499
rect 32864 19456 32916 19465
rect 33324 19456 33376 19508
rect 27896 19320 27948 19372
rect 22376 19227 22428 19236
rect 22376 19193 22385 19227
rect 22385 19193 22419 19227
rect 22419 19193 22428 19227
rect 22376 19184 22428 19193
rect 25872 19184 25924 19236
rect 23480 19159 23532 19168
rect 23480 19125 23489 19159
rect 23489 19125 23523 19159
rect 23523 19125 23532 19159
rect 23480 19116 23532 19125
rect 25136 19116 25188 19168
rect 26424 19116 26476 19168
rect 27068 19252 27120 19304
rect 27620 19252 27672 19304
rect 29368 19252 29420 19304
rect 29644 19252 29696 19304
rect 26884 19184 26936 19236
rect 29920 19363 29972 19372
rect 29920 19329 29929 19363
rect 29929 19329 29963 19363
rect 29963 19329 29972 19363
rect 29920 19320 29972 19329
rect 30840 19320 30892 19372
rect 33232 19388 33284 19440
rect 34060 19388 34112 19440
rect 31024 19320 31076 19372
rect 30288 19252 30340 19304
rect 31668 19320 31720 19372
rect 32864 19320 32916 19372
rect 33692 19320 33744 19372
rect 33876 19320 33928 19372
rect 34612 19388 34664 19440
rect 36360 19388 36412 19440
rect 34520 19320 34572 19372
rect 34888 19363 34940 19372
rect 34888 19329 34895 19363
rect 34895 19329 34940 19363
rect 34888 19320 34940 19329
rect 34981 19363 35033 19372
rect 34981 19329 34989 19363
rect 34989 19329 35023 19363
rect 35023 19329 35033 19363
rect 34981 19320 35033 19329
rect 35348 19320 35400 19372
rect 35808 19363 35860 19372
rect 35808 19329 35817 19363
rect 35817 19329 35851 19363
rect 35851 19329 35860 19363
rect 35808 19320 35860 19329
rect 33048 19295 33100 19304
rect 33048 19261 33057 19295
rect 33057 19261 33091 19295
rect 33091 19261 33100 19295
rect 33048 19252 33100 19261
rect 30472 19184 30524 19236
rect 31760 19184 31812 19236
rect 32220 19184 32272 19236
rect 32496 19184 32548 19236
rect 33508 19252 33560 19304
rect 36728 19363 36780 19372
rect 36728 19329 36737 19363
rect 36737 19329 36771 19363
rect 36771 19329 36780 19363
rect 36728 19320 36780 19329
rect 39028 19388 39080 19440
rect 37556 19320 37608 19372
rect 37924 19320 37976 19372
rect 36820 19295 36872 19304
rect 36820 19261 36829 19295
rect 36829 19261 36863 19295
rect 36863 19261 36872 19295
rect 36820 19252 36872 19261
rect 34060 19184 34112 19236
rect 34796 19184 34848 19236
rect 28724 19116 28776 19168
rect 30012 19116 30064 19168
rect 30748 19116 30800 19168
rect 31024 19116 31076 19168
rect 31668 19116 31720 19168
rect 34980 19116 35032 19168
rect 35164 19116 35216 19168
rect 35624 19116 35676 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 13544 18912 13596 18964
rect 12900 18751 12952 18760
rect 12900 18717 12909 18751
rect 12909 18717 12943 18751
rect 12943 18717 12952 18751
rect 12900 18708 12952 18717
rect 14096 18776 14148 18828
rect 14740 18844 14792 18896
rect 14832 18844 14884 18896
rect 14464 18708 14516 18760
rect 14648 18708 14700 18760
rect 15476 18776 15528 18828
rect 16212 18819 16264 18828
rect 16212 18785 16221 18819
rect 16221 18785 16255 18819
rect 16255 18785 16264 18819
rect 16212 18776 16264 18785
rect 17224 18776 17276 18828
rect 20904 18912 20956 18964
rect 21732 18955 21784 18964
rect 21732 18921 21741 18955
rect 21741 18921 21775 18955
rect 21775 18921 21784 18955
rect 21732 18912 21784 18921
rect 23112 18912 23164 18964
rect 23756 18912 23808 18964
rect 24768 18912 24820 18964
rect 25872 18955 25924 18964
rect 25872 18921 25881 18955
rect 25881 18921 25915 18955
rect 25915 18921 25924 18955
rect 25872 18912 25924 18921
rect 22376 18844 22428 18896
rect 23848 18844 23900 18896
rect 24584 18844 24636 18896
rect 28632 18912 28684 18964
rect 29920 18912 29972 18964
rect 32220 18912 32272 18964
rect 32864 18912 32916 18964
rect 33140 18912 33192 18964
rect 33508 18912 33560 18964
rect 33600 18912 33652 18964
rect 35072 18912 35124 18964
rect 35624 18912 35676 18964
rect 36452 18912 36504 18964
rect 21456 18776 21508 18828
rect 22008 18776 22060 18828
rect 15016 18751 15068 18760
rect 15016 18717 15025 18751
rect 15025 18717 15059 18751
rect 15059 18717 15068 18751
rect 15016 18708 15068 18717
rect 16764 18708 16816 18760
rect 17132 18708 17184 18760
rect 15476 18683 15528 18692
rect 15476 18649 15485 18683
rect 15485 18649 15519 18683
rect 15519 18649 15528 18683
rect 15476 18640 15528 18649
rect 11060 18572 11112 18624
rect 14740 18572 14792 18624
rect 15016 18572 15068 18624
rect 16028 18572 16080 18624
rect 18972 18708 19024 18760
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 20536 18751 20588 18760
rect 20536 18717 20545 18751
rect 20545 18717 20579 18751
rect 20579 18717 20588 18751
rect 20536 18708 20588 18717
rect 21640 18751 21692 18760
rect 21640 18717 21649 18751
rect 21649 18717 21683 18751
rect 21683 18717 21692 18751
rect 21640 18708 21692 18717
rect 22836 18708 22888 18760
rect 23296 18708 23348 18760
rect 23756 18708 23808 18760
rect 23940 18708 23992 18760
rect 26056 18844 26108 18896
rect 26976 18844 27028 18896
rect 27344 18844 27396 18896
rect 25228 18776 25280 18828
rect 27712 18776 27764 18828
rect 25872 18751 25924 18760
rect 25872 18717 25881 18751
rect 25881 18717 25915 18751
rect 25915 18717 25924 18751
rect 25872 18708 25924 18717
rect 26056 18751 26108 18760
rect 26056 18717 26065 18751
rect 26065 18717 26099 18751
rect 26099 18717 26108 18751
rect 26056 18708 26108 18717
rect 26516 18708 26568 18760
rect 26792 18708 26844 18760
rect 27068 18751 27120 18760
rect 27068 18717 27082 18751
rect 27082 18717 27116 18751
rect 27116 18717 27120 18751
rect 27068 18708 27120 18717
rect 27528 18708 27580 18760
rect 29368 18844 29420 18896
rect 17776 18640 17828 18692
rect 18328 18572 18380 18624
rect 18604 18640 18656 18692
rect 20628 18640 20680 18692
rect 23020 18640 23072 18692
rect 24400 18640 24452 18692
rect 25136 18683 25188 18692
rect 25136 18649 25145 18683
rect 25145 18649 25179 18683
rect 25179 18649 25188 18683
rect 25136 18640 25188 18649
rect 25228 18683 25280 18692
rect 25228 18649 25237 18683
rect 25237 18649 25271 18683
rect 25271 18649 25280 18683
rect 25228 18640 25280 18649
rect 28172 18751 28224 18760
rect 28172 18717 28181 18751
rect 28181 18717 28215 18751
rect 28215 18717 28224 18751
rect 28172 18708 28224 18717
rect 28356 18751 28408 18760
rect 28356 18717 28365 18751
rect 28365 18717 28399 18751
rect 28399 18717 28408 18751
rect 28356 18708 28408 18717
rect 28540 18776 28592 18828
rect 29460 18776 29512 18828
rect 27712 18640 27764 18692
rect 29828 18708 29880 18760
rect 30012 18844 30064 18896
rect 30840 18844 30892 18896
rect 31576 18844 31628 18896
rect 30012 18708 30064 18760
rect 31300 18776 31352 18828
rect 31208 18751 31260 18760
rect 31208 18717 31217 18751
rect 31217 18717 31251 18751
rect 31251 18717 31260 18751
rect 31208 18708 31260 18717
rect 31668 18751 31720 18760
rect 31668 18717 31677 18751
rect 31677 18717 31711 18751
rect 31711 18717 31720 18751
rect 31668 18708 31720 18717
rect 32404 18708 32456 18760
rect 32864 18751 32916 18760
rect 32864 18717 32873 18751
rect 32873 18717 32907 18751
rect 32907 18717 32916 18751
rect 32864 18708 32916 18717
rect 22744 18615 22796 18624
rect 22744 18581 22753 18615
rect 22753 18581 22787 18615
rect 22787 18581 22796 18615
rect 22744 18572 22796 18581
rect 23388 18572 23440 18624
rect 24584 18572 24636 18624
rect 27344 18572 27396 18624
rect 27528 18572 27580 18624
rect 29368 18640 29420 18692
rect 30472 18640 30524 18692
rect 32312 18640 32364 18692
rect 29000 18615 29052 18624
rect 29000 18581 29015 18615
rect 29015 18581 29049 18615
rect 29049 18581 29052 18615
rect 29000 18572 29052 18581
rect 30564 18572 30616 18624
rect 31208 18572 31260 18624
rect 31300 18572 31352 18624
rect 32496 18572 32548 18624
rect 32588 18615 32640 18624
rect 32588 18581 32597 18615
rect 32597 18581 32631 18615
rect 32631 18581 32640 18615
rect 32588 18572 32640 18581
rect 33232 18819 33284 18828
rect 33232 18785 33241 18819
rect 33241 18785 33275 18819
rect 33275 18785 33284 18819
rect 33232 18776 33284 18785
rect 33968 18844 34020 18896
rect 33140 18683 33192 18692
rect 33140 18649 33149 18683
rect 33149 18649 33183 18683
rect 33183 18649 33192 18683
rect 33140 18640 33192 18649
rect 36268 18776 36320 18828
rect 34520 18708 34572 18760
rect 34980 18751 35032 18760
rect 34980 18717 34990 18751
rect 34990 18717 35024 18751
rect 35024 18717 35032 18751
rect 34980 18708 35032 18717
rect 35164 18751 35216 18760
rect 35164 18717 35173 18751
rect 35173 18717 35207 18751
rect 35207 18717 35216 18751
rect 35164 18708 35216 18717
rect 35348 18751 35400 18760
rect 35348 18717 35362 18751
rect 35362 18717 35396 18751
rect 35396 18717 35400 18751
rect 35348 18708 35400 18717
rect 36544 18751 36596 18760
rect 36544 18717 36553 18751
rect 36553 18717 36587 18751
rect 36587 18717 36596 18751
rect 36544 18708 36596 18717
rect 33692 18572 33744 18624
rect 33968 18615 34020 18624
rect 33968 18581 33977 18615
rect 33977 18581 34011 18615
rect 34011 18581 34020 18615
rect 33968 18572 34020 18581
rect 36452 18640 36504 18692
rect 35348 18572 35400 18624
rect 37832 18572 37884 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 14372 18411 14424 18420
rect 14372 18377 14381 18411
rect 14381 18377 14415 18411
rect 14415 18377 14424 18411
rect 14372 18368 14424 18377
rect 15384 18368 15436 18420
rect 12900 18300 12952 18352
rect 16948 18368 17000 18420
rect 16028 18343 16080 18352
rect 16028 18309 16037 18343
rect 16037 18309 16071 18343
rect 16071 18309 16080 18343
rect 16028 18300 16080 18309
rect 14096 18275 14148 18284
rect 14096 18241 14105 18275
rect 14105 18241 14139 18275
rect 14139 18241 14148 18275
rect 14096 18232 14148 18241
rect 14832 18232 14884 18284
rect 15016 18164 15068 18216
rect 16212 18275 16264 18284
rect 16212 18241 16221 18275
rect 16221 18241 16255 18275
rect 16255 18241 16264 18275
rect 16212 18232 16264 18241
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 18328 18275 18380 18284
rect 18328 18241 18337 18275
rect 18337 18241 18371 18275
rect 18371 18241 18380 18275
rect 18328 18232 18380 18241
rect 19340 18368 19392 18420
rect 20076 18368 20128 18420
rect 20168 18368 20220 18420
rect 23204 18368 23256 18420
rect 23480 18368 23532 18420
rect 24308 18368 24360 18420
rect 18512 18164 18564 18216
rect 20444 18300 20496 18352
rect 20628 18300 20680 18352
rect 22744 18300 22796 18352
rect 22284 18275 22336 18284
rect 22284 18241 22293 18275
rect 22293 18241 22327 18275
rect 22327 18241 22336 18275
rect 22284 18232 22336 18241
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 22468 18232 22520 18284
rect 25228 18300 25280 18352
rect 19800 18207 19852 18216
rect 19800 18173 19809 18207
rect 19809 18173 19843 18207
rect 19843 18173 19852 18207
rect 19800 18164 19852 18173
rect 20076 18164 20128 18216
rect 20812 18207 20864 18216
rect 20812 18173 20821 18207
rect 20821 18173 20855 18207
rect 20855 18173 20864 18207
rect 20812 18164 20864 18173
rect 22192 18164 22244 18216
rect 24032 18232 24084 18284
rect 24308 18232 24360 18284
rect 25688 18275 25740 18284
rect 25688 18241 25697 18275
rect 25697 18241 25731 18275
rect 25731 18241 25740 18275
rect 25688 18232 25740 18241
rect 25872 18275 25924 18284
rect 25872 18241 25881 18275
rect 25881 18241 25915 18275
rect 25915 18241 25924 18275
rect 25872 18232 25924 18241
rect 26240 18232 26292 18284
rect 26608 18275 26660 18284
rect 26608 18241 26617 18275
rect 26617 18241 26651 18275
rect 26651 18241 26660 18275
rect 26608 18232 26660 18241
rect 29920 18368 29972 18420
rect 30840 18368 30892 18420
rect 32220 18368 32272 18420
rect 27620 18300 27672 18352
rect 23572 18164 23624 18216
rect 24400 18207 24452 18216
rect 24400 18173 24409 18207
rect 24409 18173 24443 18207
rect 24443 18173 24452 18207
rect 24400 18164 24452 18173
rect 25964 18207 26016 18216
rect 25964 18173 25973 18207
rect 25973 18173 26007 18207
rect 26007 18173 26016 18207
rect 25964 18164 26016 18173
rect 26056 18164 26108 18216
rect 27252 18232 27304 18284
rect 29092 18275 29144 18284
rect 29092 18241 29101 18275
rect 29101 18241 29135 18275
rect 29135 18241 29144 18275
rect 29092 18232 29144 18241
rect 32404 18300 32456 18352
rect 35256 18368 35308 18420
rect 35532 18368 35584 18420
rect 29460 18232 29512 18284
rect 30288 18232 30340 18284
rect 30380 18275 30432 18284
rect 30380 18241 30389 18275
rect 30389 18241 30423 18275
rect 30423 18241 30432 18275
rect 30380 18232 30432 18241
rect 30564 18232 30616 18284
rect 23388 18096 23440 18148
rect 24584 18096 24636 18148
rect 30012 18139 30064 18148
rect 30012 18105 30021 18139
rect 30021 18105 30055 18139
rect 30055 18105 30064 18139
rect 30012 18096 30064 18105
rect 31760 18232 31812 18284
rect 31576 18207 31628 18216
rect 31576 18173 31585 18207
rect 31585 18173 31619 18207
rect 31619 18173 31628 18207
rect 31576 18164 31628 18173
rect 32220 18164 32272 18216
rect 32496 18207 32548 18216
rect 32496 18173 32505 18207
rect 32505 18173 32539 18207
rect 32539 18173 32548 18207
rect 32496 18164 32548 18173
rect 32588 18164 32640 18216
rect 33232 18232 33284 18284
rect 33416 18275 33468 18284
rect 33416 18241 33425 18275
rect 33425 18241 33459 18275
rect 33459 18241 33468 18275
rect 33416 18232 33468 18241
rect 32864 18207 32916 18216
rect 32864 18173 32873 18207
rect 32873 18173 32907 18207
rect 32907 18173 32916 18207
rect 32864 18164 32916 18173
rect 30748 18096 30800 18148
rect 30840 18096 30892 18148
rect 33600 18232 33652 18284
rect 33876 18275 33928 18284
rect 33876 18241 33890 18275
rect 33890 18241 33924 18275
rect 33924 18241 33928 18275
rect 33876 18232 33928 18241
rect 34796 18275 34848 18284
rect 34796 18241 34805 18275
rect 34805 18241 34839 18275
rect 34839 18241 34848 18275
rect 34796 18232 34848 18241
rect 34980 18300 35032 18352
rect 35348 18300 35400 18352
rect 35808 18300 35860 18352
rect 35072 18275 35124 18284
rect 35072 18241 35081 18275
rect 35081 18241 35115 18275
rect 35115 18241 35124 18275
rect 35072 18232 35124 18241
rect 35256 18275 35308 18284
rect 35256 18241 35270 18275
rect 35270 18241 35304 18275
rect 35304 18241 35308 18275
rect 35256 18232 35308 18241
rect 33692 18096 33744 18148
rect 17408 18028 17460 18080
rect 18144 18071 18196 18080
rect 18144 18037 18153 18071
rect 18153 18037 18187 18071
rect 18187 18037 18196 18071
rect 18144 18028 18196 18037
rect 19156 18071 19208 18080
rect 19156 18037 19165 18071
rect 19165 18037 19199 18071
rect 19199 18037 19208 18071
rect 19156 18028 19208 18037
rect 20536 18028 20588 18080
rect 21640 18028 21692 18080
rect 23480 18028 23532 18080
rect 24216 18071 24268 18080
rect 24216 18037 24225 18071
rect 24225 18037 24259 18071
rect 24259 18037 24268 18071
rect 24216 18028 24268 18037
rect 25504 18071 25556 18080
rect 25504 18037 25513 18071
rect 25513 18037 25547 18071
rect 25547 18037 25556 18071
rect 25504 18028 25556 18037
rect 26516 18071 26568 18080
rect 26516 18037 26525 18071
rect 26525 18037 26559 18071
rect 26559 18037 26568 18071
rect 26516 18028 26568 18037
rect 28264 18028 28316 18080
rect 29092 18028 29144 18080
rect 31300 18028 31352 18080
rect 34612 18096 34664 18148
rect 36268 18232 36320 18284
rect 37832 18275 37884 18284
rect 37832 18241 37841 18275
rect 37841 18241 37875 18275
rect 37875 18241 37884 18275
rect 37832 18232 37884 18241
rect 36360 18164 36412 18216
rect 38108 18207 38160 18216
rect 38108 18173 38117 18207
rect 38117 18173 38151 18207
rect 38151 18173 38160 18207
rect 38108 18164 38160 18173
rect 34520 18028 34572 18080
rect 35348 18028 35400 18080
rect 36084 18028 36136 18080
rect 37464 18071 37516 18080
rect 37464 18037 37473 18071
rect 37473 18037 37507 18071
rect 37507 18037 37516 18071
rect 37464 18028 37516 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 15016 17867 15068 17876
rect 15016 17833 15025 17867
rect 15025 17833 15059 17867
rect 15059 17833 15068 17867
rect 15016 17824 15068 17833
rect 15384 17824 15436 17876
rect 15936 17824 15988 17876
rect 16304 17824 16356 17876
rect 16488 17824 16540 17876
rect 18512 17824 18564 17876
rect 19524 17824 19576 17876
rect 22008 17824 22060 17876
rect 22376 17824 22428 17876
rect 23572 17867 23624 17876
rect 23572 17833 23581 17867
rect 23581 17833 23615 17867
rect 23615 17833 23624 17867
rect 23572 17824 23624 17833
rect 26516 17824 26568 17876
rect 16028 17688 16080 17740
rect 15384 17663 15436 17672
rect 15384 17629 15393 17663
rect 15393 17629 15427 17663
rect 15427 17629 15436 17663
rect 15384 17620 15436 17629
rect 15844 17552 15896 17604
rect 17500 17620 17552 17672
rect 17776 17663 17828 17672
rect 17776 17629 17785 17663
rect 17785 17629 17819 17663
rect 17819 17629 17828 17663
rect 17776 17620 17828 17629
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 21272 17756 21324 17808
rect 23296 17756 23348 17808
rect 24676 17756 24728 17808
rect 25504 17756 25556 17808
rect 27528 17824 27580 17876
rect 31392 17824 31444 17876
rect 31944 17824 31996 17876
rect 32496 17824 32548 17876
rect 34152 17824 34204 17876
rect 35348 17867 35400 17876
rect 35348 17833 35357 17867
rect 35357 17833 35391 17867
rect 35391 17833 35400 17867
rect 35348 17824 35400 17833
rect 36452 17867 36504 17876
rect 36452 17833 36461 17867
rect 36461 17833 36495 17867
rect 36495 17833 36504 17867
rect 36452 17824 36504 17833
rect 37832 17824 37884 17876
rect 27160 17756 27212 17808
rect 28172 17756 28224 17808
rect 30748 17756 30800 17808
rect 32588 17756 32640 17808
rect 18880 17663 18932 17672
rect 18880 17629 18889 17663
rect 18889 17629 18923 17663
rect 18923 17629 18932 17663
rect 18880 17620 18932 17629
rect 19064 17620 19116 17672
rect 19524 17663 19576 17672
rect 19524 17629 19533 17663
rect 19533 17629 19567 17663
rect 19567 17629 19576 17663
rect 19524 17620 19576 17629
rect 19156 17552 19208 17604
rect 20720 17620 20772 17672
rect 20904 17663 20956 17672
rect 20904 17629 20913 17663
rect 20913 17629 20947 17663
rect 20947 17629 20956 17663
rect 20904 17620 20956 17629
rect 20812 17595 20864 17604
rect 20812 17561 20821 17595
rect 20821 17561 20855 17595
rect 20855 17561 20864 17595
rect 20812 17552 20864 17561
rect 21272 17552 21324 17604
rect 22008 17552 22060 17604
rect 22836 17663 22888 17672
rect 22836 17629 22845 17663
rect 22845 17629 22879 17663
rect 22879 17629 22888 17663
rect 22836 17620 22888 17629
rect 23204 17620 23256 17672
rect 24584 17663 24636 17672
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 24676 17663 24728 17672
rect 24676 17629 24685 17663
rect 24685 17629 24719 17663
rect 24719 17629 24728 17663
rect 24676 17620 24728 17629
rect 24768 17620 24820 17672
rect 25780 17663 25832 17672
rect 25780 17629 25789 17663
rect 25789 17629 25823 17663
rect 25823 17629 25832 17663
rect 25780 17620 25832 17629
rect 26332 17620 26384 17672
rect 30840 17688 30892 17740
rect 30932 17688 30984 17740
rect 31668 17688 31720 17740
rect 32956 17688 33008 17740
rect 33600 17688 33652 17740
rect 23940 17552 23992 17604
rect 26608 17595 26660 17604
rect 26608 17561 26617 17595
rect 26617 17561 26651 17595
rect 26651 17561 26660 17595
rect 26608 17552 26660 17561
rect 27620 17663 27672 17672
rect 27344 17595 27396 17604
rect 27344 17561 27353 17595
rect 27353 17561 27387 17595
rect 27387 17561 27396 17595
rect 27344 17552 27396 17561
rect 27620 17629 27623 17663
rect 27623 17629 27672 17663
rect 27620 17620 27672 17629
rect 27988 17552 28040 17604
rect 28632 17595 28684 17604
rect 28632 17561 28641 17595
rect 28641 17561 28675 17595
rect 28675 17561 28684 17595
rect 28632 17552 28684 17561
rect 29736 17663 29788 17672
rect 29736 17629 29745 17663
rect 29745 17629 29779 17663
rect 29779 17629 29788 17663
rect 29736 17620 29788 17629
rect 30564 17663 30616 17672
rect 30564 17629 30573 17663
rect 30573 17629 30607 17663
rect 30607 17629 30616 17663
rect 30564 17620 30616 17629
rect 31392 17663 31444 17672
rect 31392 17629 31401 17663
rect 31401 17629 31435 17663
rect 31435 17629 31444 17663
rect 31392 17620 31444 17629
rect 31484 17620 31536 17672
rect 32036 17620 32088 17672
rect 32220 17620 32272 17672
rect 32864 17620 32916 17672
rect 33324 17663 33376 17672
rect 33324 17629 33333 17663
rect 33333 17629 33367 17663
rect 33367 17629 33376 17663
rect 33324 17620 33376 17629
rect 33416 17663 33468 17672
rect 33416 17629 33426 17663
rect 33426 17629 33460 17663
rect 33460 17629 33468 17663
rect 33416 17620 33468 17629
rect 33508 17620 33560 17672
rect 15476 17484 15528 17536
rect 16212 17484 16264 17536
rect 16304 17484 16356 17536
rect 20904 17484 20956 17536
rect 26976 17484 27028 17536
rect 28356 17484 28408 17536
rect 28540 17484 28592 17536
rect 29276 17552 29328 17604
rect 31300 17552 31352 17604
rect 33784 17663 33836 17672
rect 33784 17629 33798 17663
rect 33798 17629 33832 17663
rect 33832 17629 33836 17663
rect 34060 17756 34112 17808
rect 34704 17688 34756 17740
rect 36728 17688 36780 17740
rect 33784 17620 33836 17629
rect 35164 17663 35216 17672
rect 35164 17629 35173 17663
rect 35173 17629 35207 17663
rect 35207 17629 35216 17663
rect 35164 17620 35216 17629
rect 29644 17484 29696 17536
rect 30564 17484 30616 17536
rect 33416 17484 33468 17536
rect 33692 17595 33744 17604
rect 33692 17561 33701 17595
rect 33701 17561 33735 17595
rect 33735 17561 33744 17595
rect 33692 17552 33744 17561
rect 36084 17663 36136 17672
rect 36084 17629 36093 17663
rect 36093 17629 36127 17663
rect 36127 17629 36136 17663
rect 36084 17620 36136 17629
rect 36544 17620 36596 17672
rect 36820 17620 36872 17672
rect 37464 17620 37516 17672
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 15200 17323 15252 17332
rect 15200 17289 15209 17323
rect 15209 17289 15243 17323
rect 15243 17289 15252 17323
rect 15200 17280 15252 17289
rect 15476 17212 15528 17264
rect 15844 17187 15896 17196
rect 15844 17153 15853 17187
rect 15853 17153 15887 17187
rect 15887 17153 15896 17187
rect 15844 17144 15896 17153
rect 15936 17187 15988 17196
rect 15936 17153 15945 17187
rect 15945 17153 15979 17187
rect 15979 17153 15988 17187
rect 15936 17144 15988 17153
rect 16120 17187 16172 17196
rect 16120 17153 16129 17187
rect 16129 17153 16163 17187
rect 16163 17153 16172 17187
rect 16120 17144 16172 17153
rect 16028 17076 16080 17128
rect 16304 17144 16356 17196
rect 19064 17280 19116 17332
rect 22284 17280 22336 17332
rect 24492 17280 24544 17332
rect 26700 17280 26752 17332
rect 18052 17212 18104 17264
rect 18972 17212 19024 17264
rect 17408 17144 17460 17196
rect 18512 17144 18564 17196
rect 19432 17144 19484 17196
rect 20260 17212 20312 17264
rect 21916 17212 21968 17264
rect 22192 17255 22244 17264
rect 22192 17221 22201 17255
rect 22201 17221 22235 17255
rect 22235 17221 22244 17255
rect 22192 17212 22244 17221
rect 22376 17212 22428 17264
rect 17500 17119 17552 17128
rect 17500 17085 17509 17119
rect 17509 17085 17543 17119
rect 17543 17085 17552 17119
rect 17500 17076 17552 17085
rect 18144 17076 18196 17128
rect 19340 17076 19392 17128
rect 20168 17187 20220 17196
rect 20168 17153 20177 17187
rect 20177 17153 20211 17187
rect 20211 17153 20220 17187
rect 20168 17144 20220 17153
rect 20444 17144 20496 17196
rect 20536 17144 20588 17196
rect 21640 17144 21692 17196
rect 22652 17144 22704 17196
rect 23388 17144 23440 17196
rect 26608 17212 26660 17264
rect 29920 17280 29972 17332
rect 30104 17280 30156 17332
rect 35164 17280 35216 17332
rect 37832 17323 37884 17332
rect 37832 17289 37841 17323
rect 37841 17289 37875 17323
rect 37875 17289 37884 17323
rect 37832 17280 37884 17289
rect 29184 17212 29236 17264
rect 29736 17212 29788 17264
rect 23112 17076 23164 17128
rect 23204 17076 23256 17128
rect 15016 17008 15068 17060
rect 18052 17008 18104 17060
rect 18880 17008 18932 17060
rect 21272 17008 21324 17060
rect 17040 16983 17092 16992
rect 17040 16949 17049 16983
rect 17049 16949 17083 16983
rect 17083 16949 17092 16983
rect 17040 16940 17092 16949
rect 19156 16940 19208 16992
rect 20812 16940 20864 16992
rect 23020 16940 23072 16992
rect 23848 16940 23900 16992
rect 26056 17119 26108 17128
rect 26056 17085 26065 17119
rect 26065 17085 26099 17119
rect 26099 17085 26108 17119
rect 26056 17076 26108 17085
rect 27344 17187 27396 17196
rect 27344 17153 27353 17187
rect 27353 17153 27387 17187
rect 27387 17153 27396 17187
rect 27344 17144 27396 17153
rect 27712 17144 27764 17196
rect 28540 17144 28592 17196
rect 27528 17119 27580 17128
rect 27528 17085 27537 17119
rect 27537 17085 27571 17119
rect 27571 17085 27580 17119
rect 27528 17076 27580 17085
rect 27620 17119 27672 17128
rect 27620 17085 27629 17119
rect 27629 17085 27663 17119
rect 27663 17085 27672 17119
rect 27620 17076 27672 17085
rect 26148 17008 26200 17060
rect 30656 17187 30708 17196
rect 30656 17153 30665 17187
rect 30665 17153 30699 17187
rect 30699 17153 30708 17187
rect 30656 17144 30708 17153
rect 30748 17187 30800 17196
rect 30748 17153 30758 17187
rect 30758 17153 30792 17187
rect 30792 17153 30800 17187
rect 30748 17144 30800 17153
rect 30932 17187 30984 17196
rect 30932 17153 30941 17187
rect 30941 17153 30975 17187
rect 30975 17153 30984 17187
rect 30932 17144 30984 17153
rect 31300 17212 31352 17264
rect 32680 17212 32732 17264
rect 31208 17144 31260 17196
rect 31852 17144 31904 17196
rect 32312 17144 32364 17196
rect 33232 17212 33284 17264
rect 33600 17255 33652 17264
rect 33600 17221 33609 17255
rect 33609 17221 33643 17255
rect 33643 17221 33652 17255
rect 33600 17212 33652 17221
rect 34244 17144 34296 17196
rect 34520 17187 34572 17196
rect 34520 17153 34529 17187
rect 34529 17153 34563 17187
rect 34563 17153 34572 17187
rect 34520 17144 34572 17153
rect 34612 17187 34664 17196
rect 34612 17153 34621 17187
rect 34621 17153 34655 17187
rect 34655 17153 34664 17187
rect 34612 17144 34664 17153
rect 31668 17076 31720 17128
rect 32588 17076 32640 17128
rect 36360 17144 36412 17196
rect 38844 17144 38896 17196
rect 31852 17008 31904 17060
rect 35348 17008 35400 17060
rect 38108 17119 38160 17128
rect 38108 17085 38117 17119
rect 38117 17085 38151 17119
rect 38151 17085 38160 17119
rect 38108 17076 38160 17085
rect 39028 17008 39080 17060
rect 29006 16940 29058 16992
rect 31484 16940 31536 16992
rect 31668 16940 31720 16992
rect 37096 16940 37148 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 15016 16779 15068 16788
rect 15016 16745 15025 16779
rect 15025 16745 15059 16779
rect 15059 16745 15068 16779
rect 15016 16736 15068 16745
rect 16212 16736 16264 16788
rect 15844 16668 15896 16720
rect 16856 16736 16908 16788
rect 17500 16736 17552 16788
rect 22008 16736 22060 16788
rect 22652 16736 22704 16788
rect 16028 16532 16080 16584
rect 16120 16532 16172 16584
rect 19432 16668 19484 16720
rect 16672 16600 16724 16652
rect 18420 16643 18472 16652
rect 18420 16609 18429 16643
rect 18429 16609 18463 16643
rect 18463 16609 18472 16643
rect 18420 16600 18472 16609
rect 21364 16600 21416 16652
rect 25504 16600 25556 16652
rect 17592 16575 17644 16584
rect 17592 16541 17601 16575
rect 17601 16541 17635 16575
rect 17635 16541 17644 16575
rect 17592 16532 17644 16541
rect 18052 16532 18104 16584
rect 16580 16464 16632 16516
rect 20444 16532 20496 16584
rect 21732 16575 21784 16584
rect 21732 16541 21741 16575
rect 21741 16541 21775 16575
rect 21775 16541 21784 16575
rect 21732 16532 21784 16541
rect 22376 16532 22428 16584
rect 23940 16532 23992 16584
rect 24400 16532 24452 16584
rect 25688 16532 25740 16584
rect 27712 16736 27764 16788
rect 28632 16736 28684 16788
rect 29092 16736 29144 16788
rect 30104 16736 30156 16788
rect 27528 16600 27580 16652
rect 27804 16600 27856 16652
rect 31576 16736 31628 16788
rect 32588 16668 32640 16720
rect 33692 16736 33744 16788
rect 34796 16736 34848 16788
rect 26148 16532 26200 16584
rect 27252 16532 27304 16584
rect 20904 16464 20956 16516
rect 15016 16439 15068 16448
rect 15016 16405 15041 16439
rect 15041 16405 15068 16439
rect 15016 16396 15068 16405
rect 15292 16396 15344 16448
rect 20260 16396 20312 16448
rect 23480 16464 23532 16516
rect 24124 16464 24176 16516
rect 22744 16396 22796 16448
rect 27344 16396 27396 16448
rect 28264 16532 28316 16584
rect 32956 16643 33008 16652
rect 32956 16609 32965 16643
rect 32965 16609 32999 16643
rect 32999 16609 33008 16643
rect 32956 16600 33008 16609
rect 33968 16600 34020 16652
rect 35256 16643 35308 16652
rect 35256 16609 35265 16643
rect 35265 16609 35299 16643
rect 35299 16609 35308 16643
rect 35256 16600 35308 16609
rect 28356 16464 28408 16516
rect 31668 16532 31720 16584
rect 33508 16532 33560 16584
rect 34152 16532 34204 16584
rect 35808 16532 35860 16584
rect 37004 16736 37056 16788
rect 37832 16736 37884 16788
rect 36820 16643 36872 16652
rect 29552 16464 29604 16516
rect 33600 16464 33652 16516
rect 34796 16464 34848 16516
rect 36820 16609 36829 16643
rect 36829 16609 36863 16643
rect 36863 16609 36872 16643
rect 36820 16600 36872 16609
rect 37096 16575 37148 16584
rect 37096 16541 37130 16575
rect 37130 16541 37148 16575
rect 37096 16532 37148 16541
rect 30288 16396 30340 16448
rect 32128 16396 32180 16448
rect 34336 16396 34388 16448
rect 36268 16439 36320 16448
rect 36268 16405 36277 16439
rect 36277 16405 36311 16439
rect 36311 16405 36320 16439
rect 36268 16396 36320 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 19432 16192 19484 16244
rect 21364 16235 21416 16244
rect 21364 16201 21373 16235
rect 21373 16201 21407 16235
rect 21407 16201 21416 16235
rect 21364 16192 21416 16201
rect 21548 16192 21600 16244
rect 24032 16192 24084 16244
rect 17040 16124 17092 16176
rect 21824 16124 21876 16176
rect 15292 16099 15344 16108
rect 15292 16065 15301 16099
rect 15301 16065 15335 16099
rect 15335 16065 15344 16099
rect 15292 16056 15344 16065
rect 16028 16056 16080 16108
rect 15936 15988 15988 16040
rect 16856 16099 16908 16108
rect 16856 16065 16865 16099
rect 16865 16065 16899 16099
rect 16899 16065 16908 16099
rect 16856 16056 16908 16065
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 18512 16099 18564 16108
rect 18512 16065 18521 16099
rect 18521 16065 18555 16099
rect 18555 16065 18564 16099
rect 18512 16056 18564 16065
rect 18604 16099 18656 16108
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 20352 16099 20404 16108
rect 20352 16065 20361 16099
rect 20361 16065 20395 16099
rect 20395 16065 20404 16099
rect 20352 16056 20404 16065
rect 20812 16099 20864 16108
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 21272 16099 21324 16108
rect 21272 16065 21281 16099
rect 21281 16065 21315 16099
rect 21315 16065 21324 16099
rect 21272 16056 21324 16065
rect 21732 16056 21784 16108
rect 23756 16124 23808 16176
rect 23940 16124 23992 16176
rect 24308 16099 24360 16108
rect 24308 16065 24317 16099
rect 24317 16065 24351 16099
rect 24351 16065 24360 16099
rect 24308 16056 24360 16065
rect 25596 16192 25648 16244
rect 27712 16235 27764 16244
rect 27712 16201 27721 16235
rect 27721 16201 27755 16235
rect 27755 16201 27764 16235
rect 27712 16192 27764 16201
rect 30748 16192 30800 16244
rect 31760 16192 31812 16244
rect 26424 16124 26476 16176
rect 26056 16056 26108 16108
rect 26516 16056 26568 16108
rect 16580 15988 16632 16040
rect 17592 15988 17644 16040
rect 19156 15988 19208 16040
rect 23020 15988 23072 16040
rect 15016 15920 15068 15972
rect 18420 15920 18472 15972
rect 23112 15920 23164 15972
rect 25964 16031 26016 16040
rect 25964 15997 25973 16031
rect 25973 15997 26007 16031
rect 26007 15997 26016 16031
rect 25964 15988 26016 15997
rect 28448 16056 28500 16108
rect 28540 16099 28592 16108
rect 28540 16065 28549 16099
rect 28549 16065 28583 16099
rect 28583 16065 28592 16099
rect 28540 16056 28592 16065
rect 28816 16099 28868 16108
rect 28816 16065 28850 16099
rect 28850 16065 28868 16099
rect 28816 16056 28868 16065
rect 30748 16099 30800 16108
rect 30748 16065 30757 16099
rect 30757 16065 30791 16099
rect 30791 16065 30800 16099
rect 30748 16056 30800 16065
rect 31116 16124 31168 16176
rect 33600 16235 33652 16244
rect 33600 16201 33609 16235
rect 33609 16201 33643 16235
rect 33643 16201 33652 16235
rect 33600 16192 33652 16201
rect 33692 16192 33744 16244
rect 34520 16192 34572 16244
rect 35256 16167 35308 16176
rect 35256 16133 35290 16167
rect 35290 16133 35308 16167
rect 35256 16124 35308 16133
rect 36360 16235 36412 16244
rect 36360 16201 36369 16235
rect 36369 16201 36403 16235
rect 36403 16201 36412 16235
rect 36360 16192 36412 16201
rect 37924 16167 37976 16176
rect 37924 16133 37933 16167
rect 37933 16133 37967 16167
rect 37967 16133 37976 16167
rect 37924 16124 37976 16133
rect 29552 15988 29604 16040
rect 31116 15988 31168 16040
rect 32404 16056 32456 16108
rect 32680 16099 32732 16108
rect 32680 16065 32689 16099
rect 32689 16065 32723 16099
rect 32723 16065 32732 16099
rect 32680 16056 32732 16065
rect 32956 16099 33008 16108
rect 32956 16065 32965 16099
rect 32965 16065 32999 16099
rect 32999 16065 33008 16099
rect 32956 16056 33008 16065
rect 34704 16056 34756 16108
rect 36360 16056 36412 16108
rect 37832 16099 37884 16108
rect 37832 16065 37841 16099
rect 37841 16065 37875 16099
rect 37875 16065 37884 16099
rect 37832 16056 37884 16065
rect 32588 16031 32640 16040
rect 32588 15997 32597 16031
rect 32597 15997 32631 16031
rect 32631 15997 32640 16031
rect 32588 15988 32640 15997
rect 20076 15852 20128 15904
rect 25412 15895 25464 15904
rect 25412 15861 25421 15895
rect 25421 15861 25455 15895
rect 25455 15861 25464 15895
rect 25412 15852 25464 15861
rect 27344 15852 27396 15904
rect 29920 15895 29972 15904
rect 29920 15861 29929 15895
rect 29929 15861 29963 15895
rect 29963 15861 29972 15895
rect 29920 15852 29972 15861
rect 30380 15895 30432 15904
rect 30380 15861 30389 15895
rect 30389 15861 30423 15895
rect 30423 15861 30432 15895
rect 30380 15852 30432 15861
rect 34796 15988 34848 16040
rect 38108 15988 38160 16040
rect 37464 15895 37516 15904
rect 37464 15861 37473 15895
rect 37473 15861 37507 15895
rect 37507 15861 37516 15895
rect 37464 15852 37516 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 16764 15648 16816 15700
rect 19340 15648 19392 15700
rect 19984 15648 20036 15700
rect 22560 15648 22612 15700
rect 27252 15648 27304 15700
rect 28448 15691 28500 15700
rect 28448 15657 28457 15691
rect 28457 15657 28491 15691
rect 28491 15657 28500 15691
rect 28448 15648 28500 15657
rect 29000 15691 29052 15700
rect 29000 15657 29009 15691
rect 29009 15657 29043 15691
rect 29043 15657 29052 15691
rect 29000 15648 29052 15657
rect 33140 15648 33192 15700
rect 37832 15648 37884 15700
rect 20168 15623 20220 15632
rect 20168 15589 20177 15623
rect 20177 15589 20211 15623
rect 20211 15589 20220 15623
rect 20168 15580 20220 15589
rect 20352 15580 20404 15632
rect 31944 15623 31996 15632
rect 31944 15589 31953 15623
rect 31953 15589 31987 15623
rect 31987 15589 31996 15623
rect 31944 15580 31996 15589
rect 18696 15512 18748 15564
rect 18512 15444 18564 15496
rect 18880 15487 18932 15496
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 19432 15444 19484 15496
rect 20536 15512 20588 15564
rect 20076 15444 20128 15496
rect 20260 15487 20312 15496
rect 20260 15453 20269 15487
rect 20269 15453 20303 15487
rect 20303 15453 20312 15487
rect 20260 15444 20312 15453
rect 20812 15444 20864 15496
rect 22008 15512 22060 15564
rect 26516 15512 26568 15564
rect 26608 15512 26660 15564
rect 28540 15512 28592 15564
rect 21640 15444 21692 15496
rect 23388 15487 23440 15496
rect 23388 15453 23397 15487
rect 23397 15453 23431 15487
rect 23431 15453 23440 15487
rect 23388 15444 23440 15453
rect 24952 15444 25004 15496
rect 27344 15487 27396 15496
rect 27344 15453 27378 15487
rect 27378 15453 27396 15487
rect 27344 15444 27396 15453
rect 29552 15444 29604 15496
rect 31484 15512 31536 15564
rect 38936 15512 38988 15564
rect 29828 15444 29880 15496
rect 31392 15444 31444 15496
rect 34704 15444 34756 15496
rect 37464 15444 37516 15496
rect 38016 15444 38068 15496
rect 23756 15376 23808 15428
rect 24584 15419 24636 15428
rect 24584 15385 24593 15419
rect 24593 15385 24627 15419
rect 24627 15385 24636 15419
rect 24584 15376 24636 15385
rect 22928 15351 22980 15360
rect 22928 15317 22937 15351
rect 22937 15317 22971 15351
rect 22971 15317 22980 15351
rect 22928 15308 22980 15317
rect 25504 15308 25556 15360
rect 27436 15376 27488 15428
rect 30380 15376 30432 15428
rect 32220 15376 32272 15428
rect 29552 15308 29604 15360
rect 30748 15308 30800 15360
rect 33600 15308 33652 15360
rect 33876 15351 33928 15360
rect 33876 15317 33885 15351
rect 33885 15317 33919 15351
rect 33919 15317 33928 15351
rect 33876 15308 33928 15317
rect 35716 15376 35768 15428
rect 35440 15308 35492 15360
rect 36268 15308 36320 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 22468 15104 22520 15156
rect 23388 15104 23440 15156
rect 23664 15104 23716 15156
rect 18604 15036 18656 15088
rect 17408 14968 17460 15020
rect 18144 15011 18196 15020
rect 18144 14977 18153 15011
rect 18153 14977 18187 15011
rect 18187 14977 18196 15011
rect 18144 14968 18196 14977
rect 19156 15011 19208 15020
rect 19156 14977 19165 15011
rect 19165 14977 19199 15011
rect 19199 14977 19208 15011
rect 19156 14968 19208 14977
rect 20444 14968 20496 15020
rect 21088 15011 21140 15020
rect 21088 14977 21097 15011
rect 21097 14977 21131 15011
rect 21131 14977 21140 15011
rect 21088 14968 21140 14977
rect 22376 15011 22428 15020
rect 22376 14977 22385 15011
rect 22385 14977 22419 15011
rect 22419 14977 22428 15011
rect 22376 14968 22428 14977
rect 22928 14968 22980 15020
rect 25412 14968 25464 15020
rect 27344 15011 27396 15020
rect 27344 14977 27353 15011
rect 27353 14977 27387 15011
rect 27387 14977 27396 15011
rect 27344 14968 27396 14977
rect 27436 14968 27488 15020
rect 28816 15104 28868 15156
rect 29920 15104 29972 15156
rect 30104 15147 30156 15156
rect 30104 15113 30113 15147
rect 30113 15113 30147 15147
rect 30147 15113 30156 15147
rect 30104 15104 30156 15113
rect 32220 15104 32272 15156
rect 33784 15104 33836 15156
rect 29736 15036 29788 15088
rect 27988 14968 28040 15020
rect 28448 14968 28500 15020
rect 19248 14943 19300 14952
rect 19248 14909 19257 14943
rect 19257 14909 19291 14943
rect 19291 14909 19300 14943
rect 19248 14900 19300 14909
rect 19524 14943 19576 14952
rect 19524 14909 19533 14943
rect 19533 14909 19567 14943
rect 19567 14909 19576 14943
rect 19524 14900 19576 14909
rect 20168 14900 20220 14952
rect 22284 14900 22336 14952
rect 23388 14900 23440 14952
rect 18420 14832 18472 14884
rect 18788 14832 18840 14884
rect 28356 14943 28408 14952
rect 28356 14909 28365 14943
rect 28365 14909 28399 14943
rect 28399 14909 28408 14943
rect 28356 14900 28408 14909
rect 30196 14943 30248 14952
rect 30196 14909 30205 14943
rect 30205 14909 30239 14943
rect 30239 14909 30248 14943
rect 30196 14900 30248 14909
rect 30472 14968 30524 15020
rect 32496 14968 32548 15020
rect 33508 15011 33560 15020
rect 31484 14943 31536 14952
rect 31484 14909 31493 14943
rect 31493 14909 31527 14943
rect 31527 14909 31536 14943
rect 31484 14900 31536 14909
rect 31668 14943 31720 14952
rect 31668 14909 31677 14943
rect 31677 14909 31711 14943
rect 31711 14909 31720 14943
rect 31668 14900 31720 14909
rect 33508 14977 33517 15011
rect 33517 14977 33551 15011
rect 33551 14977 33560 15011
rect 33508 14968 33560 14977
rect 33876 15036 33928 15088
rect 34612 15104 34664 15156
rect 35992 15104 36044 15156
rect 33324 14943 33376 14952
rect 33324 14909 33333 14943
rect 33333 14909 33367 14943
rect 33367 14909 33376 14943
rect 33324 14900 33376 14909
rect 22100 14764 22152 14816
rect 23756 14807 23808 14816
rect 23756 14773 23765 14807
rect 23765 14773 23799 14807
rect 23799 14773 23808 14807
rect 23756 14764 23808 14773
rect 24768 14764 24820 14816
rect 26056 14764 26108 14816
rect 29460 14764 29512 14816
rect 31576 14764 31628 14816
rect 35900 15036 35952 15088
rect 36268 15079 36320 15088
rect 36268 15045 36277 15079
rect 36277 15045 36311 15079
rect 36311 15045 36320 15079
rect 36268 15036 36320 15045
rect 36912 15036 36964 15088
rect 39028 15036 39080 15088
rect 36176 14968 36228 15020
rect 36360 14968 36412 15020
rect 35992 14900 36044 14952
rect 36360 14764 36412 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 18512 14560 18564 14612
rect 21088 14560 21140 14612
rect 19524 14492 19576 14544
rect 19432 14356 19484 14408
rect 20076 14399 20128 14408
rect 20076 14365 20085 14399
rect 20085 14365 20119 14399
rect 20119 14365 20128 14399
rect 20076 14356 20128 14365
rect 22376 14356 22428 14408
rect 22652 14356 22704 14408
rect 19340 14288 19392 14340
rect 19248 14220 19300 14272
rect 22100 14331 22152 14340
rect 22100 14297 22134 14331
rect 22134 14297 22152 14331
rect 22100 14288 22152 14297
rect 23940 14560 23992 14612
rect 24676 14560 24728 14612
rect 27344 14560 27396 14612
rect 32312 14560 32364 14612
rect 33784 14560 33836 14612
rect 35808 14560 35860 14612
rect 28356 14492 28408 14544
rect 24032 14356 24084 14408
rect 24952 14356 25004 14408
rect 26056 14424 26108 14476
rect 27712 14424 27764 14476
rect 28540 14467 28592 14476
rect 28540 14433 28549 14467
rect 28549 14433 28583 14467
rect 28583 14433 28592 14467
rect 28540 14424 28592 14433
rect 30656 14424 30708 14476
rect 24860 14288 24912 14340
rect 25504 14399 25556 14408
rect 25504 14365 25513 14399
rect 25513 14365 25547 14399
rect 25547 14365 25556 14399
rect 25504 14356 25556 14365
rect 22376 14220 22428 14272
rect 23480 14220 23532 14272
rect 24032 14263 24084 14272
rect 24032 14229 24041 14263
rect 24041 14229 24075 14263
rect 24075 14229 24084 14263
rect 24032 14220 24084 14229
rect 27988 14356 28040 14408
rect 26332 14220 26384 14272
rect 26608 14288 26660 14340
rect 28356 14399 28408 14408
rect 28356 14365 28365 14399
rect 28365 14365 28399 14399
rect 28399 14365 28408 14399
rect 28356 14356 28408 14365
rect 38108 14467 38160 14476
rect 38108 14433 38117 14467
rect 38117 14433 38151 14467
rect 38151 14433 38160 14467
rect 38108 14424 38160 14433
rect 31024 14356 31076 14408
rect 33048 14356 33100 14408
rect 34796 14356 34848 14408
rect 30932 14288 30984 14340
rect 32036 14288 32088 14340
rect 33968 14331 34020 14340
rect 33968 14297 33977 14331
rect 33977 14297 34011 14331
rect 34011 14297 34020 14331
rect 33968 14288 34020 14297
rect 34152 14331 34204 14340
rect 34152 14297 34161 14331
rect 34161 14297 34195 14331
rect 34195 14297 34204 14331
rect 34152 14288 34204 14297
rect 36084 14356 36136 14408
rect 37924 14356 37976 14408
rect 32496 14220 32548 14272
rect 33232 14220 33284 14272
rect 33324 14263 33376 14272
rect 33324 14229 33333 14263
rect 33333 14229 33367 14263
rect 33367 14229 33376 14263
rect 33324 14220 33376 14229
rect 34796 14220 34848 14272
rect 36728 14331 36780 14340
rect 36728 14297 36737 14331
rect 36737 14297 36771 14331
rect 36771 14297 36780 14331
rect 36728 14288 36780 14297
rect 37556 14331 37608 14340
rect 37556 14297 37565 14331
rect 37565 14297 37599 14331
rect 37599 14297 37608 14331
rect 37556 14288 37608 14297
rect 35348 14220 35400 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 22376 14016 22428 14068
rect 22468 14059 22520 14068
rect 22468 14025 22477 14059
rect 22477 14025 22511 14059
rect 22511 14025 22520 14059
rect 22468 14016 22520 14025
rect 22928 14016 22980 14068
rect 23020 14016 23072 14068
rect 23204 13948 23256 14000
rect 23572 13948 23624 14000
rect 25504 14016 25556 14068
rect 26148 14016 26200 14068
rect 27436 14016 27488 14068
rect 28908 14016 28960 14068
rect 32772 14016 32824 14068
rect 33968 14016 34020 14068
rect 18788 13923 18840 13932
rect 18788 13889 18797 13923
rect 18797 13889 18831 13923
rect 18831 13889 18840 13923
rect 18788 13880 18840 13889
rect 18972 13923 19024 13932
rect 18972 13889 18981 13923
rect 18981 13889 19015 13923
rect 19015 13889 19024 13923
rect 18972 13880 19024 13889
rect 19248 13880 19300 13932
rect 22376 13923 22428 13932
rect 22376 13889 22385 13923
rect 22385 13889 22419 13923
rect 22419 13889 22428 13923
rect 22376 13880 22428 13889
rect 23388 13880 23440 13932
rect 27528 13948 27580 14000
rect 29644 13991 29696 14000
rect 29644 13957 29653 13991
rect 29653 13957 29687 13991
rect 29687 13957 29696 13991
rect 29644 13948 29696 13957
rect 29920 13948 29972 14000
rect 25320 13880 25372 13932
rect 28356 13923 28408 13932
rect 28356 13889 28365 13923
rect 28365 13889 28399 13923
rect 28399 13889 28408 13923
rect 28356 13880 28408 13889
rect 18696 13812 18748 13864
rect 19432 13812 19484 13864
rect 22744 13812 22796 13864
rect 23940 13855 23992 13864
rect 23940 13821 23949 13855
rect 23949 13821 23983 13855
rect 23983 13821 23992 13855
rect 23940 13812 23992 13821
rect 20720 13744 20772 13796
rect 23112 13744 23164 13796
rect 22008 13719 22060 13728
rect 22008 13685 22017 13719
rect 22017 13685 22051 13719
rect 22051 13685 22060 13719
rect 22008 13676 22060 13685
rect 22836 13676 22888 13728
rect 23204 13676 23256 13728
rect 27620 13812 27672 13864
rect 30656 13880 30708 13932
rect 30748 13923 30800 13932
rect 30748 13889 30757 13923
rect 30757 13889 30791 13923
rect 30791 13889 30800 13923
rect 30748 13880 30800 13889
rect 29000 13812 29052 13864
rect 31024 13880 31076 13932
rect 34520 13948 34572 14000
rect 36820 14059 36872 14068
rect 36820 14025 36829 14059
rect 36829 14025 36863 14059
rect 36863 14025 36872 14059
rect 36820 14016 36872 14025
rect 37556 14016 37608 14068
rect 39488 14016 39540 14068
rect 37740 13948 37792 14000
rect 31576 13923 31628 13932
rect 31576 13889 31585 13923
rect 31585 13889 31619 13923
rect 31619 13889 31628 13923
rect 31576 13880 31628 13889
rect 31668 13880 31720 13932
rect 33232 13923 33284 13932
rect 33232 13889 33241 13923
rect 33241 13889 33275 13923
rect 33275 13889 33284 13923
rect 33232 13880 33284 13889
rect 33508 13880 33560 13932
rect 34704 13923 34756 13932
rect 34704 13889 34713 13923
rect 34713 13889 34747 13923
rect 34747 13889 34756 13923
rect 34704 13880 34756 13889
rect 35348 13880 35400 13932
rect 35532 13880 35584 13932
rect 39396 13948 39448 14000
rect 27896 13744 27948 13796
rect 28816 13744 28868 13796
rect 30472 13787 30524 13796
rect 30472 13753 30481 13787
rect 30481 13753 30515 13787
rect 30515 13753 30524 13787
rect 30472 13744 30524 13753
rect 33968 13744 34020 13796
rect 36820 13744 36872 13796
rect 26148 13719 26200 13728
rect 26148 13685 26157 13719
rect 26157 13685 26191 13719
rect 26191 13685 26200 13719
rect 26148 13676 26200 13685
rect 32956 13676 33008 13728
rect 36268 13676 36320 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19340 13472 19392 13524
rect 22376 13472 22428 13524
rect 23572 13472 23624 13524
rect 23940 13472 23992 13524
rect 25320 13515 25372 13524
rect 25320 13481 25329 13515
rect 25329 13481 25363 13515
rect 25363 13481 25372 13515
rect 25320 13472 25372 13481
rect 24308 13404 24360 13456
rect 19984 13336 20036 13388
rect 20720 13336 20772 13388
rect 22652 13379 22704 13388
rect 22652 13345 22661 13379
rect 22661 13345 22695 13379
rect 22695 13345 22704 13379
rect 22652 13336 22704 13345
rect 24216 13336 24268 13388
rect 27344 13472 27396 13524
rect 32036 13472 32088 13524
rect 34520 13472 34572 13524
rect 34796 13472 34848 13524
rect 37280 13472 37332 13524
rect 39028 13472 39080 13524
rect 31484 13404 31536 13456
rect 20536 13268 20588 13320
rect 23388 13268 23440 13320
rect 24032 13268 24084 13320
rect 24768 13311 24820 13320
rect 24768 13277 24777 13311
rect 24777 13277 24811 13311
rect 24811 13277 24820 13311
rect 24768 13268 24820 13277
rect 24860 13311 24912 13320
rect 24860 13277 24869 13311
rect 24869 13277 24903 13311
rect 24903 13277 24912 13311
rect 24860 13268 24912 13277
rect 25688 13311 25740 13320
rect 25688 13277 25697 13311
rect 25697 13277 25731 13311
rect 25731 13277 25740 13311
rect 25688 13268 25740 13277
rect 26148 13268 26200 13320
rect 26332 13268 26384 13320
rect 27528 13336 27580 13388
rect 27804 13379 27856 13388
rect 27804 13345 27813 13379
rect 27813 13345 27847 13379
rect 27847 13345 27856 13379
rect 27804 13336 27856 13345
rect 29828 13379 29880 13388
rect 29828 13345 29837 13379
rect 29837 13345 29871 13379
rect 29871 13345 29880 13379
rect 29828 13336 29880 13345
rect 34244 13404 34296 13456
rect 32496 13379 32548 13388
rect 32496 13345 32505 13379
rect 32505 13345 32539 13379
rect 32539 13345 32548 13379
rect 32496 13336 32548 13345
rect 35164 13336 35216 13388
rect 35440 13379 35492 13388
rect 35440 13345 35449 13379
rect 35449 13345 35483 13379
rect 35483 13345 35492 13379
rect 35440 13336 35492 13345
rect 36084 13447 36136 13456
rect 36084 13413 36093 13447
rect 36093 13413 36127 13447
rect 36127 13413 36136 13447
rect 36084 13404 36136 13413
rect 20260 13132 20312 13184
rect 22008 13200 22060 13252
rect 23572 13200 23624 13252
rect 27896 13268 27948 13320
rect 28816 13268 28868 13320
rect 32128 13268 32180 13320
rect 22376 13132 22428 13184
rect 25596 13132 25648 13184
rect 26240 13132 26292 13184
rect 27344 13243 27396 13252
rect 27344 13209 27353 13243
rect 27353 13209 27387 13243
rect 27387 13209 27396 13243
rect 27344 13200 27396 13209
rect 28632 13200 28684 13252
rect 30288 13200 30340 13252
rect 26884 13132 26936 13184
rect 27620 13132 27672 13184
rect 29276 13132 29328 13184
rect 29460 13132 29512 13184
rect 30748 13200 30800 13252
rect 35992 13268 36044 13320
rect 36268 13311 36320 13320
rect 36268 13277 36277 13311
rect 36277 13277 36311 13311
rect 36311 13277 36320 13311
rect 36268 13268 36320 13277
rect 38660 13336 38712 13388
rect 36912 13311 36964 13320
rect 36912 13277 36921 13311
rect 36921 13277 36955 13311
rect 36955 13277 36964 13311
rect 36912 13268 36964 13277
rect 37372 13311 37424 13320
rect 37372 13277 37381 13311
rect 37381 13277 37415 13311
rect 37415 13277 37424 13311
rect 37372 13268 37424 13277
rect 37648 13268 37700 13320
rect 30656 13132 30708 13184
rect 33324 13132 33376 13184
rect 33968 13175 34020 13184
rect 33968 13141 33977 13175
rect 33977 13141 34011 13175
rect 34011 13141 34020 13175
rect 33968 13132 34020 13141
rect 35348 13132 35400 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 20904 12860 20956 12912
rect 23204 12928 23256 12980
rect 23572 12971 23624 12980
rect 23572 12937 23581 12971
rect 23581 12937 23615 12971
rect 23615 12937 23624 12971
rect 23572 12928 23624 12937
rect 24308 12928 24360 12980
rect 24676 12928 24728 12980
rect 22928 12860 22980 12912
rect 20352 12792 20404 12844
rect 20536 12835 20588 12844
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 22100 12792 22152 12844
rect 22744 12792 22796 12844
rect 23664 12656 23716 12708
rect 24216 12767 24268 12776
rect 24216 12733 24225 12767
rect 24225 12733 24259 12767
rect 24259 12733 24268 12767
rect 24216 12724 24268 12733
rect 24952 12792 25004 12844
rect 25964 12928 26016 12980
rect 27896 12928 27948 12980
rect 28632 12971 28684 12980
rect 28632 12937 28641 12971
rect 28641 12937 28675 12971
rect 28675 12937 28684 12971
rect 28632 12928 28684 12937
rect 29092 12971 29144 12980
rect 29092 12937 29101 12971
rect 29101 12937 29135 12971
rect 29135 12937 29144 12971
rect 29092 12928 29144 12937
rect 29460 12928 29512 12980
rect 30288 12971 30340 12980
rect 30288 12937 30297 12971
rect 30297 12937 30331 12971
rect 30331 12937 30340 12971
rect 30288 12928 30340 12937
rect 30656 12971 30708 12980
rect 30656 12937 30665 12971
rect 30665 12937 30699 12971
rect 30699 12937 30708 12971
rect 30656 12928 30708 12937
rect 30748 12971 30800 12980
rect 30748 12937 30757 12971
rect 30757 12937 30791 12971
rect 30791 12937 30800 12971
rect 30748 12928 30800 12937
rect 30840 12928 30892 12980
rect 35624 12928 35676 12980
rect 38568 12928 38620 12980
rect 26056 12860 26108 12912
rect 26332 12792 26384 12844
rect 26608 12835 26660 12844
rect 26608 12801 26617 12835
rect 26617 12801 26651 12835
rect 26651 12801 26660 12835
rect 26608 12792 26660 12801
rect 27068 12792 27120 12844
rect 28356 12860 28408 12912
rect 29368 12860 29420 12912
rect 27620 12835 27672 12844
rect 27620 12801 27629 12835
rect 27629 12801 27663 12835
rect 27663 12801 27672 12835
rect 27620 12792 27672 12801
rect 28080 12792 28132 12844
rect 29276 12792 29328 12844
rect 29920 12792 29972 12844
rect 30564 12792 30616 12844
rect 32128 12860 32180 12912
rect 27436 12724 27488 12776
rect 28264 12724 28316 12776
rect 29092 12724 29144 12776
rect 30196 12724 30248 12776
rect 22008 12588 22060 12640
rect 22284 12588 22336 12640
rect 23848 12588 23900 12640
rect 26332 12588 26384 12640
rect 26792 12588 26844 12640
rect 27436 12588 27488 12640
rect 27896 12631 27948 12640
rect 27896 12597 27905 12631
rect 27905 12597 27939 12631
rect 27939 12597 27948 12631
rect 31116 12724 31168 12776
rect 32312 12835 32364 12844
rect 32312 12801 32321 12835
rect 32321 12801 32355 12835
rect 32355 12801 32364 12835
rect 32312 12792 32364 12801
rect 32864 12835 32916 12844
rect 32864 12801 32873 12835
rect 32873 12801 32907 12835
rect 32907 12801 32916 12835
rect 32864 12792 32916 12801
rect 33324 12792 33376 12844
rect 33508 12835 33560 12844
rect 33508 12801 33517 12835
rect 33517 12801 33551 12835
rect 33551 12801 33560 12835
rect 33508 12792 33560 12801
rect 33692 12835 33744 12844
rect 33692 12801 33701 12835
rect 33701 12801 33735 12835
rect 33735 12801 33744 12835
rect 33692 12792 33744 12801
rect 34796 12792 34848 12844
rect 34520 12724 34572 12776
rect 35164 12767 35216 12776
rect 35164 12733 35173 12767
rect 35173 12733 35207 12767
rect 35207 12733 35216 12767
rect 35164 12724 35216 12733
rect 35532 12724 35584 12776
rect 36360 12792 36412 12844
rect 36636 12835 36688 12844
rect 36636 12801 36645 12835
rect 36645 12801 36679 12835
rect 36679 12801 36688 12835
rect 36636 12792 36688 12801
rect 36912 12724 36964 12776
rect 33140 12656 33192 12708
rect 27896 12588 27948 12597
rect 34612 12631 34664 12640
rect 34612 12597 34621 12631
rect 34621 12597 34655 12631
rect 34655 12597 34664 12631
rect 34612 12588 34664 12597
rect 38292 12631 38344 12640
rect 38292 12597 38301 12631
rect 38301 12597 38335 12631
rect 38335 12597 38344 12631
rect 38292 12588 38344 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 20352 12384 20404 12436
rect 19432 12291 19484 12300
rect 19432 12257 19441 12291
rect 19441 12257 19475 12291
rect 19475 12257 19484 12291
rect 19432 12248 19484 12257
rect 22284 12316 22336 12368
rect 23112 12384 23164 12436
rect 24584 12384 24636 12436
rect 22008 12180 22060 12232
rect 23020 12248 23072 12300
rect 23848 12248 23900 12300
rect 26608 12384 26660 12436
rect 32312 12384 32364 12436
rect 34796 12384 34848 12436
rect 26976 12316 27028 12368
rect 26332 12248 26384 12300
rect 28632 12248 28684 12300
rect 29000 12316 29052 12368
rect 31668 12316 31720 12368
rect 32680 12359 32732 12368
rect 32680 12325 32689 12359
rect 32689 12325 32723 12359
rect 32723 12325 32732 12359
rect 32680 12316 32732 12325
rect 26608 12223 26660 12232
rect 26608 12189 26617 12223
rect 26617 12189 26651 12223
rect 26651 12189 26660 12223
rect 26608 12180 26660 12189
rect 23848 12155 23900 12164
rect 23848 12121 23889 12155
rect 23889 12121 23900 12155
rect 23848 12112 23900 12121
rect 25044 12112 25096 12164
rect 26424 12112 26476 12164
rect 26884 12223 26936 12232
rect 26884 12189 26893 12223
rect 26893 12189 26927 12223
rect 26927 12189 26936 12223
rect 26884 12180 26936 12189
rect 26976 12180 27028 12232
rect 28540 12180 28592 12232
rect 29552 12248 29604 12300
rect 27252 12112 27304 12164
rect 29000 12223 29052 12232
rect 29000 12189 29009 12223
rect 29009 12189 29043 12223
rect 29043 12189 29052 12223
rect 29000 12180 29052 12189
rect 29184 12223 29236 12232
rect 29184 12189 29193 12223
rect 29193 12189 29227 12223
rect 29227 12189 29236 12223
rect 29184 12180 29236 12189
rect 29920 12223 29972 12232
rect 29920 12189 29929 12223
rect 29929 12189 29963 12223
rect 29963 12189 29972 12223
rect 29920 12180 29972 12189
rect 30656 12180 30708 12232
rect 30932 12223 30984 12232
rect 30932 12189 30941 12223
rect 30941 12189 30975 12223
rect 30975 12189 30984 12223
rect 30932 12180 30984 12189
rect 31024 12223 31076 12232
rect 31024 12189 31033 12223
rect 31033 12189 31067 12223
rect 31067 12189 31076 12223
rect 31024 12180 31076 12189
rect 31760 12248 31812 12300
rect 32956 12248 33008 12300
rect 33508 12248 33560 12300
rect 34612 12248 34664 12300
rect 29644 12112 29696 12164
rect 29736 12155 29788 12164
rect 29736 12121 29745 12155
rect 29745 12121 29779 12155
rect 29779 12121 29788 12155
rect 29736 12112 29788 12121
rect 30472 12112 30524 12164
rect 21732 12087 21784 12096
rect 21732 12053 21741 12087
rect 21741 12053 21775 12087
rect 21775 12053 21784 12087
rect 21732 12044 21784 12053
rect 23020 12087 23072 12096
rect 23020 12053 23029 12087
rect 23029 12053 23063 12087
rect 23063 12053 23072 12087
rect 23020 12044 23072 12053
rect 24952 12087 25004 12096
rect 24952 12053 24961 12087
rect 24961 12053 24995 12087
rect 24995 12053 25004 12087
rect 24952 12044 25004 12053
rect 25320 12087 25372 12096
rect 25320 12053 25329 12087
rect 25329 12053 25363 12087
rect 25363 12053 25372 12087
rect 25320 12044 25372 12053
rect 25780 12044 25832 12096
rect 31944 12180 31996 12232
rect 31392 12112 31444 12164
rect 33324 12223 33376 12232
rect 33324 12189 33333 12223
rect 33333 12189 33367 12223
rect 33367 12189 33376 12223
rect 33324 12180 33376 12189
rect 34796 12180 34848 12232
rect 33048 12112 33100 12164
rect 31760 12087 31812 12096
rect 31760 12053 31769 12087
rect 31769 12053 31803 12087
rect 31803 12053 31812 12087
rect 31760 12044 31812 12053
rect 32312 12044 32364 12096
rect 34520 12044 34572 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 20904 11840 20956 11892
rect 21732 11840 21784 11892
rect 22652 11840 22704 11892
rect 24308 11840 24360 11892
rect 25320 11840 25372 11892
rect 23756 11772 23808 11824
rect 24952 11772 25004 11824
rect 26056 11772 26108 11824
rect 26516 11883 26568 11892
rect 26516 11849 26525 11883
rect 26525 11849 26559 11883
rect 26559 11849 26568 11883
rect 26516 11840 26568 11849
rect 26608 11840 26660 11892
rect 27252 11840 27304 11892
rect 28540 11840 28592 11892
rect 22376 11747 22428 11756
rect 22376 11713 22385 11747
rect 22385 11713 22419 11747
rect 22419 11713 22428 11747
rect 22376 11704 22428 11713
rect 23204 11747 23256 11756
rect 23204 11713 23213 11747
rect 23213 11713 23247 11747
rect 23247 11713 23256 11747
rect 23204 11704 23256 11713
rect 20628 11543 20680 11552
rect 20628 11509 20637 11543
rect 20637 11509 20671 11543
rect 20671 11509 20680 11543
rect 20628 11500 20680 11509
rect 22008 11543 22060 11552
rect 22008 11509 22017 11543
rect 22017 11509 22051 11543
rect 22051 11509 22060 11543
rect 22008 11500 22060 11509
rect 22744 11636 22796 11688
rect 24860 11704 24912 11756
rect 22192 11568 22244 11620
rect 24308 11679 24360 11688
rect 24308 11645 24317 11679
rect 24317 11645 24351 11679
rect 24351 11645 24360 11679
rect 24308 11636 24360 11645
rect 25688 11704 25740 11756
rect 26792 11636 26844 11688
rect 28632 11772 28684 11824
rect 30012 11840 30064 11892
rect 31760 11840 31812 11892
rect 31852 11840 31904 11892
rect 34796 11840 34848 11892
rect 35348 11840 35400 11892
rect 28724 11747 28776 11756
rect 28724 11713 28733 11747
rect 28733 11713 28767 11747
rect 28767 11713 28776 11747
rect 28724 11704 28776 11713
rect 30380 11704 30432 11756
rect 31024 11704 31076 11756
rect 27528 11568 27580 11620
rect 27068 11500 27120 11552
rect 28172 11500 28224 11552
rect 30196 11679 30248 11688
rect 30196 11645 30205 11679
rect 30205 11645 30239 11679
rect 30239 11645 30248 11679
rect 30196 11636 30248 11645
rect 32312 11704 32364 11756
rect 31300 11679 31352 11688
rect 31300 11645 31309 11679
rect 31309 11645 31343 11679
rect 31343 11645 31352 11679
rect 31300 11636 31352 11645
rect 32496 11772 32548 11824
rect 33140 11704 33192 11756
rect 33600 11747 33652 11756
rect 33600 11713 33609 11747
rect 33609 11713 33643 11747
rect 33643 11713 33652 11747
rect 33600 11704 33652 11713
rect 33784 11747 33836 11756
rect 33784 11713 33793 11747
rect 33793 11713 33827 11747
rect 33827 11713 33836 11747
rect 33784 11704 33836 11713
rect 34796 11704 34848 11756
rect 32864 11679 32916 11688
rect 32864 11645 32873 11679
rect 32873 11645 32907 11679
rect 32907 11645 32916 11679
rect 32864 11636 32916 11645
rect 29552 11543 29604 11552
rect 29552 11509 29561 11543
rect 29561 11509 29595 11543
rect 29595 11509 29604 11543
rect 29552 11500 29604 11509
rect 30656 11500 30708 11552
rect 30840 11500 30892 11552
rect 31392 11500 31444 11552
rect 32404 11543 32456 11552
rect 32404 11509 32413 11543
rect 32413 11509 32447 11543
rect 32447 11509 32456 11543
rect 32404 11500 32456 11509
rect 32496 11500 32548 11552
rect 33048 11500 33100 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 22376 11339 22428 11348
rect 22376 11305 22385 11339
rect 22385 11305 22419 11339
rect 22419 11305 22428 11339
rect 22376 11296 22428 11305
rect 23204 11296 23256 11348
rect 26792 11296 26844 11348
rect 27068 11296 27120 11348
rect 30380 11296 30432 11348
rect 31024 11296 31076 11348
rect 19432 11160 19484 11212
rect 23756 11203 23808 11212
rect 23756 11169 23765 11203
rect 23765 11169 23799 11203
rect 23799 11169 23808 11203
rect 23756 11160 23808 11169
rect 24216 11160 24268 11212
rect 24308 11160 24360 11212
rect 26424 11160 26476 11212
rect 22008 11092 22060 11144
rect 23296 10999 23348 11008
rect 23296 10965 23305 10999
rect 23305 10965 23339 10999
rect 23339 10965 23348 10999
rect 23296 10956 23348 10965
rect 23480 10956 23532 11008
rect 26792 11135 26844 11144
rect 26792 11101 26801 11135
rect 26801 11101 26835 11135
rect 26835 11101 26844 11135
rect 26792 11092 26844 11101
rect 27068 11203 27120 11212
rect 27068 11169 27077 11203
rect 27077 11169 27111 11203
rect 27111 11169 27120 11203
rect 27068 11160 27120 11169
rect 27160 11092 27212 11144
rect 27804 11203 27856 11212
rect 27804 11169 27813 11203
rect 27813 11169 27847 11203
rect 27847 11169 27856 11203
rect 27804 11160 27856 11169
rect 29552 11092 29604 11144
rect 29828 11160 29880 11212
rect 32496 11296 32548 11348
rect 33140 11296 33192 11348
rect 34796 11296 34848 11348
rect 35440 11203 35492 11212
rect 30472 11024 30524 11076
rect 30656 11067 30708 11076
rect 30656 11033 30679 11067
rect 30679 11033 30708 11067
rect 30656 11024 30708 11033
rect 32404 11024 32456 11076
rect 32956 11024 33008 11076
rect 35440 11169 35449 11203
rect 35449 11169 35483 11203
rect 35483 11169 35492 11203
rect 35440 11160 35492 11169
rect 35348 11092 35400 11144
rect 39212 11092 39264 11144
rect 34520 11024 34572 11076
rect 38108 11067 38160 11076
rect 38108 11033 38117 11067
rect 38117 11033 38151 11067
rect 38151 11033 38160 11067
rect 38108 11024 38160 11033
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 20904 10752 20956 10804
rect 23020 10752 23072 10804
rect 28724 10752 28776 10804
rect 29644 10752 29696 10804
rect 30288 10752 30340 10804
rect 33692 10795 33744 10804
rect 33692 10761 33701 10795
rect 33701 10761 33735 10795
rect 33735 10761 33744 10795
rect 33692 10752 33744 10761
rect 20628 10684 20680 10736
rect 19432 10616 19484 10668
rect 20536 10616 20588 10668
rect 22376 10616 22428 10668
rect 22652 10616 22704 10668
rect 23296 10616 23348 10668
rect 27712 10616 27764 10668
rect 27804 10616 27856 10668
rect 28356 10659 28408 10668
rect 28356 10625 28390 10659
rect 28390 10625 28408 10659
rect 28356 10616 28408 10625
rect 29828 10616 29880 10668
rect 30196 10659 30248 10668
rect 30196 10625 30230 10659
rect 30230 10625 30248 10659
rect 30196 10616 30248 10625
rect 32404 10616 32456 10668
rect 22192 10548 22244 10600
rect 22284 10591 22336 10600
rect 22284 10557 22293 10591
rect 22293 10557 22327 10591
rect 22327 10557 22336 10591
rect 22284 10548 22336 10557
rect 23480 10412 23532 10464
rect 29460 10455 29512 10464
rect 29460 10421 29469 10455
rect 29469 10421 29503 10455
rect 29503 10421 29512 10455
rect 29460 10412 29512 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 22100 10251 22152 10260
rect 22100 10217 22109 10251
rect 22109 10217 22143 10251
rect 22143 10217 22152 10251
rect 22100 10208 22152 10217
rect 22284 10208 22336 10260
rect 27528 10251 27580 10260
rect 27528 10217 27537 10251
rect 27537 10217 27571 10251
rect 27571 10217 27580 10251
rect 27528 10208 27580 10217
rect 27712 10208 27764 10260
rect 30196 10251 30248 10260
rect 30196 10217 30205 10251
rect 30205 10217 30239 10251
rect 30239 10217 30248 10251
rect 30196 10208 30248 10217
rect 30380 10208 30432 10260
rect 30288 10140 30340 10192
rect 23112 10004 23164 10056
rect 23480 10004 23532 10056
rect 27252 10072 27304 10124
rect 30472 10072 30524 10124
rect 23848 10004 23900 10056
rect 27804 10004 27856 10056
rect 28724 10004 28776 10056
rect 30656 10072 30708 10124
rect 31300 10072 31352 10124
rect 32404 10251 32456 10260
rect 32404 10217 32413 10251
rect 32413 10217 32447 10251
rect 32447 10217 32456 10251
rect 32404 10208 32456 10217
rect 32864 10115 32916 10124
rect 27160 9936 27212 9988
rect 29736 9868 29788 9920
rect 32864 10081 32873 10115
rect 32873 10081 32907 10115
rect 32907 10081 32916 10115
rect 32864 10072 32916 10081
rect 32956 10115 33008 10124
rect 32956 10081 32965 10115
rect 32965 10081 32999 10115
rect 32999 10081 33008 10115
rect 32956 10072 33008 10081
rect 33692 10004 33744 10056
rect 34336 10004 34388 10056
rect 30656 9911 30708 9920
rect 30656 9877 30665 9911
rect 30665 9877 30699 9911
rect 30699 9877 30708 9911
rect 38108 9979 38160 9988
rect 38108 9945 38117 9979
rect 38117 9945 38151 9979
rect 38151 9945 38160 9979
rect 38108 9936 38160 9945
rect 30656 9868 30708 9877
rect 31760 9911 31812 9920
rect 31760 9877 31769 9911
rect 31769 9877 31803 9911
rect 31803 9877 31812 9911
rect 31760 9868 31812 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 27160 9707 27212 9716
rect 27160 9673 27169 9707
rect 27169 9673 27203 9707
rect 27203 9673 27212 9707
rect 27160 9664 27212 9673
rect 27528 9707 27580 9716
rect 27528 9673 27537 9707
rect 27537 9673 27571 9707
rect 27571 9673 27580 9707
rect 27528 9664 27580 9673
rect 27252 9596 27304 9648
rect 28356 9664 28408 9716
rect 28816 9664 28868 9716
rect 30656 9664 30708 9716
rect 29460 9596 29512 9648
rect 30840 9596 30892 9648
rect 27436 9528 27488 9580
rect 29736 9571 29788 9580
rect 29736 9537 29745 9571
rect 29745 9537 29779 9571
rect 29779 9537 29788 9571
rect 29736 9528 29788 9537
rect 31024 9571 31076 9580
rect 31024 9537 31033 9571
rect 31033 9537 31067 9571
rect 31067 9537 31076 9571
rect 31024 9528 31076 9537
rect 29184 9460 29236 9512
rect 30748 9460 30800 9512
rect 29000 9324 29052 9376
rect 31760 9528 31812 9580
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 32588 8984 32640 9036
rect 37280 8984 37332 9036
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 38200 8440 38252 8492
rect 38108 8415 38160 8424
rect 38108 8381 38117 8415
rect 38117 8381 38151 8415
rect 38151 8381 38160 8415
rect 38108 8372 38160 8381
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 37832 7395 37884 7404
rect 37832 7361 37841 7395
rect 37841 7361 37875 7395
rect 37875 7361 37884 7395
rect 37832 7352 37884 7361
rect 38108 7327 38160 7336
rect 38108 7293 38117 7327
rect 38117 7293 38151 7327
rect 38151 7293 38160 7327
rect 38108 7284 38160 7293
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 37280 5652 37332 5704
rect 38108 5627 38160 5636
rect 38108 5593 38117 5627
rect 38117 5593 38151 5627
rect 38151 5593 38160 5627
rect 38108 5584 38160 5593
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 37832 4607 37884 4616
rect 37832 4573 37841 4607
rect 37841 4573 37875 4607
rect 37875 4573 37884 4607
rect 37832 4564 37884 4573
rect 38108 4539 38160 4548
rect 38108 4505 38117 4539
rect 38117 4505 38151 4539
rect 38151 4505 38160 4539
rect 38108 4496 38160 4505
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 37372 3000 37424 3052
rect 38108 2975 38160 2984
rect 38108 2941 38117 2975
rect 38117 2941 38151 2975
rect 38151 2941 38160 2975
rect 38108 2932 38160 2941
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 37832 2431 37884 2440
rect 37832 2397 37841 2431
rect 37841 2397 37875 2431
rect 37875 2397 37884 2431
rect 37832 2388 37884 2397
rect 38108 2363 38160 2372
rect 38108 2329 38117 2363
rect 38117 2329 38151 2363
rect 38151 2329 38160 2363
rect 38108 2320 38160 2329
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 1766 39200 1822 40000
rect 4988 39296 5040 39302
rect 4988 39238 5040 39244
rect 1780 37262 1808 39200
rect 3976 39024 4028 39030
rect 3976 38966 4028 38972
rect 3332 38888 3384 38894
rect 3332 38830 3384 38836
rect 3056 38548 3108 38554
rect 3056 38490 3108 38496
rect 2596 38004 2648 38010
rect 2596 37946 2648 37952
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1676 36780 1728 36786
rect 1676 36722 1728 36728
rect 1688 36281 1716 36722
rect 1768 36576 1820 36582
rect 1768 36518 1820 36524
rect 2412 36576 2464 36582
rect 2412 36518 2464 36524
rect 1674 36272 1730 36281
rect 1674 36207 1730 36216
rect 1780 27985 1808 36518
rect 1766 27976 1822 27985
rect 1766 27911 1822 27920
rect 2424 26042 2452 36518
rect 2608 36378 2636 37946
rect 3068 36922 3096 38490
rect 3056 36916 3108 36922
rect 3056 36858 3108 36864
rect 3240 36576 3292 36582
rect 3240 36518 3292 36524
rect 2596 36372 2648 36378
rect 2596 36314 2648 36320
rect 3252 36174 3280 36518
rect 3344 36378 3372 38830
rect 3606 38312 3662 38321
rect 3606 38247 3662 38256
rect 3424 37256 3476 37262
rect 3424 37198 3476 37204
rect 3332 36372 3384 36378
rect 3332 36314 3384 36320
rect 3240 36168 3292 36174
rect 3240 36110 3292 36116
rect 3436 35766 3464 37198
rect 3516 37120 3568 37126
rect 3516 37062 3568 37068
rect 3528 36038 3556 37062
rect 3516 36032 3568 36038
rect 3516 35974 3568 35980
rect 3424 35760 3476 35766
rect 3424 35702 3476 35708
rect 3620 34746 3648 38247
rect 3700 37664 3752 37670
rect 3700 37606 3752 37612
rect 3712 36922 3740 37606
rect 3792 37120 3844 37126
rect 3792 37062 3844 37068
rect 3700 36916 3752 36922
rect 3700 36858 3752 36864
rect 3700 35488 3752 35494
rect 3700 35430 3752 35436
rect 3608 34740 3660 34746
rect 3608 34682 3660 34688
rect 3516 34604 3568 34610
rect 3516 34546 3568 34552
rect 2688 32360 2740 32366
rect 2688 32302 2740 32308
rect 2412 26036 2464 26042
rect 2412 25978 2464 25984
rect 2700 24410 2728 32302
rect 3528 27606 3556 34546
rect 3516 27600 3568 27606
rect 3516 27542 3568 27548
rect 2688 24404 2740 24410
rect 2688 24346 2740 24352
rect 3712 22681 3740 35430
rect 3804 25129 3832 37062
rect 3988 33590 4016 38966
rect 4894 38720 4950 38729
rect 4894 38655 4950 38664
rect 4068 38072 4120 38078
rect 4068 38014 4120 38020
rect 4080 33998 4108 38014
rect 4804 37868 4856 37874
rect 4804 37810 4856 37816
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4528 37256 4580 37262
rect 4528 37198 4580 37204
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 4540 36650 4568 37198
rect 4632 37126 4660 37198
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 4712 37120 4764 37126
rect 4712 37062 4764 37068
rect 4528 36644 4580 36650
rect 4528 36586 4580 36592
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4342 35728 4398 35737
rect 4342 35663 4344 35672
rect 4396 35663 4398 35672
rect 4528 35692 4580 35698
rect 4344 35634 4396 35640
rect 4528 35634 4580 35640
rect 4540 35494 4568 35634
rect 4528 35488 4580 35494
rect 4528 35430 4580 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4344 35284 4396 35290
rect 4344 35226 4396 35232
rect 4356 35086 4384 35226
rect 4344 35080 4396 35086
rect 4344 35022 4396 35028
rect 4356 34649 4384 35022
rect 4620 34944 4672 34950
rect 4620 34886 4672 34892
rect 4342 34640 4398 34649
rect 4160 34604 4212 34610
rect 4342 34575 4398 34584
rect 4160 34546 4212 34552
rect 4172 34406 4200 34546
rect 4160 34400 4212 34406
rect 4632 34377 4660 34886
rect 4160 34342 4212 34348
rect 4618 34368 4674 34377
rect 4214 34300 4522 34309
rect 4618 34303 4674 34312
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4068 33992 4120 33998
rect 4068 33934 4120 33940
rect 4068 33856 4120 33862
rect 4068 33798 4120 33804
rect 3976 33584 4028 33590
rect 3976 33526 4028 33532
rect 3884 33312 3936 33318
rect 3884 33254 3936 33260
rect 3790 25120 3846 25129
rect 3790 25055 3846 25064
rect 3698 22672 3754 22681
rect 3698 22607 3754 22616
rect 3896 17105 3924 33254
rect 4080 32960 4108 33798
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4620 33040 4672 33046
rect 4620 32982 4672 32988
rect 3988 32932 4108 32960
rect 3988 29850 4016 32932
rect 4526 32600 4582 32609
rect 4526 32535 4582 32544
rect 4540 32434 4568 32535
rect 4528 32428 4580 32434
rect 4528 32370 4580 32376
rect 4632 32230 4660 32982
rect 4724 32337 4752 37062
rect 4816 36922 4844 37810
rect 4804 36916 4856 36922
rect 4804 36858 4856 36864
rect 4908 36530 4936 38655
rect 5000 36854 5028 39238
rect 5078 39200 5134 40000
rect 6826 39264 6882 39273
rect 5908 39228 5960 39234
rect 5092 37262 5120 39200
rect 6826 39199 6882 39208
rect 8390 39200 8446 40000
rect 11702 39200 11758 40000
rect 15014 39200 15070 40000
rect 18326 39200 18382 40000
rect 21638 39200 21694 40000
rect 24950 39200 25006 40000
rect 28262 39200 28318 40000
rect 31574 39200 31630 40000
rect 34886 39200 34942 40000
rect 35806 39400 35862 39409
rect 35806 39335 35862 39344
rect 5908 39170 5960 39176
rect 5354 38992 5410 39001
rect 5264 38956 5316 38962
rect 5354 38927 5410 38936
rect 5264 38898 5316 38904
rect 5170 37768 5226 37777
rect 5170 37703 5226 37712
rect 5080 37256 5132 37262
rect 5080 37198 5132 37204
rect 5078 36952 5134 36961
rect 5078 36887 5134 36896
rect 4988 36848 5040 36854
rect 4988 36790 5040 36796
rect 4988 36644 5040 36650
rect 4988 36586 5040 36592
rect 4816 36502 4936 36530
rect 4816 35834 4844 36502
rect 4894 36408 4950 36417
rect 4894 36343 4950 36352
rect 4804 35828 4856 35834
rect 4804 35770 4856 35776
rect 4804 35692 4856 35698
rect 4804 35634 4856 35640
rect 4816 34950 4844 35634
rect 4804 34944 4856 34950
rect 4804 34886 4856 34892
rect 4802 34776 4858 34785
rect 4908 34746 4936 36343
rect 5000 35873 5028 36586
rect 5092 36174 5120 36887
rect 5080 36168 5132 36174
rect 5080 36110 5132 36116
rect 5184 35986 5212 37703
rect 5276 36378 5304 38898
rect 5368 37369 5396 38927
rect 5540 38820 5592 38826
rect 5540 38762 5592 38768
rect 5354 37360 5410 37369
rect 5354 37295 5410 37304
rect 5448 36916 5500 36922
rect 5448 36858 5500 36864
rect 5356 36848 5408 36854
rect 5356 36790 5408 36796
rect 5264 36372 5316 36378
rect 5264 36314 5316 36320
rect 5092 35958 5212 35986
rect 4986 35864 5042 35873
rect 4986 35799 5042 35808
rect 4988 35692 5040 35698
rect 4988 35634 5040 35640
rect 5000 35290 5028 35634
rect 4988 35284 5040 35290
rect 4988 35226 5040 35232
rect 5092 35034 5120 35958
rect 5170 35864 5226 35873
rect 5170 35799 5226 35808
rect 5000 35006 5120 35034
rect 4802 34711 4858 34720
rect 4896 34740 4948 34746
rect 4816 33658 4844 34711
rect 4896 34682 4948 34688
rect 5000 34202 5028 35006
rect 5080 34944 5132 34950
rect 5184 34921 5212 35799
rect 5368 35766 5396 36790
rect 5460 36689 5488 36858
rect 5446 36680 5502 36689
rect 5446 36615 5502 36624
rect 5448 36576 5500 36582
rect 5448 36518 5500 36524
rect 5460 36174 5488 36518
rect 5448 36168 5500 36174
rect 5448 36110 5500 36116
rect 5460 35766 5488 36110
rect 5356 35760 5408 35766
rect 5356 35702 5408 35708
rect 5448 35760 5500 35766
rect 5448 35702 5500 35708
rect 5264 35692 5316 35698
rect 5264 35634 5316 35640
rect 5276 35290 5304 35634
rect 5264 35284 5316 35290
rect 5264 35226 5316 35232
rect 5080 34886 5132 34892
rect 5170 34912 5226 34921
rect 5092 34785 5120 34886
rect 5170 34847 5226 34856
rect 5078 34776 5134 34785
rect 5078 34711 5134 34720
rect 5172 34740 5224 34746
rect 5172 34682 5224 34688
rect 5078 34640 5134 34649
rect 5078 34575 5134 34584
rect 4988 34196 5040 34202
rect 4988 34138 5040 34144
rect 4988 33992 5040 33998
rect 4988 33934 5040 33940
rect 4896 33924 4948 33930
rect 4896 33866 4948 33872
rect 4804 33652 4856 33658
rect 4804 33594 4856 33600
rect 4804 33516 4856 33522
rect 4804 33458 4856 33464
rect 4816 33318 4844 33458
rect 4908 33454 4936 33866
rect 5000 33658 5028 33934
rect 4988 33652 5040 33658
rect 4988 33594 5040 33600
rect 4896 33448 4948 33454
rect 4896 33390 4948 33396
rect 4804 33312 4856 33318
rect 4804 33254 4856 33260
rect 4896 33312 4948 33318
rect 4896 33254 4948 33260
rect 4710 32328 4766 32337
rect 4710 32263 4766 32272
rect 4068 32224 4120 32230
rect 4068 32166 4120 32172
rect 4620 32224 4672 32230
rect 4620 32166 4672 32172
rect 4712 32224 4764 32230
rect 4712 32166 4764 32172
rect 3976 29844 4028 29850
rect 3976 29786 4028 29792
rect 4080 24857 4108 32166
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4434 31920 4490 31929
rect 4434 31855 4436 31864
rect 4488 31855 4490 31864
rect 4436 31826 4488 31832
rect 4620 31680 4672 31686
rect 4620 31622 4672 31628
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4528 29844 4580 29850
rect 4528 29786 4580 29792
rect 4540 28966 4568 29786
rect 4632 29034 4660 31622
rect 4620 29028 4672 29034
rect 4620 28970 4672 28976
rect 4528 28960 4580 28966
rect 4528 28902 4580 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4724 27674 4752 32166
rect 4712 27668 4764 27674
rect 4712 27610 4764 27616
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4816 25401 4844 33254
rect 4908 31686 4936 33254
rect 4988 32904 5040 32910
rect 4986 32872 4988 32881
rect 5040 32872 5042 32881
rect 4986 32807 5042 32816
rect 4988 31816 5040 31822
rect 4988 31758 5040 31764
rect 4896 31680 4948 31686
rect 4896 31622 4948 31628
rect 4894 31512 4950 31521
rect 4894 31447 4950 31456
rect 4908 26761 4936 31447
rect 4894 26752 4950 26761
rect 4894 26687 4950 26696
rect 5000 26217 5028 31758
rect 5092 31278 5120 34575
rect 5184 34066 5212 34682
rect 5172 34060 5224 34066
rect 5172 34002 5224 34008
rect 5172 32768 5224 32774
rect 5172 32710 5224 32716
rect 5184 32298 5212 32710
rect 5172 32292 5224 32298
rect 5172 32234 5224 32240
rect 5172 31340 5224 31346
rect 5172 31282 5224 31288
rect 5080 31272 5132 31278
rect 5080 31214 5132 31220
rect 5080 30592 5132 30598
rect 5080 30534 5132 30540
rect 4986 26208 5042 26217
rect 4986 26143 5042 26152
rect 4802 25392 4858 25401
rect 4802 25327 4858 25336
rect 4066 24848 4122 24857
rect 4066 24783 4122 24792
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 5092 22001 5120 30534
rect 5078 21992 5134 22001
rect 5078 21927 5134 21936
rect 5184 21418 5212 31282
rect 5276 31113 5304 35226
rect 5368 34950 5396 35702
rect 5448 35488 5500 35494
rect 5448 35430 5500 35436
rect 5356 34944 5408 34950
rect 5356 34886 5408 34892
rect 5460 33833 5488 35430
rect 5552 35222 5580 38762
rect 5816 38208 5868 38214
rect 5816 38150 5868 38156
rect 5724 37188 5776 37194
rect 5724 37130 5776 37136
rect 5736 36825 5764 37130
rect 5722 36816 5778 36825
rect 5632 36780 5684 36786
rect 5722 36751 5724 36760
rect 5632 36722 5684 36728
rect 5776 36751 5778 36760
rect 5724 36722 5776 36728
rect 5540 35216 5592 35222
rect 5540 35158 5592 35164
rect 5540 35080 5592 35086
rect 5540 35022 5592 35028
rect 5552 34610 5580 35022
rect 5540 34604 5592 34610
rect 5540 34546 5592 34552
rect 5540 34468 5592 34474
rect 5540 34410 5592 34416
rect 5552 34066 5580 34410
rect 5540 34060 5592 34066
rect 5540 34002 5592 34008
rect 5446 33824 5502 33833
rect 5446 33759 5502 33768
rect 5356 33516 5408 33522
rect 5356 33458 5408 33464
rect 5368 31822 5396 33458
rect 5644 33454 5672 36722
rect 5828 36106 5856 38150
rect 5920 36174 5948 39170
rect 6644 38752 6696 38758
rect 6644 38694 6696 38700
rect 6184 38616 6236 38622
rect 6184 38558 6236 38564
rect 6458 38584 6514 38593
rect 6000 38276 6052 38282
rect 6000 38218 6052 38224
rect 6012 36922 6040 38218
rect 6000 36916 6052 36922
rect 6000 36858 6052 36864
rect 5908 36168 5960 36174
rect 5908 36110 5960 36116
rect 5816 36100 5868 36106
rect 5816 36042 5868 36048
rect 6092 36100 6144 36106
rect 6092 36042 6144 36048
rect 5828 35698 5856 36042
rect 6104 36009 6132 36042
rect 6090 36000 6146 36009
rect 6090 35935 6146 35944
rect 6196 35834 6224 38558
rect 6458 38519 6514 38528
rect 6276 38480 6328 38486
rect 6276 38422 6328 38428
rect 6184 35828 6236 35834
rect 6184 35770 6236 35776
rect 5816 35692 5868 35698
rect 5816 35634 5868 35640
rect 5908 35488 5960 35494
rect 5908 35430 5960 35436
rect 5920 35086 5948 35430
rect 5908 35080 5960 35086
rect 5908 35022 5960 35028
rect 5920 34678 5948 35022
rect 6000 34944 6052 34950
rect 6000 34886 6052 34892
rect 6092 34944 6144 34950
rect 6092 34886 6144 34892
rect 5908 34672 5960 34678
rect 5908 34614 5960 34620
rect 5724 34604 5776 34610
rect 5724 34546 5776 34552
rect 5632 33448 5684 33454
rect 5632 33390 5684 33396
rect 5736 33130 5764 34546
rect 5908 34536 5960 34542
rect 5908 34478 5960 34484
rect 5814 34096 5870 34105
rect 5814 34031 5870 34040
rect 5828 33522 5856 34031
rect 5816 33516 5868 33522
rect 5816 33458 5868 33464
rect 5816 33312 5868 33318
rect 5814 33280 5816 33289
rect 5868 33280 5870 33289
rect 5814 33215 5870 33224
rect 5644 33102 5764 33130
rect 5644 32910 5672 33102
rect 5632 32904 5684 32910
rect 5632 32846 5684 32852
rect 5724 32904 5776 32910
rect 5724 32846 5776 32852
rect 5448 32768 5500 32774
rect 5448 32710 5500 32716
rect 5460 31890 5488 32710
rect 5632 32292 5684 32298
rect 5632 32234 5684 32240
rect 5448 31884 5500 31890
rect 5448 31826 5500 31832
rect 5356 31816 5408 31822
rect 5356 31758 5408 31764
rect 5262 31104 5318 31113
rect 5262 31039 5318 31048
rect 5368 30954 5396 31758
rect 5540 31680 5592 31686
rect 5540 31622 5592 31628
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 5276 30926 5396 30954
rect 5276 26246 5304 30926
rect 5356 30728 5408 30734
rect 5354 30696 5356 30705
rect 5408 30696 5410 30705
rect 5354 30631 5410 30640
rect 5356 27600 5408 27606
rect 5356 27542 5408 27548
rect 5264 26240 5316 26246
rect 5264 26182 5316 26188
rect 5368 24818 5396 27542
rect 5460 26081 5488 31078
rect 5552 29481 5580 31622
rect 5644 31385 5672 32234
rect 5630 31376 5686 31385
rect 5736 31346 5764 32846
rect 5816 32428 5868 32434
rect 5816 32370 5868 32376
rect 5828 32337 5856 32370
rect 5814 32328 5870 32337
rect 5814 32263 5870 32272
rect 5816 32224 5868 32230
rect 5816 32166 5868 32172
rect 5828 31958 5856 32166
rect 5816 31952 5868 31958
rect 5816 31894 5868 31900
rect 5828 31822 5856 31894
rect 5816 31816 5868 31822
rect 5816 31758 5868 31764
rect 5920 31362 5948 34478
rect 6012 32434 6040 34886
rect 6104 34066 6132 34886
rect 6092 34060 6144 34066
rect 6092 34002 6144 34008
rect 6184 33992 6236 33998
rect 6184 33934 6236 33940
rect 6196 33862 6224 33934
rect 6092 33856 6144 33862
rect 6092 33798 6144 33804
rect 6184 33856 6236 33862
rect 6184 33798 6236 33804
rect 6000 32428 6052 32434
rect 6000 32370 6052 32376
rect 6012 32337 6040 32370
rect 5998 32328 6054 32337
rect 5998 32263 6054 32272
rect 6000 31816 6052 31822
rect 6104 31793 6132 33798
rect 6184 33040 6236 33046
rect 6184 32982 6236 32988
rect 6000 31758 6052 31764
rect 6090 31784 6146 31793
rect 5630 31311 5686 31320
rect 5724 31340 5776 31346
rect 5724 31282 5776 31288
rect 5828 31334 5948 31362
rect 5736 30569 5764 31282
rect 5722 30560 5778 30569
rect 5722 30495 5778 30504
rect 5538 29472 5594 29481
rect 5538 29407 5594 29416
rect 5828 28762 5856 31334
rect 5908 31272 5960 31278
rect 5906 31240 5908 31249
rect 5960 31240 5962 31249
rect 5906 31175 5962 31184
rect 6012 30938 6040 31758
rect 6196 31754 6224 32982
rect 6288 32450 6316 38422
rect 6368 38140 6420 38146
rect 6368 38082 6420 38088
rect 6380 32910 6408 38082
rect 6472 33046 6500 38519
rect 6552 37188 6604 37194
rect 6552 37130 6604 37136
rect 6564 35873 6592 37130
rect 6550 35864 6606 35873
rect 6656 35834 6684 38694
rect 6736 37800 6788 37806
rect 6736 37742 6788 37748
rect 6748 36378 6776 37742
rect 6736 36372 6788 36378
rect 6736 36314 6788 36320
rect 6840 36088 6868 39199
rect 8404 39114 8432 39200
rect 11716 39166 11744 39200
rect 8220 39086 8432 39114
rect 10508 39160 10560 39166
rect 11704 39160 11756 39166
rect 10508 39102 10560 39108
rect 11242 39128 11298 39137
rect 7748 38412 7800 38418
rect 7748 38354 7800 38360
rect 7012 38344 7064 38350
rect 7012 38286 7064 38292
rect 6920 37732 6972 37738
rect 6920 37674 6972 37680
rect 6748 36060 6868 36088
rect 6550 35799 6606 35808
rect 6644 35828 6696 35834
rect 6644 35770 6696 35776
rect 6748 35086 6776 36060
rect 6932 35986 6960 37674
rect 7024 37330 7052 38286
rect 7288 37936 7340 37942
rect 7288 37878 7340 37884
rect 7378 37904 7434 37913
rect 7102 37360 7158 37369
rect 7012 37324 7064 37330
rect 7102 37295 7158 37304
rect 7012 37266 7064 37272
rect 7012 36780 7064 36786
rect 7012 36722 7064 36728
rect 7024 36553 7052 36722
rect 7010 36544 7066 36553
rect 7010 36479 7066 36488
rect 7024 36038 7052 36479
rect 6840 35958 6960 35986
rect 7012 36032 7064 36038
rect 7012 35974 7064 35980
rect 6840 35630 6868 35958
rect 6920 35760 6972 35766
rect 6920 35702 6972 35708
rect 6828 35624 6880 35630
rect 6828 35566 6880 35572
rect 6826 35184 6882 35193
rect 6932 35154 6960 35702
rect 7116 35698 7144 37295
rect 7196 37256 7248 37262
rect 7196 37198 7248 37204
rect 7208 36310 7236 37198
rect 7300 37126 7328 37878
rect 7378 37839 7434 37848
rect 7288 37120 7340 37126
rect 7288 37062 7340 37068
rect 7196 36304 7248 36310
rect 7196 36246 7248 36252
rect 7208 36106 7236 36246
rect 7196 36100 7248 36106
rect 7196 36042 7248 36048
rect 7300 35986 7328 37062
rect 7208 35958 7328 35986
rect 7104 35692 7156 35698
rect 7104 35634 7156 35640
rect 6826 35119 6882 35128
rect 6920 35148 6972 35154
rect 6840 35086 6868 35119
rect 6920 35090 6972 35096
rect 6736 35080 6788 35086
rect 6656 35040 6736 35068
rect 6552 34944 6604 34950
rect 6552 34886 6604 34892
rect 6564 34746 6592 34886
rect 6552 34740 6604 34746
rect 6552 34682 6604 34688
rect 6552 34060 6604 34066
rect 6552 34002 6604 34008
rect 6564 33930 6592 34002
rect 6656 33998 6684 35040
rect 6736 35022 6788 35028
rect 6828 35080 6880 35086
rect 6828 35022 6880 35028
rect 6840 34202 6868 35022
rect 6932 34610 6960 35090
rect 7208 34950 7236 35958
rect 7392 35816 7420 37839
rect 7656 36712 7708 36718
rect 7656 36654 7708 36660
rect 7472 36576 7524 36582
rect 7472 36518 7524 36524
rect 7484 36174 7512 36518
rect 7472 36168 7524 36174
rect 7472 36110 7524 36116
rect 7564 36032 7616 36038
rect 7564 35974 7616 35980
rect 7392 35788 7512 35816
rect 7380 35692 7432 35698
rect 7380 35634 7432 35640
rect 7392 35154 7420 35634
rect 7380 35148 7432 35154
rect 7380 35090 7432 35096
rect 7484 35086 7512 35788
rect 7472 35080 7524 35086
rect 7472 35022 7524 35028
rect 7288 35012 7340 35018
rect 7288 34954 7340 34960
rect 7196 34944 7248 34950
rect 7196 34886 7248 34892
rect 7196 34672 7248 34678
rect 7010 34640 7066 34649
rect 6920 34604 6972 34610
rect 7196 34614 7248 34620
rect 7010 34575 7012 34584
rect 6920 34546 6972 34552
rect 7064 34575 7066 34584
rect 7012 34546 7064 34552
rect 6828 34196 6880 34202
rect 6828 34138 6880 34144
rect 6644 33992 6696 33998
rect 6644 33934 6696 33940
rect 6552 33924 6604 33930
rect 6552 33866 6604 33872
rect 6564 33697 6592 33866
rect 6550 33688 6606 33697
rect 6550 33623 6606 33632
rect 6656 33561 6684 33934
rect 6736 33924 6788 33930
rect 6736 33866 6788 33872
rect 6920 33924 6972 33930
rect 6920 33866 6972 33872
rect 6642 33552 6698 33561
rect 6642 33487 6698 33496
rect 6552 33448 6604 33454
rect 6552 33390 6604 33396
rect 6564 33318 6592 33390
rect 6552 33312 6604 33318
rect 6552 33254 6604 33260
rect 6642 33144 6698 33153
rect 6642 33079 6698 33088
rect 6460 33040 6512 33046
rect 6460 32982 6512 32988
rect 6368 32904 6420 32910
rect 6368 32846 6420 32852
rect 6460 32904 6512 32910
rect 6460 32846 6512 32852
rect 6380 32609 6408 32846
rect 6366 32600 6422 32609
rect 6366 32535 6422 32544
rect 6288 32422 6408 32450
rect 6380 32366 6408 32422
rect 6368 32360 6420 32366
rect 6368 32302 6420 32308
rect 6274 32192 6330 32201
rect 6274 32127 6330 32136
rect 6090 31719 6146 31728
rect 6184 31748 6236 31754
rect 6184 31690 6236 31696
rect 6288 31634 6316 32127
rect 6368 32020 6420 32026
rect 6368 31962 6420 31968
rect 6380 31822 6408 31962
rect 6368 31816 6420 31822
rect 6368 31758 6420 31764
rect 6472 31634 6500 32846
rect 6550 32600 6606 32609
rect 6550 32535 6606 32544
rect 6564 31822 6592 32535
rect 6656 31822 6684 33079
rect 6748 32910 6776 33866
rect 6828 33312 6880 33318
rect 6828 33254 6880 33260
rect 6736 32904 6788 32910
rect 6736 32846 6788 32852
rect 6736 32428 6788 32434
rect 6736 32370 6788 32376
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6644 31816 6696 31822
rect 6644 31758 6696 31764
rect 6748 31686 6776 32370
rect 6644 31680 6696 31686
rect 6288 31606 6408 31634
rect 6472 31606 6592 31634
rect 6644 31622 6696 31628
rect 6736 31680 6788 31686
rect 6736 31622 6788 31628
rect 6274 31512 6330 31521
rect 6274 31447 6330 31456
rect 6000 30932 6052 30938
rect 6000 30874 6052 30880
rect 6012 30394 6040 30874
rect 6000 30388 6052 30394
rect 6000 30330 6052 30336
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 6288 28665 6316 31447
rect 6274 28656 6330 28665
rect 6274 28591 6330 28600
rect 6380 27305 6408 31606
rect 6564 29209 6592 31606
rect 6656 30734 6684 31622
rect 6736 31340 6788 31346
rect 6736 31282 6788 31288
rect 6644 30728 6696 30734
rect 6644 30670 6696 30676
rect 6644 30048 6696 30054
rect 6644 29990 6696 29996
rect 6656 29617 6684 29990
rect 6642 29608 6698 29617
rect 6642 29543 6698 29552
rect 6550 29200 6606 29209
rect 6550 29135 6606 29144
rect 6748 27849 6776 31282
rect 6840 28937 6868 33254
rect 6932 33017 6960 33866
rect 6918 33008 6974 33017
rect 6918 32943 6974 32952
rect 6920 32836 6972 32842
rect 6920 32778 6972 32784
rect 6932 32434 6960 32778
rect 6920 32428 6972 32434
rect 6920 32370 6972 32376
rect 7024 32366 7052 34546
rect 7208 34542 7236 34614
rect 7196 34536 7248 34542
rect 7196 34478 7248 34484
rect 7104 34400 7156 34406
rect 7104 34342 7156 34348
rect 7116 33930 7144 34342
rect 7104 33924 7156 33930
rect 7104 33866 7156 33872
rect 7102 33552 7158 33561
rect 7102 33487 7104 33496
rect 7156 33487 7158 33496
rect 7104 33458 7156 33464
rect 7208 32910 7236 34478
rect 7300 33998 7328 34954
rect 7380 34468 7432 34474
rect 7380 34410 7432 34416
rect 7288 33992 7340 33998
rect 7286 33960 7288 33969
rect 7340 33960 7342 33969
rect 7286 33895 7342 33904
rect 7392 33504 7420 34410
rect 7484 33998 7512 35022
rect 7576 34474 7604 35974
rect 7668 35630 7696 36654
rect 7760 36378 7788 38354
rect 8114 37632 8170 37641
rect 8114 37567 8170 37576
rect 7840 36644 7892 36650
rect 7840 36586 7892 36592
rect 7852 36378 7880 36586
rect 7748 36372 7800 36378
rect 7748 36314 7800 36320
rect 7840 36372 7892 36378
rect 7840 36314 7892 36320
rect 8128 36106 8156 37567
rect 8220 37262 8248 39086
rect 8758 38856 8814 38865
rect 8758 38791 8814 38800
rect 8666 38448 8722 38457
rect 8666 38383 8722 38392
rect 8576 37392 8628 37398
rect 8576 37334 8628 37340
rect 8208 37256 8260 37262
rect 8208 37198 8260 37204
rect 8484 37188 8536 37194
rect 8484 37130 8536 37136
rect 8390 36544 8446 36553
rect 8390 36479 8446 36488
rect 8116 36100 8168 36106
rect 8116 36042 8168 36048
rect 8300 36100 8352 36106
rect 8300 36042 8352 36048
rect 8116 35692 8168 35698
rect 8116 35634 8168 35640
rect 7656 35624 7708 35630
rect 7656 35566 7708 35572
rect 7564 34468 7616 34474
rect 7564 34410 7616 34416
rect 7564 34196 7616 34202
rect 7564 34138 7616 34144
rect 7472 33992 7524 33998
rect 7472 33934 7524 33940
rect 7484 33862 7512 33934
rect 7472 33856 7524 33862
rect 7472 33798 7524 33804
rect 7300 33476 7420 33504
rect 7300 33386 7328 33476
rect 7576 33425 7604 34138
rect 7668 33454 7696 35566
rect 7932 35556 7984 35562
rect 7932 35498 7984 35504
rect 7838 35456 7894 35465
rect 7838 35391 7894 35400
rect 7852 35086 7880 35391
rect 7840 35080 7892 35086
rect 7840 35022 7892 35028
rect 7748 35012 7800 35018
rect 7748 34954 7800 34960
rect 7760 34785 7788 34954
rect 7746 34776 7802 34785
rect 7746 34711 7802 34720
rect 7838 34640 7894 34649
rect 7838 34575 7840 34584
rect 7892 34575 7894 34584
rect 7840 34546 7892 34552
rect 7746 34232 7802 34241
rect 7746 34167 7802 34176
rect 7760 33862 7788 34167
rect 7944 34134 7972 35498
rect 8024 35216 8076 35222
rect 8024 35158 8076 35164
rect 8036 34610 8064 35158
rect 8024 34604 8076 34610
rect 8024 34546 8076 34552
rect 7932 34128 7984 34134
rect 7932 34070 7984 34076
rect 8024 34128 8076 34134
rect 8024 34070 8076 34076
rect 7840 33992 7892 33998
rect 7840 33934 7892 33940
rect 7748 33856 7800 33862
rect 7748 33798 7800 33804
rect 7748 33584 7800 33590
rect 7748 33526 7800 33532
rect 7656 33448 7708 33454
rect 7562 33416 7618 33425
rect 7288 33380 7340 33386
rect 7288 33322 7340 33328
rect 7380 33380 7432 33386
rect 7656 33390 7708 33396
rect 7562 33351 7618 33360
rect 7380 33322 7432 33328
rect 7196 32904 7248 32910
rect 7196 32846 7248 32852
rect 7104 32496 7156 32502
rect 7104 32438 7156 32444
rect 7012 32360 7064 32366
rect 7012 32302 7064 32308
rect 7116 32298 7144 32438
rect 7392 32366 7420 33322
rect 7380 32360 7432 32366
rect 7380 32302 7432 32308
rect 7104 32292 7156 32298
rect 7104 32234 7156 32240
rect 7012 32020 7064 32026
rect 7012 31962 7064 31968
rect 6920 30728 6972 30734
rect 6920 30670 6972 30676
rect 6932 29345 6960 30670
rect 7024 29646 7052 31962
rect 7116 30977 7144 32234
rect 7196 31340 7248 31346
rect 7196 31282 7248 31288
rect 7102 30968 7158 30977
rect 7102 30903 7158 30912
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 7116 29646 7144 30738
rect 7208 29714 7236 31282
rect 7288 30728 7340 30734
rect 7392 30716 7420 32302
rect 7564 31748 7616 31754
rect 7564 31690 7616 31696
rect 7656 31748 7708 31754
rect 7656 31690 7708 31696
rect 7340 30688 7420 30716
rect 7288 30670 7340 30676
rect 7392 30190 7420 30688
rect 7472 30592 7524 30598
rect 7472 30534 7524 30540
rect 7380 30184 7432 30190
rect 7380 30126 7432 30132
rect 7196 29708 7248 29714
rect 7196 29650 7248 29656
rect 7012 29640 7064 29646
rect 7012 29582 7064 29588
rect 7104 29640 7156 29646
rect 7104 29582 7156 29588
rect 6918 29336 6974 29345
rect 6918 29271 6974 29280
rect 7392 29238 7420 30126
rect 7484 29306 7512 30534
rect 7576 30161 7604 31690
rect 7668 31346 7696 31690
rect 7656 31340 7708 31346
rect 7656 31282 7708 31288
rect 7760 31278 7788 33526
rect 7852 33114 7880 33934
rect 7944 33862 7972 34070
rect 7932 33856 7984 33862
rect 7932 33798 7984 33804
rect 7840 33108 7892 33114
rect 7840 33050 7892 33056
rect 8036 33046 8064 34070
rect 8024 33040 8076 33046
rect 8024 32982 8076 32988
rect 7840 32904 7892 32910
rect 7840 32846 7892 32852
rect 7852 32201 7880 32846
rect 7932 32836 7984 32842
rect 7932 32778 7984 32784
rect 7838 32192 7894 32201
rect 7838 32127 7894 32136
rect 7852 31414 7880 32127
rect 7944 31890 7972 32778
rect 7932 31884 7984 31890
rect 7932 31826 7984 31832
rect 8036 31822 8064 32982
rect 8128 32473 8156 35634
rect 8208 35080 8260 35086
rect 8208 35022 8260 35028
rect 8220 34649 8248 35022
rect 8206 34640 8262 34649
rect 8206 34575 8262 34584
rect 8312 34490 8340 36042
rect 8404 35086 8432 36479
rect 8496 36106 8524 37130
rect 8588 36310 8616 37334
rect 8576 36304 8628 36310
rect 8576 36246 8628 36252
rect 8484 36100 8536 36106
rect 8484 36042 8536 36048
rect 8680 35290 8708 38383
rect 8668 35284 8720 35290
rect 8668 35226 8720 35232
rect 8392 35080 8444 35086
rect 8392 35022 8444 35028
rect 8220 34462 8340 34490
rect 8576 34468 8628 34474
rect 8220 34202 8248 34462
rect 8576 34410 8628 34416
rect 8588 34202 8616 34410
rect 8208 34196 8260 34202
rect 8208 34138 8260 34144
rect 8576 34196 8628 34202
rect 8576 34138 8628 34144
rect 8392 33992 8444 33998
rect 8392 33934 8444 33940
rect 8404 32994 8432 33934
rect 8482 33688 8538 33697
rect 8482 33623 8538 33632
rect 8576 33652 8628 33658
rect 8496 33046 8524 33623
rect 8576 33594 8628 33600
rect 8588 33318 8616 33594
rect 8772 33522 8800 38791
rect 9496 37324 9548 37330
rect 9496 37266 9548 37272
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 9140 36786 9168 37062
rect 9128 36780 9180 36786
rect 9128 36722 9180 36728
rect 9220 36644 9272 36650
rect 9220 36586 9272 36592
rect 9232 36242 9260 36586
rect 9220 36236 9272 36242
rect 9220 36178 9272 36184
rect 9402 35864 9458 35873
rect 9402 35799 9458 35808
rect 9128 35692 9180 35698
rect 9128 35634 9180 35640
rect 9140 35290 9168 35634
rect 9128 35284 9180 35290
rect 9128 35226 9180 35232
rect 9416 34950 9444 35799
rect 9508 35086 9536 37266
rect 10520 37262 10548 39102
rect 11704 39102 11756 39108
rect 11242 39063 11298 39072
rect 11058 38176 11114 38185
rect 11058 38111 11114 38120
rect 11072 37466 11100 38111
rect 11060 37460 11112 37466
rect 11060 37402 11112 37408
rect 10968 37324 11020 37330
rect 10968 37266 11020 37272
rect 10508 37256 10560 37262
rect 10508 37198 10560 37204
rect 9680 37188 9732 37194
rect 9680 37130 9732 37136
rect 9772 37188 9824 37194
rect 9772 37130 9824 37136
rect 9588 37120 9640 37126
rect 9588 37062 9640 37068
rect 9600 36922 9628 37062
rect 9588 36916 9640 36922
rect 9588 36858 9640 36864
rect 9600 36242 9628 36858
rect 9588 36236 9640 36242
rect 9588 36178 9640 36184
rect 9692 36038 9720 37130
rect 9784 36650 9812 37130
rect 10508 36780 10560 36786
rect 10508 36722 10560 36728
rect 9772 36644 9824 36650
rect 9772 36586 9824 36592
rect 10520 36378 10548 36722
rect 9864 36372 9916 36378
rect 9864 36314 9916 36320
rect 10508 36372 10560 36378
rect 10508 36314 10560 36320
rect 9876 36242 9904 36314
rect 10416 36304 10468 36310
rect 10416 36246 10468 36252
rect 9864 36236 9916 36242
rect 9864 36178 9916 36184
rect 9680 36032 9732 36038
rect 9678 36000 9680 36009
rect 9732 36000 9734 36009
rect 9678 35935 9734 35944
rect 9588 35828 9640 35834
rect 9588 35770 9640 35776
rect 9600 35154 9628 35770
rect 9772 35760 9824 35766
rect 9772 35702 9824 35708
rect 9588 35148 9640 35154
rect 9588 35090 9640 35096
rect 9784 35086 9812 35702
rect 9876 35630 9904 36178
rect 10230 35864 10286 35873
rect 10230 35799 10286 35808
rect 10244 35766 10272 35799
rect 10232 35760 10284 35766
rect 10232 35702 10284 35708
rect 9864 35624 9916 35630
rect 9864 35566 9916 35572
rect 10048 35148 10100 35154
rect 10048 35090 10100 35096
rect 9496 35080 9548 35086
rect 9496 35022 9548 35028
rect 9772 35080 9824 35086
rect 9772 35022 9824 35028
rect 9680 35012 9732 35018
rect 9680 34954 9732 34960
rect 9404 34944 9456 34950
rect 9588 34944 9640 34950
rect 9404 34886 9456 34892
rect 9508 34904 9588 34932
rect 9036 34604 9088 34610
rect 9036 34546 9088 34552
rect 9404 34604 9456 34610
rect 9404 34546 9456 34552
rect 8944 34060 8996 34066
rect 8944 34002 8996 34008
rect 8956 33590 8984 34002
rect 9048 33930 9076 34546
rect 9036 33924 9088 33930
rect 9036 33866 9088 33872
rect 8944 33584 8996 33590
rect 8944 33526 8996 33532
rect 8760 33516 8812 33522
rect 8760 33458 8812 33464
rect 8668 33448 8720 33454
rect 8668 33390 8720 33396
rect 8576 33312 8628 33318
rect 8576 33254 8628 33260
rect 8208 32972 8260 32978
rect 8208 32914 8260 32920
rect 8312 32966 8432 32994
rect 8484 33040 8536 33046
rect 8484 32982 8536 32988
rect 8588 32978 8616 33254
rect 8680 32978 8708 33390
rect 8576 32972 8628 32978
rect 8114 32464 8170 32473
rect 8114 32399 8170 32408
rect 8220 31929 8248 32914
rect 8312 32434 8340 32966
rect 8576 32914 8628 32920
rect 8668 32972 8720 32978
rect 8668 32914 8720 32920
rect 8484 32904 8536 32910
rect 8484 32846 8536 32852
rect 8852 32904 8904 32910
rect 8852 32846 8904 32852
rect 8496 32570 8524 32846
rect 8484 32564 8536 32570
rect 8484 32506 8536 32512
rect 8300 32428 8352 32434
rect 8300 32370 8352 32376
rect 8206 31920 8262 31929
rect 8206 31855 8262 31864
rect 8312 31822 8340 32370
rect 8760 32360 8812 32366
rect 8760 32302 8812 32308
rect 8772 32230 8800 32302
rect 8576 32224 8628 32230
rect 8576 32166 8628 32172
rect 8760 32224 8812 32230
rect 8760 32166 8812 32172
rect 8588 32042 8616 32166
rect 8496 32026 8616 32042
rect 8484 32020 8616 32026
rect 8536 32014 8616 32020
rect 8484 31962 8536 31968
rect 8772 31906 8800 32166
rect 8864 32008 8892 32846
rect 9048 32745 9076 33866
rect 9220 32972 9272 32978
rect 9220 32914 9272 32920
rect 9128 32768 9180 32774
rect 9034 32736 9090 32745
rect 9128 32710 9180 32716
rect 9034 32671 9090 32680
rect 8942 32600 8998 32609
rect 8942 32535 8998 32544
rect 8956 32230 8984 32535
rect 9140 32502 9168 32710
rect 9128 32496 9180 32502
rect 9128 32438 9180 32444
rect 9036 32428 9088 32434
rect 9036 32370 9088 32376
rect 9048 32230 9076 32370
rect 8944 32224 8996 32230
rect 8944 32166 8996 32172
rect 9036 32224 9088 32230
rect 9036 32166 9088 32172
rect 8864 31980 8984 32008
rect 8772 31878 8892 31906
rect 8024 31816 8076 31822
rect 8024 31758 8076 31764
rect 8300 31816 8352 31822
rect 8576 31816 8628 31822
rect 8352 31776 8524 31804
rect 8300 31758 8352 31764
rect 7932 31680 7984 31686
rect 7932 31622 7984 31628
rect 7840 31408 7892 31414
rect 7840 31350 7892 31356
rect 7944 31346 7972 31622
rect 8036 31346 8064 31758
rect 8208 31680 8260 31686
rect 8128 31640 8208 31668
rect 7932 31340 7984 31346
rect 7932 31282 7984 31288
rect 8024 31340 8076 31346
rect 8024 31282 8076 31288
rect 7748 31272 7800 31278
rect 7748 31214 7800 31220
rect 7656 31204 7708 31210
rect 7656 31146 7708 31152
rect 7840 31204 7892 31210
rect 7840 31146 7892 31152
rect 7562 30152 7618 30161
rect 7562 30087 7618 30096
rect 7564 29708 7616 29714
rect 7564 29650 7616 29656
rect 7472 29300 7524 29306
rect 7472 29242 7524 29248
rect 7380 29232 7432 29238
rect 7380 29174 7432 29180
rect 7576 29170 7604 29650
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 7012 29028 7064 29034
rect 7012 28970 7064 28976
rect 6826 28928 6882 28937
rect 6826 28863 6882 28872
rect 6734 27840 6790 27849
rect 6734 27775 6790 27784
rect 6920 27668 6972 27674
rect 6920 27610 6972 27616
rect 6366 27296 6422 27305
rect 6366 27231 6422 27240
rect 5446 26072 5502 26081
rect 5446 26007 5502 26016
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5172 21412 5224 21418
rect 5172 21354 5224 21360
rect 6932 21350 6960 27610
rect 7024 23225 7052 28970
rect 7196 28960 7248 28966
rect 7196 28902 7248 28908
rect 7104 28552 7156 28558
rect 7104 28494 7156 28500
rect 7116 27538 7144 28494
rect 7104 27532 7156 27538
rect 7104 27474 7156 27480
rect 7208 23322 7236 28902
rect 7576 27946 7604 29106
rect 7564 27940 7616 27946
rect 7564 27882 7616 27888
rect 7668 27713 7696 31146
rect 7748 30048 7800 30054
rect 7748 29990 7800 29996
rect 7760 29889 7788 29990
rect 7746 29880 7802 29889
rect 7746 29815 7802 29824
rect 7852 28966 7880 31146
rect 7944 30036 7972 31282
rect 8036 30326 8064 31282
rect 8128 30841 8156 31640
rect 8208 31622 8260 31628
rect 8390 31512 8446 31521
rect 8390 31447 8446 31456
rect 8300 31136 8352 31142
rect 8300 31078 8352 31084
rect 8208 30932 8260 30938
rect 8208 30874 8260 30880
rect 8114 30832 8170 30841
rect 8114 30767 8170 30776
rect 8024 30320 8076 30326
rect 8024 30262 8076 30268
rect 8116 30252 8168 30258
rect 8116 30194 8168 30200
rect 8024 30048 8076 30054
rect 7944 30008 8024 30036
rect 8024 29990 8076 29996
rect 8128 29850 8156 30194
rect 8220 29850 8248 30874
rect 8116 29844 8168 29850
rect 8116 29786 8168 29792
rect 8208 29844 8260 29850
rect 8208 29786 8260 29792
rect 7930 29744 7986 29753
rect 7930 29679 7986 29688
rect 7944 29170 7972 29679
rect 8312 29646 8340 31078
rect 8404 30598 8432 31447
rect 8496 30802 8524 31776
rect 8576 31758 8628 31764
rect 8484 30796 8536 30802
rect 8484 30738 8536 30744
rect 8484 30660 8536 30666
rect 8484 30602 8536 30608
rect 8392 30592 8444 30598
rect 8392 30534 8444 30540
rect 8496 30326 8524 30602
rect 8484 30320 8536 30326
rect 8484 30262 8536 30268
rect 8588 30190 8616 31758
rect 8668 31748 8720 31754
rect 8668 31690 8720 31696
rect 8576 30184 8628 30190
rect 8576 30126 8628 30132
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 8208 29504 8260 29510
rect 8208 29446 8260 29452
rect 8114 29336 8170 29345
rect 8114 29271 8116 29280
rect 8168 29271 8170 29280
rect 8116 29242 8168 29248
rect 8220 29170 8248 29446
rect 8392 29300 8444 29306
rect 8392 29242 8444 29248
rect 7932 29164 7984 29170
rect 7932 29106 7984 29112
rect 8208 29164 8260 29170
rect 8208 29106 8260 29112
rect 8220 28994 8248 29106
rect 8404 29102 8432 29242
rect 8392 29096 8444 29102
rect 8392 29038 8444 29044
rect 8220 28966 8432 28994
rect 7840 28960 7892 28966
rect 8404 28914 8432 28966
rect 7840 28902 7892 28908
rect 8312 28886 8432 28914
rect 8024 28484 8076 28490
rect 8024 28426 8076 28432
rect 8036 28218 8064 28426
rect 8024 28212 8076 28218
rect 8024 28154 8076 28160
rect 8312 28150 8340 28886
rect 8392 28416 8444 28422
rect 8392 28358 8444 28364
rect 8300 28144 8352 28150
rect 8300 28086 8352 28092
rect 8404 28082 8432 28358
rect 8392 28076 8444 28082
rect 8392 28018 8444 28024
rect 7654 27704 7710 27713
rect 7654 27639 7710 27648
rect 8208 27464 8260 27470
rect 8208 27406 8260 27412
rect 8024 27396 8076 27402
rect 8024 27338 8076 27344
rect 8036 27130 8064 27338
rect 8024 27124 8076 27130
rect 8024 27066 8076 27072
rect 8220 26450 8248 27406
rect 8208 26444 8260 26450
rect 8208 26386 8260 26392
rect 8220 25922 8248 26386
rect 8220 25906 8340 25922
rect 8220 25900 8352 25906
rect 8220 25894 8300 25900
rect 8300 25842 8352 25848
rect 8208 24744 8260 24750
rect 8208 24686 8260 24692
rect 8220 24206 8248 24686
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8220 23730 8248 24142
rect 8208 23724 8260 23730
rect 8208 23666 8260 23672
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7010 23216 7066 23225
rect 7010 23151 7066 23160
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 8404 19145 8432 28018
rect 8496 28014 8524 29582
rect 8484 28008 8536 28014
rect 8484 27950 8536 27956
rect 8588 27470 8616 30126
rect 8680 29510 8708 31690
rect 8760 31272 8812 31278
rect 8760 31214 8812 31220
rect 8772 30666 8800 31214
rect 8760 30660 8812 30666
rect 8760 30602 8812 30608
rect 8760 30048 8812 30054
rect 8758 30016 8760 30025
rect 8812 30016 8814 30025
rect 8758 29951 8814 29960
rect 8772 29714 8800 29951
rect 8760 29708 8812 29714
rect 8760 29650 8812 29656
rect 8668 29504 8720 29510
rect 8668 29446 8720 29452
rect 8758 29472 8814 29481
rect 8758 29407 8814 29416
rect 8772 29170 8800 29407
rect 8864 29170 8892 31878
rect 8956 31414 8984 31980
rect 9232 31822 9260 32914
rect 9312 32768 9364 32774
rect 9312 32710 9364 32716
rect 9220 31816 9272 31822
rect 9220 31758 9272 31764
rect 9036 31680 9088 31686
rect 9036 31622 9088 31628
rect 8944 31408 8996 31414
rect 8944 31350 8996 31356
rect 8956 31210 8984 31350
rect 8944 31204 8996 31210
rect 8944 31146 8996 31152
rect 9048 31142 9076 31622
rect 9220 31408 9272 31414
rect 9220 31350 9272 31356
rect 9036 31136 9088 31142
rect 9036 31078 9088 31084
rect 9128 31136 9180 31142
rect 9128 31078 9180 31084
rect 9036 30864 9088 30870
rect 9036 30806 9088 30812
rect 8944 30796 8996 30802
rect 8944 30738 8996 30744
rect 8956 30258 8984 30738
rect 8944 30252 8996 30258
rect 8944 30194 8996 30200
rect 8760 29164 8812 29170
rect 8760 29106 8812 29112
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 8668 29028 8720 29034
rect 8668 28970 8720 28976
rect 8576 27464 8628 27470
rect 8680 27441 8708 28970
rect 8772 27577 8800 29106
rect 8956 29034 8984 30194
rect 9048 29753 9076 30806
rect 9140 30326 9168 31078
rect 9232 30326 9260 31350
rect 9324 31278 9352 32710
rect 9416 32366 9444 34546
rect 9508 34474 9536 34904
rect 9588 34886 9640 34892
rect 9692 34649 9720 34954
rect 9678 34640 9734 34649
rect 9678 34575 9734 34584
rect 9784 34542 9812 35022
rect 10060 34610 10088 35090
rect 10428 35086 10456 36246
rect 10980 36242 11008 37266
rect 11152 36576 11204 36582
rect 11152 36518 11204 36524
rect 10968 36236 11020 36242
rect 10968 36178 11020 36184
rect 11164 36038 11192 36518
rect 11152 36032 11204 36038
rect 11152 35974 11204 35980
rect 11152 35148 11204 35154
rect 11152 35090 11204 35096
rect 10324 35080 10376 35086
rect 10322 35048 10324 35057
rect 10416 35080 10468 35086
rect 10376 35048 10378 35057
rect 10416 35022 10468 35028
rect 10322 34983 10378 34992
rect 10048 34604 10100 34610
rect 9876 34564 10048 34592
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 9496 34468 9548 34474
rect 9496 34410 9548 34416
rect 9588 34400 9640 34406
rect 9588 34342 9640 34348
rect 9496 33516 9548 33522
rect 9496 33458 9548 33464
rect 9508 32910 9536 33458
rect 9600 32994 9628 34342
rect 9680 34196 9732 34202
rect 9680 34138 9732 34144
rect 9692 34066 9720 34138
rect 9680 34060 9732 34066
rect 9680 34002 9732 34008
rect 9772 33992 9824 33998
rect 9772 33934 9824 33940
rect 9600 32978 9720 32994
rect 9600 32972 9732 32978
rect 9600 32966 9680 32972
rect 9680 32914 9732 32920
rect 9496 32904 9548 32910
rect 9496 32846 9548 32852
rect 9588 32904 9640 32910
rect 9784 32881 9812 33934
rect 9876 33454 9904 34564
rect 10048 34546 10100 34552
rect 10324 34604 10376 34610
rect 10324 34546 10376 34552
rect 10140 34400 10192 34406
rect 10140 34342 10192 34348
rect 9954 33688 10010 33697
rect 9954 33623 9956 33632
rect 10008 33623 10010 33632
rect 9956 33594 10008 33600
rect 9864 33448 9916 33454
rect 9864 33390 9916 33396
rect 9968 33386 9996 33594
rect 10048 33448 10100 33454
rect 10048 33390 10100 33396
rect 9956 33380 10008 33386
rect 9956 33322 10008 33328
rect 10060 33114 10088 33390
rect 10152 33318 10180 34342
rect 10336 33998 10364 34546
rect 10782 34504 10838 34513
rect 10782 34439 10838 34448
rect 10876 34468 10928 34474
rect 10324 33992 10376 33998
rect 10324 33934 10376 33940
rect 10692 33448 10744 33454
rect 10692 33390 10744 33396
rect 10140 33312 10192 33318
rect 10140 33254 10192 33260
rect 10048 33108 10100 33114
rect 10048 33050 10100 33056
rect 10152 32994 10180 33254
rect 10060 32966 10180 32994
rect 10414 33008 10470 33017
rect 9588 32846 9640 32852
rect 9770 32872 9826 32881
rect 9494 32736 9550 32745
rect 9494 32671 9550 32680
rect 9404 32360 9456 32366
rect 9404 32302 9456 32308
rect 9402 32192 9458 32201
rect 9402 32127 9458 32136
rect 9416 32026 9444 32127
rect 9404 32020 9456 32026
rect 9404 31962 9456 31968
rect 9508 31890 9536 32671
rect 9600 31958 9628 32846
rect 9770 32807 9826 32816
rect 9956 32428 10008 32434
rect 9956 32370 10008 32376
rect 9770 32328 9826 32337
rect 9692 32298 9770 32314
rect 9680 32292 9770 32298
rect 9732 32286 9770 32292
rect 9770 32263 9826 32272
rect 9680 32234 9732 32240
rect 9588 31952 9640 31958
rect 9588 31894 9640 31900
rect 9404 31884 9456 31890
rect 9404 31826 9456 31832
rect 9496 31884 9548 31890
rect 9496 31826 9548 31832
rect 9416 31521 9444 31826
rect 9402 31512 9458 31521
rect 9402 31447 9458 31456
rect 9508 31414 9536 31826
rect 9496 31408 9548 31414
rect 9496 31350 9548 31356
rect 9404 31340 9456 31346
rect 9404 31282 9456 31288
rect 9312 31272 9364 31278
rect 9312 31214 9364 31220
rect 9128 30320 9180 30326
rect 9128 30262 9180 30268
rect 9220 30320 9272 30326
rect 9220 30262 9272 30268
rect 9128 30048 9180 30054
rect 9128 29990 9180 29996
rect 9034 29744 9090 29753
rect 9140 29714 9168 29990
rect 9034 29679 9090 29688
rect 9128 29708 9180 29714
rect 9128 29650 9180 29656
rect 9324 29646 9352 31214
rect 9416 29866 9444 31282
rect 9586 30968 9642 30977
rect 9586 30903 9642 30912
rect 9494 30832 9550 30841
rect 9494 30767 9550 30776
rect 9508 30734 9536 30767
rect 9496 30728 9548 30734
rect 9496 30670 9548 30676
rect 9600 30666 9628 30903
rect 9692 30802 9720 32234
rect 9772 32224 9824 32230
rect 9772 32166 9824 32172
rect 9864 32224 9916 32230
rect 9864 32166 9916 32172
rect 9784 31958 9812 32166
rect 9772 31952 9824 31958
rect 9772 31894 9824 31900
rect 9772 31816 9824 31822
rect 9772 31758 9824 31764
rect 9784 31210 9812 31758
rect 9876 31278 9904 32166
rect 9968 31385 9996 32370
rect 9954 31376 10010 31385
rect 9954 31311 10010 31320
rect 9864 31272 9916 31278
rect 9864 31214 9916 31220
rect 9772 31204 9824 31210
rect 9772 31146 9824 31152
rect 9956 31136 10008 31142
rect 9956 31078 10008 31084
rect 9770 30832 9826 30841
rect 9680 30796 9732 30802
rect 9770 30767 9826 30776
rect 9680 30738 9732 30744
rect 9588 30660 9640 30666
rect 9588 30602 9640 30608
rect 9496 30592 9548 30598
rect 9496 30534 9548 30540
rect 9508 30054 9536 30534
rect 9678 30288 9734 30297
rect 9784 30258 9812 30767
rect 9678 30223 9734 30232
rect 9772 30252 9824 30258
rect 9692 30054 9720 30223
rect 9772 30194 9824 30200
rect 9496 30048 9548 30054
rect 9496 29990 9548 29996
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9416 29838 9628 29866
rect 9404 29776 9456 29782
rect 9404 29718 9456 29724
rect 9496 29776 9548 29782
rect 9496 29718 9548 29724
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9416 29481 9444 29718
rect 9402 29472 9458 29481
rect 9402 29407 9458 29416
rect 9416 29102 9444 29407
rect 9220 29096 9272 29102
rect 9218 29064 9220 29073
rect 9404 29096 9456 29102
rect 9272 29064 9274 29073
rect 8852 29028 8904 29034
rect 8852 28970 8904 28976
rect 8944 29028 8996 29034
rect 9404 29038 9456 29044
rect 9218 28999 9274 29008
rect 8944 28970 8996 28976
rect 8758 27568 8814 27577
rect 8758 27503 8814 27512
rect 8576 27406 8628 27412
rect 8666 27432 8722 27441
rect 8666 27367 8722 27376
rect 8576 27328 8628 27334
rect 8576 27270 8628 27276
rect 8588 27062 8616 27270
rect 8576 27056 8628 27062
rect 8576 26998 8628 27004
rect 8864 25294 8892 28970
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 9128 28416 9180 28422
rect 9128 28358 9180 28364
rect 9140 28218 9168 28358
rect 9128 28212 9180 28218
rect 9128 28154 9180 28160
rect 9324 27674 9352 28494
rect 9312 27668 9364 27674
rect 9312 27610 9364 27616
rect 9324 27130 9352 27610
rect 9312 27124 9364 27130
rect 9312 27066 9364 27072
rect 9508 25362 9536 29718
rect 9600 29714 9628 29838
rect 9588 29708 9640 29714
rect 9588 29650 9640 29656
rect 9692 29560 9720 29990
rect 9600 29532 9720 29560
rect 9600 29306 9628 29532
rect 9772 29504 9824 29510
rect 9772 29446 9824 29452
rect 9588 29300 9640 29306
rect 9588 29242 9640 29248
rect 9680 29300 9732 29306
rect 9680 29242 9732 29248
rect 9588 29096 9640 29102
rect 9588 29038 9640 29044
rect 9600 28914 9628 29038
rect 9692 29034 9720 29242
rect 9784 29170 9812 29446
rect 9772 29164 9824 29170
rect 9772 29106 9824 29112
rect 9680 29028 9732 29034
rect 9680 28970 9732 28976
rect 9600 28886 9720 28914
rect 9588 27872 9640 27878
rect 9588 27814 9640 27820
rect 9600 26994 9628 27814
rect 9692 27470 9720 28886
rect 9784 28626 9812 29106
rect 9864 28960 9916 28966
rect 9864 28902 9916 28908
rect 9772 28620 9824 28626
rect 9772 28562 9824 28568
rect 9876 28558 9904 28902
rect 9864 28552 9916 28558
rect 9864 28494 9916 28500
rect 9772 28484 9824 28490
rect 9772 28426 9824 28432
rect 9784 27946 9812 28426
rect 9968 28064 9996 31078
rect 10060 29753 10088 32966
rect 10414 32943 10470 32952
rect 10428 32910 10456 32943
rect 10704 32910 10732 33390
rect 10416 32904 10468 32910
rect 10336 32864 10416 32892
rect 10140 32428 10192 32434
rect 10140 32370 10192 32376
rect 10152 32026 10180 32370
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 10152 31890 10180 31962
rect 10140 31884 10192 31890
rect 10140 31826 10192 31832
rect 10336 31521 10364 32864
rect 10692 32904 10744 32910
rect 10416 32846 10468 32852
rect 10690 32872 10692 32881
rect 10744 32872 10746 32881
rect 10690 32807 10746 32816
rect 10416 32768 10468 32774
rect 10416 32710 10468 32716
rect 10428 31929 10456 32710
rect 10796 32484 10824 34439
rect 10876 34410 10928 34416
rect 10888 33998 10916 34410
rect 11058 34232 11114 34241
rect 11058 34167 11114 34176
rect 10876 33992 10928 33998
rect 10876 33934 10928 33940
rect 10888 32745 10916 33934
rect 11072 33590 11100 34167
rect 11164 33998 11192 35090
rect 11152 33992 11204 33998
rect 11152 33934 11204 33940
rect 11060 33584 11112 33590
rect 11060 33526 11112 33532
rect 10968 33516 11020 33522
rect 10968 33458 11020 33464
rect 10980 33114 11008 33458
rect 11072 33130 11100 33526
rect 11164 33289 11192 33934
rect 11150 33280 11206 33289
rect 11150 33215 11206 33224
rect 10968 33108 11020 33114
rect 11072 33102 11192 33130
rect 10968 33050 11020 33056
rect 10874 32736 10930 32745
rect 10874 32671 10930 32680
rect 10796 32456 10916 32484
rect 10508 32360 10560 32366
rect 10560 32320 10640 32348
rect 10508 32302 10560 32308
rect 10414 31920 10470 31929
rect 10414 31855 10470 31864
rect 10428 31822 10456 31855
rect 10416 31816 10468 31822
rect 10416 31758 10468 31764
rect 10508 31816 10560 31822
rect 10508 31758 10560 31764
rect 10322 31512 10378 31521
rect 10322 31447 10378 31456
rect 10416 31204 10468 31210
rect 10416 31146 10468 31152
rect 10140 30796 10192 30802
rect 10140 30738 10192 30744
rect 10046 29744 10102 29753
rect 10046 29679 10102 29688
rect 10060 28558 10088 29679
rect 10152 29646 10180 30738
rect 10232 30728 10284 30734
rect 10284 30676 10364 30682
rect 10232 30670 10364 30676
rect 10244 30654 10364 30670
rect 10232 30592 10284 30598
rect 10232 30534 10284 30540
rect 10244 29646 10272 30534
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 10232 29640 10284 29646
rect 10232 29582 10284 29588
rect 10336 29345 10364 30654
rect 10428 29850 10456 31146
rect 10520 30122 10548 31758
rect 10508 30116 10560 30122
rect 10508 30058 10560 30064
rect 10416 29844 10468 29850
rect 10416 29786 10468 29792
rect 10508 29708 10560 29714
rect 10508 29650 10560 29656
rect 10322 29336 10378 29345
rect 10322 29271 10378 29280
rect 10048 28552 10100 28558
rect 10048 28494 10100 28500
rect 10140 28212 10192 28218
rect 10140 28154 10192 28160
rect 10048 28076 10100 28082
rect 9968 28036 10048 28064
rect 10048 28018 10100 28024
rect 10152 28014 10180 28154
rect 10140 28008 10192 28014
rect 10140 27950 10192 27956
rect 9772 27940 9824 27946
rect 9772 27882 9824 27888
rect 10048 27940 10100 27946
rect 10048 27882 10100 27888
rect 10060 27674 10088 27882
rect 10152 27878 10180 27950
rect 10140 27872 10192 27878
rect 10140 27814 10192 27820
rect 10048 27668 10100 27674
rect 10048 27610 10100 27616
rect 9680 27464 9732 27470
rect 9680 27406 9732 27412
rect 9862 27024 9918 27033
rect 9588 26988 9640 26994
rect 9862 26959 9864 26968
rect 9588 26930 9640 26936
rect 9916 26959 9918 26968
rect 9864 26930 9916 26936
rect 9876 25770 9904 26930
rect 10140 26920 10192 26926
rect 9968 26868 10140 26874
rect 9968 26862 10192 26868
rect 9968 26858 10180 26862
rect 9956 26852 10180 26858
rect 10008 26846 10180 26852
rect 9956 26794 10008 26800
rect 10140 26784 10192 26790
rect 10140 26726 10192 26732
rect 10152 25974 10180 26726
rect 10140 25968 10192 25974
rect 10140 25910 10192 25916
rect 9864 25764 9916 25770
rect 9864 25706 9916 25712
rect 10140 25424 10192 25430
rect 10140 25366 10192 25372
rect 9496 25356 9548 25362
rect 9496 25298 9548 25304
rect 8852 25288 8904 25294
rect 8852 25230 8904 25236
rect 9128 25152 9180 25158
rect 9128 25094 9180 25100
rect 9496 25152 9548 25158
rect 9496 25094 9548 25100
rect 9140 24886 9168 25094
rect 9508 24954 9536 25094
rect 9496 24948 9548 24954
rect 9496 24890 9548 24896
rect 9128 24880 9180 24886
rect 9128 24822 9180 24828
rect 10152 24818 10180 25366
rect 10232 25152 10284 25158
rect 10232 25094 10284 25100
rect 10244 24818 10272 25094
rect 10336 24818 10364 29271
rect 10416 29164 10468 29170
rect 10416 29106 10468 29112
rect 10428 28966 10456 29106
rect 10520 29034 10548 29650
rect 10612 29170 10640 32320
rect 10782 32056 10838 32065
rect 10782 31991 10838 32000
rect 10796 31822 10824 31991
rect 10784 31816 10836 31822
rect 10784 31758 10836 31764
rect 10692 31680 10744 31686
rect 10692 31622 10744 31628
rect 10704 31414 10732 31622
rect 10692 31408 10744 31414
rect 10692 31350 10744 31356
rect 10704 29646 10732 31350
rect 10692 29640 10744 29646
rect 10692 29582 10744 29588
rect 10796 29170 10824 31758
rect 10888 31482 10916 32456
rect 11060 32224 11112 32230
rect 11060 32166 11112 32172
rect 11072 31498 11100 32166
rect 11164 31754 11192 33102
rect 11256 32434 11284 39063
rect 13728 38684 13780 38690
rect 13728 38626 13780 38632
rect 13740 38010 13768 38626
rect 13728 38004 13780 38010
rect 13728 37946 13780 37952
rect 12254 37496 12310 37505
rect 12254 37431 12310 37440
rect 11796 37120 11848 37126
rect 11796 37062 11848 37068
rect 11704 36848 11756 36854
rect 11704 36790 11756 36796
rect 11716 36718 11744 36790
rect 11704 36712 11756 36718
rect 11704 36654 11756 36660
rect 11716 36242 11744 36654
rect 11704 36236 11756 36242
rect 11704 36178 11756 36184
rect 11808 36174 11836 37062
rect 11980 36576 12032 36582
rect 11980 36518 12032 36524
rect 11796 36168 11848 36174
rect 11796 36110 11848 36116
rect 11704 36100 11756 36106
rect 11704 36042 11756 36048
rect 11716 35698 11744 36042
rect 11704 35692 11756 35698
rect 11704 35634 11756 35640
rect 11716 35601 11744 35634
rect 11702 35592 11758 35601
rect 11702 35527 11758 35536
rect 11612 34944 11664 34950
rect 11612 34886 11664 34892
rect 11520 33992 11572 33998
rect 11520 33934 11572 33940
rect 11428 32904 11480 32910
rect 11428 32846 11480 32852
rect 11244 32428 11296 32434
rect 11244 32370 11296 32376
rect 11336 32428 11388 32434
rect 11336 32370 11388 32376
rect 11256 32298 11284 32370
rect 11244 32292 11296 32298
rect 11244 32234 11296 32240
rect 11348 31890 11376 32370
rect 11336 31884 11388 31890
rect 11336 31826 11388 31832
rect 11440 31754 11468 32846
rect 11532 32178 11560 33934
rect 11624 32910 11652 34886
rect 11886 34776 11942 34785
rect 11992 34746 12020 36518
rect 12072 36032 12124 36038
rect 12072 35974 12124 35980
rect 12084 35698 12112 35974
rect 12072 35692 12124 35698
rect 12072 35634 12124 35640
rect 12164 35080 12216 35086
rect 12164 35022 12216 35028
rect 12176 34785 12204 35022
rect 12162 34776 12218 34785
rect 11886 34711 11942 34720
rect 11980 34740 12032 34746
rect 11702 33960 11758 33969
rect 11702 33895 11758 33904
rect 11716 33561 11744 33895
rect 11702 33552 11758 33561
rect 11900 33522 11928 34711
rect 12162 34711 12218 34720
rect 11980 34682 12032 34688
rect 11980 34604 12032 34610
rect 11980 34546 12032 34552
rect 12164 34604 12216 34610
rect 12164 34546 12216 34552
rect 11992 33969 12020 34546
rect 11978 33960 12034 33969
rect 11978 33895 12034 33904
rect 11888 33516 11940 33522
rect 11702 33487 11704 33496
rect 11756 33487 11758 33496
rect 11704 33458 11756 33464
rect 11808 33476 11888 33504
rect 11704 33312 11756 33318
rect 11704 33254 11756 33260
rect 11612 32904 11664 32910
rect 11612 32846 11664 32852
rect 11612 32224 11664 32230
rect 11532 32172 11612 32178
rect 11532 32166 11664 32172
rect 11532 32150 11652 32166
rect 11518 32056 11574 32065
rect 11518 31991 11574 32000
rect 11532 31822 11560 31991
rect 11624 31929 11652 32150
rect 11610 31920 11666 31929
rect 11610 31855 11666 31864
rect 11520 31816 11572 31822
rect 11520 31758 11572 31764
rect 11164 31726 11284 31754
rect 10876 31476 10928 31482
rect 10876 31418 10928 31424
rect 10968 31476 11020 31482
rect 11072 31470 11192 31498
rect 10968 31418 11020 31424
rect 10888 31346 10916 31418
rect 10876 31340 10928 31346
rect 10876 31282 10928 31288
rect 10876 31136 10928 31142
rect 10876 31078 10928 31084
rect 10888 30977 10916 31078
rect 10874 30968 10930 30977
rect 10874 30903 10930 30912
rect 10874 30560 10930 30569
rect 10874 30495 10930 30504
rect 10888 30054 10916 30495
rect 10980 30161 11008 31418
rect 11058 31376 11114 31385
rect 11058 31311 11060 31320
rect 11112 31311 11114 31320
rect 11060 31282 11112 31288
rect 11060 31204 11112 31210
rect 11060 31146 11112 31152
rect 11072 30938 11100 31146
rect 11060 30932 11112 30938
rect 11060 30874 11112 30880
rect 10966 30152 11022 30161
rect 10966 30087 11022 30096
rect 10980 30054 11008 30087
rect 10876 30048 10928 30054
rect 10876 29990 10928 29996
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 10876 29572 10928 29578
rect 10876 29514 10928 29520
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10784 29164 10836 29170
rect 10784 29106 10836 29112
rect 10508 29028 10560 29034
rect 10508 28970 10560 28976
rect 10416 28960 10468 28966
rect 10416 28902 10468 28908
rect 10520 28150 10548 28970
rect 10598 28792 10654 28801
rect 10598 28727 10654 28736
rect 10612 28694 10640 28727
rect 10600 28688 10652 28694
rect 10600 28630 10652 28636
rect 10692 28688 10744 28694
rect 10796 28676 10824 29106
rect 10744 28648 10824 28676
rect 10692 28630 10744 28636
rect 10784 28552 10836 28558
rect 10784 28494 10836 28500
rect 10692 28484 10744 28490
rect 10612 28444 10692 28472
rect 10508 28144 10560 28150
rect 10508 28086 10560 28092
rect 10416 27328 10468 27334
rect 10416 27270 10468 27276
rect 10428 25906 10456 27270
rect 10508 26920 10560 26926
rect 10612 26908 10640 28444
rect 10692 28426 10744 28432
rect 10796 28218 10824 28494
rect 10784 28212 10836 28218
rect 10784 28154 10836 28160
rect 10888 28082 10916 29514
rect 10968 28960 11020 28966
rect 10968 28902 11020 28908
rect 10980 28558 11008 28902
rect 10968 28552 11020 28558
rect 11072 28529 11100 30874
rect 11164 30705 11192 31470
rect 11150 30696 11206 30705
rect 11150 30631 11206 30640
rect 11256 30326 11284 31726
rect 11348 31726 11468 31754
rect 11348 31414 11376 31726
rect 11336 31408 11388 31414
rect 11336 31350 11388 31356
rect 11348 30666 11376 31350
rect 11520 31272 11572 31278
rect 11520 31214 11572 31220
rect 11428 30796 11480 30802
rect 11428 30738 11480 30744
rect 11336 30660 11388 30666
rect 11336 30602 11388 30608
rect 11348 30394 11376 30602
rect 11336 30388 11388 30394
rect 11336 30330 11388 30336
rect 11152 30320 11204 30326
rect 11150 30288 11152 30297
rect 11244 30320 11296 30326
rect 11204 30288 11206 30297
rect 11244 30262 11296 30268
rect 11150 30223 11206 30232
rect 11164 29782 11192 30223
rect 11244 30048 11296 30054
rect 11244 29990 11296 29996
rect 11152 29776 11204 29782
rect 11152 29718 11204 29724
rect 11256 29578 11284 29990
rect 11334 29880 11390 29889
rect 11440 29866 11468 30738
rect 11532 30666 11560 31214
rect 11520 30660 11572 30666
rect 11520 30602 11572 30608
rect 11532 30258 11560 30602
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 11518 30152 11574 30161
rect 11518 30087 11574 30096
rect 11390 29838 11468 29866
rect 11334 29815 11390 29824
rect 11244 29572 11296 29578
rect 11244 29514 11296 29520
rect 10968 28494 11020 28500
rect 11058 28520 11114 28529
rect 10876 28076 10928 28082
rect 10876 28018 10928 28024
rect 10692 28008 10744 28014
rect 10692 27950 10744 27956
rect 10704 27538 10732 27950
rect 10692 27532 10744 27538
rect 10692 27474 10744 27480
rect 10888 27470 10916 28018
rect 10876 27464 10928 27470
rect 10876 27406 10928 27412
rect 10980 26994 11008 28494
rect 11058 28455 11114 28464
rect 11060 28416 11112 28422
rect 11060 28358 11112 28364
rect 11242 28384 11298 28393
rect 11072 27470 11100 28358
rect 11242 28319 11298 28328
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 11058 27160 11114 27169
rect 11058 27095 11114 27104
rect 11072 27062 11100 27095
rect 11060 27056 11112 27062
rect 11060 26998 11112 27004
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10560 26880 10640 26908
rect 10876 26920 10928 26926
rect 10508 26862 10560 26868
rect 10876 26862 10928 26868
rect 10416 25900 10468 25906
rect 10416 25842 10468 25848
rect 10520 25362 10548 26862
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10612 25906 10640 26726
rect 10888 25906 10916 26862
rect 10968 26308 11020 26314
rect 10968 26250 11020 26256
rect 10980 26042 11008 26250
rect 11060 26240 11112 26246
rect 11060 26182 11112 26188
rect 11072 26042 11100 26182
rect 10968 26036 11020 26042
rect 10968 25978 11020 25984
rect 11060 26036 11112 26042
rect 11060 25978 11112 25984
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10508 25356 10560 25362
rect 10508 25298 10560 25304
rect 10888 25294 10916 25842
rect 10876 25288 10928 25294
rect 10876 25230 10928 25236
rect 10888 24818 10916 25230
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 10876 24676 10928 24682
rect 10876 24618 10928 24624
rect 10048 24608 10100 24614
rect 10048 24550 10100 24556
rect 10060 23798 10088 24550
rect 10888 23866 10916 24618
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 10048 23792 10100 23798
rect 10048 23734 10100 23740
rect 11072 23662 11100 25162
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 11256 23322 11284 28319
rect 11348 26738 11376 29815
rect 11532 29617 11560 30087
rect 11518 29608 11574 29617
rect 11518 29543 11574 29552
rect 11520 29096 11572 29102
rect 11520 29038 11572 29044
rect 11426 28792 11482 28801
rect 11426 28727 11482 28736
rect 11440 28490 11468 28727
rect 11532 28558 11560 29038
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 11428 28484 11480 28490
rect 11428 28426 11480 28432
rect 11348 26710 11468 26738
rect 11336 26580 11388 26586
rect 11336 26522 11388 26528
rect 11348 25838 11376 26522
rect 11336 25832 11388 25838
rect 11336 25774 11388 25780
rect 11440 25362 11468 26710
rect 11428 25356 11480 25362
rect 11428 25298 11480 25304
rect 11624 25294 11652 31855
rect 11716 30682 11744 33254
rect 11808 33017 11836 33476
rect 11888 33458 11940 33464
rect 12070 33416 12126 33425
rect 12070 33351 12072 33360
rect 12124 33351 12126 33360
rect 12072 33322 12124 33328
rect 12070 33280 12126 33289
rect 12070 33215 12126 33224
rect 11888 33108 11940 33114
rect 11888 33050 11940 33056
rect 11794 33008 11850 33017
rect 11794 32943 11850 32952
rect 11796 32904 11848 32910
rect 11796 32846 11848 32852
rect 11808 32774 11836 32846
rect 11900 32774 11928 33050
rect 12084 32978 12112 33215
rect 12176 33046 12204 34546
rect 12164 33040 12216 33046
rect 12164 32982 12216 32988
rect 12072 32972 12124 32978
rect 12072 32914 12124 32920
rect 11796 32768 11848 32774
rect 11796 32710 11848 32716
rect 11888 32768 11940 32774
rect 11940 32728 12020 32756
rect 11888 32710 11940 32716
rect 11796 32496 11848 32502
rect 11796 32438 11848 32444
rect 11808 32366 11836 32438
rect 11796 32360 11848 32366
rect 11796 32302 11848 32308
rect 11992 31328 12020 32728
rect 12268 32026 12296 37431
rect 14832 37324 14884 37330
rect 14832 37266 14884 37272
rect 14372 37256 14424 37262
rect 14372 37198 14424 37204
rect 14648 37256 14700 37262
rect 14648 37198 14700 37204
rect 12440 37188 12492 37194
rect 12440 37130 12492 37136
rect 12452 36922 12480 37130
rect 12716 37120 12768 37126
rect 12716 37062 12768 37068
rect 13084 37120 13136 37126
rect 13360 37120 13412 37126
rect 13084 37062 13136 37068
rect 13358 37088 13360 37097
rect 14280 37120 14332 37126
rect 13412 37088 13414 37097
rect 12440 36916 12492 36922
rect 12440 36858 12492 36864
rect 12728 36854 12756 37062
rect 12716 36848 12768 36854
rect 12716 36790 12768 36796
rect 12440 36712 12492 36718
rect 12440 36654 12492 36660
rect 12452 35698 12480 36654
rect 12728 36310 12756 36790
rect 13096 36786 13124 37062
rect 14280 37062 14332 37068
rect 13358 37023 13414 37032
rect 14292 36922 14320 37062
rect 13544 36916 13596 36922
rect 13544 36858 13596 36864
rect 14280 36916 14332 36922
rect 14280 36858 14332 36864
rect 13084 36780 13136 36786
rect 13084 36722 13136 36728
rect 13266 36408 13322 36417
rect 13266 36343 13322 36352
rect 12716 36304 12768 36310
rect 12716 36246 12768 36252
rect 12440 35692 12492 35698
rect 12440 35634 12492 35640
rect 13084 35692 13136 35698
rect 13084 35634 13136 35640
rect 12716 35624 12768 35630
rect 12716 35566 12768 35572
rect 12728 35154 12756 35566
rect 13096 35222 13124 35634
rect 13084 35216 13136 35222
rect 13084 35158 13136 35164
rect 12716 35148 12768 35154
rect 12716 35090 12768 35096
rect 12530 35048 12586 35057
rect 12530 34983 12586 34992
rect 12624 35012 12676 35018
rect 12440 34536 12492 34542
rect 12440 34478 12492 34484
rect 12452 33998 12480 34478
rect 12544 33998 12572 34983
rect 12624 34954 12676 34960
rect 12440 33992 12492 33998
rect 12440 33934 12492 33940
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 12348 33856 12400 33862
rect 12348 33798 12400 33804
rect 12360 33590 12388 33798
rect 12348 33584 12400 33590
rect 12348 33526 12400 33532
rect 12452 32842 12480 33934
rect 12348 32836 12400 32842
rect 12348 32778 12400 32784
rect 12440 32836 12492 32842
rect 12440 32778 12492 32784
rect 12360 32609 12388 32778
rect 12346 32600 12402 32609
rect 12346 32535 12402 32544
rect 12256 32020 12308 32026
rect 12256 31962 12308 31968
rect 12452 31754 12480 32778
rect 12544 32366 12572 33934
rect 12636 33522 12664 34954
rect 12808 34468 12860 34474
rect 12808 34410 12860 34416
rect 12900 34468 12952 34474
rect 12900 34410 12952 34416
rect 12624 33516 12676 33522
rect 12676 33476 12756 33504
rect 12624 33458 12676 33464
rect 12624 33108 12676 33114
rect 12624 33050 12676 33056
rect 12532 32360 12584 32366
rect 12532 32302 12584 32308
rect 12544 31890 12572 32302
rect 12532 31884 12584 31890
rect 12532 31826 12584 31832
rect 12452 31726 12572 31754
rect 12348 31680 12400 31686
rect 12348 31622 12400 31628
rect 12360 31346 12388 31622
rect 12348 31340 12400 31346
rect 11992 31300 12112 31328
rect 11980 31204 12032 31210
rect 11980 31146 12032 31152
rect 11716 30654 11928 30682
rect 11796 30592 11848 30598
rect 11796 30534 11848 30540
rect 11704 30252 11756 30258
rect 11704 30194 11756 30200
rect 11716 30036 11744 30194
rect 11808 30190 11836 30534
rect 11900 30297 11928 30654
rect 11886 30288 11942 30297
rect 11886 30223 11942 30232
rect 11796 30184 11848 30190
rect 11992 30172 12020 31146
rect 12084 30666 12112 31300
rect 12176 31300 12348 31328
rect 12176 30938 12204 31300
rect 12348 31282 12400 31288
rect 12440 31340 12492 31346
rect 12440 31282 12492 31288
rect 12256 31136 12308 31142
rect 12256 31078 12308 31084
rect 12164 30932 12216 30938
rect 12164 30874 12216 30880
rect 12072 30660 12124 30666
rect 12072 30602 12124 30608
rect 11992 30144 12112 30172
rect 11796 30126 11848 30132
rect 11716 30008 11836 30036
rect 11702 29200 11758 29209
rect 11702 29135 11704 29144
rect 11756 29135 11758 29144
rect 11704 29106 11756 29112
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 11716 27538 11744 28358
rect 11704 27532 11756 27538
rect 11704 27474 11756 27480
rect 11704 26376 11756 26382
rect 11704 26318 11756 26324
rect 11716 25906 11744 26318
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11808 25786 11836 30008
rect 11980 29776 12032 29782
rect 11980 29718 12032 29724
rect 11886 29608 11942 29617
rect 11886 29543 11942 29552
rect 11900 27418 11928 29543
rect 11992 29034 12020 29718
rect 11980 29028 12032 29034
rect 11980 28970 12032 28976
rect 12084 28801 12112 30144
rect 12070 28792 12126 28801
rect 12070 28727 12126 28736
rect 12084 28082 12112 28727
rect 12176 28082 12204 30874
rect 12268 30870 12296 31078
rect 12256 30864 12308 30870
rect 12452 30841 12480 31282
rect 12256 30806 12308 30812
rect 12438 30832 12494 30841
rect 12438 30767 12494 30776
rect 12440 30252 12492 30258
rect 12440 30194 12492 30200
rect 12348 30048 12400 30054
rect 12348 29990 12400 29996
rect 12256 29572 12308 29578
rect 12256 29514 12308 29520
rect 12268 28558 12296 29514
rect 12360 28558 12388 29990
rect 12452 29782 12480 30194
rect 12440 29776 12492 29782
rect 12440 29718 12492 29724
rect 12438 29608 12494 29617
rect 12438 29543 12440 29552
rect 12492 29543 12494 29552
rect 12440 29514 12492 29520
rect 12544 28994 12572 31726
rect 12636 31278 12664 33050
rect 12728 32910 12756 33476
rect 12820 33318 12848 34410
rect 12808 33312 12860 33318
rect 12808 33254 12860 33260
rect 12716 32904 12768 32910
rect 12716 32846 12768 32852
rect 12820 32756 12848 33254
rect 12912 33114 12940 34410
rect 13096 34202 13124 35158
rect 13280 35086 13308 36343
rect 13556 35329 13584 36858
rect 13636 36032 13688 36038
rect 13634 36000 13636 36009
rect 13688 36000 13690 36009
rect 13634 35935 13690 35944
rect 14292 35562 14320 36858
rect 14280 35556 14332 35562
rect 14280 35498 14332 35504
rect 14096 35488 14148 35494
rect 14384 35465 14412 37198
rect 14556 37120 14608 37126
rect 14556 37062 14608 37068
rect 14568 36417 14596 37062
rect 14554 36408 14610 36417
rect 14554 36343 14610 36352
rect 14096 35430 14148 35436
rect 14370 35456 14426 35465
rect 13542 35320 13598 35329
rect 13542 35255 13598 35264
rect 13636 35284 13688 35290
rect 13636 35226 13688 35232
rect 13268 35080 13320 35086
rect 13268 35022 13320 35028
rect 13174 34912 13230 34921
rect 13174 34847 13230 34856
rect 13084 34196 13136 34202
rect 13084 34138 13136 34144
rect 12992 33856 13044 33862
rect 12992 33798 13044 33804
rect 12900 33108 12952 33114
rect 12900 33050 12952 33056
rect 12728 32728 12848 32756
rect 12900 32768 12952 32774
rect 12898 32736 12900 32745
rect 13004 32756 13032 33798
rect 12952 32736 13032 32756
rect 12728 31482 12756 32728
rect 12954 32728 13032 32736
rect 12898 32671 12954 32680
rect 12808 32428 12860 32434
rect 12808 32370 12860 32376
rect 12716 31476 12768 31482
rect 12716 31418 12768 31424
rect 12624 31272 12676 31278
rect 12624 31214 12676 31220
rect 12728 31142 12756 31418
rect 12820 31210 12848 32370
rect 12808 31204 12860 31210
rect 12808 31146 12860 31152
rect 12624 31136 12676 31142
rect 12624 31078 12676 31084
rect 12716 31136 12768 31142
rect 12716 31078 12768 31084
rect 12636 30802 12664 31078
rect 12624 30796 12676 30802
rect 12624 30738 12676 30744
rect 12912 30666 12940 32671
rect 12990 32600 13046 32609
rect 13096 32586 13124 34138
rect 13188 34134 13216 34847
rect 13280 34762 13308 35022
rect 13280 34734 13584 34762
rect 13556 34474 13584 34734
rect 13544 34468 13596 34474
rect 13544 34410 13596 34416
rect 13648 34406 13676 35226
rect 14108 34950 14136 35430
rect 14370 35391 14426 35400
rect 14660 35222 14688 37198
rect 14844 36174 14872 37266
rect 15028 37262 15056 39200
rect 16948 38820 17000 38826
rect 16948 38762 17000 38768
rect 18144 38820 18196 38826
rect 18144 38762 18196 38768
rect 16488 38140 16540 38146
rect 16488 38082 16540 38088
rect 16500 37777 16528 38082
rect 15382 37768 15438 37777
rect 15382 37703 15438 37712
rect 16486 37768 16542 37777
rect 16486 37703 16542 37712
rect 15200 37460 15252 37466
rect 15200 37402 15252 37408
rect 15016 37256 15068 37262
rect 15016 37198 15068 37204
rect 15016 37120 15068 37126
rect 15016 37062 15068 37068
rect 14924 36780 14976 36786
rect 14924 36722 14976 36728
rect 14936 36310 14964 36722
rect 15028 36582 15056 37062
rect 15106 36952 15162 36961
rect 15212 36938 15240 37402
rect 15162 36910 15240 36938
rect 15106 36887 15162 36896
rect 15016 36576 15068 36582
rect 15016 36518 15068 36524
rect 15200 36576 15252 36582
rect 15200 36518 15252 36524
rect 14924 36304 14976 36310
rect 14924 36246 14976 36252
rect 15212 36242 15240 36518
rect 15200 36236 15252 36242
rect 15200 36178 15252 36184
rect 14832 36168 14884 36174
rect 14832 36110 14884 36116
rect 14648 35216 14700 35222
rect 14648 35158 14700 35164
rect 14844 35154 14872 36110
rect 15212 35698 15240 36178
rect 15200 35692 15252 35698
rect 15200 35634 15252 35640
rect 15292 35488 15344 35494
rect 15014 35456 15070 35465
rect 15014 35391 15070 35400
rect 15198 35456 15254 35465
rect 15292 35430 15344 35436
rect 15198 35391 15254 35400
rect 14832 35148 14884 35154
rect 14832 35090 14884 35096
rect 14556 35080 14608 35086
rect 14556 35022 14608 35028
rect 14096 34944 14148 34950
rect 14096 34886 14148 34892
rect 14280 34672 14332 34678
rect 14280 34614 14332 34620
rect 14004 34604 14056 34610
rect 14004 34546 14056 34552
rect 14188 34604 14240 34610
rect 14188 34546 14240 34552
rect 13268 34400 13320 34406
rect 13268 34342 13320 34348
rect 13636 34400 13688 34406
rect 13636 34342 13688 34348
rect 13820 34400 13872 34406
rect 13820 34342 13872 34348
rect 13176 34128 13228 34134
rect 13176 34070 13228 34076
rect 13176 33924 13228 33930
rect 13176 33866 13228 33872
rect 13188 33454 13216 33866
rect 13280 33590 13308 34342
rect 13360 34196 13412 34202
rect 13412 34156 13676 34184
rect 13360 34138 13412 34144
rect 13542 34096 13598 34105
rect 13542 34031 13598 34040
rect 13452 33856 13504 33862
rect 13452 33798 13504 33804
rect 13464 33658 13492 33798
rect 13556 33658 13584 34031
rect 13648 33998 13676 34156
rect 13832 34105 13860 34342
rect 13818 34096 13874 34105
rect 13818 34031 13874 34040
rect 13832 33998 13860 34031
rect 13636 33992 13688 33998
rect 13820 33992 13872 33998
rect 13688 33952 13768 33980
rect 13636 33934 13688 33940
rect 13452 33652 13504 33658
rect 13452 33594 13504 33600
rect 13544 33652 13596 33658
rect 13544 33594 13596 33600
rect 13268 33584 13320 33590
rect 13268 33526 13320 33532
rect 13176 33448 13228 33454
rect 13176 33390 13228 33396
rect 13266 33144 13322 33153
rect 13266 33079 13268 33088
rect 13320 33079 13322 33088
rect 13268 33050 13320 33056
rect 13360 33040 13412 33046
rect 13360 32982 13412 32988
rect 13464 32994 13492 33594
rect 13740 33572 13768 33952
rect 13820 33934 13872 33940
rect 13910 33960 13966 33969
rect 13910 33895 13966 33904
rect 13740 33544 13860 33572
rect 13636 33516 13688 33522
rect 13688 33476 13768 33504
rect 13636 33458 13688 33464
rect 13544 33448 13596 33454
rect 13544 33390 13596 33396
rect 13556 33114 13584 33390
rect 13740 33318 13768 33476
rect 13832 33454 13860 33544
rect 13820 33448 13872 33454
rect 13820 33390 13872 33396
rect 13728 33312 13780 33318
rect 13820 33312 13872 33318
rect 13780 33260 13820 33266
rect 13728 33254 13872 33260
rect 13740 33238 13860 33254
rect 13544 33108 13596 33114
rect 13544 33050 13596 33056
rect 13096 32558 13216 32586
rect 12990 32535 13046 32544
rect 13004 32502 13032 32535
rect 12992 32496 13044 32502
rect 12992 32438 13044 32444
rect 12992 32360 13044 32366
rect 12992 32302 13044 32308
rect 13084 32360 13136 32366
rect 13084 32302 13136 32308
rect 13004 31958 13032 32302
rect 13096 32026 13124 32302
rect 13084 32020 13136 32026
rect 13084 31962 13136 31968
rect 12992 31952 13044 31958
rect 12992 31894 13044 31900
rect 12992 31816 13044 31822
rect 12992 31758 13044 31764
rect 13004 30734 13032 31758
rect 13096 31346 13124 31962
rect 13188 31822 13216 32558
rect 13372 32337 13400 32982
rect 13464 32966 13676 32994
rect 13544 32904 13596 32910
rect 13544 32846 13596 32852
rect 13358 32328 13414 32337
rect 13268 32292 13320 32298
rect 13358 32263 13414 32272
rect 13268 32234 13320 32240
rect 13280 32042 13308 32234
rect 13280 32014 13400 32042
rect 13372 31822 13400 32014
rect 13452 31952 13504 31958
rect 13452 31894 13504 31900
rect 13176 31816 13228 31822
rect 13176 31758 13228 31764
rect 13360 31816 13412 31822
rect 13360 31758 13412 31764
rect 13464 31686 13492 31894
rect 13452 31680 13504 31686
rect 13174 31648 13230 31657
rect 13452 31622 13504 31628
rect 13174 31583 13230 31592
rect 13084 31340 13136 31346
rect 13084 31282 13136 31288
rect 13082 30832 13138 30841
rect 13082 30767 13138 30776
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 12900 30660 12952 30666
rect 12900 30602 12952 30608
rect 12912 30326 12940 30602
rect 13096 30580 13124 30767
rect 13188 30734 13216 31583
rect 13556 31346 13584 32846
rect 13648 31906 13676 32966
rect 13740 32212 13768 33238
rect 13818 33144 13874 33153
rect 13818 33079 13874 33088
rect 13832 32570 13860 33079
rect 13820 32564 13872 32570
rect 13820 32506 13872 32512
rect 13740 32184 13860 32212
rect 13648 31878 13768 31906
rect 13636 31816 13688 31822
rect 13636 31758 13688 31764
rect 13648 31482 13676 31758
rect 13636 31476 13688 31482
rect 13636 31418 13688 31424
rect 13544 31340 13596 31346
rect 13544 31282 13596 31288
rect 13268 31272 13320 31278
rect 13268 31214 13320 31220
rect 13176 30728 13228 30734
rect 13176 30670 13228 30676
rect 13004 30552 13124 30580
rect 12900 30320 12952 30326
rect 12900 30262 12952 30268
rect 12624 30184 12676 30190
rect 12624 30126 12676 30132
rect 12716 30184 12768 30190
rect 12808 30184 12860 30190
rect 12716 30126 12768 30132
rect 12806 30152 12808 30161
rect 12860 30152 12862 30161
rect 12636 29730 12664 30126
rect 12728 29850 12756 30126
rect 12806 30087 12862 30096
rect 12716 29844 12768 29850
rect 12716 29786 12768 29792
rect 13004 29753 13032 30552
rect 13176 30388 13228 30394
rect 13176 30330 13228 30336
rect 13084 30048 13136 30054
rect 13084 29990 13136 29996
rect 12990 29744 13046 29753
rect 12636 29702 12756 29730
rect 12624 29572 12676 29578
rect 12624 29514 12676 29520
rect 12636 29102 12664 29514
rect 12728 29510 12756 29702
rect 12990 29679 13046 29688
rect 12992 29640 13044 29646
rect 12992 29582 13044 29588
rect 12716 29504 12768 29510
rect 12716 29446 12768 29452
rect 12728 29306 12756 29446
rect 12716 29300 12768 29306
rect 12716 29242 12768 29248
rect 12624 29096 12676 29102
rect 12624 29038 12676 29044
rect 12452 28966 12572 28994
rect 12452 28608 12480 28966
rect 12532 28620 12584 28626
rect 12452 28580 12532 28608
rect 12256 28552 12308 28558
rect 12256 28494 12308 28500
rect 12348 28552 12400 28558
rect 12348 28494 12400 28500
rect 12348 28416 12400 28422
rect 12348 28358 12400 28364
rect 12072 28076 12124 28082
rect 12072 28018 12124 28024
rect 12164 28076 12216 28082
rect 12164 28018 12216 28024
rect 12256 28076 12308 28082
rect 12256 28018 12308 28024
rect 12072 27600 12124 27606
rect 12176 27588 12204 28018
rect 12268 27674 12296 28018
rect 12256 27668 12308 27674
rect 12256 27610 12308 27616
rect 12124 27560 12204 27588
rect 12072 27542 12124 27548
rect 12360 27538 12388 28358
rect 12452 28082 12480 28580
rect 12532 28562 12584 28568
rect 12636 28132 12664 29038
rect 12716 28552 12768 28558
rect 12716 28494 12768 28500
rect 12728 28218 12756 28494
rect 12808 28484 12860 28490
rect 12808 28426 12860 28432
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 12544 28104 12664 28132
rect 12440 28076 12492 28082
rect 12440 28018 12492 28024
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 11900 27390 12112 27418
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 12084 27282 12112 27390
rect 11716 25758 11836 25786
rect 11716 25702 11744 25758
rect 11704 25696 11756 25702
rect 11704 25638 11756 25644
rect 11612 25288 11664 25294
rect 11612 25230 11664 25236
rect 11704 25152 11756 25158
rect 11704 25094 11756 25100
rect 11716 24818 11744 25094
rect 11900 24818 11928 27270
rect 11992 27033 12020 27270
rect 12084 27254 12204 27282
rect 11978 27024 12034 27033
rect 11978 26959 12034 26968
rect 11980 26240 12032 26246
rect 11980 26182 12032 26188
rect 11992 25906 12020 26182
rect 11980 25900 12032 25906
rect 11980 25842 12032 25848
rect 12072 25220 12124 25226
rect 12072 25162 12124 25168
rect 12084 24818 12112 25162
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 11428 24744 11480 24750
rect 11428 24686 11480 24692
rect 11440 24206 11468 24686
rect 11992 24274 12020 24754
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 11440 23186 11468 24142
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 11428 23180 11480 23186
rect 11428 23122 11480 23128
rect 11992 23118 12020 23462
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 11060 22024 11112 22030
rect 11112 21972 11284 21978
rect 11060 21966 11284 21972
rect 11072 21950 11284 21966
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 8390 19136 8446 19145
rect 4214 19068 4522 19077
rect 8390 19071 8446 19080
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 11072 18630 11100 21286
rect 11256 20942 11284 21950
rect 11796 21956 11848 21962
rect 11796 21898 11848 21904
rect 11808 21690 11836 21898
rect 12176 21690 12204 27254
rect 12256 26784 12308 26790
rect 12256 26726 12308 26732
rect 12268 26314 12296 26726
rect 12256 26308 12308 26314
rect 12256 26250 12308 26256
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12268 24138 12296 24550
rect 12360 24206 12388 27474
rect 12452 27470 12480 28018
rect 12544 27946 12572 28104
rect 12532 27940 12584 27946
rect 12532 27882 12584 27888
rect 12440 27464 12492 27470
rect 12440 27406 12492 27412
rect 12452 26314 12480 27406
rect 12440 26308 12492 26314
rect 12440 26250 12492 26256
rect 12544 26246 12572 27882
rect 12716 27872 12768 27878
rect 12716 27814 12768 27820
rect 12728 27674 12756 27814
rect 12716 27668 12768 27674
rect 12716 27610 12768 27616
rect 12728 27470 12756 27610
rect 12820 27470 12848 28426
rect 12900 28008 12952 28014
rect 12900 27950 12952 27956
rect 12716 27464 12768 27470
rect 12716 27406 12768 27412
rect 12808 27464 12860 27470
rect 12808 27406 12860 27412
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12728 25974 12756 27406
rect 12820 27062 12848 27406
rect 12808 27056 12860 27062
rect 12808 26998 12860 27004
rect 12912 26382 12940 27950
rect 13004 27452 13032 29582
rect 13096 29578 13124 29990
rect 13084 29572 13136 29578
rect 13084 29514 13136 29520
rect 13096 29034 13124 29514
rect 13084 29028 13136 29034
rect 13084 28970 13136 28976
rect 13188 28994 13216 30330
rect 13280 29850 13308 31214
rect 13450 30968 13506 30977
rect 13450 30903 13506 30912
rect 13358 30832 13414 30841
rect 13358 30767 13414 30776
rect 13372 30734 13400 30767
rect 13464 30734 13492 30903
rect 13360 30728 13412 30734
rect 13360 30670 13412 30676
rect 13452 30728 13504 30734
rect 13452 30670 13504 30676
rect 13452 30592 13504 30598
rect 13452 30534 13504 30540
rect 13268 29844 13320 29850
rect 13268 29786 13320 29792
rect 13280 29170 13308 29786
rect 13464 29510 13492 30534
rect 13648 30258 13676 31418
rect 13740 31414 13768 31878
rect 13832 31464 13860 32184
rect 13924 32026 13952 33895
rect 14016 33862 14044 34546
rect 14200 33930 14228 34546
rect 14188 33924 14240 33930
rect 14188 33866 14240 33872
rect 14004 33856 14056 33862
rect 14004 33798 14056 33804
rect 14004 33516 14056 33522
rect 14004 33458 14056 33464
rect 14016 33114 14044 33458
rect 14004 33108 14056 33114
rect 14004 33050 14056 33056
rect 14096 32972 14148 32978
rect 14096 32914 14148 32920
rect 14108 32745 14136 32914
rect 14200 32910 14228 33866
rect 14292 33386 14320 34614
rect 14372 34604 14424 34610
rect 14372 34546 14424 34552
rect 14384 34066 14412 34546
rect 14464 34400 14516 34406
rect 14464 34342 14516 34348
rect 14372 34060 14424 34066
rect 14372 34002 14424 34008
rect 14370 33824 14426 33833
rect 14370 33759 14426 33768
rect 14280 33380 14332 33386
rect 14280 33322 14332 33328
rect 14188 32904 14240 32910
rect 14188 32846 14240 32852
rect 14188 32768 14240 32774
rect 14094 32736 14150 32745
rect 14188 32710 14240 32716
rect 14280 32768 14332 32774
rect 14280 32710 14332 32716
rect 14094 32671 14150 32680
rect 14004 32564 14056 32570
rect 14004 32506 14056 32512
rect 14016 32337 14044 32506
rect 14096 32428 14148 32434
rect 14096 32370 14148 32376
rect 14002 32328 14058 32337
rect 14002 32263 14058 32272
rect 13912 32020 13964 32026
rect 13912 31962 13964 31968
rect 13832 31436 13952 31464
rect 13728 31408 13780 31414
rect 13728 31350 13780 31356
rect 13924 31346 13952 31436
rect 14108 31385 14136 32370
rect 14200 31890 14228 32710
rect 14188 31884 14240 31890
rect 14188 31826 14240 31832
rect 14292 31822 14320 32710
rect 14384 32609 14412 33759
rect 14370 32600 14426 32609
rect 14370 32535 14426 32544
rect 14476 32026 14504 34342
rect 14568 34202 14596 35022
rect 15028 34785 15056 35391
rect 14738 34776 14794 34785
rect 14738 34711 14794 34720
rect 15014 34776 15070 34785
rect 15212 34746 15240 35391
rect 15014 34711 15070 34720
rect 15200 34740 15252 34746
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 14660 34406 14688 34546
rect 14648 34400 14700 34406
rect 14648 34342 14700 34348
rect 14556 34196 14608 34202
rect 14556 34138 14608 34144
rect 14568 33522 14596 34138
rect 14660 33998 14688 34342
rect 14752 34202 14780 34711
rect 15200 34682 15252 34688
rect 14922 34640 14978 34649
rect 14922 34575 14978 34584
rect 15016 34604 15068 34610
rect 14740 34196 14792 34202
rect 14740 34138 14792 34144
rect 14648 33992 14700 33998
rect 14648 33934 14700 33940
rect 14648 33584 14700 33590
rect 14648 33526 14700 33532
rect 14556 33516 14608 33522
rect 14556 33458 14608 33464
rect 14660 32978 14688 33526
rect 14648 32972 14700 32978
rect 14648 32914 14700 32920
rect 14646 32600 14702 32609
rect 14646 32535 14702 32544
rect 14660 32337 14688 32535
rect 14646 32328 14702 32337
rect 14646 32263 14702 32272
rect 14464 32020 14516 32026
rect 14464 31962 14516 31968
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 14464 31816 14516 31822
rect 14464 31758 14516 31764
rect 14372 31680 14424 31686
rect 14476 31657 14504 31758
rect 14372 31622 14424 31628
rect 14462 31648 14518 31657
rect 14384 31482 14412 31622
rect 14462 31583 14518 31592
rect 14372 31476 14424 31482
rect 14372 31418 14424 31424
rect 14094 31376 14150 31385
rect 13820 31340 13872 31346
rect 13820 31282 13872 31288
rect 13912 31340 13964 31346
rect 14094 31311 14150 31320
rect 13912 31282 13964 31288
rect 13728 31272 13780 31278
rect 13728 31214 13780 31220
rect 13740 30666 13768 31214
rect 13832 30734 13860 31282
rect 13820 30728 13872 30734
rect 13820 30670 13872 30676
rect 13728 30660 13780 30666
rect 13728 30602 13780 30608
rect 13924 30569 13952 31282
rect 13910 30560 13966 30569
rect 13910 30495 13966 30504
rect 13636 30252 13688 30258
rect 13636 30194 13688 30200
rect 13648 29714 13676 30194
rect 13728 30184 13780 30190
rect 13728 30126 13780 30132
rect 13636 29708 13688 29714
rect 13636 29650 13688 29656
rect 13740 29646 13768 30126
rect 13820 30048 13872 30054
rect 13820 29990 13872 29996
rect 13728 29640 13780 29646
rect 13728 29582 13780 29588
rect 13740 29510 13768 29582
rect 13452 29504 13504 29510
rect 13452 29446 13504 29452
rect 13728 29504 13780 29510
rect 13728 29446 13780 29452
rect 13268 29164 13320 29170
rect 13268 29106 13320 29112
rect 13096 27674 13124 28970
rect 13188 28966 13676 28994
rect 13542 28656 13598 28665
rect 13542 28591 13598 28600
rect 13556 28422 13584 28591
rect 13452 28416 13504 28422
rect 13452 28358 13504 28364
rect 13544 28416 13596 28422
rect 13544 28358 13596 28364
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 13188 27674 13216 28018
rect 13084 27668 13136 27674
rect 13084 27610 13136 27616
rect 13176 27668 13228 27674
rect 13176 27610 13228 27616
rect 13360 27600 13412 27606
rect 13360 27542 13412 27548
rect 13084 27464 13136 27470
rect 13004 27424 13084 27452
rect 13004 27130 13032 27424
rect 13084 27406 13136 27412
rect 12992 27124 13044 27130
rect 12992 27066 13044 27072
rect 13372 26994 13400 27542
rect 13464 27470 13492 28358
rect 13648 28082 13676 28966
rect 13726 28792 13782 28801
rect 13726 28727 13782 28736
rect 13740 28490 13768 28727
rect 13728 28484 13780 28490
rect 13728 28426 13780 28432
rect 13636 28076 13688 28082
rect 13636 28018 13688 28024
rect 13452 27464 13504 27470
rect 13452 27406 13504 27412
rect 13464 27130 13492 27406
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 13450 27024 13506 27033
rect 13360 26988 13412 26994
rect 13450 26959 13452 26968
rect 13360 26930 13412 26936
rect 13504 26959 13506 26968
rect 13452 26930 13504 26936
rect 13176 26920 13228 26926
rect 13176 26862 13228 26868
rect 13266 26888 13322 26897
rect 13188 26518 13216 26862
rect 13266 26823 13322 26832
rect 13280 26790 13308 26823
rect 13268 26784 13320 26790
rect 13268 26726 13320 26732
rect 13176 26512 13228 26518
rect 13176 26454 13228 26460
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12992 26240 13044 26246
rect 12992 26182 13044 26188
rect 13004 26042 13032 26182
rect 12992 26036 13044 26042
rect 12992 25978 13044 25984
rect 12716 25968 12768 25974
rect 12716 25910 12768 25916
rect 12990 25800 13046 25809
rect 12990 25735 13046 25744
rect 12900 24744 12952 24750
rect 12900 24686 12952 24692
rect 12912 24274 12940 24686
rect 12900 24268 12952 24274
rect 12900 24210 12952 24216
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12360 23866 12388 24142
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12256 23656 12308 23662
rect 12256 23598 12308 23604
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12268 21486 12296 23598
rect 12820 23322 12848 23666
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12912 22642 12940 24210
rect 13004 24070 13032 25735
rect 13464 25294 13492 26930
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 13648 25140 13676 28018
rect 13740 25906 13768 28426
rect 13728 25900 13780 25906
rect 13728 25842 13780 25848
rect 13372 25112 13676 25140
rect 13372 24070 13400 25112
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 13084 24064 13136 24070
rect 13084 24006 13136 24012
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13096 23798 13124 24006
rect 13084 23792 13136 23798
rect 13084 23734 13136 23740
rect 13464 23730 13492 24210
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13452 23724 13504 23730
rect 13452 23666 13504 23672
rect 13740 23526 13768 24142
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13832 23118 13860 29990
rect 13924 29306 13952 30495
rect 13912 29300 13964 29306
rect 13912 29242 13964 29248
rect 14108 28801 14136 31311
rect 14372 31272 14424 31278
rect 14372 31214 14424 31220
rect 14280 29572 14332 29578
rect 14280 29514 14332 29520
rect 14094 28792 14150 28801
rect 14094 28727 14150 28736
rect 14292 28558 14320 29514
rect 14384 28762 14412 31214
rect 14554 30968 14610 30977
rect 14464 30932 14516 30938
rect 14554 30903 14610 30912
rect 14464 30874 14516 30880
rect 14476 30802 14504 30874
rect 14464 30796 14516 30802
rect 14464 30738 14516 30744
rect 14372 28756 14424 28762
rect 14372 28698 14424 28704
rect 14188 28552 14240 28558
rect 14188 28494 14240 28500
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 14200 28150 14228 28494
rect 14188 28144 14240 28150
rect 14188 28086 14240 28092
rect 14096 27940 14148 27946
rect 14096 27882 14148 27888
rect 14108 27402 14136 27882
rect 14096 27396 14148 27402
rect 14096 27338 14148 27344
rect 13912 26920 13964 26926
rect 13912 26862 13964 26868
rect 13924 26382 13952 26862
rect 13912 26376 13964 26382
rect 13912 26318 13964 26324
rect 13924 25838 13952 26318
rect 14200 25906 14228 28086
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 14188 25900 14240 25906
rect 14188 25842 14240 25848
rect 13912 25832 13964 25838
rect 13912 25774 13964 25780
rect 14108 25702 14136 25842
rect 14096 25696 14148 25702
rect 14096 25638 14148 25644
rect 13912 25424 13964 25430
rect 13912 25366 13964 25372
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 13096 22710 13124 22918
rect 13084 22704 13136 22710
rect 13084 22646 13136 22652
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12912 22098 12940 22578
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 12900 22092 12952 22098
rect 12900 22034 12952 22040
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 12360 21622 12388 21830
rect 12348 21616 12400 21622
rect 12348 21558 12400 21564
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 13096 21418 13124 21830
rect 13464 21486 13492 22374
rect 13924 22094 13952 25366
rect 14004 24132 14056 24138
rect 14004 24074 14056 24080
rect 14016 23730 14044 24074
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 14292 22710 14320 28494
rect 14384 24750 14412 28698
rect 14568 27606 14596 30903
rect 14556 27600 14608 27606
rect 14556 27542 14608 27548
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14568 27033 14596 27406
rect 14554 27024 14610 27033
rect 14464 26988 14516 26994
rect 14554 26959 14610 26968
rect 14464 26930 14516 26936
rect 14476 26314 14504 26930
rect 14464 26308 14516 26314
rect 14464 26250 14516 26256
rect 14476 25906 14504 26250
rect 14464 25900 14516 25906
rect 14464 25842 14516 25848
rect 14660 25294 14688 32263
rect 14752 30841 14780 34138
rect 14936 34105 14964 34575
rect 15016 34546 15068 34552
rect 14922 34096 14978 34105
rect 14922 34031 14978 34040
rect 14832 33992 14884 33998
rect 14832 33934 14884 33940
rect 14924 33992 14976 33998
rect 14924 33934 14976 33940
rect 14844 32881 14872 33934
rect 14936 33658 14964 33934
rect 14924 33652 14976 33658
rect 14924 33594 14976 33600
rect 15028 33318 15056 34546
rect 15108 34536 15160 34542
rect 15160 34496 15240 34524
rect 15304 34513 15332 35430
rect 15108 34478 15160 34484
rect 15108 33992 15160 33998
rect 15108 33934 15160 33940
rect 15120 33658 15148 33934
rect 15108 33652 15160 33658
rect 15108 33594 15160 33600
rect 15108 33516 15160 33522
rect 15108 33458 15160 33464
rect 15016 33312 15068 33318
rect 15016 33254 15068 33260
rect 15028 32978 15056 33254
rect 15016 32972 15068 32978
rect 15016 32914 15068 32920
rect 14830 32872 14886 32881
rect 14830 32807 14886 32816
rect 14832 32496 14884 32502
rect 14832 32438 14884 32444
rect 14844 31754 14872 32438
rect 15016 32360 15068 32366
rect 15016 32302 15068 32308
rect 14924 32020 14976 32026
rect 14924 31962 14976 31968
rect 14832 31748 14884 31754
rect 14832 31690 14884 31696
rect 14936 31634 14964 31962
rect 15028 31890 15056 32302
rect 15120 32230 15148 33458
rect 15212 32502 15240 34496
rect 15290 34504 15346 34513
rect 15290 34439 15346 34448
rect 15396 33946 15424 37703
rect 16488 37392 16540 37398
rect 16488 37334 16540 37340
rect 16500 37244 16528 37334
rect 16500 37216 16620 37244
rect 15752 37188 15804 37194
rect 15752 37130 15804 37136
rect 15936 37188 15988 37194
rect 15936 37130 15988 37136
rect 15764 36922 15792 37130
rect 15948 37097 15976 37130
rect 15934 37088 15990 37097
rect 15934 37023 15990 37032
rect 15752 36916 15804 36922
rect 15752 36858 15804 36864
rect 15844 36644 15896 36650
rect 15844 36586 15896 36592
rect 15856 36394 15884 36586
rect 15764 36366 15884 36394
rect 15764 36038 15792 36366
rect 15844 36304 15896 36310
rect 15844 36246 15896 36252
rect 15752 36032 15804 36038
rect 15752 35974 15804 35980
rect 15764 35698 15792 35974
rect 15752 35692 15804 35698
rect 15752 35634 15804 35640
rect 15476 35624 15528 35630
rect 15476 35566 15528 35572
rect 15750 35592 15806 35601
rect 15488 34746 15516 35566
rect 15750 35527 15806 35536
rect 15568 35080 15620 35086
rect 15764 35057 15792 35527
rect 15568 35022 15620 35028
rect 15750 35048 15806 35057
rect 15476 34740 15528 34746
rect 15476 34682 15528 34688
rect 15488 34048 15516 34682
rect 15580 34241 15608 35022
rect 15750 34983 15806 34992
rect 15660 34944 15712 34950
rect 15660 34886 15712 34892
rect 15566 34232 15622 34241
rect 15566 34167 15622 34176
rect 15568 34060 15620 34066
rect 15488 34020 15568 34048
rect 15568 34002 15620 34008
rect 15672 33998 15700 34886
rect 15856 34513 15884 36246
rect 15948 35834 15976 37023
rect 16486 36272 16542 36281
rect 16486 36207 16542 36216
rect 16396 36100 16448 36106
rect 16396 36042 16448 36048
rect 15936 35828 15988 35834
rect 15936 35770 15988 35776
rect 15948 34649 15976 35770
rect 16304 35624 16356 35630
rect 16304 35566 16356 35572
rect 16210 35320 16266 35329
rect 16210 35255 16266 35264
rect 16120 35080 16172 35086
rect 16120 35022 16172 35028
rect 15934 34640 15990 34649
rect 15934 34575 15990 34584
rect 15842 34504 15898 34513
rect 15842 34439 15898 34448
rect 16028 34468 16080 34474
rect 16028 34410 16080 34416
rect 15844 34196 15896 34202
rect 15844 34138 15896 34144
rect 15856 34066 15884 34138
rect 15752 34060 15804 34066
rect 15752 34002 15804 34008
rect 15844 34060 15896 34066
rect 15844 34002 15896 34008
rect 15660 33992 15712 33998
rect 15396 33918 15608 33946
rect 15660 33934 15712 33940
rect 15476 33856 15528 33862
rect 15476 33798 15528 33804
rect 15292 33108 15344 33114
rect 15292 33050 15344 33056
rect 15200 32496 15252 32502
rect 15200 32438 15252 32444
rect 15108 32224 15160 32230
rect 15108 32166 15160 32172
rect 15016 31884 15068 31890
rect 15016 31826 15068 31832
rect 14844 31606 14964 31634
rect 14844 30938 14872 31606
rect 14922 31512 14978 31521
rect 14922 31447 14978 31456
rect 14936 31346 14964 31447
rect 14924 31340 14976 31346
rect 14924 31282 14976 31288
rect 15016 31272 15068 31278
rect 15016 31214 15068 31220
rect 14832 30932 14884 30938
rect 14832 30874 14884 30880
rect 14738 30832 14794 30841
rect 14738 30767 14794 30776
rect 15028 30666 15056 31214
rect 15016 30660 15068 30666
rect 15016 30602 15068 30608
rect 14832 30592 14884 30598
rect 14752 30552 14832 30580
rect 14752 29646 14780 30552
rect 14832 30534 14884 30540
rect 15120 30394 15148 32166
rect 15304 32042 15332 33050
rect 15488 32910 15516 33798
rect 15580 33590 15608 33918
rect 15764 33658 15792 34002
rect 15752 33652 15804 33658
rect 15752 33594 15804 33600
rect 15568 33584 15620 33590
rect 15568 33526 15620 33532
rect 15660 33584 15712 33590
rect 15660 33526 15712 33532
rect 15672 33114 15700 33526
rect 15764 33522 15792 33594
rect 15752 33516 15804 33522
rect 15752 33458 15804 33464
rect 15856 33289 15884 34002
rect 16040 33998 16068 34410
rect 16028 33992 16080 33998
rect 16028 33934 16080 33940
rect 16040 33810 16068 33934
rect 15948 33782 16068 33810
rect 15948 33522 15976 33782
rect 15936 33516 15988 33522
rect 15936 33458 15988 33464
rect 15842 33280 15898 33289
rect 15842 33215 15898 33224
rect 16132 33114 16160 35022
rect 15660 33108 15712 33114
rect 15580 33068 15660 33096
rect 15384 32904 15436 32910
rect 15384 32846 15436 32852
rect 15476 32904 15528 32910
rect 15476 32846 15528 32852
rect 15396 32298 15424 32846
rect 15474 32600 15530 32609
rect 15474 32535 15530 32544
rect 15488 32434 15516 32535
rect 15476 32428 15528 32434
rect 15476 32370 15528 32376
rect 15384 32292 15436 32298
rect 15384 32234 15436 32240
rect 15382 32192 15438 32201
rect 15382 32127 15438 32136
rect 15212 32014 15332 32042
rect 15212 31414 15240 32014
rect 15292 31952 15344 31958
rect 15292 31894 15344 31900
rect 15304 31754 15332 31894
rect 15292 31748 15344 31754
rect 15292 31690 15344 31696
rect 15200 31408 15252 31414
rect 15200 31350 15252 31356
rect 15198 31240 15254 31249
rect 15198 31175 15200 31184
rect 15252 31175 15254 31184
rect 15200 31146 15252 31152
rect 15304 30734 15332 31690
rect 15396 30734 15424 32127
rect 15488 31822 15516 32370
rect 15476 31816 15528 31822
rect 15476 31758 15528 31764
rect 15292 30728 15344 30734
rect 15292 30670 15344 30676
rect 15384 30728 15436 30734
rect 15384 30670 15436 30676
rect 15108 30388 15160 30394
rect 15108 30330 15160 30336
rect 14832 30252 14884 30258
rect 14832 30194 14884 30200
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14752 29170 14780 29582
rect 14844 29306 14872 30194
rect 15028 29578 15056 30194
rect 15580 29866 15608 33068
rect 15660 33050 15712 33056
rect 15844 33108 15896 33114
rect 15844 33050 15896 33056
rect 16120 33108 16172 33114
rect 16120 33050 16172 33056
rect 15752 32972 15804 32978
rect 15752 32914 15804 32920
rect 15660 32224 15712 32230
rect 15660 32166 15712 32172
rect 15672 31385 15700 32166
rect 15658 31376 15714 31385
rect 15658 31311 15714 31320
rect 15764 30802 15792 32914
rect 15856 32570 15884 33050
rect 15934 32872 15990 32881
rect 15934 32807 15990 32816
rect 15844 32564 15896 32570
rect 15844 32506 15896 32512
rect 15948 31414 15976 32807
rect 16224 32722 16252 35255
rect 16316 33969 16344 35566
rect 16408 35290 16436 36042
rect 16500 35873 16528 36207
rect 16486 35864 16542 35873
rect 16486 35799 16542 35808
rect 16396 35284 16448 35290
rect 16396 35226 16448 35232
rect 16394 34504 16450 34513
rect 16394 34439 16450 34448
rect 16408 34241 16436 34439
rect 16394 34232 16450 34241
rect 16394 34167 16450 34176
rect 16302 33960 16358 33969
rect 16302 33895 16358 33904
rect 16408 32756 16436 34167
rect 16488 33516 16540 33522
rect 16488 33458 16540 33464
rect 16500 33114 16528 33458
rect 16488 33108 16540 33114
rect 16488 33050 16540 33056
rect 16040 32694 16252 32722
rect 16316 32728 16436 32756
rect 15936 31408 15988 31414
rect 15936 31350 15988 31356
rect 16040 31226 16068 32694
rect 16316 32586 16344 32728
rect 16120 32564 16172 32570
rect 16120 32506 16172 32512
rect 16224 32558 16344 32586
rect 16132 31822 16160 32506
rect 16224 32026 16252 32558
rect 16212 32020 16264 32026
rect 16212 31962 16264 31968
rect 16120 31816 16172 31822
rect 16120 31758 16172 31764
rect 16304 31816 16356 31822
rect 16304 31758 16356 31764
rect 16316 31657 16344 31758
rect 16302 31648 16358 31657
rect 16302 31583 16358 31592
rect 16040 31198 16344 31226
rect 16120 31136 16172 31142
rect 16120 31078 16172 31084
rect 15752 30796 15804 30802
rect 15752 30738 15804 30744
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15580 29838 15884 29866
rect 15384 29776 15436 29782
rect 15384 29718 15436 29724
rect 15750 29744 15806 29753
rect 15016 29572 15068 29578
rect 15016 29514 15068 29520
rect 14832 29300 14884 29306
rect 14832 29242 14884 29248
rect 15028 29238 15056 29514
rect 15016 29232 15068 29238
rect 15016 29174 15068 29180
rect 14740 29164 14792 29170
rect 14740 29106 14792 29112
rect 14752 26382 14780 29106
rect 15016 28960 15068 28966
rect 15016 28902 15068 28908
rect 15200 28960 15252 28966
rect 15200 28902 15252 28908
rect 15028 28762 15056 28902
rect 15016 28756 15068 28762
rect 15016 28698 15068 28704
rect 15212 28694 15240 28902
rect 15200 28688 15252 28694
rect 15200 28630 15252 28636
rect 15016 28076 15068 28082
rect 15016 28018 15068 28024
rect 14832 27328 14884 27334
rect 14832 27270 14884 27276
rect 14844 27062 14872 27270
rect 14832 27056 14884 27062
rect 14832 26998 14884 27004
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14832 26376 14884 26382
rect 14832 26318 14884 26324
rect 14740 25968 14792 25974
rect 14740 25910 14792 25916
rect 14752 25430 14780 25910
rect 14740 25424 14792 25430
rect 14740 25366 14792 25372
rect 14648 25288 14700 25294
rect 14462 25256 14518 25265
rect 14648 25230 14700 25236
rect 14462 25191 14464 25200
rect 14516 25191 14518 25200
rect 14464 25162 14516 25168
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14740 24336 14792 24342
rect 14740 24278 14792 24284
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 13832 22066 13952 22094
rect 13832 21622 13860 22066
rect 14292 22030 14320 22646
rect 14752 22098 14780 24278
rect 14844 24206 14872 26318
rect 14936 26314 14964 26726
rect 14924 26308 14976 26314
rect 14924 26250 14976 26256
rect 14936 25226 14964 26250
rect 15028 25294 15056 28018
rect 15108 27872 15160 27878
rect 15106 27840 15108 27849
rect 15160 27840 15162 27849
rect 15106 27775 15162 27784
rect 15212 27470 15240 28630
rect 15292 28484 15344 28490
rect 15292 28426 15344 28432
rect 15304 27470 15332 28426
rect 15396 28082 15424 29718
rect 15750 29679 15806 29688
rect 15476 29572 15528 29578
rect 15476 29514 15528 29520
rect 15384 28076 15436 28082
rect 15384 28018 15436 28024
rect 15200 27464 15252 27470
rect 15200 27406 15252 27412
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 15290 27024 15346 27033
rect 15290 26959 15346 26968
rect 15200 26852 15252 26858
rect 15200 26794 15252 26800
rect 15212 26518 15240 26794
rect 15304 26790 15332 26959
rect 15384 26920 15436 26926
rect 15384 26862 15436 26868
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15200 26512 15252 26518
rect 15200 26454 15252 26460
rect 15200 26376 15252 26382
rect 15396 26330 15424 26862
rect 15252 26324 15424 26330
rect 15200 26318 15424 26324
rect 15212 26302 15424 26318
rect 15108 25424 15160 25430
rect 15108 25366 15160 25372
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 14924 25220 14976 25226
rect 14924 25162 14976 25168
rect 15120 24954 15148 25366
rect 15200 25356 15252 25362
rect 15200 25298 15252 25304
rect 15212 24993 15240 25298
rect 15396 25294 15424 26302
rect 15488 25498 15516 29514
rect 15568 29164 15620 29170
rect 15568 29106 15620 29112
rect 15580 28150 15608 29106
rect 15568 28144 15620 28150
rect 15568 28086 15620 28092
rect 15568 27532 15620 27538
rect 15568 27474 15620 27480
rect 15580 26790 15608 27474
rect 15660 27464 15712 27470
rect 15764 27441 15792 29679
rect 15660 27406 15712 27412
rect 15750 27432 15806 27441
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15568 26512 15620 26518
rect 15568 26454 15620 26460
rect 15580 26382 15608 26454
rect 15672 26450 15700 27406
rect 15750 27367 15806 27376
rect 15856 27305 15884 29838
rect 15948 29646 15976 29990
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 16040 29646 16068 29786
rect 15936 29640 15988 29646
rect 15936 29582 15988 29588
rect 16028 29640 16080 29646
rect 16028 29582 16080 29588
rect 16040 29170 16068 29582
rect 16028 29164 16080 29170
rect 16028 29106 16080 29112
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 15948 28558 15976 28902
rect 15936 28552 15988 28558
rect 15936 28494 15988 28500
rect 16040 28082 16068 29106
rect 16132 28937 16160 31078
rect 16212 30252 16264 30258
rect 16212 30194 16264 30200
rect 16224 29850 16252 30194
rect 16212 29844 16264 29850
rect 16212 29786 16264 29792
rect 16118 28928 16174 28937
rect 16118 28863 16174 28872
rect 16118 28520 16174 28529
rect 16118 28455 16120 28464
rect 16172 28455 16174 28464
rect 16120 28426 16172 28432
rect 16028 28076 16080 28082
rect 16028 28018 16080 28024
rect 15936 27872 15988 27878
rect 15936 27814 15988 27820
rect 15948 27470 15976 27814
rect 15936 27464 15988 27470
rect 15936 27406 15988 27412
rect 15842 27296 15898 27305
rect 15842 27231 15898 27240
rect 16040 26926 16068 28018
rect 16028 26920 16080 26926
rect 16028 26862 16080 26868
rect 16120 26784 16172 26790
rect 16120 26726 16172 26732
rect 15660 26444 15712 26450
rect 15660 26386 15712 26392
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15844 26036 15896 26042
rect 15844 25978 15896 25984
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15580 25498 15608 25842
rect 15476 25492 15528 25498
rect 15476 25434 15528 25440
rect 15568 25492 15620 25498
rect 15568 25434 15620 25440
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 15198 24984 15254 24993
rect 15108 24948 15160 24954
rect 15198 24919 15254 24928
rect 15108 24890 15160 24896
rect 15016 24676 15068 24682
rect 15016 24618 15068 24624
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 15028 24138 15056 24618
rect 15304 24410 15332 25094
rect 15856 24682 15884 25978
rect 15844 24676 15896 24682
rect 15844 24618 15896 24624
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15660 24200 15712 24206
rect 15660 24142 15712 24148
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 15028 23322 15056 24074
rect 15672 23730 15700 24142
rect 15936 24132 15988 24138
rect 15936 24074 15988 24080
rect 15948 23866 15976 24074
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 16132 23798 16160 26726
rect 16212 25696 16264 25702
rect 16212 25638 16264 25644
rect 16224 25362 16252 25638
rect 16212 25356 16264 25362
rect 16212 25298 16264 25304
rect 16316 24954 16344 31198
rect 16500 30977 16528 33050
rect 16592 32881 16620 37216
rect 16856 35012 16908 35018
rect 16856 34954 16908 34960
rect 16868 34610 16896 34954
rect 16856 34604 16908 34610
rect 16856 34546 16908 34552
rect 16672 33992 16724 33998
rect 16672 33934 16724 33940
rect 16578 32872 16634 32881
rect 16578 32807 16634 32816
rect 16580 31952 16632 31958
rect 16578 31920 16580 31929
rect 16632 31920 16634 31929
rect 16578 31855 16634 31864
rect 16684 31754 16712 33934
rect 16960 33862 16988 38762
rect 17960 38480 18012 38486
rect 17960 38422 18012 38428
rect 17040 37256 17092 37262
rect 17040 37198 17092 37204
rect 17222 37224 17278 37233
rect 17052 36281 17080 37198
rect 17222 37159 17278 37168
rect 17316 37188 17368 37194
rect 17132 36780 17184 36786
rect 17132 36722 17184 36728
rect 17038 36272 17094 36281
rect 17038 36207 17094 36216
rect 17144 36174 17172 36722
rect 17236 36689 17264 37159
rect 17316 37130 17368 37136
rect 17222 36680 17278 36689
rect 17222 36615 17278 36624
rect 17132 36168 17184 36174
rect 17328 36145 17356 37130
rect 17406 36680 17462 36689
rect 17406 36615 17462 36624
rect 17420 36582 17448 36615
rect 17408 36576 17460 36582
rect 17408 36518 17460 36524
rect 17776 36576 17828 36582
rect 17776 36518 17828 36524
rect 17132 36110 17184 36116
rect 17314 36136 17370 36145
rect 17314 36071 17370 36080
rect 17316 36032 17368 36038
rect 17316 35974 17368 35980
rect 17328 35834 17356 35974
rect 17316 35828 17368 35834
rect 17316 35770 17368 35776
rect 17040 35556 17092 35562
rect 17040 35498 17092 35504
rect 16856 33856 16908 33862
rect 16856 33798 16908 33804
rect 16948 33856 17000 33862
rect 16948 33798 17000 33804
rect 16868 33289 16896 33798
rect 16960 33658 16988 33798
rect 16948 33652 17000 33658
rect 16948 33594 17000 33600
rect 16948 33448 17000 33454
rect 16948 33390 17000 33396
rect 16854 33280 16910 33289
rect 16854 33215 16910 33224
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 16868 32745 16896 32846
rect 16854 32736 16910 32745
rect 16854 32671 16910 32680
rect 16960 32434 16988 33390
rect 16948 32428 17000 32434
rect 16948 32370 17000 32376
rect 16856 32020 16908 32026
rect 16856 31962 16908 31968
rect 16868 31754 16896 31962
rect 16592 31726 16712 31754
rect 16776 31726 16896 31754
rect 16592 31210 16620 31726
rect 16580 31204 16632 31210
rect 16580 31146 16632 31152
rect 16486 30968 16542 30977
rect 16486 30903 16542 30912
rect 16488 30660 16540 30666
rect 16488 30602 16540 30608
rect 16396 30252 16448 30258
rect 16396 30194 16448 30200
rect 16408 29578 16436 30194
rect 16500 30122 16528 30602
rect 16488 30116 16540 30122
rect 16488 30058 16540 30064
rect 16486 30016 16542 30025
rect 16486 29951 16542 29960
rect 16500 29850 16528 29951
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16592 29730 16620 31146
rect 16670 30968 16726 30977
rect 16670 30903 16726 30912
rect 16500 29702 16620 29730
rect 16396 29572 16448 29578
rect 16396 29514 16448 29520
rect 16396 28960 16448 28966
rect 16396 28902 16448 28908
rect 16304 24948 16356 24954
rect 16304 24890 16356 24896
rect 16212 24812 16264 24818
rect 16212 24754 16264 24760
rect 16224 24410 16252 24754
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 16120 23792 16172 23798
rect 16120 23734 16172 23740
rect 16408 23730 16436 28902
rect 16500 27470 16528 29702
rect 16684 28966 16712 30903
rect 16672 28960 16724 28966
rect 16672 28902 16724 28908
rect 16578 28656 16634 28665
rect 16578 28591 16634 28600
rect 16592 28422 16620 28591
rect 16580 28416 16632 28422
rect 16580 28358 16632 28364
rect 16776 28257 16804 31726
rect 17052 31686 17080 35498
rect 17132 35148 17184 35154
rect 17132 35090 17184 35096
rect 17144 34746 17172 35090
rect 17328 35086 17356 35770
rect 17408 35148 17460 35154
rect 17408 35090 17460 35096
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 17420 34921 17448 35090
rect 17406 34912 17462 34921
rect 17406 34847 17462 34856
rect 17314 34776 17370 34785
rect 17132 34740 17184 34746
rect 17314 34711 17370 34720
rect 17132 34682 17184 34688
rect 17224 33108 17276 33114
rect 17224 33050 17276 33056
rect 17236 32586 17264 33050
rect 17328 33046 17356 34711
rect 17420 33658 17448 34847
rect 17788 34762 17816 36518
rect 17972 35714 18000 38422
rect 18156 38350 18184 38762
rect 18236 38480 18288 38486
rect 18236 38422 18288 38428
rect 18144 38344 18196 38350
rect 18144 38286 18196 38292
rect 18052 36032 18104 36038
rect 18050 36000 18052 36009
rect 18104 36000 18106 36009
rect 18050 35935 18106 35944
rect 17972 35686 18092 35714
rect 17960 35624 18012 35630
rect 17958 35592 17960 35601
rect 18012 35592 18014 35601
rect 17958 35527 18014 35536
rect 17972 35018 18000 35527
rect 17960 35012 18012 35018
rect 17960 34954 18012 34960
rect 17604 34734 17816 34762
rect 17500 34604 17552 34610
rect 17500 34546 17552 34552
rect 17512 34134 17540 34546
rect 17500 34128 17552 34134
rect 17500 34070 17552 34076
rect 17408 33652 17460 33658
rect 17408 33594 17460 33600
rect 17408 33380 17460 33386
rect 17408 33322 17460 33328
rect 17316 33040 17368 33046
rect 17316 32982 17368 32988
rect 17236 32558 17356 32586
rect 17132 32428 17184 32434
rect 17132 32370 17184 32376
rect 17144 31754 17172 32370
rect 17144 31726 17264 31754
rect 17040 31680 17092 31686
rect 17040 31622 17092 31628
rect 17132 31680 17184 31686
rect 17132 31622 17184 31628
rect 17144 31346 17172 31622
rect 16856 31340 16908 31346
rect 17132 31340 17184 31346
rect 16908 31300 16988 31328
rect 16856 31282 16908 31288
rect 16856 31204 16908 31210
rect 16856 31146 16908 31152
rect 16868 29510 16896 31146
rect 16960 30666 16988 31300
rect 17132 31282 17184 31288
rect 17236 31142 17264 31726
rect 17224 31136 17276 31142
rect 17224 31078 17276 31084
rect 16948 30660 17000 30666
rect 16948 30602 17000 30608
rect 17328 30376 17356 32558
rect 17420 31754 17448 33322
rect 17512 32434 17540 34070
rect 17604 33930 17632 34734
rect 17684 34604 17736 34610
rect 17684 34546 17736 34552
rect 17960 34604 18012 34610
rect 17960 34546 18012 34552
rect 17592 33924 17644 33930
rect 17592 33866 17644 33872
rect 17604 33658 17632 33866
rect 17592 33652 17644 33658
rect 17592 33594 17644 33600
rect 17592 33516 17644 33522
rect 17592 33458 17644 33464
rect 17500 32428 17552 32434
rect 17500 32370 17552 32376
rect 17500 32020 17552 32026
rect 17500 31962 17552 31968
rect 17512 31890 17540 31962
rect 17500 31884 17552 31890
rect 17500 31826 17552 31832
rect 17604 31754 17632 33458
rect 17696 33454 17724 34546
rect 17776 34536 17828 34542
rect 17776 34478 17828 34484
rect 17684 33448 17736 33454
rect 17684 33390 17736 33396
rect 17788 33318 17816 34478
rect 17972 34406 18000 34546
rect 17960 34400 18012 34406
rect 17960 34342 18012 34348
rect 17866 34096 17922 34105
rect 17866 34031 17922 34040
rect 17880 33980 17908 34031
rect 17960 33992 18012 33998
rect 17880 33952 17960 33980
rect 17960 33934 18012 33940
rect 17868 33652 17920 33658
rect 17868 33594 17920 33600
rect 17776 33312 17828 33318
rect 17776 33254 17828 33260
rect 17880 33114 17908 33594
rect 17972 33318 18000 33934
rect 17960 33312 18012 33318
rect 17960 33254 18012 33260
rect 17868 33108 17920 33114
rect 17868 33050 17920 33056
rect 17684 33040 17736 33046
rect 17684 32982 17736 32988
rect 17408 31748 17460 31754
rect 17408 31690 17460 31696
rect 17512 31726 17632 31754
rect 17420 31346 17448 31690
rect 17408 31340 17460 31346
rect 17408 31282 17460 31288
rect 17144 30348 17356 30376
rect 17040 30252 17092 30258
rect 17040 30194 17092 30200
rect 17052 29782 17080 30194
rect 17040 29776 17092 29782
rect 17144 29753 17172 30348
rect 17224 30252 17276 30258
rect 17224 30194 17276 30200
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 17040 29718 17092 29724
rect 17130 29744 17186 29753
rect 17130 29679 17186 29688
rect 16948 29640 17000 29646
rect 16948 29582 17000 29588
rect 16856 29504 16908 29510
rect 16856 29446 16908 29452
rect 16868 29170 16896 29446
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16762 28248 16818 28257
rect 16762 28183 16818 28192
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 16868 27946 16896 28018
rect 16856 27940 16908 27946
rect 16856 27882 16908 27888
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16868 26518 16896 27882
rect 16960 26994 16988 29582
rect 17040 29232 17092 29238
rect 17040 29174 17092 29180
rect 17052 28694 17080 29174
rect 17132 29164 17184 29170
rect 17132 29106 17184 29112
rect 17040 28688 17092 28694
rect 17040 28630 17092 28636
rect 17144 28150 17172 29106
rect 17236 29102 17264 30194
rect 17328 29646 17356 30194
rect 17316 29640 17368 29646
rect 17316 29582 17368 29588
rect 17420 29209 17448 31282
rect 17406 29200 17462 29209
rect 17406 29135 17462 29144
rect 17224 29096 17276 29102
rect 17224 29038 17276 29044
rect 17420 28914 17448 29135
rect 17236 28886 17448 28914
rect 17132 28144 17184 28150
rect 17132 28086 17184 28092
rect 17144 27606 17172 28086
rect 17132 27600 17184 27606
rect 17132 27542 17184 27548
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16856 26512 16908 26518
rect 16856 26454 16908 26460
rect 16580 26308 16632 26314
rect 16580 26250 16632 26256
rect 16488 26240 16540 26246
rect 16488 26182 16540 26188
rect 16500 26042 16528 26182
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 16592 25498 16620 26250
rect 17236 26246 17264 28886
rect 17512 28506 17540 31726
rect 17592 31408 17644 31414
rect 17592 31350 17644 31356
rect 17604 30938 17632 31350
rect 17592 30932 17644 30938
rect 17592 30874 17644 30880
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17604 30326 17632 30534
rect 17592 30320 17644 30326
rect 17592 30262 17644 30268
rect 17604 29578 17632 30262
rect 17592 29572 17644 29578
rect 17592 29514 17644 29520
rect 17696 28966 17724 32982
rect 17866 32600 17922 32609
rect 17866 32535 17922 32544
rect 17776 32428 17828 32434
rect 17776 32370 17828 32376
rect 17788 31822 17816 32370
rect 17880 32314 17908 32535
rect 17960 32496 18012 32502
rect 18064 32484 18092 35686
rect 18144 35284 18196 35290
rect 18144 35226 18196 35232
rect 18012 32456 18092 32484
rect 17960 32438 18012 32444
rect 17880 32286 18000 32314
rect 18064 32298 18092 32456
rect 17868 32224 17920 32230
rect 17868 32166 17920 32172
rect 17776 31816 17828 31822
rect 17776 31758 17828 31764
rect 17776 31680 17828 31686
rect 17776 31622 17828 31628
rect 17788 29306 17816 31622
rect 17880 31521 17908 32166
rect 17972 31958 18000 32286
rect 18052 32292 18104 32298
rect 18052 32234 18104 32240
rect 17960 31952 18012 31958
rect 17960 31894 18012 31900
rect 18052 31680 18104 31686
rect 18156 31668 18184 35226
rect 18248 34921 18276 38422
rect 18340 37262 18368 39200
rect 21652 39166 21680 39200
rect 21640 39160 21692 39166
rect 21640 39102 21692 39108
rect 22100 39160 22152 39166
rect 22100 39102 22152 39108
rect 18604 38956 18656 38962
rect 18604 38898 18656 38904
rect 18328 37256 18380 37262
rect 18328 37198 18380 37204
rect 18616 36854 18644 38898
rect 20168 38820 20220 38826
rect 20168 38762 20220 38768
rect 19430 37360 19486 37369
rect 19430 37295 19486 37304
rect 20076 37324 20128 37330
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 18788 37188 18840 37194
rect 18788 37130 18840 37136
rect 18512 36848 18564 36854
rect 18512 36790 18564 36796
rect 18604 36848 18656 36854
rect 18604 36790 18656 36796
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 18432 36310 18460 36722
rect 18420 36304 18472 36310
rect 18420 36246 18472 36252
rect 18524 36174 18552 36790
rect 18604 36576 18656 36582
rect 18604 36518 18656 36524
rect 18616 36242 18644 36518
rect 18604 36236 18656 36242
rect 18604 36178 18656 36184
rect 18420 36168 18472 36174
rect 18420 36110 18472 36116
rect 18512 36168 18564 36174
rect 18512 36110 18564 36116
rect 18328 35692 18380 35698
rect 18432 35680 18460 36110
rect 18380 35652 18460 35680
rect 18328 35634 18380 35640
rect 18432 35494 18460 35652
rect 18524 35630 18552 36110
rect 18604 36100 18656 36106
rect 18604 36042 18656 36048
rect 18512 35624 18564 35630
rect 18512 35566 18564 35572
rect 18420 35488 18472 35494
rect 18420 35430 18472 35436
rect 18328 35080 18380 35086
rect 18328 35022 18380 35028
rect 18234 34912 18290 34921
rect 18234 34847 18290 34856
rect 18340 34474 18368 35022
rect 18328 34468 18380 34474
rect 18328 34410 18380 34416
rect 18236 34060 18288 34066
rect 18236 34002 18288 34008
rect 18248 33153 18276 34002
rect 18234 33144 18290 33153
rect 18234 33079 18290 33088
rect 18340 32960 18368 34410
rect 18418 33688 18474 33697
rect 18418 33623 18474 33632
rect 18432 33522 18460 33623
rect 18420 33516 18472 33522
rect 18420 33458 18472 33464
rect 18432 33046 18460 33458
rect 18420 33040 18472 33046
rect 18420 32982 18472 32988
rect 18248 32932 18368 32960
rect 18248 32609 18276 32932
rect 18328 32836 18380 32842
rect 18328 32778 18380 32784
rect 18420 32836 18472 32842
rect 18420 32778 18472 32784
rect 18234 32600 18290 32609
rect 18234 32535 18290 32544
rect 18248 32434 18276 32535
rect 18340 32502 18368 32778
rect 18432 32745 18460 32778
rect 18418 32736 18474 32745
rect 18418 32671 18474 32680
rect 18328 32496 18380 32502
rect 18328 32438 18380 32444
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 18236 32224 18288 32230
rect 18236 32166 18288 32172
rect 18104 31640 18184 31668
rect 18052 31622 18104 31628
rect 17866 31512 17922 31521
rect 17866 31447 17922 31456
rect 18248 31414 18276 32166
rect 18236 31408 18288 31414
rect 18236 31350 18288 31356
rect 18144 31136 18196 31142
rect 18144 31078 18196 31084
rect 18052 30864 18104 30870
rect 18052 30806 18104 30812
rect 17960 30660 18012 30666
rect 17960 30602 18012 30608
rect 17972 29646 18000 30602
rect 18064 30433 18092 30806
rect 18156 30734 18184 31078
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 18340 30666 18368 32438
rect 18420 31952 18472 31958
rect 18420 31894 18472 31900
rect 18328 30660 18380 30666
rect 18328 30602 18380 30608
rect 18050 30424 18106 30433
rect 18050 30359 18106 30368
rect 18432 30190 18460 31894
rect 18524 31142 18552 35566
rect 18616 32201 18644 36042
rect 18800 35601 18828 37130
rect 18880 36780 18932 36786
rect 18880 36722 18932 36728
rect 19156 36780 19208 36786
rect 19156 36722 19208 36728
rect 18786 35592 18842 35601
rect 18786 35527 18842 35536
rect 18696 35148 18748 35154
rect 18696 35090 18748 35096
rect 18602 32192 18658 32201
rect 18602 32127 18658 32136
rect 18604 31816 18656 31822
rect 18604 31758 18656 31764
rect 18512 31136 18564 31142
rect 18512 31078 18564 31084
rect 18512 30660 18564 30666
rect 18512 30602 18564 30608
rect 18328 30184 18380 30190
rect 18328 30126 18380 30132
rect 18420 30184 18472 30190
rect 18420 30126 18472 30132
rect 17960 29640 18012 29646
rect 17960 29582 18012 29588
rect 18050 29472 18106 29481
rect 18050 29407 18106 29416
rect 17776 29300 17828 29306
rect 17776 29242 17828 29248
rect 17684 28960 17736 28966
rect 17684 28902 17736 28908
rect 17684 28688 17736 28694
rect 17684 28630 17736 28636
rect 17420 28478 17540 28506
rect 17316 28076 17368 28082
rect 17420 28064 17448 28478
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17368 28036 17448 28064
rect 17316 28018 17368 28024
rect 17224 26240 17276 26246
rect 17224 26182 17276 26188
rect 17328 26058 17356 28018
rect 17406 27024 17462 27033
rect 17512 26994 17540 28358
rect 17604 26994 17632 28358
rect 17696 28014 17724 28630
rect 17868 28552 17920 28558
rect 17868 28494 17920 28500
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 17880 27674 17908 28494
rect 17868 27668 17920 27674
rect 17868 27610 17920 27616
rect 17866 27568 17922 27577
rect 17866 27503 17922 27512
rect 17682 27432 17738 27441
rect 17682 27367 17738 27376
rect 17406 26959 17462 26968
rect 17500 26988 17552 26994
rect 17420 26450 17448 26959
rect 17500 26930 17552 26936
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17408 26444 17460 26450
rect 17408 26386 17460 26392
rect 17236 26030 17356 26058
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 17052 25498 17080 25842
rect 16580 25492 16632 25498
rect 16580 25434 16632 25440
rect 17040 25492 17092 25498
rect 17040 25434 17092 25440
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 16856 25288 16908 25294
rect 16856 25230 16908 25236
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 16592 24206 16620 25230
rect 16868 24818 16896 25230
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16764 24608 16816 24614
rect 16764 24550 16816 24556
rect 16580 24200 16632 24206
rect 16580 24142 16632 24148
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 16396 23724 16448 23730
rect 16396 23666 16448 23672
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15120 22778 15148 23054
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15304 22098 15332 22578
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14832 22024 14884 22030
rect 14832 21966 14884 21972
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 14292 21622 14320 21966
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13084 21412 13136 21418
rect 13084 21354 13136 21360
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 11256 19854 11284 20878
rect 12438 20632 12494 20641
rect 12438 20567 12440 20576
rect 12492 20567 12494 20576
rect 12440 20538 12492 20544
rect 12348 20324 12400 20330
rect 12348 20266 12400 20272
rect 12360 19854 12388 20266
rect 12636 20058 12664 20878
rect 13464 20398 13492 21422
rect 13648 21146 13676 21490
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13268 20392 13320 20398
rect 13268 20334 13320 20340
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13280 20058 13308 20334
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12360 19378 12388 19790
rect 13832 19514 13860 21558
rect 14844 21554 14872 21966
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 15212 21026 15240 21966
rect 15120 20998 15240 21026
rect 15292 21004 15344 21010
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 14002 20632 14058 20641
rect 15028 20602 15056 20878
rect 15120 20602 15148 20998
rect 15292 20946 15344 20952
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 14002 20567 14058 20576
rect 15016 20596 15068 20602
rect 14016 20330 14044 20567
rect 15016 20538 15068 20544
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15028 20398 15056 20538
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 14004 20324 14056 20330
rect 14004 20266 14056 20272
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 14476 19310 14504 19722
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 13556 18970 13584 19178
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 12912 18358 12940 18702
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 14108 18290 14136 18770
rect 14384 18426 14412 19246
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18766 14504 19110
rect 14660 18766 14688 20198
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14752 19854 14780 19994
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14924 19848 14976 19854
rect 15028 19836 15056 20334
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 15120 19854 15148 20198
rect 14976 19808 15056 19836
rect 15108 19848 15160 19854
rect 14924 19790 14976 19796
rect 15108 19790 15160 19796
rect 14752 19514 14780 19790
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14752 18902 14780 19450
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14844 18902 14872 19314
rect 15212 19310 15240 20878
rect 15304 20466 15332 20946
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15304 19922 15332 20198
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 15396 19310 15424 22034
rect 15488 21010 15516 23054
rect 16592 22642 16620 24142
rect 16672 23588 16724 23594
rect 16672 23530 16724 23536
rect 16684 22982 16712 23530
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16776 22710 16804 24550
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16868 23050 16896 24006
rect 16856 23044 16908 23050
rect 16856 22986 16908 22992
rect 16764 22704 16816 22710
rect 16764 22646 16816 22652
rect 16212 22636 16264 22642
rect 16212 22578 16264 22584
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15844 22568 15896 22574
rect 15844 22510 15896 22516
rect 15580 22030 15608 22510
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15856 21690 15884 22510
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15580 21350 15608 21490
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15580 20398 15608 20810
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15488 20058 15516 20334
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15672 19854 15700 21422
rect 16224 20602 16252 22578
rect 16212 20596 16264 20602
rect 16212 20538 16264 20544
rect 15752 20528 15804 20534
rect 15752 20470 15804 20476
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15764 19786 15792 20470
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16040 19990 16068 20198
rect 16028 19984 16080 19990
rect 16028 19926 16080 19932
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 16500 19718 16528 22578
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16592 20058 16620 20402
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 15936 19712 15988 19718
rect 15936 19654 15988 19660
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 14832 18896 14884 18902
rect 14832 18838 14884 18844
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3882 17096 3938 17105
rect 3882 17031 3938 17040
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 14752 15609 14780 18566
rect 14844 18290 14872 18838
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 15028 18630 15056 18702
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 15028 18222 15056 18566
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 15028 17882 15056 18158
rect 15016 17876 15068 17882
rect 15016 17818 15068 17824
rect 15212 17338 15240 19246
rect 15396 18426 15424 19246
rect 15948 19174 15976 19654
rect 16592 19378 16620 19994
rect 16684 19854 16712 22374
rect 16960 22094 16988 25230
rect 17236 24154 17264 26030
rect 17592 25764 17644 25770
rect 17696 25752 17724 27367
rect 17880 26382 17908 27503
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17972 27033 18000 27406
rect 18064 27334 18092 29407
rect 18144 28620 18196 28626
rect 18144 28562 18196 28568
rect 18052 27328 18104 27334
rect 18052 27270 18104 27276
rect 18156 27130 18184 28562
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18248 27470 18276 28494
rect 18340 28082 18368 30126
rect 18524 29170 18552 30602
rect 18616 29782 18644 31758
rect 18604 29776 18656 29782
rect 18604 29718 18656 29724
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 18328 28076 18380 28082
rect 18328 28018 18380 28024
rect 18328 27872 18380 27878
rect 18328 27814 18380 27820
rect 18420 27872 18472 27878
rect 18420 27814 18472 27820
rect 18340 27538 18368 27814
rect 18432 27538 18460 27814
rect 18328 27532 18380 27538
rect 18328 27474 18380 27480
rect 18420 27532 18472 27538
rect 18420 27474 18472 27480
rect 18236 27464 18288 27470
rect 18432 27418 18460 27474
rect 18236 27406 18288 27412
rect 18144 27124 18196 27130
rect 18144 27066 18196 27072
rect 17958 27024 18014 27033
rect 17958 26959 18014 26968
rect 18248 26790 18276 27406
rect 18340 27390 18460 27418
rect 18236 26784 18288 26790
rect 18050 26752 18106 26761
rect 18236 26726 18288 26732
rect 18050 26687 18106 26696
rect 18064 26450 18092 26687
rect 18052 26444 18104 26450
rect 18052 26386 18104 26392
rect 18248 26382 18276 26726
rect 17776 26376 17828 26382
rect 17776 26318 17828 26324
rect 17868 26376 17920 26382
rect 18236 26376 18288 26382
rect 17868 26318 17920 26324
rect 17958 26344 18014 26353
rect 17644 25724 17724 25752
rect 17592 25706 17644 25712
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17316 24948 17368 24954
rect 17316 24890 17368 24896
rect 17328 24818 17356 24890
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17328 24274 17356 24550
rect 17420 24274 17448 25638
rect 17592 25356 17644 25362
rect 17592 25298 17644 25304
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 17512 24954 17540 25094
rect 17500 24948 17552 24954
rect 17500 24890 17552 24896
rect 17316 24268 17368 24274
rect 17316 24210 17368 24216
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 17236 24126 17448 24154
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 16868 22066 16988 22094
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 16776 21486 16804 21898
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16684 19446 16712 19790
rect 16672 19440 16724 19446
rect 16672 19382 16724 19388
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16776 19242 16804 21014
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16224 18834 16252 19110
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 15488 18698 15516 18770
rect 16776 18766 16804 19178
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 16040 18358 16068 18566
rect 16028 18352 16080 18358
rect 16028 18294 16080 18300
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15396 17678 15424 17818
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15844 17604 15896 17610
rect 15844 17546 15896 17552
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15488 17270 15516 17478
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 15856 17202 15884 17546
rect 15948 17202 15976 17818
rect 16040 17746 16068 18294
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 16224 17542 16252 18226
rect 16316 17882 16344 18226
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 15016 17060 15068 17066
rect 15016 17002 15068 17008
rect 15028 16794 15056 17002
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 15856 16726 15884 17138
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 16040 16590 16068 17070
rect 16132 16590 16160 17138
rect 16224 16794 16252 17478
rect 16316 17202 16344 17478
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16500 16674 16528 17818
rect 16868 16946 16896 22066
rect 17052 20602 17080 23666
rect 17144 22982 17172 24006
rect 17316 23724 17368 23730
rect 17316 23666 17368 23672
rect 17224 23520 17276 23526
rect 17328 23497 17356 23666
rect 17224 23462 17276 23468
rect 17314 23488 17370 23497
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 17236 22098 17264 23462
rect 17314 23423 17370 23432
rect 17316 23316 17368 23322
rect 17316 23258 17368 23264
rect 17328 22574 17356 23258
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 17328 22234 17356 22510
rect 17420 22506 17448 24126
rect 17604 22658 17632 25298
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17696 23769 17724 24754
rect 17788 24449 17816 26318
rect 18236 26318 18288 26324
rect 17958 26279 18014 26288
rect 17868 26240 17920 26246
rect 17868 26182 17920 26188
rect 17880 25906 17908 26182
rect 17972 25974 18000 26279
rect 17960 25968 18012 25974
rect 17960 25910 18012 25916
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 17880 25140 17908 25842
rect 17880 25112 18092 25140
rect 18064 24721 18092 25112
rect 18340 24750 18368 27390
rect 18524 27282 18552 29106
rect 18604 29028 18656 29034
rect 18604 28970 18656 28976
rect 18432 27254 18552 27282
rect 18432 25922 18460 27254
rect 18616 26994 18644 28970
rect 18708 27878 18736 35090
rect 18892 34134 18920 36722
rect 18972 36576 19024 36582
rect 18970 36544 18972 36553
rect 19024 36544 19026 36553
rect 18970 36479 19026 36488
rect 18972 36100 19024 36106
rect 18972 36042 19024 36048
rect 18984 36009 19012 36042
rect 18970 36000 19026 36009
rect 18970 35935 19026 35944
rect 19168 35834 19196 36722
rect 19260 36582 19288 37198
rect 19338 36952 19394 36961
rect 19338 36887 19394 36896
rect 19248 36576 19300 36582
rect 19248 36518 19300 36524
rect 19260 36174 19288 36518
rect 19352 36281 19380 36887
rect 19338 36272 19394 36281
rect 19338 36207 19394 36216
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 19246 35864 19302 35873
rect 19156 35828 19208 35834
rect 19246 35799 19248 35808
rect 19156 35770 19208 35776
rect 19300 35799 19302 35808
rect 19248 35770 19300 35776
rect 19444 35748 19472 37295
rect 20076 37266 20128 37272
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19984 36712 20036 36718
rect 19984 36654 20036 36660
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19444 35720 19656 35748
rect 19628 35562 19656 35720
rect 19616 35556 19668 35562
rect 19616 35498 19668 35504
rect 19628 35086 19656 35498
rect 19996 35222 20024 36654
rect 19984 35216 20036 35222
rect 19984 35158 20036 35164
rect 19616 35080 19668 35086
rect 19616 35022 19668 35028
rect 19984 35080 20036 35086
rect 19984 35022 20036 35028
rect 19340 35012 19392 35018
rect 19340 34954 19392 34960
rect 19432 35012 19484 35018
rect 19432 34954 19484 34960
rect 19352 34474 19380 34954
rect 19340 34468 19392 34474
rect 19340 34410 19392 34416
rect 18880 34128 18932 34134
rect 19444 34105 19472 34954
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19892 34740 19944 34746
rect 19892 34682 19944 34688
rect 19904 34626 19932 34682
rect 19996 34626 20024 35022
rect 20088 34746 20116 37266
rect 20180 36417 20208 38762
rect 20904 38140 20956 38146
rect 20904 38082 20956 38088
rect 20720 37664 20772 37670
rect 20720 37606 20772 37612
rect 20534 37360 20590 37369
rect 20534 37295 20590 37304
rect 20166 36408 20222 36417
rect 20166 36343 20222 36352
rect 20444 36304 20496 36310
rect 20444 36246 20496 36252
rect 20168 36168 20220 36174
rect 20168 36110 20220 36116
rect 20076 34740 20128 34746
rect 20076 34682 20128 34688
rect 19616 34604 19668 34610
rect 19616 34546 19668 34552
rect 19708 34604 19760 34610
rect 19904 34598 20024 34626
rect 19708 34546 19760 34552
rect 19628 34513 19656 34546
rect 19614 34504 19670 34513
rect 19614 34439 19670 34448
rect 19720 34134 19748 34546
rect 19708 34128 19760 34134
rect 18880 34070 18932 34076
rect 19430 34096 19486 34105
rect 18892 33998 18920 34070
rect 19708 34070 19760 34076
rect 19430 34031 19486 34040
rect 19524 34060 19576 34066
rect 19524 34002 19576 34008
rect 18880 33992 18932 33998
rect 18880 33934 18932 33940
rect 18788 33856 18840 33862
rect 18788 33798 18840 33804
rect 18880 33856 18932 33862
rect 19536 33844 19564 34002
rect 19982 33960 20038 33969
rect 19982 33895 20038 33904
rect 18880 33798 18932 33804
rect 19352 33816 19564 33844
rect 18800 32230 18828 33798
rect 18892 33658 18920 33798
rect 18880 33652 18932 33658
rect 18880 33594 18932 33600
rect 18880 33312 18932 33318
rect 18880 33254 18932 33260
rect 18892 32978 18920 33254
rect 18972 33108 19024 33114
rect 18972 33050 19024 33056
rect 18880 32972 18932 32978
rect 18880 32914 18932 32920
rect 18880 32292 18932 32298
rect 18880 32234 18932 32240
rect 18788 32224 18840 32230
rect 18788 32166 18840 32172
rect 18788 32020 18840 32026
rect 18788 31962 18840 31968
rect 18800 31657 18828 31962
rect 18892 31958 18920 32234
rect 18880 31952 18932 31958
rect 18880 31894 18932 31900
rect 18880 31680 18932 31686
rect 18786 31648 18842 31657
rect 18880 31622 18932 31628
rect 18786 31583 18842 31592
rect 18892 31521 18920 31622
rect 18878 31512 18934 31521
rect 18878 31447 18934 31456
rect 18984 30569 19012 33050
rect 19064 32768 19116 32774
rect 19064 32710 19116 32716
rect 19156 32768 19208 32774
rect 19156 32710 19208 32716
rect 19076 31142 19104 32710
rect 19168 32570 19196 32710
rect 19156 32564 19208 32570
rect 19156 32506 19208 32512
rect 19352 32366 19380 33816
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19432 33448 19484 33454
rect 19432 33390 19484 33396
rect 19444 32910 19472 33390
rect 19996 33114 20024 33895
rect 20074 33688 20130 33697
rect 20074 33623 20130 33632
rect 20088 33590 20116 33623
rect 20076 33584 20128 33590
rect 20076 33526 20128 33532
rect 19984 33108 20036 33114
rect 19984 33050 20036 33056
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19444 32570 19472 32846
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19432 32564 19484 32570
rect 19432 32506 19484 32512
rect 19340 32360 19392 32366
rect 19340 32302 19392 32308
rect 19248 32224 19300 32230
rect 19248 32166 19300 32172
rect 19340 32224 19392 32230
rect 19340 32166 19392 32172
rect 19064 31136 19116 31142
rect 19064 31078 19116 31084
rect 18970 30560 19026 30569
rect 18970 30495 19026 30504
rect 18786 30152 18842 30161
rect 18786 30087 18842 30096
rect 18800 28393 18828 30087
rect 19156 29640 19208 29646
rect 19156 29582 19208 29588
rect 18972 29504 19024 29510
rect 18972 29446 19024 29452
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 18892 28558 18920 28698
rect 18880 28552 18932 28558
rect 18880 28494 18932 28500
rect 18786 28384 18842 28393
rect 18786 28319 18842 28328
rect 18880 28008 18932 28014
rect 18880 27950 18932 27956
rect 18696 27872 18748 27878
rect 18696 27814 18748 27820
rect 18696 27328 18748 27334
rect 18696 27270 18748 27276
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 18708 26874 18736 27270
rect 18892 26994 18920 27950
rect 18880 26988 18932 26994
rect 18880 26930 18932 26936
rect 18512 26852 18564 26858
rect 18512 26794 18564 26800
rect 18616 26846 18736 26874
rect 18524 26586 18552 26794
rect 18512 26580 18564 26586
rect 18512 26522 18564 26528
rect 18616 26353 18644 26846
rect 18880 26784 18932 26790
rect 18786 26752 18842 26761
rect 18880 26726 18932 26732
rect 18786 26687 18842 26696
rect 18696 26444 18748 26450
rect 18696 26386 18748 26392
rect 18602 26344 18658 26353
rect 18602 26279 18658 26288
rect 18512 26240 18564 26246
rect 18512 26182 18564 26188
rect 18602 26208 18658 26217
rect 18524 26042 18552 26182
rect 18602 26143 18658 26152
rect 18512 26036 18564 26042
rect 18512 25978 18564 25984
rect 18432 25894 18552 25922
rect 18616 25906 18644 26143
rect 18420 25832 18472 25838
rect 18420 25774 18472 25780
rect 18524 25786 18552 25894
rect 18604 25900 18656 25906
rect 18604 25842 18656 25848
rect 18432 25673 18460 25774
rect 18524 25758 18644 25786
rect 18418 25664 18474 25673
rect 18418 25599 18474 25608
rect 18432 25129 18460 25599
rect 18616 25362 18644 25758
rect 18604 25356 18656 25362
rect 18604 25298 18656 25304
rect 18512 25220 18564 25226
rect 18512 25162 18564 25168
rect 18418 25120 18474 25129
rect 18418 25055 18474 25064
rect 18328 24744 18380 24750
rect 18050 24712 18106 24721
rect 18328 24686 18380 24692
rect 18050 24647 18106 24656
rect 17774 24440 17830 24449
rect 17774 24375 17830 24384
rect 17682 23760 17738 23769
rect 17682 23695 17738 23704
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17788 23050 17816 23462
rect 17767 23044 17819 23050
rect 17767 22986 17819 22992
rect 17868 22976 17920 22982
rect 17868 22918 17920 22924
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 17512 22642 17632 22658
rect 17500 22636 17632 22642
rect 17552 22630 17632 22636
rect 17500 22578 17552 22584
rect 17880 22574 17908 22918
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17408 22500 17460 22506
rect 17408 22442 17460 22448
rect 17316 22228 17368 22234
rect 17316 22170 17368 22176
rect 17880 22166 17908 22510
rect 17972 22506 18000 22918
rect 18064 22545 18092 24647
rect 18420 24200 18472 24206
rect 18524 24188 18552 25162
rect 18616 24206 18644 25298
rect 18708 24410 18736 26386
rect 18800 26042 18828 26687
rect 18788 26036 18840 26042
rect 18788 25978 18840 25984
rect 18892 25922 18920 26726
rect 18800 25894 18920 25922
rect 18800 25294 18828 25894
rect 18788 25288 18840 25294
rect 18788 25230 18840 25236
rect 18800 24886 18828 25230
rect 18788 24880 18840 24886
rect 18788 24822 18840 24828
rect 18696 24404 18748 24410
rect 18696 24346 18748 24352
rect 18472 24160 18552 24188
rect 18604 24200 18656 24206
rect 18420 24142 18472 24148
rect 18604 24142 18656 24148
rect 18420 24064 18472 24070
rect 18472 24024 18644 24052
rect 18420 24006 18472 24012
rect 18616 23594 18644 24024
rect 18604 23588 18656 23594
rect 18604 23530 18656 23536
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18616 22778 18644 22986
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18708 22642 18736 24346
rect 18800 23633 18828 24822
rect 18984 24800 19012 29446
rect 19168 29050 19196 29582
rect 19260 29170 19288 32166
rect 19352 31929 19380 32166
rect 19338 31920 19394 31929
rect 19338 31855 19394 31864
rect 19444 31346 19472 32506
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 19892 32020 19944 32026
rect 19892 31962 19944 31968
rect 19904 31822 19932 31962
rect 19892 31816 19944 31822
rect 19892 31758 19944 31764
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19340 31272 19392 31278
rect 19340 31214 19392 31220
rect 19996 31226 20024 32370
rect 20180 32212 20208 36110
rect 20352 35488 20404 35494
rect 20352 35430 20404 35436
rect 20364 35290 20392 35430
rect 20352 35284 20404 35290
rect 20352 35226 20404 35232
rect 20456 35086 20484 36246
rect 20548 35680 20576 37295
rect 20732 37194 20760 37606
rect 20720 37188 20772 37194
rect 20720 37130 20772 37136
rect 20916 36174 20944 38082
rect 21272 38004 21324 38010
rect 21272 37946 21324 37952
rect 20996 37460 21048 37466
rect 20996 37402 21048 37408
rect 21008 37369 21036 37402
rect 20994 37360 21050 37369
rect 20994 37295 21050 37304
rect 20904 36168 20956 36174
rect 20904 36110 20956 36116
rect 21180 36100 21232 36106
rect 21180 36042 21232 36048
rect 20548 35652 20668 35680
rect 20536 35556 20588 35562
rect 20536 35498 20588 35504
rect 20548 35290 20576 35498
rect 20536 35284 20588 35290
rect 20536 35226 20588 35232
rect 20640 35170 20668 35652
rect 20548 35142 20668 35170
rect 20904 35216 20956 35222
rect 20904 35158 20956 35164
rect 20444 35080 20496 35086
rect 20444 35022 20496 35028
rect 20444 34944 20496 34950
rect 20444 34886 20496 34892
rect 20456 34678 20484 34886
rect 20444 34672 20496 34678
rect 20444 34614 20496 34620
rect 20352 34060 20404 34066
rect 20352 34002 20404 34008
rect 20260 33380 20312 33386
rect 20260 33322 20312 33328
rect 20088 32184 20208 32212
rect 20088 31754 20116 32184
rect 20272 32042 20300 33322
rect 20364 33114 20392 34002
rect 20444 33516 20496 33522
rect 20444 33458 20496 33464
rect 20352 33108 20404 33114
rect 20352 33050 20404 33056
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 20364 32337 20392 32370
rect 20350 32328 20406 32337
rect 20350 32263 20406 32272
rect 20180 32014 20300 32042
rect 20076 31748 20128 31754
rect 20076 31690 20128 31696
rect 19352 30258 19380 31214
rect 19996 31198 20116 31226
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 19352 29578 19380 30194
rect 19708 30048 19760 30054
rect 19708 29990 19760 29996
rect 19720 29782 19748 29990
rect 19708 29776 19760 29782
rect 19708 29718 19760 29724
rect 19340 29572 19392 29578
rect 19340 29514 19392 29520
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 19168 29022 19472 29050
rect 19156 28008 19208 28014
rect 19156 27950 19208 27956
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 19076 26994 19104 27270
rect 19064 26988 19116 26994
rect 19064 26930 19116 26936
rect 19062 26072 19118 26081
rect 19062 26007 19064 26016
rect 19116 26007 19118 26016
rect 19064 25978 19116 25984
rect 19064 25832 19116 25838
rect 19064 25774 19116 25780
rect 19076 25362 19104 25774
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 19064 24812 19116 24818
rect 18984 24772 19064 24800
rect 19064 24754 19116 24760
rect 18880 24404 18932 24410
rect 18880 24346 18932 24352
rect 18892 23866 18920 24346
rect 19062 24304 19118 24313
rect 19062 24239 19118 24248
rect 19076 24206 19104 24239
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18786 23624 18842 23633
rect 18786 23559 18842 23568
rect 18892 23254 18920 23802
rect 18972 23656 19024 23662
rect 18972 23598 19024 23604
rect 18984 23497 19012 23598
rect 18970 23488 19026 23497
rect 18970 23423 19026 23432
rect 19168 23361 19196 27950
rect 19444 27849 19472 29022
rect 19996 28778 20024 31078
rect 20088 29073 20116 31198
rect 20180 30394 20208 32014
rect 20350 31648 20406 31657
rect 20350 31583 20406 31592
rect 20260 31340 20312 31346
rect 20260 31282 20312 31288
rect 20272 30938 20300 31282
rect 20260 30932 20312 30938
rect 20260 30874 20312 30880
rect 20168 30388 20220 30394
rect 20168 30330 20220 30336
rect 20074 29064 20130 29073
rect 20074 28999 20130 29008
rect 20076 28960 20128 28966
rect 20076 28902 20128 28908
rect 20088 28778 20116 28902
rect 19996 28750 20116 28778
rect 19984 28620 20036 28626
rect 19984 28562 20036 28568
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19524 28008 19576 28014
rect 19524 27950 19576 27956
rect 19430 27840 19486 27849
rect 19430 27775 19486 27784
rect 19248 27396 19300 27402
rect 19536 27384 19564 27950
rect 19892 27940 19944 27946
rect 19892 27882 19944 27888
rect 19904 27674 19932 27882
rect 19892 27668 19944 27674
rect 19892 27610 19944 27616
rect 19248 27338 19300 27344
rect 19444 27356 19564 27384
rect 19260 27130 19288 27338
rect 19248 27124 19300 27130
rect 19248 27066 19300 27072
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 19260 25770 19288 26930
rect 19352 26518 19380 26998
rect 19340 26512 19392 26518
rect 19340 26454 19392 26460
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19352 25838 19380 26318
rect 19444 26296 19472 27356
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19892 26920 19944 26926
rect 19892 26862 19944 26868
rect 19904 26314 19932 26862
rect 19424 26268 19472 26296
rect 19892 26308 19944 26314
rect 19424 26058 19452 26268
rect 19892 26250 19944 26256
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19424 26030 19472 26058
rect 19444 25906 19472 26030
rect 19432 25900 19484 25906
rect 19616 25900 19668 25906
rect 19432 25842 19484 25848
rect 19536 25860 19616 25888
rect 19340 25832 19392 25838
rect 19444 25809 19472 25842
rect 19340 25774 19392 25780
rect 19430 25800 19486 25809
rect 19248 25764 19300 25770
rect 19430 25735 19486 25744
rect 19248 25706 19300 25712
rect 19536 25650 19564 25860
rect 19616 25842 19668 25848
rect 19892 25832 19944 25838
rect 19892 25774 19944 25780
rect 19444 25622 19564 25650
rect 19444 25401 19472 25622
rect 19904 25430 19932 25774
rect 19996 25702 20024 28562
rect 20088 28082 20116 28750
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 20180 27538 20208 30330
rect 20260 29572 20312 29578
rect 20260 29514 20312 29520
rect 20272 29238 20300 29514
rect 20260 29232 20312 29238
rect 20260 29174 20312 29180
rect 20168 27532 20220 27538
rect 20168 27474 20220 27480
rect 20076 27124 20128 27130
rect 20076 27066 20128 27072
rect 20088 26382 20116 27066
rect 20272 26586 20300 29174
rect 20260 26580 20312 26586
rect 20260 26522 20312 26528
rect 20076 26376 20128 26382
rect 20076 26318 20128 26324
rect 19984 25696 20036 25702
rect 19984 25638 20036 25644
rect 20088 25480 20116 26318
rect 20364 25906 20392 31583
rect 20456 31414 20484 33458
rect 20548 32230 20576 35142
rect 20628 35080 20680 35086
rect 20628 35022 20680 35028
rect 20720 35080 20772 35086
rect 20720 35022 20772 35028
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20640 34202 20668 35022
rect 20732 34950 20760 35022
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 20824 34626 20852 35022
rect 20916 34746 20944 35158
rect 21088 35012 21140 35018
rect 21088 34954 21140 34960
rect 20904 34740 20956 34746
rect 20904 34682 20956 34688
rect 20732 34610 21036 34626
rect 20732 34604 21048 34610
rect 20732 34598 20996 34604
rect 20732 34406 20760 34598
rect 20996 34546 21048 34552
rect 21100 34406 21128 34954
rect 21192 34746 21220 36042
rect 21284 35766 21312 37946
rect 21916 37664 21968 37670
rect 21916 37606 21968 37612
rect 21638 37088 21694 37097
rect 21638 37023 21694 37032
rect 21548 36712 21600 36718
rect 21548 36654 21600 36660
rect 21456 36576 21508 36582
rect 21456 36518 21508 36524
rect 21468 35834 21496 36518
rect 21560 36242 21588 36654
rect 21548 36236 21600 36242
rect 21548 36178 21600 36184
rect 21456 35828 21508 35834
rect 21456 35770 21508 35776
rect 21272 35760 21324 35766
rect 21272 35702 21324 35708
rect 21456 35624 21508 35630
rect 21456 35566 21508 35572
rect 21468 35222 21496 35566
rect 21456 35216 21508 35222
rect 21456 35158 21508 35164
rect 21272 35148 21324 35154
rect 21272 35090 21324 35096
rect 21180 34740 21232 34746
rect 21180 34682 21232 34688
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20812 34400 20864 34406
rect 20812 34342 20864 34348
rect 21088 34400 21140 34406
rect 21088 34342 21140 34348
rect 20628 34196 20680 34202
rect 20628 34138 20680 34144
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20640 33114 20668 33934
rect 20720 33924 20772 33930
rect 20720 33866 20772 33872
rect 20732 33833 20760 33866
rect 20718 33824 20774 33833
rect 20718 33759 20774 33768
rect 20824 33289 20852 34342
rect 20904 33856 20956 33862
rect 20904 33798 20956 33804
rect 20810 33280 20866 33289
rect 20810 33215 20866 33224
rect 20628 33108 20680 33114
rect 20628 33050 20680 33056
rect 20628 32904 20680 32910
rect 20916 32858 20944 33798
rect 21100 33454 21128 34342
rect 21284 33998 21312 35090
rect 21652 35086 21680 37023
rect 21640 35080 21692 35086
rect 21640 35022 21692 35028
rect 21732 34944 21784 34950
rect 21732 34886 21784 34892
rect 21364 34536 21416 34542
rect 21364 34478 21416 34484
rect 21456 34536 21508 34542
rect 21456 34478 21508 34484
rect 21376 34134 21404 34478
rect 21364 34128 21416 34134
rect 21364 34070 21416 34076
rect 21272 33992 21324 33998
rect 21324 33952 21404 33980
rect 21272 33934 21324 33940
rect 21272 33652 21324 33658
rect 21272 33594 21324 33600
rect 21088 33448 21140 33454
rect 21088 33390 21140 33396
rect 21284 33318 21312 33594
rect 21180 33312 21232 33318
rect 20628 32846 20680 32852
rect 20536 32224 20588 32230
rect 20536 32166 20588 32172
rect 20640 31958 20668 32846
rect 20824 32830 20944 32858
rect 21008 33272 21180 33300
rect 20824 32774 20852 32830
rect 20812 32768 20864 32774
rect 20812 32710 20864 32716
rect 20904 32768 20956 32774
rect 20904 32710 20956 32716
rect 20720 32496 20772 32502
rect 20720 32438 20772 32444
rect 20812 32496 20864 32502
rect 20812 32438 20864 32444
rect 20628 31952 20680 31958
rect 20628 31894 20680 31900
rect 20536 31748 20588 31754
rect 20536 31690 20588 31696
rect 20444 31408 20496 31414
rect 20444 31350 20496 31356
rect 20548 31226 20576 31690
rect 20456 31198 20576 31226
rect 20456 28121 20484 31198
rect 20628 31136 20680 31142
rect 20548 31084 20628 31090
rect 20548 31078 20680 31084
rect 20548 31062 20668 31078
rect 20548 30734 20576 31062
rect 20536 30728 20588 30734
rect 20536 30670 20588 30676
rect 20628 30660 20680 30666
rect 20628 30602 20680 30608
rect 20640 30326 20668 30602
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20732 29306 20760 32438
rect 20824 32201 20852 32438
rect 20810 32192 20866 32201
rect 20810 32127 20866 32136
rect 20810 31920 20866 31929
rect 20810 31855 20812 31864
rect 20864 31855 20866 31864
rect 20812 31826 20864 31832
rect 20916 30682 20944 32710
rect 21008 32230 21036 33272
rect 21180 33254 21232 33260
rect 21272 33312 21324 33318
rect 21272 33254 21324 33260
rect 21088 32904 21140 32910
rect 21088 32846 21140 32852
rect 21180 32904 21232 32910
rect 21180 32846 21232 32852
rect 20996 32224 21048 32230
rect 20996 32166 21048 32172
rect 21008 32026 21036 32166
rect 20996 32020 21048 32026
rect 20996 31962 21048 31968
rect 20996 31816 21048 31822
rect 20996 31758 21048 31764
rect 21008 31482 21036 31758
rect 20996 31476 21048 31482
rect 20996 31418 21048 31424
rect 21100 30938 21128 32846
rect 21192 31929 21220 32846
rect 21272 32836 21324 32842
rect 21272 32778 21324 32784
rect 21284 32337 21312 32778
rect 21270 32328 21326 32337
rect 21270 32263 21326 32272
rect 21376 31958 21404 33952
rect 21468 33658 21496 34478
rect 21640 34196 21692 34202
rect 21640 34138 21692 34144
rect 21548 33992 21600 33998
rect 21548 33934 21600 33940
rect 21456 33652 21508 33658
rect 21456 33594 21508 33600
rect 21456 33516 21508 33522
rect 21456 33458 21508 33464
rect 21468 32774 21496 33458
rect 21456 32768 21508 32774
rect 21456 32710 21508 32716
rect 21272 31952 21324 31958
rect 21178 31920 21234 31929
rect 21272 31894 21324 31900
rect 21364 31952 21416 31958
rect 21364 31894 21416 31900
rect 21178 31855 21234 31864
rect 21180 31476 21232 31482
rect 21180 31418 21232 31424
rect 21088 30932 21140 30938
rect 21088 30874 21140 30880
rect 20916 30654 21036 30682
rect 20904 30592 20956 30598
rect 20904 30534 20956 30540
rect 20916 30258 20944 30534
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 20904 29776 20956 29782
rect 20904 29718 20956 29724
rect 20720 29300 20772 29306
rect 20720 29242 20772 29248
rect 20916 28914 20944 29718
rect 21008 29102 21036 30654
rect 21192 30394 21220 31418
rect 21284 31210 21312 31894
rect 21468 31754 21496 32710
rect 21456 31748 21508 31754
rect 21456 31690 21508 31696
rect 21272 31204 21324 31210
rect 21272 31146 21324 31152
rect 21560 30705 21588 33934
rect 21652 32609 21680 34138
rect 21638 32600 21694 32609
rect 21638 32535 21694 32544
rect 21638 32464 21694 32473
rect 21638 32399 21640 32408
rect 21692 32399 21694 32408
rect 21640 32370 21692 32376
rect 21546 30696 21602 30705
rect 21546 30631 21602 30640
rect 21180 30388 21232 30394
rect 21180 30330 21232 30336
rect 21456 30320 21508 30326
rect 21456 30262 21508 30268
rect 21088 30252 21140 30258
rect 21088 30194 21140 30200
rect 21272 30252 21324 30258
rect 21272 30194 21324 30200
rect 21100 30054 21128 30194
rect 21180 30184 21232 30190
rect 21180 30126 21232 30132
rect 21088 30048 21140 30054
rect 21088 29990 21140 29996
rect 20996 29096 21048 29102
rect 20996 29038 21048 29044
rect 20916 28886 21036 28914
rect 20536 28416 20588 28422
rect 20536 28358 20588 28364
rect 20812 28416 20864 28422
rect 20812 28358 20864 28364
rect 20442 28112 20498 28121
rect 20442 28047 20498 28056
rect 20444 27396 20496 27402
rect 20444 27338 20496 27344
rect 20168 25900 20220 25906
rect 20168 25842 20220 25848
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20180 25809 20208 25842
rect 20166 25800 20222 25809
rect 20166 25735 20222 25744
rect 20352 25764 20404 25770
rect 20352 25706 20404 25712
rect 20168 25696 20220 25702
rect 20168 25638 20220 25644
rect 19996 25452 20116 25480
rect 19800 25424 19852 25430
rect 19430 25392 19486 25401
rect 19800 25366 19852 25372
rect 19892 25424 19944 25430
rect 19892 25366 19944 25372
rect 19430 25327 19486 25336
rect 19812 25254 19840 25366
rect 19996 25344 20024 25452
rect 19996 25316 20116 25344
rect 19812 25226 20024 25254
rect 19996 25129 20024 25226
rect 20088 25158 20116 25316
rect 20076 25152 20128 25158
rect 19430 25120 19486 25129
rect 19430 25055 19486 25064
rect 19982 25120 20038 25129
rect 20076 25094 20128 25100
rect 19444 24970 19472 25055
rect 19574 25052 19882 25061
rect 19982 25055 20038 25064
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 20088 24970 20116 25094
rect 19424 24942 19472 24970
rect 19524 24948 19576 24954
rect 19424 24868 19452 24942
rect 19524 24890 19576 24896
rect 19996 24942 20116 24970
rect 19352 24840 19452 24868
rect 19352 24834 19380 24840
rect 19260 24806 19380 24834
rect 19260 23497 19288 24806
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 19246 23488 19302 23497
rect 19246 23423 19302 23432
rect 19154 23352 19210 23361
rect 19154 23287 19210 23296
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 19156 23112 19208 23118
rect 19156 23054 19208 23060
rect 19168 22642 19196 23054
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 18788 22568 18840 22574
rect 18050 22536 18106 22545
rect 17960 22500 18012 22506
rect 18788 22510 18840 22516
rect 18050 22471 18106 22480
rect 17960 22442 18012 22448
rect 18800 22234 18828 22510
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 17776 21344 17828 21350
rect 17776 21286 17828 21292
rect 17130 20904 17186 20913
rect 17130 20839 17132 20848
rect 17184 20839 17186 20848
rect 17132 20810 17184 20816
rect 17788 20806 17816 21286
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 17788 20618 17816 20742
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 17040 20596 17092 20602
rect 17040 20538 17092 20544
rect 17696 20590 17816 20618
rect 16960 20466 16988 20538
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 17052 19242 17080 20538
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17512 20262 17540 20402
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17040 19236 17092 19242
rect 17040 19178 17092 19184
rect 17144 18766 17172 19314
rect 17236 18834 17264 20198
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16776 16918 16896 16946
rect 16500 16658 16712 16674
rect 16500 16652 16724 16658
rect 16500 16646 16672 16652
rect 16672 16594 16724 16600
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15028 15978 15056 16390
rect 15304 16114 15332 16390
rect 16040 16266 16068 16526
rect 15948 16238 16068 16266
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15948 16046 15976 16238
rect 16132 16130 16160 16526
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16040 16114 16160 16130
rect 16028 16108 16160 16114
rect 16080 16102 16160 16108
rect 16028 16050 16080 16056
rect 16592 16046 16620 16458
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 16776 15706 16804 16918
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16868 16114 16896 16730
rect 16960 16114 16988 18362
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17420 17202 17448 18022
rect 17512 17678 17540 20198
rect 17696 19378 17724 20590
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17788 19378 17816 20402
rect 17972 19854 18000 21558
rect 18050 20496 18106 20505
rect 18050 20431 18106 20440
rect 18064 19922 18092 20431
rect 18156 20369 18184 21830
rect 18248 21690 18276 21966
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 18512 21480 18564 21486
rect 18512 21422 18564 21428
rect 18234 21040 18290 21049
rect 18234 20975 18290 20984
rect 18142 20360 18198 20369
rect 18142 20295 18198 20304
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18064 19378 18092 19654
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 17788 17678 17816 18634
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 17052 16182 17080 16934
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 14738 15600 14794 15609
rect 14738 15535 14794 15544
rect 17420 15026 17448 17138
rect 17512 17134 17540 17614
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17512 16794 17540 17070
rect 18064 17066 18092 17206
rect 18156 17134 18184 18022
rect 18248 17678 18276 20975
rect 18524 20806 18552 21422
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18524 20534 18552 20742
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18524 19174 18552 19246
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18616 18698 18644 21830
rect 19168 21622 19196 22578
rect 19260 21690 19288 23423
rect 19352 23186 19380 24278
rect 19536 24177 19564 24890
rect 19800 24880 19852 24886
rect 19800 24822 19852 24828
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 19628 24410 19656 24754
rect 19812 24750 19840 24822
rect 19800 24744 19852 24750
rect 19800 24686 19852 24692
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 19522 24168 19578 24177
rect 19522 24103 19578 24112
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19616 23860 19668 23866
rect 19996 23848 20024 24942
rect 20180 24682 20208 25638
rect 20364 25362 20392 25706
rect 20456 25498 20484 27338
rect 20548 27044 20576 28358
rect 20718 28248 20774 28257
rect 20718 28183 20720 28192
rect 20772 28183 20774 28192
rect 20720 28154 20772 28160
rect 20720 27328 20772 27334
rect 20720 27270 20772 27276
rect 20628 27056 20680 27062
rect 20548 27016 20628 27044
rect 20548 26926 20576 27016
rect 20628 26998 20680 27004
rect 20536 26920 20588 26926
rect 20536 26862 20588 26868
rect 20628 26784 20680 26790
rect 20628 26726 20680 26732
rect 20536 26376 20588 26382
rect 20534 26344 20536 26353
rect 20588 26344 20590 26353
rect 20534 26279 20590 26288
rect 20534 26208 20590 26217
rect 20534 26143 20590 26152
rect 20548 25974 20576 26143
rect 20536 25968 20588 25974
rect 20536 25910 20588 25916
rect 20640 25906 20668 26726
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20536 25764 20588 25770
rect 20536 25706 20588 25712
rect 20444 25492 20496 25498
rect 20444 25434 20496 25440
rect 20548 25378 20576 25706
rect 20626 25528 20682 25537
rect 20626 25463 20628 25472
rect 20680 25463 20682 25472
rect 20628 25434 20680 25440
rect 20352 25356 20404 25362
rect 20548 25350 20668 25378
rect 20352 25298 20404 25304
rect 20640 25226 20668 25350
rect 20352 25220 20404 25226
rect 20352 25162 20404 25168
rect 20628 25220 20680 25226
rect 20628 25162 20680 25168
rect 20260 24812 20312 24818
rect 20260 24754 20312 24760
rect 20168 24676 20220 24682
rect 20168 24618 20220 24624
rect 20272 24070 20300 24754
rect 20364 24721 20392 25162
rect 20536 24744 20588 24750
rect 20350 24712 20406 24721
rect 20350 24647 20406 24656
rect 20456 24692 20536 24698
rect 20456 24686 20588 24692
rect 20456 24670 20576 24686
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 19616 23802 19668 23808
rect 19812 23820 20024 23848
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19352 22098 19380 22714
rect 19444 22234 19472 23666
rect 19628 23594 19656 23802
rect 19708 23724 19760 23730
rect 19708 23666 19760 23672
rect 19720 23594 19748 23666
rect 19616 23588 19668 23594
rect 19616 23530 19668 23536
rect 19708 23588 19760 23594
rect 19708 23530 19760 23536
rect 19812 23474 19840 23820
rect 20088 23662 20116 24006
rect 20456 23866 20484 24670
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20548 24138 20576 24550
rect 20536 24132 20588 24138
rect 20536 24074 20588 24080
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 19892 23656 19944 23662
rect 19892 23598 19944 23604
rect 20076 23656 20128 23662
rect 20076 23598 20128 23604
rect 19628 23446 19840 23474
rect 19628 23118 19656 23446
rect 19904 23254 19932 23598
rect 19892 23248 19944 23254
rect 19892 23190 19944 23196
rect 20168 23180 20220 23186
rect 20168 23122 20220 23128
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19720 22982 19748 23054
rect 19708 22976 19760 22982
rect 19708 22918 19760 22924
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19798 22536 19854 22545
rect 19798 22471 19854 22480
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19536 22030 19564 22374
rect 19812 22166 19840 22471
rect 20180 22409 20208 23122
rect 20272 22953 20300 23802
rect 20548 23730 20576 23802
rect 20640 23730 20668 25162
rect 20732 24698 20760 27270
rect 20824 26790 20852 28358
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20916 25702 20944 26862
rect 21008 26081 21036 28886
rect 21100 28558 21128 29990
rect 21088 28552 21140 28558
rect 21088 28494 21140 28500
rect 21088 28212 21140 28218
rect 21088 28154 21140 28160
rect 21100 28082 21128 28154
rect 21088 28076 21140 28082
rect 21088 28018 21140 28024
rect 20994 26072 21050 26081
rect 20994 26007 21050 26016
rect 20996 25832 21048 25838
rect 20996 25774 21048 25780
rect 21008 25702 21036 25774
rect 20904 25696 20956 25702
rect 20904 25638 20956 25644
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 20996 25152 21048 25158
rect 20996 25094 21048 25100
rect 21008 24954 21036 25094
rect 20996 24948 21048 24954
rect 20996 24890 21048 24896
rect 20904 24812 20956 24818
rect 20904 24754 20956 24760
rect 20916 24721 20944 24754
rect 20902 24712 20958 24721
rect 20732 24670 20852 24698
rect 20720 24608 20772 24614
rect 20718 24576 20720 24585
rect 20772 24576 20774 24585
rect 20718 24511 20774 24520
rect 20824 24342 20852 24670
rect 20902 24647 20958 24656
rect 20916 24410 20944 24647
rect 20904 24404 20956 24410
rect 20904 24346 20956 24352
rect 20812 24336 20864 24342
rect 20812 24278 20864 24284
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20628 23724 20680 23730
rect 20824 23712 20852 24278
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 20904 23724 20956 23730
rect 20824 23684 20904 23712
rect 20628 23666 20680 23672
rect 20904 23666 20956 23672
rect 20718 23624 20774 23633
rect 20718 23559 20774 23568
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 20628 23520 20680 23526
rect 20628 23462 20680 23468
rect 20442 23352 20498 23361
rect 20442 23287 20498 23296
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 20258 22944 20314 22953
rect 20258 22879 20314 22888
rect 20364 22710 20392 23054
rect 20456 22778 20484 23287
rect 20444 22772 20496 22778
rect 20444 22714 20496 22720
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 20166 22400 20222 22409
rect 20166 22335 20222 22344
rect 19800 22160 19852 22166
rect 19800 22102 19852 22108
rect 19996 22080 20392 22094
rect 20456 22080 20484 22714
rect 19996 22066 20484 22080
rect 19524 22024 19576 22030
rect 19892 22024 19944 22030
rect 19524 21966 19576 21972
rect 19890 21992 19892 22001
rect 19944 21992 19946 22001
rect 19890 21927 19946 21936
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19248 21684 19300 21690
rect 19996 21672 20024 22066
rect 20364 22052 20484 22066
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 19248 21626 19300 21632
rect 19904 21644 20024 21672
rect 20074 21720 20130 21729
rect 20074 21655 20130 21664
rect 19156 21616 19208 21622
rect 19156 21558 19208 21564
rect 19156 21480 19208 21486
rect 19904 21457 19932 21644
rect 20088 21554 20116 21655
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 19156 21422 19208 21428
rect 19890 21448 19946 21457
rect 18696 21412 18748 21418
rect 18696 21354 18748 21360
rect 18708 20466 18736 21354
rect 19168 21078 19196 21422
rect 20088 21434 20116 21490
rect 19890 21383 19946 21392
rect 19996 21406 20116 21434
rect 19996 21350 20024 21406
rect 20180 21350 20208 21966
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 19156 21072 19208 21078
rect 19156 21014 19208 21020
rect 19248 21072 19300 21078
rect 19248 21014 19300 21020
rect 19984 21072 20036 21078
rect 19984 21014 20036 21020
rect 19260 20942 19288 21014
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 19352 20262 19380 20878
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 18880 19780 18932 19786
rect 18880 19722 18932 19728
rect 18604 18692 18656 18698
rect 18604 18634 18656 18640
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 18290 18368 18566
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18524 17882 18552 18158
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18052 17060 18104 17066
rect 18052 17002 18104 17008
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 18064 16590 18092 17002
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 17604 16046 17632 16526
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 18156 15026 18184 17070
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18432 15978 18460 16594
rect 18524 16114 18552 17138
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18420 15972 18472 15978
rect 18420 15914 18472 15920
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18432 14890 18460 15914
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 18524 14618 18552 15438
rect 18616 15094 18644 16050
rect 18708 15570 18736 19722
rect 18892 17678 18920 19722
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18984 18766 19012 19110
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 19352 18426 19380 19246
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 19076 17338 19104 17614
rect 19168 17610 19196 18022
rect 19156 17604 19208 17610
rect 19156 17546 19208 17552
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18972 17264 19024 17270
rect 18972 17206 19024 17212
rect 18880 17060 18932 17066
rect 18880 17002 18932 17008
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18708 13870 18736 15506
rect 18892 15502 18920 17002
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18800 13938 18828 14826
rect 18984 13938 19012 17206
rect 19168 16998 19196 17546
rect 19444 17202 19472 20266
rect 19996 19990 20024 21014
rect 20088 20398 20116 21286
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 20180 20330 20208 20878
rect 20272 20466 20300 21626
rect 20548 21536 20576 23462
rect 20640 23254 20668 23462
rect 20732 23361 20760 23559
rect 20718 23352 20774 23361
rect 20718 23287 20774 23296
rect 20628 23248 20680 23254
rect 20628 23190 20680 23196
rect 20640 21690 20668 23190
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20732 22642 20760 23054
rect 20812 22976 20864 22982
rect 20812 22918 20864 22924
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20824 22094 20852 22918
rect 20824 22066 20944 22094
rect 20628 21684 20680 21690
rect 20628 21626 20680 21632
rect 20364 21508 20576 21536
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 20088 20097 20116 20198
rect 20074 20088 20130 20097
rect 20074 20023 20130 20032
rect 19984 19984 20036 19990
rect 19984 19926 20036 19932
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 19628 18766 19656 19382
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20088 18426 20116 20023
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 20272 19514 20300 19926
rect 20364 19718 20392 21508
rect 20444 21412 20496 21418
rect 20444 21354 20496 21360
rect 20456 21010 20484 21354
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20548 20602 20576 21286
rect 20640 21078 20668 21286
rect 20628 21072 20680 21078
rect 20628 21014 20680 21020
rect 20536 20596 20588 20602
rect 20720 20596 20772 20602
rect 20588 20556 20668 20584
rect 20536 20538 20588 20544
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 19798 18320 19854 18329
rect 19798 18255 19854 18264
rect 19812 18222 19840 18255
rect 20088 18222 20116 18362
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19536 17678 19564 17818
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20180 17202 20208 18362
rect 20272 17354 20300 19450
rect 20456 18358 20484 19994
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20548 19446 20576 19790
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 20548 18766 20576 19382
rect 20640 19378 20668 20556
rect 20720 20538 20772 20544
rect 20732 19854 20760 20538
rect 20916 20482 20944 22066
rect 21008 21622 21036 23802
rect 21100 23730 21128 28018
rect 21192 25514 21220 30126
rect 21284 29306 21312 30194
rect 21468 30054 21496 30262
rect 21456 30048 21508 30054
rect 21456 29990 21508 29996
rect 21652 29889 21680 32370
rect 21744 32298 21772 34886
rect 21824 34400 21876 34406
rect 21824 34342 21876 34348
rect 21836 34202 21864 34342
rect 21824 34196 21876 34202
rect 21824 34138 21876 34144
rect 21928 33522 21956 37606
rect 22112 37262 22140 39102
rect 23296 39024 23348 39030
rect 22374 38992 22430 39001
rect 23296 38966 23348 38972
rect 22374 38927 22430 38936
rect 22284 38752 22336 38758
rect 22284 38694 22336 38700
rect 22100 37256 22152 37262
rect 22100 37198 22152 37204
rect 22098 36136 22154 36145
rect 22296 36106 22324 38694
rect 22098 36071 22154 36080
rect 22284 36100 22336 36106
rect 22006 36000 22062 36009
rect 22006 35935 22062 35944
rect 22020 35698 22048 35935
rect 22008 35692 22060 35698
rect 22008 35634 22060 35640
rect 22112 34406 22140 36071
rect 22284 36042 22336 36048
rect 22388 35766 22416 38927
rect 23204 38752 23256 38758
rect 23204 38694 23256 38700
rect 23020 38072 23072 38078
rect 23020 38014 23072 38020
rect 22560 37460 22612 37466
rect 22560 37402 22612 37408
rect 22468 37188 22520 37194
rect 22468 37130 22520 37136
rect 22376 35760 22428 35766
rect 22376 35702 22428 35708
rect 22480 35018 22508 37130
rect 22572 36854 22600 37402
rect 22652 37188 22704 37194
rect 22652 37130 22704 37136
rect 22560 36848 22612 36854
rect 22560 36790 22612 36796
rect 22560 36712 22612 36718
rect 22664 36689 22692 37130
rect 22560 36654 22612 36660
rect 22650 36680 22706 36689
rect 22572 35086 22600 36654
rect 22650 36615 22706 36624
rect 22652 36236 22704 36242
rect 22652 36178 22704 36184
rect 22560 35080 22612 35086
rect 22560 35022 22612 35028
rect 22468 35012 22520 35018
rect 22468 34954 22520 34960
rect 22560 34944 22612 34950
rect 22560 34886 22612 34892
rect 22100 34400 22152 34406
rect 22100 34342 22152 34348
rect 22100 34196 22152 34202
rect 22152 34156 22416 34184
rect 22100 34138 22152 34144
rect 22100 34060 22152 34066
rect 22100 34002 22152 34008
rect 22112 33969 22140 34002
rect 22098 33960 22154 33969
rect 22098 33895 22154 33904
rect 22388 33862 22416 34156
rect 22466 33960 22522 33969
rect 22466 33895 22522 33904
rect 22376 33856 22428 33862
rect 22376 33798 22428 33804
rect 22282 33688 22338 33697
rect 22192 33652 22244 33658
rect 22112 33612 22192 33640
rect 21916 33516 21968 33522
rect 21916 33458 21968 33464
rect 22008 33380 22060 33386
rect 22008 33322 22060 33328
rect 22020 33130 22048 33322
rect 22112 33318 22140 33612
rect 22282 33623 22338 33632
rect 22192 33594 22244 33600
rect 22296 33522 22324 33623
rect 22284 33516 22336 33522
rect 22284 33458 22336 33464
rect 22480 33386 22508 33895
rect 22572 33862 22600 34886
rect 22664 34746 22692 36178
rect 23032 36145 23060 38014
rect 23110 36544 23166 36553
rect 23110 36479 23166 36488
rect 23018 36136 23074 36145
rect 23018 36071 23074 36080
rect 22928 35624 22980 35630
rect 22928 35566 22980 35572
rect 22652 34740 22704 34746
rect 22652 34682 22704 34688
rect 22652 34400 22704 34406
rect 22652 34342 22704 34348
rect 22742 34368 22798 34377
rect 22664 33998 22692 34342
rect 22742 34303 22798 34312
rect 22652 33992 22704 33998
rect 22652 33934 22704 33940
rect 22560 33856 22612 33862
rect 22560 33798 22612 33804
rect 22560 33516 22612 33522
rect 22560 33458 22612 33464
rect 22284 33380 22336 33386
rect 22284 33322 22336 33328
rect 22468 33380 22520 33386
rect 22468 33322 22520 33328
rect 22100 33312 22152 33318
rect 22100 33254 22152 33260
rect 22020 33102 22232 33130
rect 21824 33040 21876 33046
rect 21824 32982 21876 32988
rect 22100 33040 22152 33046
rect 22204 33017 22232 33102
rect 22100 32982 22152 32988
rect 22190 33008 22246 33017
rect 21836 32473 21864 32982
rect 22112 32858 22140 32982
rect 22190 32943 22246 32952
rect 22112 32830 22232 32858
rect 22100 32768 22152 32774
rect 21914 32736 21970 32745
rect 22100 32710 22152 32716
rect 21914 32671 21970 32680
rect 21822 32464 21878 32473
rect 21822 32399 21878 32408
rect 21732 32292 21784 32298
rect 21732 32234 21784 32240
rect 21744 31890 21772 32234
rect 21732 31884 21784 31890
rect 21732 31826 21784 31832
rect 21928 31822 21956 32671
rect 22112 32570 22140 32710
rect 22204 32570 22232 32830
rect 22100 32564 22152 32570
rect 22100 32506 22152 32512
rect 22192 32564 22244 32570
rect 22192 32506 22244 32512
rect 22192 32428 22244 32434
rect 22192 32370 22244 32376
rect 22098 32192 22154 32201
rect 22098 32127 22154 32136
rect 22112 31822 22140 32127
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 21928 31142 21956 31758
rect 22204 31482 22232 32370
rect 22192 31476 22244 31482
rect 22192 31418 22244 31424
rect 21824 31136 21876 31142
rect 21824 31078 21876 31084
rect 21916 31136 21968 31142
rect 21916 31078 21968 31084
rect 21732 30932 21784 30938
rect 21732 30874 21784 30880
rect 21638 29880 21694 29889
rect 21638 29815 21694 29824
rect 21548 29776 21600 29782
rect 21548 29718 21600 29724
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 21272 29300 21324 29306
rect 21272 29242 21324 29248
rect 21272 29164 21324 29170
rect 21272 29106 21324 29112
rect 21284 27606 21312 29106
rect 21362 28928 21418 28937
rect 21362 28863 21418 28872
rect 21376 28082 21404 28863
rect 21468 28422 21496 29582
rect 21456 28416 21508 28422
rect 21456 28358 21508 28364
rect 21560 28218 21588 29718
rect 21640 29572 21692 29578
rect 21640 29514 21692 29520
rect 21652 28422 21680 29514
rect 21744 28694 21772 30874
rect 21836 30818 21864 31078
rect 22296 30954 22324 33322
rect 22376 33108 22428 33114
rect 22376 33050 22428 33056
rect 22388 32026 22416 33050
rect 22572 32858 22600 33458
rect 22480 32830 22600 32858
rect 22480 32434 22508 32830
rect 22560 32768 22612 32774
rect 22560 32710 22612 32716
rect 22468 32428 22520 32434
rect 22468 32370 22520 32376
rect 22468 32292 22520 32298
rect 22468 32234 22520 32240
rect 22480 32026 22508 32234
rect 22376 32020 22428 32026
rect 22376 31962 22428 31968
rect 22468 32020 22520 32026
rect 22468 31962 22520 31968
rect 22480 31906 22508 31962
rect 22204 30926 22324 30954
rect 22388 31878 22508 31906
rect 21836 30790 22140 30818
rect 22112 30734 22140 30790
rect 22008 30728 22060 30734
rect 22008 30670 22060 30676
rect 22100 30728 22152 30734
rect 22100 30670 22152 30676
rect 22020 30258 22048 30670
rect 22204 30598 22232 30926
rect 22284 30864 22336 30870
rect 22284 30806 22336 30812
rect 22192 30592 22244 30598
rect 22192 30534 22244 30540
rect 22204 30410 22232 30534
rect 22112 30382 22232 30410
rect 22008 30252 22060 30258
rect 21836 30212 22008 30240
rect 21732 28688 21784 28694
rect 21732 28630 21784 28636
rect 21836 28626 21864 30212
rect 22008 30194 22060 30200
rect 22008 30116 22060 30122
rect 22008 30058 22060 30064
rect 22020 29714 22048 30058
rect 21916 29708 21968 29714
rect 21916 29650 21968 29656
rect 22008 29708 22060 29714
rect 22008 29650 22060 29656
rect 21824 28620 21876 28626
rect 21824 28562 21876 28568
rect 21732 28552 21784 28558
rect 21732 28494 21784 28500
rect 21640 28416 21692 28422
rect 21640 28358 21692 28364
rect 21548 28212 21600 28218
rect 21548 28154 21600 28160
rect 21454 28112 21510 28121
rect 21364 28076 21416 28082
rect 21454 28047 21510 28056
rect 21364 28018 21416 28024
rect 21364 27940 21416 27946
rect 21364 27882 21416 27888
rect 21272 27600 21324 27606
rect 21272 27542 21324 27548
rect 21284 25702 21312 27542
rect 21376 27130 21404 27882
rect 21364 27124 21416 27130
rect 21364 27066 21416 27072
rect 21376 26926 21404 27066
rect 21364 26920 21416 26926
rect 21364 26862 21416 26868
rect 21468 26246 21496 28047
rect 21638 27976 21694 27985
rect 21638 27911 21694 27920
rect 21548 27396 21600 27402
rect 21548 27338 21600 27344
rect 21456 26240 21508 26246
rect 21456 26182 21508 26188
rect 21272 25696 21324 25702
rect 21272 25638 21324 25644
rect 21560 25650 21588 27338
rect 21652 26382 21680 27911
rect 21744 26450 21772 28494
rect 21824 27328 21876 27334
rect 21824 27270 21876 27276
rect 21836 27062 21864 27270
rect 21824 27056 21876 27062
rect 21824 26998 21876 27004
rect 21732 26444 21784 26450
rect 21732 26386 21784 26392
rect 21640 26376 21692 26382
rect 21640 26318 21692 26324
rect 21732 25900 21784 25906
rect 21732 25842 21784 25848
rect 21560 25622 21680 25650
rect 21192 25486 21588 25514
rect 21456 25356 21508 25362
rect 21456 25298 21508 25304
rect 21468 25158 21496 25298
rect 21364 25152 21416 25158
rect 21364 25094 21416 25100
rect 21456 25152 21508 25158
rect 21456 25094 21508 25100
rect 21376 24886 21404 25094
rect 21364 24880 21416 24886
rect 21364 24822 21416 24828
rect 21088 23724 21140 23730
rect 21088 23666 21140 23672
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 20996 21616 21048 21622
rect 20996 21558 21048 21564
rect 21100 21486 21128 21898
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21088 21480 21140 21486
rect 21088 21422 21140 21428
rect 21468 20942 21496 21490
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 20824 20454 20944 20482
rect 20824 19990 20852 20454
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20916 19990 20944 20334
rect 20812 19984 20864 19990
rect 20812 19926 20864 19932
rect 20904 19984 20956 19990
rect 20904 19926 20956 19932
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20824 19514 20852 19790
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20536 18760 20588 18766
rect 20536 18702 20588 18708
rect 20640 18698 20668 19314
rect 20916 18970 20944 19790
rect 21008 19310 21036 20334
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 21100 19242 21128 20878
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21284 20262 21312 20402
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21284 19514 21312 20198
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21468 19378 21496 20402
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21088 19236 21140 19242
rect 21088 19178 21140 19184
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 21468 18834 21496 19314
rect 21456 18828 21508 18834
rect 21456 18770 21508 18776
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20640 18358 20668 18634
rect 20444 18352 20496 18358
rect 20444 18294 20496 18300
rect 20628 18352 20680 18358
rect 20680 18300 20760 18306
rect 20628 18294 20760 18300
rect 20640 18278 20760 18294
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20272 17326 20392 17354
rect 20260 17264 20312 17270
rect 20260 17206 20312 17212
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 19168 15026 19196 15982
rect 19352 15706 19380 17070
rect 19432 16720 19484 16726
rect 19432 16662 19484 16668
rect 19444 16250 19472 16662
rect 20272 16454 20300 17206
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19260 14278 19288 14894
rect 19444 14414 19472 15438
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19536 14550 19564 14894
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19260 13938 19288 14214
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 19352 13530 19380 14282
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 19444 12306 19472 13806
rect 19996 13394 20024 15642
rect 20088 15502 20116 15846
rect 20168 15632 20220 15638
rect 20168 15574 20220 15580
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 20088 14414 20116 15438
rect 20180 14958 20208 15574
rect 20272 15502 20300 16390
rect 20364 16266 20392 17326
rect 20548 17202 20576 18022
rect 20732 17678 20760 18278
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20902 18184 20958 18193
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20824 17610 20852 18158
rect 20902 18119 20958 18128
rect 20916 17678 20944 18119
rect 21272 17808 21324 17814
rect 21272 17750 21324 17756
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 21284 17610 21312 17750
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20456 16590 20484 17138
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20364 16238 20484 16266
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20364 15638 20392 16050
rect 20352 15632 20404 15638
rect 20352 15574 20404 15580
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 20272 13190 20300 15438
rect 20456 15026 20484 16238
rect 20548 15570 20576 17138
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20824 16114 20852 16934
rect 20916 16522 20944 17478
rect 21284 17066 21312 17546
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 20904 16516 20956 16522
rect 20904 16458 20956 16464
rect 21284 16114 21312 17002
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21376 16250 21404 16594
rect 21560 16250 21588 25486
rect 21652 23526 21680 25622
rect 21744 24993 21772 25842
rect 21730 24984 21786 24993
rect 21730 24919 21786 24928
rect 21744 24313 21772 24919
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21836 24410 21864 24754
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21730 24304 21786 24313
rect 21730 24239 21786 24248
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21928 22094 21956 29650
rect 22112 29170 22140 30382
rect 22192 30320 22244 30326
rect 22192 30262 22244 30268
rect 22204 29646 22232 30262
rect 22296 30258 22324 30806
rect 22388 30734 22416 31878
rect 22572 31822 22600 32710
rect 22664 32026 22692 33934
rect 22756 33930 22784 34303
rect 22940 34066 22968 35566
rect 23032 34610 23060 36071
rect 23124 36038 23152 36479
rect 23112 36032 23164 36038
rect 23112 35974 23164 35980
rect 23110 35456 23166 35465
rect 23110 35391 23166 35400
rect 23020 34604 23072 34610
rect 23020 34546 23072 34552
rect 23020 34196 23072 34202
rect 23020 34138 23072 34144
rect 22928 34060 22980 34066
rect 22848 34020 22928 34048
rect 22744 33924 22796 33930
rect 22744 33866 22796 33872
rect 22744 33516 22796 33522
rect 22744 33458 22796 33464
rect 22756 32978 22784 33458
rect 22744 32972 22796 32978
rect 22744 32914 22796 32920
rect 22756 32473 22784 32914
rect 22848 32745 22876 34020
rect 22928 34002 22980 34008
rect 23032 33998 23060 34138
rect 23124 34066 23152 35391
rect 23112 34060 23164 34066
rect 23112 34002 23164 34008
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 23020 33856 23072 33862
rect 23020 33798 23072 33804
rect 22928 33312 22980 33318
rect 22928 33254 22980 33260
rect 22940 32842 22968 33254
rect 22928 32836 22980 32842
rect 22928 32778 22980 32784
rect 22834 32736 22890 32745
rect 22834 32671 22890 32680
rect 22926 32600 22982 32609
rect 22926 32535 22982 32544
rect 22742 32464 22798 32473
rect 22742 32399 22798 32408
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 22744 32360 22796 32366
rect 22744 32302 22796 32308
rect 22756 32201 22784 32302
rect 22848 32298 22876 32370
rect 22836 32292 22888 32298
rect 22836 32234 22888 32240
rect 22742 32192 22798 32201
rect 22798 32150 22876 32178
rect 22742 32127 22798 32136
rect 22652 32020 22704 32026
rect 22652 31962 22704 31968
rect 22560 31816 22612 31822
rect 22560 31758 22612 31764
rect 22468 31340 22520 31346
rect 22468 31282 22520 31288
rect 22652 31340 22704 31346
rect 22652 31282 22704 31288
rect 22376 30728 22428 30734
rect 22376 30670 22428 30676
rect 22480 30666 22508 31282
rect 22560 31136 22612 31142
rect 22560 31078 22612 31084
rect 22572 30666 22600 31078
rect 22664 30870 22692 31282
rect 22744 31136 22796 31142
rect 22744 31078 22796 31084
rect 22652 30864 22704 30870
rect 22652 30806 22704 30812
rect 22652 30728 22704 30734
rect 22652 30670 22704 30676
rect 22468 30660 22520 30666
rect 22468 30602 22520 30608
rect 22560 30660 22612 30666
rect 22560 30602 22612 30608
rect 22480 30258 22508 30602
rect 22560 30320 22612 30326
rect 22560 30262 22612 30268
rect 22284 30252 22336 30258
rect 22284 30194 22336 30200
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22572 30122 22600 30262
rect 22560 30116 22612 30122
rect 22560 30058 22612 30064
rect 22468 30048 22520 30054
rect 22468 29990 22520 29996
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 22480 29306 22508 29990
rect 22468 29300 22520 29306
rect 22468 29242 22520 29248
rect 22190 29200 22246 29209
rect 22100 29164 22152 29170
rect 22190 29135 22246 29144
rect 22376 29164 22428 29170
rect 22100 29106 22152 29112
rect 22008 28960 22060 28966
rect 22008 28902 22060 28908
rect 22020 28218 22048 28902
rect 22098 28792 22154 28801
rect 22098 28727 22154 28736
rect 22008 28212 22060 28218
rect 22008 28154 22060 28160
rect 22112 28014 22140 28727
rect 22204 28558 22232 29135
rect 22376 29106 22428 29112
rect 22388 29073 22416 29106
rect 22374 29064 22430 29073
rect 22374 28999 22430 29008
rect 22284 28960 22336 28966
rect 22284 28902 22336 28908
rect 22192 28552 22244 28558
rect 22192 28494 22244 28500
rect 22100 28008 22152 28014
rect 22100 27950 22152 27956
rect 22008 27872 22060 27878
rect 22008 27814 22060 27820
rect 22020 27538 22048 27814
rect 22192 27668 22244 27674
rect 22192 27610 22244 27616
rect 22008 27532 22060 27538
rect 22008 27474 22060 27480
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 22008 27124 22060 27130
rect 22008 27066 22060 27072
rect 22020 25974 22048 27066
rect 22008 25968 22060 25974
rect 22008 25910 22060 25916
rect 22112 25770 22140 27406
rect 22204 26042 22232 27610
rect 22192 26036 22244 26042
rect 22192 25978 22244 25984
rect 22100 25764 22152 25770
rect 22100 25706 22152 25712
rect 22192 25764 22244 25770
rect 22192 25706 22244 25712
rect 22008 24744 22060 24750
rect 22008 24686 22060 24692
rect 22020 24206 22048 24686
rect 22008 24200 22060 24206
rect 22204 24177 22232 25706
rect 22008 24142 22060 24148
rect 22190 24168 22246 24177
rect 22020 23118 22048 24142
rect 22190 24103 22246 24112
rect 22296 23730 22324 28902
rect 22572 28490 22600 30058
rect 22664 29782 22692 30670
rect 22652 29776 22704 29782
rect 22652 29718 22704 29724
rect 22650 29608 22706 29617
rect 22650 29543 22706 29552
rect 22664 28642 22692 29543
rect 22756 29209 22784 31078
rect 22848 30802 22876 32150
rect 22836 30796 22888 30802
rect 22836 30738 22888 30744
rect 22940 29306 22968 32535
rect 23032 32008 23060 33798
rect 23124 32473 23152 34002
rect 23216 33454 23244 38694
rect 23308 35834 23336 38966
rect 23388 38888 23440 38894
rect 23388 38830 23440 38836
rect 23400 36961 23428 38830
rect 23664 38548 23716 38554
rect 23664 38490 23716 38496
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 23480 37120 23532 37126
rect 23480 37062 23532 37068
rect 23386 36952 23442 36961
rect 23386 36887 23442 36896
rect 23296 35828 23348 35834
rect 23296 35770 23348 35776
rect 23308 34610 23336 35770
rect 23388 35148 23440 35154
rect 23388 35090 23440 35096
rect 23400 35057 23428 35090
rect 23492 35086 23520 37062
rect 23584 36378 23612 37198
rect 23676 36786 23704 38490
rect 24674 38176 24730 38185
rect 24674 38111 24730 38120
rect 24308 37392 24360 37398
rect 24308 37334 24360 37340
rect 24490 37360 24546 37369
rect 23848 37188 23900 37194
rect 23848 37130 23900 37136
rect 24124 37188 24176 37194
rect 24124 37130 24176 37136
rect 23860 36922 23888 37130
rect 23848 36916 23900 36922
rect 23900 36876 23980 36904
rect 23848 36858 23900 36864
rect 23664 36780 23716 36786
rect 23664 36722 23716 36728
rect 23664 36576 23716 36582
rect 23664 36518 23716 36524
rect 23572 36372 23624 36378
rect 23572 36314 23624 36320
rect 23572 36032 23624 36038
rect 23572 35974 23624 35980
rect 23480 35080 23532 35086
rect 23386 35048 23442 35057
rect 23480 35022 23532 35028
rect 23386 34983 23442 34992
rect 23388 34672 23440 34678
rect 23386 34640 23388 34649
rect 23440 34640 23442 34649
rect 23296 34604 23348 34610
rect 23386 34575 23442 34584
rect 23296 34546 23348 34552
rect 23294 34504 23350 34513
rect 23294 34439 23350 34448
rect 23308 33522 23336 34439
rect 23584 33538 23612 35974
rect 23296 33516 23348 33522
rect 23296 33458 23348 33464
rect 23400 33510 23612 33538
rect 23204 33448 23256 33454
rect 23204 33390 23256 33396
rect 23296 32904 23348 32910
rect 23296 32846 23348 32852
rect 23204 32768 23256 32774
rect 23204 32710 23256 32716
rect 23110 32464 23166 32473
rect 23110 32399 23166 32408
rect 23032 31980 23152 32008
rect 23020 31884 23072 31890
rect 23020 31826 23072 31832
rect 22928 29300 22980 29306
rect 22928 29242 22980 29248
rect 22742 29200 22798 29209
rect 22742 29135 22798 29144
rect 22664 28614 22784 28642
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 22664 27713 22692 28494
rect 22756 28014 22784 28614
rect 22928 28552 22980 28558
rect 22928 28494 22980 28500
rect 22940 28234 22968 28494
rect 22848 28206 22968 28234
rect 22744 28008 22796 28014
rect 22744 27950 22796 27956
rect 22650 27704 22706 27713
rect 22650 27639 22706 27648
rect 22376 27600 22428 27606
rect 22376 27542 22428 27548
rect 22388 23798 22416 27542
rect 22848 27146 22876 28206
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 22940 27713 22968 28018
rect 23032 27946 23060 31826
rect 23124 31482 23152 31980
rect 23112 31476 23164 31482
rect 23112 31418 23164 31424
rect 23216 31346 23244 32710
rect 23308 31929 23336 32846
rect 23400 32337 23428 33510
rect 23572 33448 23624 33454
rect 23572 33390 23624 33396
rect 23480 33380 23532 33386
rect 23480 33322 23532 33328
rect 23492 33017 23520 33322
rect 23478 33008 23534 33017
rect 23478 32943 23534 32952
rect 23480 32836 23532 32842
rect 23480 32778 23532 32784
rect 23492 32502 23520 32778
rect 23480 32496 23532 32502
rect 23480 32438 23532 32444
rect 23386 32328 23442 32337
rect 23386 32263 23442 32272
rect 23294 31920 23350 31929
rect 23294 31855 23350 31864
rect 23204 31340 23256 31346
rect 23204 31282 23256 31288
rect 23112 31272 23164 31278
rect 23112 31214 23164 31220
rect 23124 30326 23152 31214
rect 23308 30954 23336 31855
rect 23400 31822 23428 32263
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 23388 31680 23440 31686
rect 23388 31622 23440 31628
rect 23400 31346 23428 31622
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 23216 30926 23336 30954
rect 23112 30320 23164 30326
rect 23112 30262 23164 30268
rect 23112 30116 23164 30122
rect 23112 30058 23164 30064
rect 23020 27940 23072 27946
rect 23020 27882 23072 27888
rect 22926 27704 22982 27713
rect 22926 27639 22982 27648
rect 23032 27470 23060 27882
rect 23124 27674 23152 30058
rect 23216 28218 23244 30926
rect 23492 30802 23520 32438
rect 23480 30796 23532 30802
rect 23480 30738 23532 30744
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 23492 29646 23520 30194
rect 23584 30190 23612 33390
rect 23676 32910 23704 36518
rect 23848 36168 23900 36174
rect 23848 36110 23900 36116
rect 23860 35737 23888 36110
rect 23952 35766 23980 36876
rect 23940 35760 23992 35766
rect 23846 35728 23902 35737
rect 23756 35692 23808 35698
rect 23940 35702 23992 35708
rect 23846 35663 23902 35672
rect 24032 35692 24084 35698
rect 23756 35634 23808 35640
rect 24032 35634 24084 35640
rect 23768 35494 23796 35634
rect 23756 35488 23808 35494
rect 23756 35430 23808 35436
rect 23768 35086 23796 35430
rect 23848 35216 23900 35222
rect 23848 35158 23900 35164
rect 23756 35080 23808 35086
rect 23756 35022 23808 35028
rect 23860 34746 23888 35158
rect 24044 35018 24072 35634
rect 24032 35012 24084 35018
rect 24032 34954 24084 34960
rect 23848 34740 23900 34746
rect 23848 34682 23900 34688
rect 23940 34196 23992 34202
rect 23940 34138 23992 34144
rect 23952 34066 23980 34138
rect 23756 34060 23808 34066
rect 23756 34002 23808 34008
rect 23940 34060 23992 34066
rect 23940 34002 23992 34008
rect 23768 33114 23796 34002
rect 24136 33930 24164 37130
rect 24320 36854 24348 37334
rect 24490 37295 24546 37304
rect 24308 36848 24360 36854
rect 24308 36790 24360 36796
rect 24400 36712 24452 36718
rect 24400 36654 24452 36660
rect 24216 36168 24268 36174
rect 24216 36110 24268 36116
rect 24228 34610 24256 36110
rect 24306 35320 24362 35329
rect 24306 35255 24362 35264
rect 24216 34604 24268 34610
rect 24216 34546 24268 34552
rect 24228 34406 24256 34546
rect 24216 34400 24268 34406
rect 24216 34342 24268 34348
rect 24124 33924 24176 33930
rect 24124 33866 24176 33872
rect 24124 33652 24176 33658
rect 24124 33594 24176 33600
rect 24032 33516 24084 33522
rect 24032 33458 24084 33464
rect 23848 33448 23900 33454
rect 24044 33402 24072 33458
rect 24136 33454 24164 33594
rect 23848 33390 23900 33396
rect 23756 33108 23808 33114
rect 23756 33050 23808 33056
rect 23756 32972 23808 32978
rect 23756 32914 23808 32920
rect 23664 32904 23716 32910
rect 23664 32846 23716 32852
rect 23768 32570 23796 32914
rect 23860 32910 23888 33390
rect 23952 33374 24072 33402
rect 24124 33448 24176 33454
rect 24124 33390 24176 33396
rect 24214 33416 24270 33425
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23756 32564 23808 32570
rect 23756 32506 23808 32512
rect 23754 32328 23810 32337
rect 23754 32263 23810 32272
rect 23848 32292 23900 32298
rect 23662 31648 23718 31657
rect 23662 31583 23718 31592
rect 23676 31414 23704 31583
rect 23664 31408 23716 31414
rect 23664 31350 23716 31356
rect 23768 31113 23796 32263
rect 23848 32234 23900 32240
rect 23754 31104 23810 31113
rect 23754 31039 23810 31048
rect 23756 30932 23808 30938
rect 23756 30874 23808 30880
rect 23768 30394 23796 30874
rect 23756 30388 23808 30394
rect 23756 30330 23808 30336
rect 23860 30274 23888 32234
rect 23952 31754 23980 33374
rect 24214 33351 24270 33360
rect 24032 33312 24084 33318
rect 24228 33300 24256 33351
rect 24084 33272 24256 33300
rect 24032 33254 24084 33260
rect 24030 32736 24086 32745
rect 24030 32671 24086 32680
rect 24044 32434 24072 32671
rect 24032 32428 24084 32434
rect 24032 32370 24084 32376
rect 24124 32360 24176 32366
rect 24124 32302 24176 32308
rect 24136 32065 24164 32302
rect 24122 32056 24178 32065
rect 24122 31991 24178 32000
rect 23952 31748 24084 31754
rect 23952 31726 24032 31748
rect 24032 31690 24084 31696
rect 23940 31680 23992 31686
rect 23940 31622 23992 31628
rect 23952 30938 23980 31622
rect 24122 31104 24178 31113
rect 24122 31039 24178 31048
rect 23940 30932 23992 30938
rect 23940 30874 23992 30880
rect 23676 30246 23888 30274
rect 23572 30184 23624 30190
rect 23572 30126 23624 30132
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23584 29510 23612 30126
rect 23676 29646 23704 30246
rect 23952 29646 23980 30874
rect 24032 30592 24084 30598
rect 24032 30534 24084 30540
rect 23664 29640 23716 29646
rect 23664 29582 23716 29588
rect 23756 29640 23808 29646
rect 23756 29582 23808 29588
rect 23940 29640 23992 29646
rect 23940 29582 23992 29588
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 23572 29504 23624 29510
rect 23572 29446 23624 29452
rect 23204 28212 23256 28218
rect 23204 28154 23256 28160
rect 23308 28150 23336 29446
rect 23480 29096 23532 29102
rect 23480 29038 23532 29044
rect 23492 28490 23520 29038
rect 23676 28966 23704 29582
rect 23768 29034 23796 29582
rect 23756 29028 23808 29034
rect 23756 28970 23808 28976
rect 23664 28960 23716 28966
rect 23664 28902 23716 28908
rect 24044 28642 24072 30534
rect 23768 28626 24072 28642
rect 23768 28620 24084 28626
rect 23768 28614 24032 28620
rect 23388 28484 23440 28490
rect 23388 28426 23440 28432
rect 23480 28484 23532 28490
rect 23480 28426 23532 28432
rect 23296 28144 23348 28150
rect 23296 28086 23348 28092
rect 23204 27872 23256 27878
rect 23204 27814 23256 27820
rect 23112 27668 23164 27674
rect 23112 27610 23164 27616
rect 23216 27538 23244 27814
rect 23296 27668 23348 27674
rect 23296 27610 23348 27616
rect 23204 27532 23256 27538
rect 23204 27474 23256 27480
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 23124 27305 23152 27406
rect 23110 27296 23166 27305
rect 23110 27231 23166 27240
rect 23308 27146 23336 27610
rect 22848 27118 23336 27146
rect 22468 26988 22520 26994
rect 22520 26948 22692 26976
rect 22468 26930 22520 26936
rect 22664 26586 22692 26948
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 22480 26217 22508 26250
rect 22466 26208 22522 26217
rect 22466 26143 22522 26152
rect 22744 25696 22796 25702
rect 22744 25638 22796 25644
rect 22650 25528 22706 25537
rect 22650 25463 22706 25472
rect 22664 25362 22692 25463
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 22480 25129 22508 25230
rect 22560 25220 22612 25226
rect 22560 25162 22612 25168
rect 22466 25120 22522 25129
rect 22466 25055 22522 25064
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 22480 24274 22508 24346
rect 22572 24274 22600 25162
rect 22756 24993 22784 25638
rect 22848 25106 22876 27118
rect 23296 26988 23348 26994
rect 23296 26930 23348 26936
rect 22926 26888 22982 26897
rect 22926 26823 22982 26832
rect 22940 25265 22968 26823
rect 23308 26353 23336 26930
rect 23294 26344 23350 26353
rect 23294 26279 23350 26288
rect 23204 25832 23256 25838
rect 23204 25774 23256 25780
rect 23216 25378 23244 25774
rect 23032 25350 23244 25378
rect 22926 25256 22982 25265
rect 22926 25191 22982 25200
rect 22848 25078 22968 25106
rect 22742 24984 22798 24993
rect 22652 24948 22704 24954
rect 22742 24919 22798 24928
rect 22652 24890 22704 24896
rect 22664 24614 22692 24890
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 22468 24268 22520 24274
rect 22468 24210 22520 24216
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22376 23792 22428 23798
rect 22376 23734 22428 23740
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22836 23724 22888 23730
rect 22836 23666 22888 23672
rect 22192 23588 22244 23594
rect 22192 23530 22244 23536
rect 22008 23112 22060 23118
rect 22008 23054 22060 23060
rect 22204 22642 22232 23530
rect 22742 23080 22798 23089
rect 22742 23015 22798 23024
rect 22756 22982 22784 23015
rect 22744 22976 22796 22982
rect 22282 22944 22338 22953
rect 22848 22953 22876 23666
rect 22940 23118 22968 25078
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 22744 22918 22796 22924
rect 22834 22944 22890 22953
rect 22282 22879 22338 22888
rect 22834 22879 22890 22888
rect 22296 22642 22324 22879
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 21836 22066 21956 22094
rect 21638 21720 21694 21729
rect 21638 21655 21694 21664
rect 21652 21418 21680 21655
rect 21640 21412 21692 21418
rect 21640 21354 21692 21360
rect 21640 19984 21692 19990
rect 21640 19926 21692 19932
rect 21652 18766 21680 19926
rect 21732 19916 21784 19922
rect 21732 19858 21784 19864
rect 21744 19310 21772 19858
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21744 18970 21772 19246
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21652 17202 21680 18022
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20824 15502 20852 16050
rect 21652 15502 21680 17138
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 21744 16114 21772 16526
rect 21836 16182 21864 22066
rect 22204 21962 22232 22578
rect 22284 22500 22336 22506
rect 22284 22442 22336 22448
rect 22296 22166 22324 22442
rect 22572 22234 22600 22714
rect 22744 22636 22796 22642
rect 22744 22578 22796 22584
rect 22468 22228 22520 22234
rect 22468 22170 22520 22176
rect 22560 22228 22612 22234
rect 22560 22170 22612 22176
rect 22284 22160 22336 22166
rect 22284 22102 22336 22108
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 22284 21956 22336 21962
rect 22284 21898 22336 21904
rect 22296 21842 22324 21898
rect 22112 21814 22324 21842
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 22020 21146 22048 21286
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 22112 21010 22140 21814
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22204 21010 22232 21626
rect 22388 21554 22416 21830
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 22192 21004 22244 21010
rect 22192 20946 22244 20952
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 22112 20330 22140 20810
rect 22204 20466 22232 20946
rect 22296 20602 22324 21490
rect 22480 21350 22508 22170
rect 22756 22030 22784 22578
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 22848 22098 22876 22510
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22744 21616 22796 21622
rect 22664 21576 22744 21604
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22466 21176 22522 21185
rect 22572 21146 22600 21490
rect 22466 21111 22522 21120
rect 22560 21140 22612 21146
rect 22480 21026 22508 21111
rect 22560 21082 22612 21088
rect 22480 20998 22600 21026
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22468 20460 22520 20466
rect 22468 20402 22520 20408
rect 22100 20324 22152 20330
rect 22100 20266 22152 20272
rect 22480 20262 22508 20402
rect 22192 20256 22244 20262
rect 22468 20256 22520 20262
rect 22192 20198 22244 20204
rect 22388 20216 22468 20244
rect 22204 19961 22232 20198
rect 22190 19952 22246 19961
rect 22008 19916 22060 19922
rect 22190 19887 22246 19896
rect 22008 19858 22060 19864
rect 22020 19310 22048 19858
rect 22204 19854 22232 19887
rect 22388 19854 22416 20216
rect 22468 20198 22520 20204
rect 22192 19848 22244 19854
rect 22098 19816 22154 19825
rect 22192 19790 22244 19796
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22098 19751 22154 19760
rect 22284 19780 22336 19786
rect 22112 19446 22140 19751
rect 22284 19722 22336 19728
rect 22296 19666 22324 19722
rect 22296 19638 22508 19666
rect 22100 19440 22152 19446
rect 22100 19382 22152 19388
rect 22008 19304 22060 19310
rect 22480 19281 22508 19638
rect 22008 19246 22060 19252
rect 22466 19272 22522 19281
rect 21916 19236 21968 19242
rect 21916 19178 21968 19184
rect 22376 19236 22428 19242
rect 22466 19207 22522 19216
rect 22376 19178 22428 19184
rect 21928 17270 21956 19178
rect 22388 18902 22416 19178
rect 22376 18896 22428 18902
rect 22376 18838 22428 18844
rect 22008 18828 22060 18834
rect 22008 18770 22060 18776
rect 22020 17882 22048 18770
rect 22480 18290 22508 19207
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22192 18216 22244 18222
rect 22192 18158 22244 18164
rect 22008 17876 22060 17882
rect 22008 17818 22060 17824
rect 22008 17604 22060 17610
rect 22008 17546 22060 17552
rect 21916 17264 21968 17270
rect 21916 17206 21968 17212
rect 22020 16794 22048 17546
rect 22204 17270 22232 18158
rect 22296 17338 22324 18226
rect 22388 17882 22416 18226
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22192 17264 22244 17270
rect 22190 17232 22192 17241
rect 22376 17264 22428 17270
rect 22244 17232 22246 17241
rect 22376 17206 22428 17212
rect 22190 17167 22246 17176
rect 22008 16788 22060 16794
rect 22008 16730 22060 16736
rect 21824 16176 21876 16182
rect 21824 16118 21876 16124
rect 21732 16108 21784 16114
rect 21732 16050 21784 16056
rect 22020 15570 22048 16730
rect 22388 16590 22416 17206
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 22388 15026 22416 16526
rect 22572 15706 22600 20998
rect 22664 20874 22692 21576
rect 22744 21558 22796 21564
rect 22744 21412 22796 21418
rect 22744 21354 22796 21360
rect 22836 21412 22888 21418
rect 22836 21354 22888 21360
rect 22652 20868 22704 20874
rect 22652 20810 22704 20816
rect 22650 20632 22706 20641
rect 22756 20618 22784 21354
rect 22848 21049 22876 21354
rect 22834 21040 22890 21049
rect 22834 20975 22890 20984
rect 22928 21004 22980 21010
rect 22928 20946 22980 20952
rect 22940 20806 22968 20946
rect 22928 20800 22980 20806
rect 22928 20742 22980 20748
rect 22756 20590 22876 20618
rect 22650 20567 22706 20576
rect 22664 18170 22692 20567
rect 22848 20466 22876 20590
rect 22940 20505 22968 20742
rect 22926 20496 22982 20505
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22836 20460 22888 20466
rect 22926 20431 22982 20440
rect 22836 20402 22888 20408
rect 22756 19990 22784 20402
rect 22744 19984 22796 19990
rect 22744 19926 22796 19932
rect 22848 18766 22876 20402
rect 23032 19938 23060 25350
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23124 20641 23152 25230
rect 23308 23866 23336 26279
rect 23400 25770 23428 28426
rect 23492 28082 23520 28426
rect 23572 28416 23624 28422
rect 23572 28358 23624 28364
rect 23584 28082 23612 28358
rect 23768 28257 23796 28614
rect 24032 28562 24084 28568
rect 23848 28552 23900 28558
rect 23846 28520 23848 28529
rect 23900 28520 23902 28529
rect 24136 28506 24164 31039
rect 24228 30161 24256 33272
rect 24320 30802 24348 35255
rect 24412 34202 24440 36654
rect 24400 34196 24452 34202
rect 24400 34138 24452 34144
rect 24400 33924 24452 33930
rect 24400 33866 24452 33872
rect 24412 33318 24440 33866
rect 24400 33312 24452 33318
rect 24400 33254 24452 33260
rect 24504 33114 24532 37295
rect 24688 36242 24716 38111
rect 24964 37262 24992 39200
rect 28276 39166 28304 39200
rect 31588 39166 31616 39200
rect 28264 39160 28316 39166
rect 28264 39102 28316 39108
rect 31576 39160 31628 39166
rect 31576 39102 31628 39108
rect 30010 38856 30066 38865
rect 26884 38820 26936 38826
rect 30010 38791 30066 38800
rect 26884 38762 26936 38768
rect 26422 38720 26478 38729
rect 26422 38655 26478 38664
rect 26792 38684 26844 38690
rect 25964 38412 26016 38418
rect 25964 38354 26016 38360
rect 25870 38176 25926 38185
rect 25870 38111 25926 38120
rect 25504 38072 25556 38078
rect 25504 38014 25556 38020
rect 25516 37670 25544 38014
rect 25504 37664 25556 37670
rect 25504 37606 25556 37612
rect 25780 37460 25832 37466
rect 25780 37402 25832 37408
rect 24952 37256 25004 37262
rect 24952 37198 25004 37204
rect 25320 37188 25372 37194
rect 25320 37130 25372 37136
rect 25332 36553 25360 37130
rect 25502 36952 25558 36961
rect 25502 36887 25558 36896
rect 25516 36854 25544 36887
rect 25504 36848 25556 36854
rect 25504 36790 25556 36796
rect 25318 36544 25374 36553
rect 25318 36479 25374 36488
rect 24676 36236 24728 36242
rect 25412 36236 25464 36242
rect 24676 36178 24728 36184
rect 25240 36196 25412 36224
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 24596 35737 24624 36110
rect 24676 36100 24728 36106
rect 24676 36042 24728 36048
rect 25044 36100 25096 36106
rect 25044 36042 25096 36048
rect 24582 35728 24638 35737
rect 24582 35663 24638 35672
rect 24688 35018 24716 36042
rect 24860 36032 24912 36038
rect 24860 35974 24912 35980
rect 24872 35873 24900 35974
rect 24858 35864 24914 35873
rect 24858 35799 24914 35808
rect 24768 35624 24820 35630
rect 24768 35566 24820 35572
rect 24676 35012 24728 35018
rect 24676 34954 24728 34960
rect 24584 33924 24636 33930
rect 24584 33866 24636 33872
rect 24596 33522 24624 33866
rect 24584 33516 24636 33522
rect 24584 33458 24636 33464
rect 24582 33144 24638 33153
rect 24492 33108 24544 33114
rect 24582 33079 24638 33088
rect 24492 33050 24544 33056
rect 24400 32904 24452 32910
rect 24400 32846 24452 32852
rect 24490 32872 24546 32881
rect 24308 30796 24360 30802
rect 24308 30738 24360 30744
rect 24214 30152 24270 30161
rect 24214 30087 24270 30096
rect 24214 29336 24270 29345
rect 24214 29271 24270 29280
rect 24228 29170 24256 29271
rect 24216 29164 24268 29170
rect 24216 29106 24268 29112
rect 24228 28762 24256 29106
rect 24216 28756 24268 28762
rect 24216 28698 24268 28704
rect 24308 28756 24360 28762
rect 24308 28698 24360 28704
rect 23846 28455 23902 28464
rect 24044 28478 24164 28506
rect 23754 28248 23810 28257
rect 23754 28183 23810 28192
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23572 28076 23624 28082
rect 23624 28036 23704 28064
rect 23572 28018 23624 28024
rect 23480 27940 23532 27946
rect 23480 27882 23532 27888
rect 23492 27674 23520 27882
rect 23480 27668 23532 27674
rect 23480 27610 23532 27616
rect 23572 27396 23624 27402
rect 23572 27338 23624 27344
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23388 25764 23440 25770
rect 23388 25706 23440 25712
rect 23492 24206 23520 27270
rect 23584 26518 23612 27338
rect 23572 26512 23624 26518
rect 23572 26454 23624 26460
rect 23572 26308 23624 26314
rect 23572 26250 23624 26256
rect 23584 25498 23612 26250
rect 23572 25492 23624 25498
rect 23572 25434 23624 25440
rect 23676 25430 23704 28036
rect 23768 26926 23796 28183
rect 23860 28150 23888 28455
rect 23938 28248 23994 28257
rect 23938 28183 23994 28192
rect 23848 28144 23900 28150
rect 23848 28086 23900 28092
rect 23846 27296 23902 27305
rect 23846 27231 23902 27240
rect 23860 27062 23888 27231
rect 23848 27056 23900 27062
rect 23848 26998 23900 27004
rect 23756 26920 23808 26926
rect 23756 26862 23808 26868
rect 23756 26784 23808 26790
rect 23756 26726 23808 26732
rect 23768 26382 23796 26726
rect 23848 26512 23900 26518
rect 23848 26454 23900 26460
rect 23756 26376 23808 26382
rect 23860 26353 23888 26454
rect 23756 26318 23808 26324
rect 23846 26344 23902 26353
rect 23846 26279 23902 26288
rect 23952 25673 23980 28183
rect 24044 27849 24072 28478
rect 24124 28212 24176 28218
rect 24124 28154 24176 28160
rect 24030 27840 24086 27849
rect 24030 27775 24086 27784
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 23938 25664 23994 25673
rect 23938 25599 23994 25608
rect 24044 25430 24072 27406
rect 24136 27062 24164 28154
rect 24124 27056 24176 27062
rect 24124 26998 24176 27004
rect 24214 26208 24270 26217
rect 24214 26143 24270 26152
rect 24124 25764 24176 25770
rect 24124 25706 24176 25712
rect 23664 25424 23716 25430
rect 23664 25366 23716 25372
rect 24032 25424 24084 25430
rect 24032 25366 24084 25372
rect 23572 25356 23624 25362
rect 23572 25298 23624 25304
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23584 24154 23612 25298
rect 23938 24848 23994 24857
rect 23938 24783 23940 24792
rect 23992 24783 23994 24792
rect 23940 24754 23992 24760
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 23584 24126 23704 24154
rect 23860 24138 23888 24550
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23308 23730 23336 23802
rect 23296 23724 23348 23730
rect 23296 23666 23348 23672
rect 23202 23624 23258 23633
rect 23202 23559 23258 23568
rect 23216 22681 23244 23559
rect 23202 22672 23258 22681
rect 23202 22607 23258 22616
rect 23308 22574 23336 23666
rect 23584 23322 23612 24006
rect 23572 23316 23624 23322
rect 23572 23258 23624 23264
rect 23676 23186 23704 24126
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 23940 24132 23992 24138
rect 23940 24074 23992 24080
rect 23756 23316 23808 23322
rect 23756 23258 23808 23264
rect 23664 23180 23716 23186
rect 23664 23122 23716 23128
rect 23768 23118 23796 23258
rect 23756 23112 23808 23118
rect 23662 23080 23718 23089
rect 23756 23054 23808 23060
rect 23662 23015 23664 23024
rect 23716 23015 23718 23024
rect 23664 22986 23716 22992
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 23296 22432 23348 22438
rect 23296 22374 23348 22380
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23204 22160 23256 22166
rect 23204 22102 23256 22108
rect 23216 21894 23244 22102
rect 23204 21888 23256 21894
rect 23204 21830 23256 21836
rect 23110 20632 23166 20641
rect 23110 20567 23166 20576
rect 23112 20460 23164 20466
rect 23112 20402 23164 20408
rect 22940 19910 23060 19938
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22756 18358 22784 18566
rect 22744 18352 22796 18358
rect 22744 18294 22796 18300
rect 22664 18142 22784 18170
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22664 16794 22692 17138
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22756 16454 22784 18142
rect 22848 17678 22876 18702
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22940 15450 22968 19910
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 23032 19718 23060 19790
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 23032 18698 23060 19654
rect 23124 18970 23152 20402
rect 23216 19961 23244 21830
rect 23308 21078 23336 22374
rect 23676 22094 23704 22374
rect 23860 22234 23888 24074
rect 23952 22982 23980 24074
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 23400 22066 23704 22094
rect 23400 22030 23428 22066
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23400 21690 23428 21966
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 23296 21072 23348 21078
rect 23296 21014 23348 21020
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23308 20058 23336 20402
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23202 19952 23258 19961
rect 23202 19887 23258 19896
rect 23400 19718 23428 20878
rect 23492 20058 23520 20878
rect 23480 20052 23532 20058
rect 23480 19994 23532 20000
rect 23584 19922 23612 21490
rect 23676 20466 23704 22066
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 23952 21690 23980 21966
rect 23848 21684 23900 21690
rect 23848 21626 23900 21632
rect 23940 21684 23992 21690
rect 23940 21626 23992 21632
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23768 21146 23796 21490
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 23860 20602 23888 21626
rect 23848 20596 23900 20602
rect 23848 20538 23900 20544
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 23572 19916 23624 19922
rect 23572 19858 23624 19864
rect 23676 19854 23704 20402
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 23952 19802 23980 21626
rect 24044 20505 24072 22578
rect 24136 22001 24164 25706
rect 24228 23202 24256 26143
rect 24320 25809 24348 28698
rect 24412 27554 24440 32846
rect 24490 32807 24546 32816
rect 24504 31686 24532 32807
rect 24596 32609 24624 33079
rect 24688 32842 24716 34954
rect 24780 32910 24808 35566
rect 25056 35086 25084 36042
rect 25136 36032 25188 36038
rect 25136 35974 25188 35980
rect 25148 35698 25176 35974
rect 25240 35873 25268 36196
rect 25412 36178 25464 36184
rect 25504 36236 25556 36242
rect 25504 36178 25556 36184
rect 25226 35864 25282 35873
rect 25226 35799 25282 35808
rect 25136 35692 25188 35698
rect 25136 35634 25188 35640
rect 25148 35222 25176 35634
rect 25240 35630 25268 35799
rect 25516 35698 25544 36178
rect 25792 35737 25820 37402
rect 25778 35728 25834 35737
rect 25504 35692 25556 35698
rect 25778 35663 25834 35672
rect 25504 35634 25556 35640
rect 25228 35624 25280 35630
rect 25228 35566 25280 35572
rect 25596 35624 25648 35630
rect 25596 35566 25648 35572
rect 25136 35216 25188 35222
rect 25136 35158 25188 35164
rect 25044 35080 25096 35086
rect 25044 35022 25096 35028
rect 25148 34950 25176 35158
rect 25240 35154 25268 35566
rect 25504 35556 25556 35562
rect 25504 35498 25556 35504
rect 25516 35154 25544 35498
rect 25228 35148 25280 35154
rect 25228 35090 25280 35096
rect 25504 35148 25556 35154
rect 25504 35090 25556 35096
rect 25412 35012 25464 35018
rect 25412 34954 25464 34960
rect 25136 34944 25188 34950
rect 25136 34886 25188 34892
rect 25134 34776 25190 34785
rect 25134 34711 25190 34720
rect 24860 34196 24912 34202
rect 24860 34138 24912 34144
rect 24952 34196 25004 34202
rect 24952 34138 25004 34144
rect 24872 33590 24900 34138
rect 24964 33998 24992 34138
rect 24952 33992 25004 33998
rect 24952 33934 25004 33940
rect 24860 33584 24912 33590
rect 24860 33526 24912 33532
rect 24768 32904 24820 32910
rect 24768 32846 24820 32852
rect 24676 32836 24728 32842
rect 24676 32778 24728 32784
rect 24582 32600 24638 32609
rect 24780 32570 24808 32846
rect 24582 32535 24638 32544
rect 24768 32564 24820 32570
rect 24768 32506 24820 32512
rect 24768 32360 24820 32366
rect 24768 32302 24820 32308
rect 24584 32292 24636 32298
rect 24584 32234 24636 32240
rect 24676 32292 24728 32298
rect 24676 32234 24728 32240
rect 24596 31754 24624 32234
rect 24584 31748 24636 31754
rect 24584 31690 24636 31696
rect 24492 31680 24544 31686
rect 24492 31622 24544 31628
rect 24688 31385 24716 32234
rect 24780 32026 24808 32302
rect 24768 32020 24820 32026
rect 24768 31962 24820 31968
rect 24674 31376 24730 31385
rect 24674 31311 24730 31320
rect 24766 30968 24822 30977
rect 24766 30903 24822 30912
rect 24780 30802 24808 30903
rect 24768 30796 24820 30802
rect 24768 30738 24820 30744
rect 24768 30660 24820 30666
rect 24768 30602 24820 30608
rect 24584 30320 24636 30326
rect 24584 30262 24636 30268
rect 24492 30252 24544 30258
rect 24492 30194 24544 30200
rect 24504 29850 24532 30194
rect 24596 30054 24624 30262
rect 24780 30138 24808 30602
rect 24872 30258 24900 33526
rect 25044 33516 25096 33522
rect 25044 33458 25096 33464
rect 25056 33114 25084 33458
rect 25148 33318 25176 34711
rect 25228 34468 25280 34474
rect 25228 34410 25280 34416
rect 25240 33318 25268 34410
rect 25320 34128 25372 34134
rect 25320 34070 25372 34076
rect 25332 33998 25360 34070
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 25424 33930 25452 34954
rect 25608 34678 25636 35566
rect 25688 34944 25740 34950
rect 25688 34886 25740 34892
rect 25596 34672 25648 34678
rect 25596 34614 25648 34620
rect 25596 34468 25648 34474
rect 25596 34410 25648 34416
rect 25504 34400 25556 34406
rect 25504 34342 25556 34348
rect 25516 34241 25544 34342
rect 25502 34232 25558 34241
rect 25502 34167 25558 34176
rect 25608 33946 25636 34410
rect 25412 33924 25464 33930
rect 25412 33866 25464 33872
rect 25516 33918 25636 33946
rect 25700 33946 25728 34886
rect 25792 34202 25820 35663
rect 25884 35290 25912 38111
rect 25976 35766 26004 38354
rect 26148 38344 26200 38350
rect 26148 38286 26200 38292
rect 26160 37233 26188 38286
rect 26332 37868 26384 37874
rect 26332 37810 26384 37816
rect 26240 37664 26292 37670
rect 26240 37606 26292 37612
rect 26146 37224 26202 37233
rect 26146 37159 26202 37168
rect 26252 37126 26280 37606
rect 26240 37120 26292 37126
rect 26240 37062 26292 37068
rect 26240 36712 26292 36718
rect 26240 36654 26292 36660
rect 26148 36644 26200 36650
rect 26148 36586 26200 36592
rect 26056 36168 26108 36174
rect 26056 36110 26108 36116
rect 26068 36038 26096 36110
rect 26056 36032 26108 36038
rect 26056 35974 26108 35980
rect 25964 35760 26016 35766
rect 26016 35720 26096 35748
rect 25964 35702 26016 35708
rect 25964 35488 26016 35494
rect 26068 35465 26096 35720
rect 25964 35430 26016 35436
rect 26054 35456 26110 35465
rect 25872 35284 25924 35290
rect 25872 35226 25924 35232
rect 25884 35018 25912 35226
rect 25872 35012 25924 35018
rect 25872 34954 25924 34960
rect 25872 34468 25924 34474
rect 25872 34410 25924 34416
rect 25780 34196 25832 34202
rect 25780 34138 25832 34144
rect 25700 33918 25820 33946
rect 25410 33552 25466 33561
rect 25332 33510 25410 33538
rect 25136 33312 25188 33318
rect 25136 33254 25188 33260
rect 25228 33312 25280 33318
rect 25228 33254 25280 33260
rect 25332 33153 25360 33510
rect 25410 33487 25466 33496
rect 25318 33144 25374 33153
rect 25044 33108 25096 33114
rect 25318 33079 25374 33088
rect 25044 33050 25096 33056
rect 25332 33046 25360 33079
rect 25228 33040 25280 33046
rect 25042 33008 25098 33017
rect 25228 32982 25280 32988
rect 25320 33040 25372 33046
rect 25320 32982 25372 32988
rect 25042 32943 25098 32952
rect 25056 32910 25084 32943
rect 25240 32910 25268 32982
rect 24952 32904 25004 32910
rect 24950 32872 24952 32881
rect 25044 32904 25096 32910
rect 25004 32872 25006 32881
rect 25044 32846 25096 32852
rect 25228 32904 25280 32910
rect 25228 32846 25280 32852
rect 24950 32807 25006 32816
rect 25056 32298 25084 32846
rect 25136 32428 25188 32434
rect 25136 32370 25188 32376
rect 25044 32292 25096 32298
rect 25044 32234 25096 32240
rect 24952 31884 25004 31890
rect 24952 31826 25004 31832
rect 25044 31884 25096 31890
rect 25044 31826 25096 31832
rect 24964 31793 24992 31826
rect 24950 31784 25006 31793
rect 25056 31754 25084 31826
rect 24950 31719 25006 31728
rect 25044 31748 25096 31754
rect 25044 31690 25096 31696
rect 24952 31204 25004 31210
rect 24952 31146 25004 31152
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24780 30110 24900 30138
rect 24584 30048 24636 30054
rect 24584 29990 24636 29996
rect 24492 29844 24544 29850
rect 24492 29786 24544 29792
rect 24504 28994 24532 29786
rect 24768 29708 24820 29714
rect 24768 29650 24820 29656
rect 24780 29306 24808 29650
rect 24872 29646 24900 30110
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24584 29300 24636 29306
rect 24768 29300 24820 29306
rect 24636 29260 24716 29288
rect 24584 29242 24636 29248
rect 24504 28966 24624 28994
rect 24596 28694 24624 28966
rect 24584 28688 24636 28694
rect 24584 28630 24636 28636
rect 24596 28558 24624 28630
rect 24584 28552 24636 28558
rect 24490 28520 24546 28529
rect 24584 28494 24636 28500
rect 24490 28455 24546 28464
rect 24504 27985 24532 28455
rect 24490 27976 24546 27985
rect 24490 27911 24546 27920
rect 24688 27878 24716 29260
rect 24768 29242 24820 29248
rect 24872 29170 24900 29582
rect 24964 29306 24992 31146
rect 25044 30320 25096 30326
rect 25044 30262 25096 30268
rect 25056 29617 25084 30262
rect 25148 29714 25176 32370
rect 25240 30977 25268 32846
rect 25320 32836 25372 32842
rect 25320 32778 25372 32784
rect 25332 32434 25360 32778
rect 25516 32570 25544 33918
rect 25596 33856 25648 33862
rect 25596 33798 25648 33804
rect 25688 33856 25740 33862
rect 25688 33798 25740 33804
rect 25608 33522 25636 33798
rect 25700 33590 25728 33798
rect 25688 33584 25740 33590
rect 25688 33526 25740 33532
rect 25596 33516 25648 33522
rect 25596 33458 25648 33464
rect 25688 33448 25740 33454
rect 25688 33390 25740 33396
rect 25700 33318 25728 33390
rect 25688 33312 25740 33318
rect 25688 33254 25740 33260
rect 25686 33008 25742 33017
rect 25608 32966 25686 32994
rect 25412 32564 25464 32570
rect 25412 32506 25464 32512
rect 25504 32564 25556 32570
rect 25504 32506 25556 32512
rect 25320 32428 25372 32434
rect 25320 32370 25372 32376
rect 25332 32337 25360 32370
rect 25424 32366 25452 32506
rect 25412 32360 25464 32366
rect 25318 32328 25374 32337
rect 25412 32302 25464 32308
rect 25318 32263 25374 32272
rect 25412 32224 25464 32230
rect 25318 32192 25374 32201
rect 25412 32166 25464 32172
rect 25318 32127 25374 32136
rect 25332 31958 25360 32127
rect 25320 31952 25372 31958
rect 25424 31929 25452 32166
rect 25320 31894 25372 31900
rect 25410 31920 25466 31929
rect 25410 31855 25412 31864
rect 25464 31855 25466 31864
rect 25412 31826 25464 31832
rect 25608 31521 25636 32966
rect 25686 32943 25742 32952
rect 25792 32450 25820 33918
rect 25884 33454 25912 34410
rect 25872 33448 25924 33454
rect 25872 33390 25924 33396
rect 25872 33040 25924 33046
rect 25872 32982 25924 32988
rect 25700 32422 25820 32450
rect 25700 31958 25728 32422
rect 25780 32360 25832 32366
rect 25780 32302 25832 32308
rect 25688 31952 25740 31958
rect 25688 31894 25740 31900
rect 25792 31890 25820 32302
rect 25780 31884 25832 31890
rect 25780 31826 25832 31832
rect 25594 31512 25650 31521
rect 25594 31447 25650 31456
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25226 30968 25282 30977
rect 25226 30903 25282 30912
rect 25516 30734 25544 31282
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 25608 30326 25636 31282
rect 25686 31240 25742 31249
rect 25686 31175 25742 31184
rect 25700 30705 25728 31175
rect 25792 30802 25820 31826
rect 25780 30796 25832 30802
rect 25780 30738 25832 30744
rect 25686 30696 25742 30705
rect 25686 30631 25742 30640
rect 25596 30320 25648 30326
rect 25596 30262 25648 30268
rect 25596 30184 25648 30190
rect 25594 30152 25596 30161
rect 25648 30152 25650 30161
rect 25228 30116 25280 30122
rect 25228 30058 25280 30064
rect 25320 30116 25372 30122
rect 25594 30087 25650 30096
rect 25320 30058 25372 30064
rect 25240 29714 25268 30058
rect 25136 29708 25188 29714
rect 25136 29650 25188 29656
rect 25228 29708 25280 29714
rect 25228 29650 25280 29656
rect 25042 29608 25098 29617
rect 25042 29543 25098 29552
rect 25042 29336 25098 29345
rect 24952 29300 25004 29306
rect 25042 29271 25098 29280
rect 24952 29242 25004 29248
rect 25056 29170 25084 29271
rect 24860 29164 24912 29170
rect 24860 29106 24912 29112
rect 25044 29164 25096 29170
rect 25044 29106 25096 29112
rect 24766 29064 24822 29073
rect 25042 29064 25098 29073
rect 24822 29022 24900 29050
rect 24766 28999 24822 29008
rect 24872 28994 24900 29022
rect 25042 28999 25098 29008
rect 24872 28966 24992 28994
rect 24768 28484 24820 28490
rect 24768 28426 24820 28432
rect 24492 27872 24544 27878
rect 24492 27814 24544 27820
rect 24676 27872 24728 27878
rect 24676 27814 24728 27820
rect 24504 27674 24532 27814
rect 24492 27668 24544 27674
rect 24492 27610 24544 27616
rect 24412 27538 24532 27554
rect 24412 27532 24544 27538
rect 24412 27526 24492 27532
rect 24492 27474 24544 27480
rect 24400 27396 24452 27402
rect 24400 27338 24452 27344
rect 24306 25800 24362 25809
rect 24306 25735 24362 25744
rect 24308 23588 24360 23594
rect 24308 23530 24360 23536
rect 24320 23497 24348 23530
rect 24306 23488 24362 23497
rect 24306 23423 24362 23432
rect 24228 23174 24348 23202
rect 24320 23118 24348 23174
rect 24216 23112 24268 23118
rect 24216 23054 24268 23060
rect 24308 23112 24360 23118
rect 24308 23054 24360 23060
rect 24228 22710 24256 23054
rect 24308 22976 24360 22982
rect 24308 22918 24360 22924
rect 24216 22704 24268 22710
rect 24216 22646 24268 22652
rect 24122 21992 24178 22001
rect 24122 21927 24178 21936
rect 24124 21888 24176 21894
rect 24124 21830 24176 21836
rect 24216 21888 24268 21894
rect 24216 21830 24268 21836
rect 24136 21622 24164 21830
rect 24124 21616 24176 21622
rect 24124 21558 24176 21564
rect 24228 21010 24256 21830
rect 24320 21570 24348 22918
rect 24412 21690 24440 27338
rect 24504 27062 24532 27474
rect 24584 27396 24636 27402
rect 24584 27338 24636 27344
rect 24492 27056 24544 27062
rect 24492 26998 24544 27004
rect 24492 26784 24544 26790
rect 24596 26761 24624 27338
rect 24492 26726 24544 26732
rect 24582 26752 24638 26761
rect 24504 25344 24532 26726
rect 24582 26687 24638 26696
rect 24596 26518 24624 26687
rect 24584 26512 24636 26518
rect 24584 26454 24636 26460
rect 24688 26382 24716 27814
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24584 25356 24636 25362
rect 24504 25316 24584 25344
rect 24584 25298 24636 25304
rect 24596 24698 24624 25298
rect 24688 24818 24716 26318
rect 24780 25838 24808 28426
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 24872 26790 24900 28018
rect 24860 26784 24912 26790
rect 24860 26726 24912 26732
rect 24858 26480 24914 26489
rect 24858 26415 24914 26424
rect 24872 26382 24900 26415
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24768 25832 24820 25838
rect 24768 25774 24820 25780
rect 24780 25242 24808 25774
rect 24872 25362 24900 26318
rect 24964 25673 24992 28966
rect 24950 25664 25006 25673
rect 24950 25599 25006 25608
rect 25056 25430 25084 28999
rect 25332 28082 25360 30058
rect 25412 30048 25464 30054
rect 25412 29990 25464 29996
rect 25424 28558 25452 29990
rect 25596 29640 25648 29646
rect 25596 29582 25648 29588
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 25412 28552 25464 28558
rect 25412 28494 25464 28500
rect 25412 28416 25464 28422
rect 25412 28358 25464 28364
rect 25424 28082 25452 28358
rect 25320 28076 25372 28082
rect 25320 28018 25372 28024
rect 25412 28076 25464 28082
rect 25412 28018 25464 28024
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 25228 27328 25280 27334
rect 25228 27270 25280 27276
rect 25240 27130 25268 27270
rect 25228 27124 25280 27130
rect 25228 27066 25280 27072
rect 25228 26988 25280 26994
rect 25228 26930 25280 26936
rect 25240 26761 25268 26930
rect 25226 26752 25282 26761
rect 25226 26687 25282 26696
rect 25134 26480 25190 26489
rect 25134 26415 25190 26424
rect 25148 26314 25176 26415
rect 25136 26308 25188 26314
rect 25136 26250 25188 26256
rect 25228 26308 25280 26314
rect 25332 26296 25360 27406
rect 25280 26268 25360 26296
rect 25228 26250 25280 26256
rect 24952 25424 25004 25430
rect 24952 25366 25004 25372
rect 25044 25424 25096 25430
rect 25044 25366 25096 25372
rect 24860 25356 24912 25362
rect 24860 25298 24912 25304
rect 24780 25226 24900 25242
rect 24780 25220 24912 25226
rect 24780 25214 24860 25220
rect 24860 25162 24912 25168
rect 24858 24984 24914 24993
rect 24858 24919 24914 24928
rect 24676 24812 24728 24818
rect 24676 24754 24728 24760
rect 24596 24670 24716 24698
rect 24584 23792 24636 23798
rect 24584 23734 24636 23740
rect 24596 23089 24624 23734
rect 24582 23080 24638 23089
rect 24582 23015 24638 23024
rect 24492 22976 24544 22982
rect 24492 22918 24544 22924
rect 24504 22778 24532 22918
rect 24492 22772 24544 22778
rect 24492 22714 24544 22720
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24320 21542 24440 21570
rect 24308 21480 24360 21486
rect 24308 21422 24360 21428
rect 24320 21321 24348 21422
rect 24306 21312 24362 21321
rect 24306 21247 24362 21256
rect 24216 21004 24268 21010
rect 24216 20946 24268 20952
rect 24030 20496 24086 20505
rect 24030 20431 24086 20440
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 24044 19961 24072 19994
rect 24030 19952 24086 19961
rect 24030 19887 24086 19896
rect 24228 19854 24256 20946
rect 24216 19848 24268 19854
rect 23480 19780 23532 19786
rect 23480 19722 23532 19728
rect 23388 19712 23440 19718
rect 23388 19654 23440 19660
rect 23204 19508 23256 19514
rect 23204 19450 23256 19456
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23020 18692 23072 18698
rect 23020 18634 23072 18640
rect 23216 18578 23244 19450
rect 23492 19378 23520 19722
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23032 18550 23244 18578
rect 23032 16998 23060 18550
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 23216 17678 23244 18362
rect 23308 17814 23336 18702
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23400 18154 23428 18566
rect 23492 18426 23520 19110
rect 23676 18748 23704 19790
rect 23952 19774 24072 19802
rect 24216 19790 24268 19796
rect 23754 19408 23810 19417
rect 23754 19343 23756 19352
rect 23808 19343 23810 19352
rect 23756 19314 23808 19320
rect 23768 18970 23796 19314
rect 23940 19304 23992 19310
rect 23940 19246 23992 19252
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23848 18896 23900 18902
rect 23848 18838 23900 18844
rect 23756 18760 23808 18766
rect 23676 18720 23756 18748
rect 23756 18702 23808 18708
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23572 18216 23624 18222
rect 23572 18158 23624 18164
rect 23388 18148 23440 18154
rect 23388 18090 23440 18096
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23296 17808 23348 17814
rect 23296 17750 23348 17756
rect 23204 17672 23256 17678
rect 23110 17640 23166 17649
rect 23204 17614 23256 17620
rect 23110 17575 23166 17584
rect 23124 17134 23152 17575
rect 23216 17377 23244 17614
rect 23202 17368 23258 17377
rect 23202 17303 23258 17312
rect 23388 17196 23440 17202
rect 23492 17184 23520 18022
rect 23584 17882 23612 18158
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23860 17184 23888 18838
rect 23952 18766 23980 19246
rect 24044 19145 24072 19774
rect 24320 19666 24348 21247
rect 24136 19638 24348 19666
rect 24030 19136 24086 19145
rect 24030 19071 24086 19080
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 23952 17610 23980 18702
rect 24044 18290 24072 19071
rect 24136 18873 24164 19638
rect 24412 19446 24440 21542
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 24504 21185 24532 21490
rect 24596 21350 24624 23015
rect 24688 22506 24716 24670
rect 24872 24274 24900 24919
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24964 24206 24992 25366
rect 25044 25152 25096 25158
rect 25044 25094 25096 25100
rect 25136 25152 25188 25158
rect 25136 25094 25188 25100
rect 25056 24313 25084 25094
rect 25042 24304 25098 24313
rect 25042 24239 25098 24248
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24780 23118 24808 23258
rect 24860 23180 24912 23186
rect 24964 23168 24992 24142
rect 25148 23798 25176 25094
rect 25240 24993 25268 26250
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25226 24984 25282 24993
rect 25226 24919 25282 24928
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 24912 23140 24992 23168
rect 24860 23122 24912 23128
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24676 22500 24728 22506
rect 24676 22442 24728 22448
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 24490 21176 24546 21185
rect 24490 21111 24546 21120
rect 24400 19440 24452 19446
rect 24400 19382 24452 19388
rect 24308 19372 24360 19378
rect 24308 19314 24360 19320
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 24216 19304 24268 19310
rect 24216 19246 24268 19252
rect 24122 18864 24178 18873
rect 24122 18799 24178 18808
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 23940 17604 23992 17610
rect 23940 17546 23992 17552
rect 23440 17156 23520 17184
rect 23768 17156 23888 17184
rect 23388 17138 23440 17144
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 23204 17128 23256 17134
rect 23204 17070 23256 17076
rect 23020 16992 23072 16998
rect 23020 16934 23072 16940
rect 23032 16046 23060 16934
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 23112 15972 23164 15978
rect 23112 15914 23164 15920
rect 22848 15422 22968 15450
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 21100 14618 21128 14962
rect 22284 14952 22336 14958
rect 22284 14894 22336 14900
rect 22100 14816 22152 14822
rect 22100 14758 22152 14764
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 22112 14346 22140 14758
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 20720 13796 20772 13802
rect 20720 13738 20772 13744
rect 20732 13394 20760 13738
rect 22008 13728 22060 13734
rect 22008 13670 22060 13676
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 20548 12850 20576 13262
rect 22020 13258 22048 13670
rect 22008 13252 22060 13258
rect 22008 13194 22060 13200
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20364 12442 20392 12786
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 19444 11218 19472 12242
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19444 10674 19472 11154
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 20548 10674 20576 12786
rect 20916 11898 20944 12854
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22008 12640 22060 12646
rect 22008 12582 22060 12588
rect 22020 12238 22048 12582
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21744 11898 21772 12038
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20640 10742 20668 11494
rect 20916 10810 20944 11834
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22020 11150 22048 11494
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20628 10736 20680 10742
rect 20628 10678 20680 10684
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 22112 10266 22140 12786
rect 22296 12646 22324 14894
rect 22388 14414 22416 14962
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 22376 14272 22428 14278
rect 22376 14214 22428 14220
rect 22388 14074 22416 14214
rect 22480 14074 22508 15098
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22388 13530 22416 13874
rect 22376 13524 22428 13530
rect 22376 13466 22428 13472
rect 22388 13190 22416 13466
rect 22664 13394 22692 14350
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22296 12374 22324 12582
rect 22284 12368 22336 12374
rect 22284 12310 22336 12316
rect 22664 11898 22692 13330
rect 22756 12850 22784 13806
rect 22848 13734 22876 15422
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22940 15026 22968 15302
rect 22928 15020 22980 15026
rect 22928 14962 22980 14968
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22940 12918 22968 14010
rect 22928 12912 22980 12918
rect 22928 12854 22980 12860
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22192 11620 22244 11626
rect 22192 11562 22244 11568
rect 22204 10606 22232 11562
rect 22388 11354 22416 11698
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22388 10674 22416 11290
rect 22664 10674 22692 11834
rect 22756 11694 22784 12786
rect 23032 12306 23060 14010
rect 23124 13802 23152 15914
rect 23216 14006 23244 17070
rect 23480 16516 23532 16522
rect 23480 16458 23532 16464
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23400 15162 23428 15438
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23388 14952 23440 14958
rect 23388 14894 23440 14900
rect 23204 14000 23256 14006
rect 23204 13942 23256 13948
rect 23400 13938 23428 14894
rect 23492 14278 23520 16458
rect 23768 16182 23796 17156
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23756 16176 23808 16182
rect 23756 16118 23808 16124
rect 23756 15428 23808 15434
rect 23756 15370 23808 15376
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23480 14272 23532 14278
rect 23480 14214 23532 14220
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23112 13796 23164 13802
rect 23112 13738 23164 13744
rect 23204 13728 23256 13734
rect 23204 13670 23256 13676
rect 23216 12986 23244 13670
rect 23400 13326 23428 13874
rect 23584 13530 23612 13942
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23572 13252 23624 13258
rect 23572 13194 23624 13200
rect 23584 12986 23612 13194
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23112 12436 23164 12442
rect 23112 12378 23164 12384
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 23032 10810 23060 12038
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 22284 10600 22336 10606
rect 22284 10542 22336 10548
rect 22296 10266 22324 10542
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 23124 10062 23152 12378
rect 23216 11762 23244 12922
rect 23676 12714 23704 15098
rect 23768 14822 23796 15370
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23860 13240 23888 16934
rect 23952 16590 23980 17546
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 24136 16522 24164 18799
rect 24228 18086 24256 19246
rect 24320 18426 24348 19314
rect 24400 18692 24452 18698
rect 24400 18634 24452 18640
rect 24308 18420 24360 18426
rect 24308 18362 24360 18368
rect 24306 18320 24362 18329
rect 24306 18255 24308 18264
rect 24360 18255 24362 18264
rect 24308 18226 24360 18232
rect 24412 18222 24440 18634
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 24216 18080 24268 18086
rect 24216 18022 24268 18028
rect 24412 16590 24440 18158
rect 24504 17338 24532 19314
rect 24596 19145 24624 21286
rect 24688 20874 24716 22442
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 24872 22166 24900 22374
rect 24768 22160 24820 22166
rect 24768 22102 24820 22108
rect 24860 22160 24912 22166
rect 24860 22102 24912 22108
rect 24780 22030 24808 22102
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24676 20868 24728 20874
rect 24676 20810 24728 20816
rect 24872 20806 24900 22102
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 25056 21457 25084 21490
rect 25042 21448 25098 21457
rect 25042 21383 25098 21392
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 25044 20800 25096 20806
rect 25044 20742 25096 20748
rect 24860 19984 24912 19990
rect 24860 19926 24912 19932
rect 24768 19712 24820 19718
rect 24768 19654 24820 19660
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24688 19378 24716 19450
rect 24780 19378 24808 19654
rect 24676 19372 24728 19378
rect 24676 19314 24728 19320
rect 24768 19372 24820 19378
rect 24768 19314 24820 19320
rect 24582 19136 24638 19145
rect 24582 19071 24638 19080
rect 24596 18902 24624 19071
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24584 18896 24636 18902
rect 24584 18838 24636 18844
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 18154 24624 18566
rect 24584 18148 24636 18154
rect 24584 18090 24636 18096
rect 24596 17678 24624 18090
rect 24676 17808 24728 17814
rect 24676 17750 24728 17756
rect 24688 17678 24716 17750
rect 24780 17678 24808 18906
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24676 17672 24728 17678
rect 24768 17672 24820 17678
rect 24676 17614 24728 17620
rect 24766 17640 24768 17649
rect 24820 17640 24822 17649
rect 24688 17524 24716 17614
rect 24766 17575 24822 17584
rect 24872 17592 24900 19926
rect 24964 19417 24992 20742
rect 25056 19514 25084 20742
rect 25148 20097 25176 23462
rect 25240 23050 25268 24919
rect 25332 24614 25360 25230
rect 25424 25129 25452 28018
rect 25516 28014 25544 29106
rect 25608 28218 25636 29582
rect 25700 29238 25728 30631
rect 25780 30592 25832 30598
rect 25780 30534 25832 30540
rect 25792 30002 25820 30534
rect 25884 30122 25912 32982
rect 25872 30116 25924 30122
rect 25872 30058 25924 30064
rect 25792 29974 25912 30002
rect 25780 29776 25832 29782
rect 25780 29718 25832 29724
rect 25688 29232 25740 29238
rect 25688 29174 25740 29180
rect 25688 29028 25740 29034
rect 25688 28970 25740 28976
rect 25700 28490 25728 28970
rect 25688 28484 25740 28490
rect 25688 28426 25740 28432
rect 25596 28212 25648 28218
rect 25596 28154 25648 28160
rect 25504 28008 25556 28014
rect 25504 27950 25556 27956
rect 25608 27946 25636 28154
rect 25596 27940 25648 27946
rect 25596 27882 25648 27888
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25504 26240 25556 26246
rect 25504 26182 25556 26188
rect 25410 25120 25466 25129
rect 25410 25055 25466 25064
rect 25516 24970 25544 26182
rect 25608 25945 25636 26930
rect 25594 25936 25650 25945
rect 25594 25871 25650 25880
rect 25688 25492 25740 25498
rect 25688 25434 25740 25440
rect 25594 25256 25650 25265
rect 25594 25191 25650 25200
rect 25424 24942 25544 24970
rect 25320 24608 25372 24614
rect 25320 24550 25372 24556
rect 25424 23225 25452 24942
rect 25502 24712 25558 24721
rect 25502 24647 25504 24656
rect 25556 24647 25558 24656
rect 25504 24618 25556 24624
rect 25608 24120 25636 25191
rect 25700 24274 25728 25434
rect 25792 24886 25820 29718
rect 25884 28914 25912 29974
rect 25976 29714 26004 35430
rect 26054 35391 26110 35400
rect 26160 35306 26188 36586
rect 26252 36378 26280 36654
rect 26240 36372 26292 36378
rect 26240 36314 26292 36320
rect 26240 36100 26292 36106
rect 26240 36042 26292 36048
rect 26252 35562 26280 36042
rect 26240 35556 26292 35562
rect 26240 35498 26292 35504
rect 26068 35278 26188 35306
rect 26068 33318 26096 35278
rect 26344 35086 26372 37810
rect 26332 35080 26384 35086
rect 26332 35022 26384 35028
rect 26332 34944 26384 34950
rect 26332 34886 26384 34892
rect 26146 34368 26202 34377
rect 26146 34303 26202 34312
rect 26160 33998 26188 34303
rect 26238 34232 26294 34241
rect 26238 34167 26294 34176
rect 26252 33998 26280 34167
rect 26344 34105 26372 34886
rect 26436 34610 26464 38655
rect 26792 38626 26844 38632
rect 26608 37256 26660 37262
rect 26608 37198 26660 37204
rect 26516 37120 26568 37126
rect 26516 37062 26568 37068
rect 26528 34785 26556 37062
rect 26620 36650 26648 37198
rect 26608 36644 26660 36650
rect 26608 36586 26660 36592
rect 26608 36168 26660 36174
rect 26608 36110 26660 36116
rect 26620 35630 26648 36110
rect 26698 35728 26754 35737
rect 26698 35663 26754 35672
rect 26608 35624 26660 35630
rect 26608 35566 26660 35572
rect 26514 34776 26570 34785
rect 26514 34711 26570 34720
rect 26620 34678 26648 35566
rect 26712 35562 26740 35663
rect 26804 35630 26832 38626
rect 26896 37126 26924 38762
rect 27894 38584 27950 38593
rect 27894 38519 27950 38528
rect 27528 37936 27580 37942
rect 27528 37878 27580 37884
rect 26976 37868 27028 37874
rect 26976 37810 27028 37816
rect 26988 37330 27016 37810
rect 26976 37324 27028 37330
rect 26976 37266 27028 37272
rect 27252 37256 27304 37262
rect 27252 37198 27304 37204
rect 26884 37120 26936 37126
rect 26884 37062 26936 37068
rect 26896 36174 26924 37062
rect 26884 36168 26936 36174
rect 26884 36110 26936 36116
rect 26976 36032 27028 36038
rect 26976 35974 27028 35980
rect 26792 35624 26844 35630
rect 26792 35566 26844 35572
rect 26700 35556 26752 35562
rect 26700 35498 26752 35504
rect 26804 35290 26832 35566
rect 26884 35488 26936 35494
rect 26884 35430 26936 35436
rect 26896 35329 26924 35430
rect 26882 35320 26938 35329
rect 26792 35284 26844 35290
rect 26882 35255 26938 35264
rect 26792 35226 26844 35232
rect 26896 35086 26924 35255
rect 26884 35080 26936 35086
rect 26884 35022 26936 35028
rect 26608 34672 26660 34678
rect 26608 34614 26660 34620
rect 26424 34604 26476 34610
rect 26424 34546 26476 34552
rect 26792 34604 26844 34610
rect 26792 34546 26844 34552
rect 26330 34096 26386 34105
rect 26330 34031 26386 34040
rect 26148 33992 26200 33998
rect 26148 33934 26200 33940
rect 26240 33992 26292 33998
rect 26240 33934 26292 33940
rect 26148 33516 26200 33522
rect 26148 33458 26200 33464
rect 26056 33312 26108 33318
rect 26056 33254 26108 33260
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 26068 31890 26096 32846
rect 26160 32774 26188 33458
rect 26344 33402 26372 34031
rect 26424 33992 26476 33998
rect 26804 33946 26832 34546
rect 26882 34096 26938 34105
rect 26882 34031 26938 34040
rect 26424 33934 26476 33940
rect 26436 33425 26464 33934
rect 26516 33924 26568 33930
rect 26516 33866 26568 33872
rect 26620 33918 26832 33946
rect 26252 33374 26372 33402
rect 26422 33416 26478 33425
rect 26148 32768 26200 32774
rect 26148 32710 26200 32716
rect 26056 31884 26108 31890
rect 26252 31872 26280 33374
rect 26422 33351 26478 33360
rect 26332 33312 26384 33318
rect 26330 33280 26332 33289
rect 26384 33280 26386 33289
rect 26330 33215 26386 33224
rect 26528 32230 26556 33866
rect 26516 32224 26568 32230
rect 26330 32192 26386 32201
rect 26516 32166 26568 32172
rect 26330 32127 26386 32136
rect 26056 31826 26108 31832
rect 26160 31844 26280 31872
rect 26056 31680 26108 31686
rect 26056 31622 26108 31628
rect 26068 30870 26096 31622
rect 26160 31249 26188 31844
rect 26344 31804 26372 32127
rect 26516 32020 26568 32026
rect 26516 31962 26568 31968
rect 26528 31890 26556 31962
rect 26424 31884 26476 31890
rect 26424 31826 26476 31832
rect 26516 31884 26568 31890
rect 26516 31826 26568 31832
rect 26252 31776 26372 31804
rect 26146 31240 26202 31249
rect 26146 31175 26202 31184
rect 26148 31136 26200 31142
rect 26148 31078 26200 31084
rect 26056 30864 26108 30870
rect 26056 30806 26108 30812
rect 26068 30433 26096 30806
rect 26054 30424 26110 30433
rect 26054 30359 26110 30368
rect 26056 30320 26108 30326
rect 26056 30262 26108 30268
rect 25964 29708 26016 29714
rect 25964 29650 26016 29656
rect 25884 28886 26004 28914
rect 25872 28484 25924 28490
rect 25872 28426 25924 28432
rect 25884 27606 25912 28426
rect 25976 28422 26004 28886
rect 26068 28762 26096 30262
rect 26056 28756 26108 28762
rect 26056 28698 26108 28704
rect 26160 28558 26188 31078
rect 26252 30394 26280 31776
rect 26330 31240 26386 31249
rect 26330 31175 26386 31184
rect 26344 30598 26372 31175
rect 26436 30666 26464 31826
rect 26620 31754 26648 33918
rect 26792 33516 26844 33522
rect 26792 33458 26844 33464
rect 26700 33108 26752 33114
rect 26700 33050 26752 33056
rect 26528 31726 26648 31754
rect 26424 30660 26476 30666
rect 26424 30602 26476 30608
rect 26332 30592 26384 30598
rect 26332 30534 26384 30540
rect 26240 30388 26292 30394
rect 26240 30330 26292 30336
rect 26332 30116 26384 30122
rect 26332 30058 26384 30064
rect 26238 29200 26294 29209
rect 26238 29135 26294 29144
rect 26252 29102 26280 29135
rect 26240 29096 26292 29102
rect 26240 29038 26292 29044
rect 26240 28620 26292 28626
rect 26240 28562 26292 28568
rect 26148 28552 26200 28558
rect 26054 28520 26110 28529
rect 26252 28529 26280 28562
rect 26148 28494 26200 28500
rect 26238 28520 26294 28529
rect 26054 28455 26110 28464
rect 25964 28416 26016 28422
rect 25964 28358 26016 28364
rect 26068 28150 26096 28455
rect 26056 28144 26108 28150
rect 26056 28086 26108 28092
rect 26160 28014 26188 28494
rect 26238 28455 26294 28464
rect 26344 28370 26372 30058
rect 26424 29300 26476 29306
rect 26424 29242 26476 29248
rect 26436 29073 26464 29242
rect 26422 29064 26478 29073
rect 26422 28999 26478 29008
rect 26528 28966 26556 31726
rect 26608 30728 26660 30734
rect 26608 30670 26660 30676
rect 26620 29578 26648 30670
rect 26608 29572 26660 29578
rect 26608 29514 26660 29520
rect 26606 29336 26662 29345
rect 26606 29271 26608 29280
rect 26660 29271 26662 29280
rect 26608 29242 26660 29248
rect 26516 28960 26568 28966
rect 26516 28902 26568 28908
rect 26424 28620 26476 28626
rect 26424 28562 26476 28568
rect 26252 28342 26372 28370
rect 26056 28008 26108 28014
rect 26056 27950 26108 27956
rect 26148 28008 26200 28014
rect 26148 27950 26200 27956
rect 26068 27674 26096 27950
rect 26148 27872 26200 27878
rect 26148 27814 26200 27820
rect 26056 27668 26108 27674
rect 26056 27610 26108 27616
rect 25872 27600 25924 27606
rect 25872 27542 25924 27548
rect 26054 27568 26110 27577
rect 26054 27503 26056 27512
rect 26108 27503 26110 27512
rect 26056 27474 26108 27480
rect 26056 27056 26108 27062
rect 26056 26998 26108 27004
rect 25872 26852 25924 26858
rect 25872 26794 25924 26800
rect 25884 26314 25912 26794
rect 25964 26580 26016 26586
rect 25964 26522 26016 26528
rect 25872 26308 25924 26314
rect 25872 26250 25924 26256
rect 25976 26194 26004 26522
rect 25884 26166 26004 26194
rect 25884 25498 25912 26166
rect 25964 25900 26016 25906
rect 25964 25842 26016 25848
rect 25976 25809 26004 25842
rect 25962 25800 26018 25809
rect 25962 25735 26018 25744
rect 25962 25664 26018 25673
rect 25962 25599 26018 25608
rect 25872 25492 25924 25498
rect 25872 25434 25924 25440
rect 25872 25356 25924 25362
rect 25872 25298 25924 25304
rect 25780 24880 25832 24886
rect 25780 24822 25832 24828
rect 25688 24268 25740 24274
rect 25688 24210 25740 24216
rect 25884 24206 25912 25298
rect 25976 24818 26004 25599
rect 26068 24818 26096 26998
rect 26160 26450 26188 27814
rect 26252 27402 26280 28342
rect 26332 27872 26384 27878
rect 26332 27814 26384 27820
rect 26344 27713 26372 27814
rect 26330 27704 26386 27713
rect 26330 27639 26386 27648
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 26332 27396 26384 27402
rect 26332 27338 26384 27344
rect 26148 26444 26200 26450
rect 26148 26386 26200 26392
rect 26146 26344 26202 26353
rect 26344 26314 26372 27338
rect 26436 27130 26464 28562
rect 26514 27704 26570 27713
rect 26514 27639 26570 27648
rect 26424 27124 26476 27130
rect 26424 27066 26476 27072
rect 26528 26314 26556 27639
rect 26608 27464 26660 27470
rect 26608 27406 26660 27412
rect 26146 26279 26202 26288
rect 26240 26308 26292 26314
rect 26160 24954 26188 26279
rect 26240 26250 26292 26256
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26516 26308 26568 26314
rect 26516 26250 26568 26256
rect 26252 25430 26280 26250
rect 26344 25770 26372 26250
rect 26514 25936 26570 25945
rect 26514 25871 26570 25880
rect 26332 25764 26384 25770
rect 26332 25706 26384 25712
rect 26240 25424 26292 25430
rect 26240 25366 26292 25372
rect 26528 25294 26556 25871
rect 26620 25294 26648 27406
rect 26712 26994 26740 33050
rect 26804 33046 26832 33458
rect 26792 33040 26844 33046
rect 26792 32982 26844 32988
rect 26896 32978 26924 34031
rect 26884 32972 26936 32978
rect 26884 32914 26936 32920
rect 26884 32020 26936 32026
rect 26884 31962 26936 31968
rect 26790 31512 26846 31521
rect 26790 31447 26846 31456
rect 26804 30326 26832 31447
rect 26896 30598 26924 31962
rect 26988 31958 27016 35974
rect 27066 35456 27122 35465
rect 27066 35391 27122 35400
rect 27080 35086 27108 35391
rect 27160 35284 27212 35290
rect 27160 35226 27212 35232
rect 27068 35080 27120 35086
rect 27068 35022 27120 35028
rect 27172 34932 27200 35226
rect 27264 35154 27292 37198
rect 27434 36544 27490 36553
rect 27434 36479 27490 36488
rect 27342 35864 27398 35873
rect 27342 35799 27344 35808
rect 27396 35799 27398 35808
rect 27344 35770 27396 35776
rect 27342 35320 27398 35329
rect 27342 35255 27398 35264
rect 27252 35148 27304 35154
rect 27252 35090 27304 35096
rect 27250 35048 27306 35057
rect 27250 34983 27252 34992
rect 27304 34983 27306 34992
rect 27252 34954 27304 34960
rect 27080 34904 27200 34932
rect 27356 34921 27384 35255
rect 27342 34912 27398 34921
rect 26976 31952 27028 31958
rect 26976 31894 27028 31900
rect 27080 31657 27108 34904
rect 27342 34847 27398 34856
rect 27160 34672 27212 34678
rect 27160 34614 27212 34620
rect 27172 33998 27200 34614
rect 27252 34400 27304 34406
rect 27252 34342 27304 34348
rect 27160 33992 27212 33998
rect 27160 33934 27212 33940
rect 27160 33856 27212 33862
rect 27160 33798 27212 33804
rect 27172 33318 27200 33798
rect 27264 33658 27292 34342
rect 27448 34134 27476 36479
rect 27540 35057 27568 37878
rect 27620 37460 27672 37466
rect 27620 37402 27672 37408
rect 27632 36825 27660 37402
rect 27712 36848 27764 36854
rect 27618 36816 27674 36825
rect 27712 36790 27764 36796
rect 27618 36751 27674 36760
rect 27620 36712 27672 36718
rect 27620 36654 27672 36660
rect 27632 36242 27660 36654
rect 27724 36378 27752 36790
rect 27712 36372 27764 36378
rect 27712 36314 27764 36320
rect 27620 36236 27672 36242
rect 27620 36178 27672 36184
rect 27804 36168 27856 36174
rect 27804 36110 27856 36116
rect 27620 36100 27672 36106
rect 27620 36042 27672 36048
rect 27526 35048 27582 35057
rect 27526 34983 27582 34992
rect 27540 34610 27568 34983
rect 27528 34604 27580 34610
rect 27528 34546 27580 34552
rect 27436 34128 27488 34134
rect 27632 34082 27660 36042
rect 27816 35834 27844 36110
rect 27804 35828 27856 35834
rect 27804 35770 27856 35776
rect 27816 35630 27844 35770
rect 27804 35624 27856 35630
rect 27804 35566 27856 35572
rect 27804 34944 27856 34950
rect 27908 34921 27936 38519
rect 28998 37496 29054 37505
rect 28998 37431 29054 37440
rect 28448 37392 28500 37398
rect 28448 37334 28500 37340
rect 28080 37324 28132 37330
rect 28080 37266 28132 37272
rect 28092 36786 28120 37266
rect 28264 37256 28316 37262
rect 28264 37198 28316 37204
rect 28080 36780 28132 36786
rect 28080 36722 28132 36728
rect 28276 36122 28304 37198
rect 28356 37120 28408 37126
rect 28356 37062 28408 37068
rect 28000 36094 28304 36122
rect 27804 34886 27856 34892
rect 27894 34912 27950 34921
rect 27816 34678 27844 34886
rect 27894 34847 27950 34856
rect 27894 34776 27950 34785
rect 27894 34711 27950 34720
rect 27908 34678 27936 34711
rect 27804 34672 27856 34678
rect 27804 34614 27856 34620
rect 27896 34672 27948 34678
rect 27896 34614 27948 34620
rect 27804 34536 27856 34542
rect 27804 34478 27856 34484
rect 27712 34196 27764 34202
rect 27712 34138 27764 34144
rect 27436 34070 27488 34076
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 27344 33652 27396 33658
rect 27344 33594 27396 33600
rect 27356 33561 27384 33594
rect 27342 33552 27398 33561
rect 27264 33510 27342 33538
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 27066 31648 27122 31657
rect 27066 31583 27122 31592
rect 26976 31340 27028 31346
rect 26976 31282 27028 31288
rect 26884 30592 26936 30598
rect 26884 30534 26936 30540
rect 26792 30320 26844 30326
rect 26792 30262 26844 30268
rect 26988 30025 27016 31282
rect 27080 31113 27108 31583
rect 27172 31210 27200 33254
rect 27264 31906 27292 33510
rect 27448 33522 27476 34070
rect 27540 34054 27660 34082
rect 27540 33998 27568 34054
rect 27528 33992 27580 33998
rect 27528 33934 27580 33940
rect 27620 33992 27672 33998
rect 27620 33934 27672 33940
rect 27526 33688 27582 33697
rect 27526 33623 27582 33632
rect 27540 33522 27568 33623
rect 27342 33487 27398 33496
rect 27436 33516 27488 33522
rect 27436 33458 27488 33464
rect 27528 33516 27580 33522
rect 27528 33458 27580 33464
rect 27344 33312 27396 33318
rect 27344 33254 27396 33260
rect 27356 32502 27384 33254
rect 27540 32994 27568 33458
rect 27448 32966 27568 32994
rect 27448 32910 27476 32966
rect 27436 32904 27488 32910
rect 27436 32846 27488 32852
rect 27528 32904 27580 32910
rect 27528 32846 27580 32852
rect 27540 32609 27568 32846
rect 27526 32600 27582 32609
rect 27526 32535 27582 32544
rect 27344 32496 27396 32502
rect 27344 32438 27396 32444
rect 27528 32428 27580 32434
rect 27528 32370 27580 32376
rect 27540 31958 27568 32370
rect 27632 32026 27660 33934
rect 27620 32020 27672 32026
rect 27620 31962 27672 31968
rect 27528 31952 27580 31958
rect 27264 31878 27384 31906
rect 27528 31894 27580 31900
rect 27252 31680 27304 31686
rect 27252 31622 27304 31628
rect 27160 31204 27212 31210
rect 27160 31146 27212 31152
rect 27066 31104 27122 31113
rect 27066 31039 27122 31048
rect 27068 30796 27120 30802
rect 27068 30738 27120 30744
rect 27080 30326 27108 30738
rect 27068 30320 27120 30326
rect 27068 30262 27120 30268
rect 26974 30016 27030 30025
rect 26974 29951 27030 29960
rect 27080 29850 27108 30262
rect 27160 30048 27212 30054
rect 27160 29990 27212 29996
rect 27068 29844 27120 29850
rect 27068 29786 27120 29792
rect 26976 29640 27028 29646
rect 26976 29582 27028 29588
rect 26884 29164 26936 29170
rect 26884 29106 26936 29112
rect 26792 27668 26844 27674
rect 26792 27610 26844 27616
rect 26700 26988 26752 26994
rect 26700 26930 26752 26936
rect 26712 25974 26740 26930
rect 26804 26217 26832 27610
rect 26896 26858 26924 29106
rect 26988 28762 27016 29582
rect 27080 29170 27108 29786
rect 27172 29753 27200 29990
rect 27158 29744 27214 29753
rect 27264 29730 27292 31622
rect 27356 30870 27384 31878
rect 27724 31754 27752 34138
rect 27816 33930 27844 34478
rect 27908 34406 27936 34614
rect 27896 34400 27948 34406
rect 27896 34342 27948 34348
rect 27804 33924 27856 33930
rect 27804 33866 27856 33872
rect 27896 33924 27948 33930
rect 27896 33866 27948 33872
rect 27908 33454 27936 33866
rect 27896 33448 27948 33454
rect 27896 33390 27948 33396
rect 27908 33318 27936 33390
rect 27896 33312 27948 33318
rect 27896 33254 27948 33260
rect 27896 33040 27948 33046
rect 27896 32982 27948 32988
rect 27908 32881 27936 32982
rect 27894 32872 27950 32881
rect 27894 32807 27950 32816
rect 27804 32428 27856 32434
rect 27804 32370 27856 32376
rect 27712 31748 27764 31754
rect 27712 31690 27764 31696
rect 27620 31408 27672 31414
rect 27620 31350 27672 31356
rect 27528 31272 27580 31278
rect 27528 31214 27580 31220
rect 27540 30938 27568 31214
rect 27528 30932 27580 30938
rect 27528 30874 27580 30880
rect 27344 30864 27396 30870
rect 27632 30841 27660 31350
rect 27344 30806 27396 30812
rect 27618 30832 27674 30841
rect 27618 30767 27674 30776
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27344 30388 27396 30394
rect 27344 30330 27396 30336
rect 27356 30190 27384 30330
rect 27344 30184 27396 30190
rect 27344 30126 27396 30132
rect 27448 30054 27476 30670
rect 27620 30592 27672 30598
rect 27620 30534 27672 30540
rect 27712 30592 27764 30598
rect 27712 30534 27764 30540
rect 27526 30288 27582 30297
rect 27526 30223 27582 30232
rect 27344 30048 27396 30054
rect 27344 29990 27396 29996
rect 27436 30048 27488 30054
rect 27436 29990 27488 29996
rect 27356 29850 27384 29990
rect 27434 29880 27490 29889
rect 27344 29844 27396 29850
rect 27434 29815 27490 29824
rect 27344 29786 27396 29792
rect 27264 29702 27384 29730
rect 27158 29679 27214 29688
rect 27252 29640 27304 29646
rect 27252 29582 27304 29588
rect 27160 29572 27212 29578
rect 27160 29514 27212 29520
rect 27172 29345 27200 29514
rect 27158 29336 27214 29345
rect 27158 29271 27214 29280
rect 27158 29200 27214 29209
rect 27068 29164 27120 29170
rect 27158 29135 27214 29144
rect 27068 29106 27120 29112
rect 27068 28960 27120 28966
rect 27068 28902 27120 28908
rect 27080 28762 27108 28902
rect 27172 28801 27200 29135
rect 27158 28792 27214 28801
rect 26976 28756 27028 28762
rect 26976 28698 27028 28704
rect 27068 28756 27120 28762
rect 27158 28727 27214 28736
rect 27068 28698 27120 28704
rect 27080 27577 27108 28698
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27172 28082 27200 28494
rect 27160 28076 27212 28082
rect 27160 28018 27212 28024
rect 27066 27568 27122 27577
rect 27066 27503 27122 27512
rect 27264 27418 27292 29582
rect 27356 29170 27384 29702
rect 27448 29578 27476 29815
rect 27436 29572 27488 29578
rect 27436 29514 27488 29520
rect 27344 29164 27396 29170
rect 27344 29106 27396 29112
rect 27344 28960 27396 28966
rect 27344 28902 27396 28908
rect 27356 27538 27384 28902
rect 27344 27532 27396 27538
rect 27344 27474 27396 27480
rect 27172 27390 27292 27418
rect 27172 27305 27200 27390
rect 27252 27328 27304 27334
rect 27158 27296 27214 27305
rect 27252 27270 27304 27276
rect 27158 27231 27214 27240
rect 27264 26994 27292 27270
rect 27252 26988 27304 26994
rect 27252 26930 27304 26936
rect 27448 26926 27476 29514
rect 27540 28558 27568 30223
rect 27528 28552 27580 28558
rect 27528 28494 27580 28500
rect 27528 28212 27580 28218
rect 27528 28154 27580 28160
rect 27540 27577 27568 28154
rect 27526 27568 27582 27577
rect 27526 27503 27582 27512
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 26884 26852 26936 26858
rect 26884 26794 26936 26800
rect 26790 26208 26846 26217
rect 26790 26143 26846 26152
rect 26700 25968 26752 25974
rect 26700 25910 26752 25916
rect 26700 25832 26752 25838
rect 26700 25774 26752 25780
rect 26516 25288 26568 25294
rect 26516 25230 26568 25236
rect 26608 25288 26660 25294
rect 26608 25230 26660 25236
rect 26148 24948 26200 24954
rect 26148 24890 26200 24896
rect 25964 24812 26016 24818
rect 25964 24754 26016 24760
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 26240 24812 26292 24818
rect 26292 24772 26372 24800
rect 26240 24754 26292 24760
rect 25976 24721 26004 24754
rect 25962 24712 26018 24721
rect 25962 24647 26018 24656
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25872 24200 25924 24206
rect 25872 24142 25924 24148
rect 25688 24132 25740 24138
rect 25608 24092 25688 24120
rect 25688 24074 25740 24080
rect 25872 24064 25924 24070
rect 25872 24006 25924 24012
rect 25504 23724 25556 23730
rect 25504 23666 25556 23672
rect 25410 23216 25466 23225
rect 25320 23180 25372 23186
rect 25410 23151 25466 23160
rect 25320 23122 25372 23128
rect 25228 23044 25280 23050
rect 25228 22986 25280 22992
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25240 22545 25268 22578
rect 25226 22536 25282 22545
rect 25226 22471 25282 22480
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25240 20602 25268 20946
rect 25332 20806 25360 23122
rect 25516 23118 25544 23666
rect 25780 23520 25832 23526
rect 25780 23462 25832 23468
rect 25504 23112 25556 23118
rect 25504 23054 25556 23060
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25700 22574 25728 23054
rect 25688 22568 25740 22574
rect 25688 22510 25740 22516
rect 25412 22500 25464 22506
rect 25412 22442 25464 22448
rect 25596 22500 25648 22506
rect 25596 22442 25648 22448
rect 25424 21962 25452 22442
rect 25412 21956 25464 21962
rect 25412 21898 25464 21904
rect 25608 21622 25636 22442
rect 25686 22400 25742 22409
rect 25686 22335 25742 22344
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25424 20534 25452 21490
rect 25596 21480 25648 21486
rect 25596 21422 25648 21428
rect 25412 20528 25464 20534
rect 25412 20470 25464 20476
rect 25228 20392 25280 20398
rect 25228 20334 25280 20340
rect 25134 20088 25190 20097
rect 25134 20023 25190 20032
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 24950 19408 25006 19417
rect 24950 19343 25006 19352
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 25148 18698 25176 19110
rect 25240 18834 25268 20334
rect 25424 19854 25452 20470
rect 25412 19848 25464 19854
rect 25412 19790 25464 19796
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 25228 18692 25280 18698
rect 25228 18634 25280 18640
rect 25240 18358 25268 18634
rect 25228 18352 25280 18358
rect 25228 18294 25280 18300
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 25516 17814 25544 18022
rect 25504 17808 25556 17814
rect 25504 17750 25556 17756
rect 24872 17564 24992 17592
rect 24688 17496 24900 17524
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 24872 16833 24900 17496
rect 24858 16824 24914 16833
rect 24858 16759 24914 16768
rect 24400 16584 24452 16590
rect 24400 16526 24452 16532
rect 24582 16552 24638 16561
rect 24124 16516 24176 16522
rect 24582 16487 24638 16496
rect 24124 16458 24176 16464
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 23940 16176 23992 16182
rect 23940 16118 23992 16124
rect 23952 14618 23980 16118
rect 23940 14612 23992 14618
rect 23940 14554 23992 14560
rect 24044 14414 24072 16186
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 23952 13530 23980 13806
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 24044 13326 24072 14214
rect 24320 13462 24348 16050
rect 24596 15434 24624 16487
rect 24964 15502 24992 17564
rect 25516 16658 25544 17750
rect 25504 16652 25556 16658
rect 25504 16594 25556 16600
rect 25608 16250 25636 21422
rect 25700 21146 25728 22335
rect 25688 21140 25740 21146
rect 25688 21082 25740 21088
rect 25700 20466 25728 21082
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25686 19136 25742 19145
rect 25686 19071 25742 19080
rect 25700 18465 25728 19071
rect 25686 18456 25742 18465
rect 25686 18391 25742 18400
rect 25700 18290 25728 18391
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25792 17678 25820 23462
rect 25884 21486 25912 24006
rect 25976 23798 26004 24550
rect 25964 23792 26016 23798
rect 25964 23734 26016 23740
rect 26068 22642 26096 24754
rect 26238 24712 26294 24721
rect 26238 24647 26294 24656
rect 26252 24206 26280 24647
rect 26240 24200 26292 24206
rect 26146 24168 26202 24177
rect 26240 24142 26292 24148
rect 26146 24103 26202 24112
rect 26160 23730 26188 24103
rect 26344 23866 26372 24772
rect 26424 24608 26476 24614
rect 26424 24550 26476 24556
rect 26332 23860 26384 23866
rect 26332 23802 26384 23808
rect 26148 23724 26200 23730
rect 26148 23666 26200 23672
rect 26148 22976 26200 22982
rect 26148 22918 26200 22924
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 26056 22636 26108 22642
rect 26056 22578 26108 22584
rect 25976 22545 26004 22578
rect 25962 22536 26018 22545
rect 26068 22506 26096 22578
rect 25962 22471 26018 22480
rect 26056 22500 26108 22506
rect 26056 22442 26108 22448
rect 26160 21706 26188 22918
rect 26068 21678 26188 21706
rect 26068 21486 26096 21678
rect 26148 21616 26200 21622
rect 26148 21558 26200 21564
rect 25872 21480 25924 21486
rect 25872 21422 25924 21428
rect 26056 21480 26108 21486
rect 26056 21422 26108 21428
rect 25872 21140 25924 21146
rect 26056 21140 26108 21146
rect 25872 21082 25924 21088
rect 25976 21100 26056 21128
rect 25884 20874 25912 21082
rect 25872 20868 25924 20874
rect 25872 20810 25924 20816
rect 25976 20806 26004 21100
rect 26056 21082 26108 21088
rect 25964 20800 26016 20806
rect 25964 20742 26016 20748
rect 25976 20534 26004 20742
rect 25964 20528 26016 20534
rect 25964 20470 26016 20476
rect 26054 20088 26110 20097
rect 26054 20023 26110 20032
rect 26068 19854 26096 20023
rect 26056 19848 26108 19854
rect 26056 19790 26108 19796
rect 26160 19802 26188 21558
rect 26240 21004 26292 21010
rect 26240 20946 26292 20952
rect 26252 20534 26280 20946
rect 26240 20528 26292 20534
rect 26240 20470 26292 20476
rect 26344 20398 26372 22918
rect 26436 21894 26464 24550
rect 26712 24342 26740 25774
rect 26896 25702 26924 26794
rect 27436 26784 27488 26790
rect 27436 26726 27488 26732
rect 26976 26308 27028 26314
rect 26976 26250 27028 26256
rect 27068 26308 27120 26314
rect 27068 26250 27120 26256
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 26884 24744 26936 24750
rect 26884 24686 26936 24692
rect 26700 24336 26752 24342
rect 26700 24278 26752 24284
rect 26608 24200 26660 24206
rect 26608 24142 26660 24148
rect 26516 24064 26568 24070
rect 26514 24032 26516 24041
rect 26568 24032 26570 24041
rect 26514 23967 26570 23976
rect 26620 23866 26648 24142
rect 26700 24132 26752 24138
rect 26700 24074 26752 24080
rect 26608 23860 26660 23866
rect 26608 23802 26660 23808
rect 26516 23656 26568 23662
rect 26516 23598 26568 23604
rect 26528 22166 26556 23598
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 26516 22160 26568 22166
rect 26516 22102 26568 22108
rect 26424 21888 26476 21894
rect 26424 21830 26476 21836
rect 26620 21690 26648 22578
rect 26608 21684 26660 21690
rect 26608 21626 26660 21632
rect 26516 21344 26568 21350
rect 26516 21286 26568 21292
rect 26332 20392 26384 20398
rect 26332 20334 26384 20340
rect 26528 20330 26556 21286
rect 26620 20913 26648 21626
rect 26712 20942 26740 24074
rect 26790 23216 26846 23225
rect 26790 23151 26846 23160
rect 26804 23118 26832 23151
rect 26792 23112 26844 23118
rect 26792 23054 26844 23060
rect 26896 22574 26924 24686
rect 26884 22568 26936 22574
rect 26884 22510 26936 22516
rect 26896 21554 26924 22510
rect 26884 21548 26936 21554
rect 26884 21490 26936 21496
rect 26700 20936 26752 20942
rect 26606 20904 26662 20913
rect 26700 20878 26752 20884
rect 26606 20839 26662 20848
rect 26700 20800 26752 20806
rect 26700 20742 26752 20748
rect 26608 20392 26660 20398
rect 26608 20334 26660 20340
rect 26516 20324 26568 20330
rect 26516 20266 26568 20272
rect 26620 20210 26648 20334
rect 26528 20182 26648 20210
rect 26332 19848 26384 19854
rect 26160 19796 26332 19802
rect 26160 19790 26384 19796
rect 26160 19774 26372 19790
rect 26528 19786 26556 20182
rect 26608 20052 26660 20058
rect 26608 19994 26660 20000
rect 26516 19780 26568 19786
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 25962 19544 26018 19553
rect 25962 19479 26018 19488
rect 25976 19378 26004 19479
rect 25964 19372 26016 19378
rect 25964 19314 26016 19320
rect 26068 19258 26096 19654
rect 26160 19378 26188 19774
rect 26516 19722 26568 19728
rect 26240 19712 26292 19718
rect 26240 19654 26292 19660
rect 26252 19378 26280 19654
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26148 19372 26200 19378
rect 26148 19314 26200 19320
rect 26240 19372 26292 19378
rect 26436 19334 26464 19450
rect 26240 19314 26292 19320
rect 26344 19306 26464 19334
rect 25872 19236 25924 19242
rect 26068 19230 26188 19258
rect 25872 19178 25924 19184
rect 25884 19145 25912 19178
rect 25870 19136 25926 19145
rect 25870 19071 25926 19080
rect 25872 18964 25924 18970
rect 25924 18924 26004 18952
rect 25872 18906 25924 18912
rect 25976 18850 26004 18924
rect 26056 18896 26108 18902
rect 25976 18844 26056 18850
rect 25976 18838 26108 18844
rect 25976 18822 26096 18838
rect 25872 18760 25924 18766
rect 25872 18702 25924 18708
rect 25884 18290 25912 18702
rect 25872 18284 25924 18290
rect 25872 18226 25924 18232
rect 25976 18222 26004 18822
rect 26056 18760 26108 18766
rect 26056 18702 26108 18708
rect 26068 18465 26096 18702
rect 26054 18456 26110 18465
rect 26054 18391 26110 18400
rect 25964 18216 26016 18222
rect 25964 18158 26016 18164
rect 26056 18216 26108 18222
rect 26056 18158 26108 18164
rect 25780 17672 25832 17678
rect 25778 17640 25780 17649
rect 25832 17640 25834 17649
rect 25778 17575 25834 17584
rect 25792 16697 25820 17575
rect 25778 16688 25834 16697
rect 25778 16623 25834 16632
rect 25688 16584 25740 16590
rect 25976 16572 26004 18158
rect 26068 17134 26096 18158
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 26160 17066 26188 19230
rect 26238 18728 26294 18737
rect 26238 18663 26294 18672
rect 26252 18290 26280 18663
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 26252 18193 26280 18226
rect 26238 18184 26294 18193
rect 26238 18119 26294 18128
rect 26344 17678 26372 19306
rect 26514 19272 26570 19281
rect 26514 19207 26570 19216
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 26436 18329 26464 19110
rect 26528 18766 26556 19207
rect 26516 18760 26568 18766
rect 26516 18702 26568 18708
rect 26422 18320 26478 18329
rect 26422 18255 26478 18264
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 26146 16688 26202 16697
rect 26146 16623 26202 16632
rect 26160 16590 26188 16623
rect 25740 16544 26004 16572
rect 26148 16584 26200 16590
rect 25688 16526 25740 16532
rect 25596 16244 25648 16250
rect 25596 16186 25648 16192
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24584 15428 24636 15434
rect 24584 15370 24636 15376
rect 25424 15026 25452 15846
rect 25504 15360 25556 15366
rect 25504 15302 25556 15308
rect 25412 15020 25464 15026
rect 25412 14962 25464 14968
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 24308 13456 24360 13462
rect 24308 13398 24360 13404
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 23768 13212 23888 13240
rect 23664 12708 23716 12714
rect 23664 12650 23716 12656
rect 23768 11830 23796 13212
rect 24228 12782 24256 13330
rect 24320 12986 24348 13398
rect 24688 12986 24716 14554
rect 24780 13326 24808 14758
rect 25516 14414 25544 15302
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 25504 14408 25556 14414
rect 25504 14350 25556 14356
rect 24860 14340 24912 14346
rect 24860 14282 24912 14288
rect 24872 13326 24900 14282
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24308 12980 24360 12986
rect 24676 12980 24728 12986
rect 24308 12922 24360 12928
rect 24596 12940 24676 12968
rect 24216 12776 24268 12782
rect 24216 12718 24268 12724
rect 23848 12640 23900 12646
rect 23848 12582 23900 12588
rect 23860 12306 23888 12582
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23848 12164 23900 12170
rect 23848 12106 23900 12112
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23204 11756 23256 11762
rect 23204 11698 23256 11704
rect 23216 11354 23244 11698
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23768 11218 23796 11766
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 23296 11008 23348 11014
rect 23296 10950 23348 10956
rect 23480 11008 23532 11014
rect 23480 10950 23532 10956
rect 23308 10674 23336 10950
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 23492 10470 23520 10950
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23492 10062 23520 10406
rect 23860 10062 23888 12106
rect 24228 11218 24256 12718
rect 24596 12442 24624 12940
rect 24676 12922 24728 12928
rect 24584 12436 24636 12442
rect 24584 12378 24636 12384
rect 24308 11892 24360 11898
rect 24308 11834 24360 11840
rect 24320 11694 24348 11834
rect 24872 11762 24900 13262
rect 24964 12850 24992 14350
rect 25516 14074 25544 14350
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25332 13530 25360 13874
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25608 13190 25636 16186
rect 25688 13320 25740 13326
rect 25688 13262 25740 13268
rect 25596 13184 25648 13190
rect 25596 13126 25648 13132
rect 24952 12844 25004 12850
rect 25004 12804 25084 12832
rect 24952 12786 25004 12792
rect 25056 12170 25084 12804
rect 25044 12164 25096 12170
rect 25044 12106 25096 12112
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 25320 12096 25372 12102
rect 25320 12038 25372 12044
rect 24964 11830 24992 12038
rect 25332 11898 25360 12038
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 24952 11824 25004 11830
rect 24952 11766 25004 11772
rect 25700 11762 25728 13262
rect 25792 12102 25820 16544
rect 26148 16526 26200 16532
rect 26436 16182 26464 18255
rect 26528 18193 26556 18702
rect 26620 18290 26648 19994
rect 26608 18284 26660 18290
rect 26608 18226 26660 18232
rect 26514 18184 26570 18193
rect 26514 18119 26570 18128
rect 26516 18080 26568 18086
rect 26516 18022 26568 18028
rect 26528 17882 26556 18022
rect 26516 17876 26568 17882
rect 26516 17818 26568 17824
rect 26608 17604 26660 17610
rect 26608 17546 26660 17552
rect 26620 17270 26648 17546
rect 26712 17338 26740 20742
rect 26896 19922 26924 21490
rect 26988 21434 27016 26250
rect 27080 24206 27108 26250
rect 27252 25152 27304 25158
rect 27252 25094 27304 25100
rect 27160 24268 27212 24274
rect 27160 24210 27212 24216
rect 27068 24200 27120 24206
rect 27068 24142 27120 24148
rect 27172 23769 27200 24210
rect 27158 23760 27214 23769
rect 27158 23695 27214 23704
rect 27068 22772 27120 22778
rect 27068 22714 27120 22720
rect 27080 22574 27108 22714
rect 27172 22642 27200 23695
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 27068 22568 27120 22574
rect 27068 22510 27120 22516
rect 27068 22432 27120 22438
rect 27068 22374 27120 22380
rect 27080 22098 27108 22374
rect 27068 22092 27120 22098
rect 27068 22034 27120 22040
rect 27080 21554 27108 22034
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 27068 21548 27120 21554
rect 27068 21490 27120 21496
rect 27172 21486 27200 21626
rect 27160 21480 27212 21486
rect 26988 21406 27108 21434
rect 27160 21422 27212 21428
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 26988 21146 27016 21286
rect 26976 21140 27028 21146
rect 26976 21082 27028 21088
rect 26976 20800 27028 20806
rect 26976 20742 27028 20748
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 26792 19780 26844 19786
rect 26792 19722 26844 19728
rect 26804 18766 26832 19722
rect 26896 19378 26924 19858
rect 26884 19372 26936 19378
rect 26884 19314 26936 19320
rect 26884 19236 26936 19242
rect 26884 19178 26936 19184
rect 26896 19145 26924 19178
rect 26882 19136 26938 19145
rect 26882 19071 26938 19080
rect 26988 18902 27016 20742
rect 27080 20466 27108 21406
rect 27172 21185 27200 21422
rect 27158 21176 27214 21185
rect 27158 21111 27214 21120
rect 27068 20460 27120 20466
rect 27068 20402 27120 20408
rect 27264 19922 27292 25094
rect 27344 24880 27396 24886
rect 27344 24822 27396 24828
rect 27356 23526 27384 24822
rect 27448 24041 27476 26726
rect 27632 25906 27660 30534
rect 27724 30326 27752 30534
rect 27712 30320 27764 30326
rect 27712 30262 27764 30268
rect 27724 30190 27752 30262
rect 27712 30184 27764 30190
rect 27712 30126 27764 30132
rect 27816 30122 27844 32370
rect 27908 31793 27936 32807
rect 27894 31784 27950 31793
rect 27894 31719 27896 31728
rect 27948 31719 27950 31728
rect 27896 31690 27948 31696
rect 27894 30968 27950 30977
rect 27894 30903 27950 30912
rect 27804 30116 27856 30122
rect 27804 30058 27856 30064
rect 27712 29504 27764 29510
rect 27712 29446 27764 29452
rect 27804 29504 27856 29510
rect 27804 29446 27856 29452
rect 27724 28098 27752 29446
rect 27816 28694 27844 29446
rect 27908 29238 27936 30903
rect 27896 29232 27948 29238
rect 27896 29174 27948 29180
rect 27908 28966 27936 29174
rect 27896 28960 27948 28966
rect 27896 28902 27948 28908
rect 27804 28688 27856 28694
rect 27804 28630 27856 28636
rect 27804 28484 27856 28490
rect 27804 28426 27856 28432
rect 27816 28393 27844 28426
rect 27802 28384 27858 28393
rect 27802 28319 27858 28328
rect 27724 28070 27844 28098
rect 27712 28008 27764 28014
rect 27712 27950 27764 27956
rect 27724 27062 27752 27950
rect 27816 27538 27844 28070
rect 27896 27600 27948 27606
rect 27896 27542 27948 27548
rect 27804 27532 27856 27538
rect 27804 27474 27856 27480
rect 27802 27296 27858 27305
rect 27802 27231 27858 27240
rect 27712 27056 27764 27062
rect 27712 26998 27764 27004
rect 27712 26240 27764 26246
rect 27710 26208 27712 26217
rect 27764 26208 27766 26217
rect 27710 26143 27766 26152
rect 27620 25900 27672 25906
rect 27620 25842 27672 25848
rect 27712 25832 27764 25838
rect 27712 25774 27764 25780
rect 27526 25392 27582 25401
rect 27526 25327 27582 25336
rect 27434 24032 27490 24041
rect 27434 23967 27490 23976
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 27344 23520 27396 23526
rect 27344 23462 27396 23468
rect 27344 23112 27396 23118
rect 27344 23054 27396 23060
rect 27356 22778 27384 23054
rect 27448 23050 27476 23666
rect 27540 23633 27568 25327
rect 27620 25288 27672 25294
rect 27618 25256 27620 25265
rect 27672 25256 27674 25265
rect 27618 25191 27674 25200
rect 27620 24948 27672 24954
rect 27620 24890 27672 24896
rect 27632 24818 27660 24890
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 27632 24177 27660 24754
rect 27618 24168 27674 24177
rect 27618 24103 27674 24112
rect 27526 23624 27582 23633
rect 27526 23559 27582 23568
rect 27724 23526 27752 25774
rect 27816 24857 27844 27231
rect 27908 27062 27936 27542
rect 28000 27130 28028 36094
rect 28080 36032 28132 36038
rect 28080 35974 28132 35980
rect 28172 36032 28224 36038
rect 28172 35974 28224 35980
rect 28092 35630 28120 35974
rect 28080 35624 28132 35630
rect 28080 35566 28132 35572
rect 28080 34128 28132 34134
rect 28080 34070 28132 34076
rect 28092 30433 28120 34070
rect 28184 33998 28212 35974
rect 28262 35864 28318 35873
rect 28262 35799 28318 35808
rect 28276 35494 28304 35799
rect 28264 35488 28316 35494
rect 28264 35430 28316 35436
rect 28276 35222 28304 35430
rect 28264 35216 28316 35222
rect 28264 35158 28316 35164
rect 28368 34785 28396 37062
rect 28460 35290 28488 37334
rect 29012 36854 29040 37431
rect 29184 37256 29236 37262
rect 29184 37198 29236 37204
rect 29642 37224 29698 37233
rect 29092 37120 29144 37126
rect 29092 37062 29144 37068
rect 28724 36848 28776 36854
rect 28724 36790 28776 36796
rect 29000 36848 29052 36854
rect 29000 36790 29052 36796
rect 28736 36689 28764 36790
rect 28722 36680 28778 36689
rect 28722 36615 28778 36624
rect 29104 36582 29132 37062
rect 29092 36576 29144 36582
rect 29092 36518 29144 36524
rect 29196 36281 29224 37198
rect 29460 37188 29512 37194
rect 29642 37159 29698 37168
rect 29460 37130 29512 37136
rect 29368 36576 29420 36582
rect 29368 36518 29420 36524
rect 29276 36372 29328 36378
rect 29276 36314 29328 36320
rect 29182 36272 29238 36281
rect 28540 36236 28592 36242
rect 29182 36207 29238 36216
rect 28540 36178 28592 36184
rect 28552 35986 28580 36178
rect 28816 36168 28868 36174
rect 28816 36110 28868 36116
rect 28908 36168 28960 36174
rect 28908 36110 28960 36116
rect 29092 36168 29144 36174
rect 29092 36110 29144 36116
rect 28552 35958 28764 35986
rect 28632 35692 28684 35698
rect 28632 35634 28684 35640
rect 28448 35284 28500 35290
rect 28448 35226 28500 35232
rect 28644 35154 28672 35634
rect 28632 35148 28684 35154
rect 28632 35090 28684 35096
rect 28538 34912 28594 34921
rect 28538 34847 28594 34856
rect 28354 34776 28410 34785
rect 28354 34711 28410 34720
rect 28264 34604 28316 34610
rect 28264 34546 28316 34552
rect 28172 33992 28224 33998
rect 28172 33934 28224 33940
rect 28172 33856 28224 33862
rect 28172 33798 28224 33804
rect 28184 33318 28212 33798
rect 28172 33312 28224 33318
rect 28172 33254 28224 33260
rect 28184 32910 28212 33254
rect 28172 32904 28224 32910
rect 28172 32846 28224 32852
rect 28276 32552 28304 34546
rect 28368 33930 28396 34711
rect 28446 34096 28502 34105
rect 28446 34031 28502 34040
rect 28356 33924 28408 33930
rect 28356 33866 28408 33872
rect 28460 33810 28488 34031
rect 28368 33782 28488 33810
rect 28368 33114 28396 33782
rect 28552 33402 28580 34847
rect 28644 33930 28672 35090
rect 28632 33924 28684 33930
rect 28632 33866 28684 33872
rect 28736 33862 28764 35958
rect 28828 35834 28856 36110
rect 28816 35828 28868 35834
rect 28816 35770 28868 35776
rect 28828 34950 28856 35770
rect 28920 35494 28948 36110
rect 29000 35624 29052 35630
rect 29104 35612 29132 36110
rect 29052 35584 29132 35612
rect 29000 35566 29052 35572
rect 28908 35488 28960 35494
rect 28908 35430 28960 35436
rect 29012 35222 29040 35566
rect 29000 35216 29052 35222
rect 29000 35158 29052 35164
rect 29184 35148 29236 35154
rect 29184 35090 29236 35096
rect 29196 35018 29224 35090
rect 29288 35086 29316 36314
rect 29276 35080 29328 35086
rect 29276 35022 29328 35028
rect 29184 35012 29236 35018
rect 29184 34954 29236 34960
rect 28816 34944 28868 34950
rect 28816 34886 28868 34892
rect 28906 34912 28962 34921
rect 28906 34847 28962 34856
rect 28816 34400 28868 34406
rect 28816 34342 28868 34348
rect 28828 33998 28856 34342
rect 28816 33992 28868 33998
rect 28816 33934 28868 33940
rect 28724 33856 28776 33862
rect 28920 33844 28948 34847
rect 29000 34672 29052 34678
rect 28998 34640 29000 34649
rect 29052 34640 29054 34649
rect 28998 34575 29054 34584
rect 28998 34096 29054 34105
rect 28998 34031 29054 34040
rect 28724 33798 28776 33804
rect 28828 33816 28948 33844
rect 29012 33833 29040 34031
rect 29288 33998 29316 35022
rect 29092 33992 29144 33998
rect 29276 33992 29328 33998
rect 29144 33952 29224 33980
rect 29092 33934 29144 33940
rect 29092 33856 29144 33862
rect 28998 33824 29054 33833
rect 28552 33374 28764 33402
rect 28632 33312 28684 33318
rect 28538 33280 28594 33289
rect 28632 33254 28684 33260
rect 28538 33215 28594 33224
rect 28356 33108 28408 33114
rect 28356 33050 28408 33056
rect 28448 33040 28500 33046
rect 28354 33008 28410 33017
rect 28448 32982 28500 32988
rect 28354 32943 28410 32952
rect 28368 32910 28396 32943
rect 28356 32904 28408 32910
rect 28356 32846 28408 32852
rect 28276 32524 28396 32552
rect 28264 32428 28316 32434
rect 28264 32370 28316 32376
rect 28172 32292 28224 32298
rect 28172 32234 28224 32240
rect 28184 30870 28212 32234
rect 28276 31906 28304 32370
rect 28368 32026 28396 32524
rect 28356 32020 28408 32026
rect 28356 31962 28408 31968
rect 28276 31878 28396 31906
rect 28264 31680 28316 31686
rect 28264 31622 28316 31628
rect 28172 30864 28224 30870
rect 28172 30806 28224 30812
rect 28172 30660 28224 30666
rect 28172 30602 28224 30608
rect 28078 30424 28134 30433
rect 28078 30359 28134 30368
rect 28184 30190 28212 30602
rect 28080 30184 28132 30190
rect 28080 30126 28132 30132
rect 28172 30184 28224 30190
rect 28172 30126 28224 30132
rect 28092 27606 28120 30126
rect 28184 29850 28212 30126
rect 28172 29844 28224 29850
rect 28172 29786 28224 29792
rect 28172 29640 28224 29646
rect 28172 29582 28224 29588
rect 28184 29170 28212 29582
rect 28276 29170 28304 31622
rect 28368 31362 28396 31878
rect 28460 31822 28488 32982
rect 28552 32609 28580 33215
rect 28644 33017 28672 33254
rect 28630 33008 28686 33017
rect 28630 32943 28686 32952
rect 28538 32600 28594 32609
rect 28538 32535 28594 32544
rect 28736 32434 28764 33374
rect 28828 32910 28856 33816
rect 29092 33798 29144 33804
rect 28998 33759 29054 33768
rect 28908 33584 28960 33590
rect 28906 33552 28908 33561
rect 28960 33552 28962 33561
rect 28906 33487 28962 33496
rect 29012 33130 29040 33759
rect 29104 33289 29132 33798
rect 29090 33280 29146 33289
rect 29090 33215 29146 33224
rect 29012 33102 29132 33130
rect 28816 32904 28868 32910
rect 28816 32846 28868 32852
rect 28828 32745 28856 32846
rect 29104 32824 29132 33102
rect 29012 32796 29132 32824
rect 28908 32768 28960 32774
rect 28814 32736 28870 32745
rect 28908 32710 28960 32716
rect 28814 32671 28870 32680
rect 28724 32428 28776 32434
rect 28644 32388 28724 32416
rect 28644 32178 28672 32388
rect 28724 32370 28776 32376
rect 28920 32366 28948 32710
rect 29012 32366 29040 32796
rect 29090 32736 29146 32745
rect 29090 32671 29146 32680
rect 29104 32473 29132 32671
rect 29090 32464 29146 32473
rect 29090 32399 29146 32408
rect 28908 32360 28960 32366
rect 28814 32328 28870 32337
rect 28908 32302 28960 32308
rect 29000 32360 29052 32366
rect 29000 32302 29052 32308
rect 29090 32328 29146 32337
rect 28814 32263 28870 32272
rect 29090 32263 29146 32272
rect 28552 32150 28672 32178
rect 28448 31816 28500 31822
rect 28448 31758 28500 31764
rect 28552 31754 28580 32150
rect 28630 32056 28686 32065
rect 28630 31991 28686 32000
rect 28644 31822 28672 31991
rect 28828 31929 28856 32263
rect 29000 31952 29052 31958
rect 28814 31920 28870 31929
rect 29000 31894 29052 31900
rect 28814 31855 28870 31864
rect 28632 31816 28684 31822
rect 28632 31758 28684 31764
rect 28722 31784 28778 31793
rect 28540 31748 28592 31754
rect 28722 31719 28778 31728
rect 28540 31690 28592 31696
rect 28446 31376 28502 31385
rect 28368 31334 28446 31362
rect 28446 31311 28502 31320
rect 28632 31340 28684 31346
rect 28356 30864 28408 30870
rect 28356 30806 28408 30812
rect 28172 29164 28224 29170
rect 28172 29106 28224 29112
rect 28264 29164 28316 29170
rect 28264 29106 28316 29112
rect 28170 29064 28226 29073
rect 28170 28999 28226 29008
rect 28184 28082 28212 28999
rect 28276 28626 28304 29106
rect 28264 28620 28316 28626
rect 28264 28562 28316 28568
rect 28172 28076 28224 28082
rect 28172 28018 28224 28024
rect 28276 28014 28304 28562
rect 28264 28008 28316 28014
rect 28264 27950 28316 27956
rect 28368 27674 28396 30806
rect 28460 30433 28488 31311
rect 28632 31282 28684 31288
rect 28540 31272 28592 31278
rect 28540 31214 28592 31220
rect 28552 30598 28580 31214
rect 28644 30938 28672 31282
rect 28632 30932 28684 30938
rect 28632 30874 28684 30880
rect 28632 30728 28684 30734
rect 28632 30670 28684 30676
rect 28540 30592 28592 30598
rect 28540 30534 28592 30540
rect 28446 30424 28502 30433
rect 28446 30359 28502 30368
rect 28448 30252 28500 30258
rect 28448 30194 28500 30200
rect 28460 29646 28488 30194
rect 28644 30122 28672 30670
rect 28736 30598 28764 31719
rect 29012 30870 29040 31894
rect 29104 31414 29132 32263
rect 29092 31408 29144 31414
rect 29092 31350 29144 31356
rect 29196 31226 29224 33952
rect 29380 33969 29408 36518
rect 29472 36310 29500 37130
rect 29460 36304 29512 36310
rect 29460 36246 29512 36252
rect 29460 35488 29512 35494
rect 29460 35430 29512 35436
rect 29472 34649 29500 35430
rect 29458 34640 29514 34649
rect 29458 34575 29514 34584
rect 29552 34536 29604 34542
rect 29552 34478 29604 34484
rect 29564 33969 29592 34478
rect 29276 33934 29328 33940
rect 29366 33960 29422 33969
rect 29288 33318 29316 33934
rect 29366 33895 29422 33904
rect 29550 33960 29606 33969
rect 29550 33895 29606 33904
rect 29460 33856 29512 33862
rect 29460 33798 29512 33804
rect 29276 33312 29328 33318
rect 29276 33254 29328 33260
rect 29368 32972 29420 32978
rect 29368 32914 29420 32920
rect 29276 32836 29328 32842
rect 29276 32778 29328 32784
rect 29288 32366 29316 32778
rect 29276 32360 29328 32366
rect 29276 32302 29328 32308
rect 29276 32224 29328 32230
rect 29276 32166 29328 32172
rect 29288 31346 29316 32166
rect 29276 31340 29328 31346
rect 29276 31282 29328 31288
rect 29104 31198 29224 31226
rect 28816 30864 28868 30870
rect 28816 30806 28868 30812
rect 29000 30864 29052 30870
rect 29000 30806 29052 30812
rect 28828 30734 28856 30806
rect 28816 30728 28868 30734
rect 28816 30670 28868 30676
rect 28724 30592 28776 30598
rect 28724 30534 28776 30540
rect 28908 30592 28960 30598
rect 28908 30534 28960 30540
rect 28632 30116 28684 30122
rect 28632 30058 28684 30064
rect 28920 29646 28948 30534
rect 28998 30424 29054 30433
rect 28998 30359 29054 30368
rect 28448 29640 28500 29646
rect 28448 29582 28500 29588
rect 28724 29640 28776 29646
rect 28724 29582 28776 29588
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 28632 29572 28684 29578
rect 28632 29514 28684 29520
rect 28446 29336 28502 29345
rect 28446 29271 28502 29280
rect 28356 27668 28408 27674
rect 28356 27610 28408 27616
rect 28080 27600 28132 27606
rect 28080 27542 28132 27548
rect 28092 27470 28120 27542
rect 28080 27464 28132 27470
rect 28132 27424 28212 27452
rect 28080 27406 28132 27412
rect 27988 27124 28040 27130
rect 27988 27066 28040 27072
rect 28080 27124 28132 27130
rect 28080 27066 28132 27072
rect 27896 27056 27948 27062
rect 27896 26998 27948 27004
rect 27896 26240 27948 26246
rect 27896 26182 27948 26188
rect 27908 25838 27936 26182
rect 28000 25906 28028 27066
rect 28092 26586 28120 27066
rect 28184 26994 28212 27424
rect 28172 26988 28224 26994
rect 28172 26930 28224 26936
rect 28080 26580 28132 26586
rect 28080 26522 28132 26528
rect 28264 26580 28316 26586
rect 28264 26522 28316 26528
rect 28276 26450 28304 26522
rect 28460 26466 28488 29271
rect 28644 28218 28672 29514
rect 28632 28212 28684 28218
rect 28632 28154 28684 28160
rect 28736 28150 28764 29582
rect 28908 28484 28960 28490
rect 28908 28426 28960 28432
rect 28816 28416 28868 28422
rect 28816 28358 28868 28364
rect 28724 28144 28776 28150
rect 28724 28086 28776 28092
rect 28540 28076 28592 28082
rect 28540 28018 28592 28024
rect 28552 27674 28580 28018
rect 28540 27668 28592 27674
rect 28540 27610 28592 27616
rect 28724 27532 28776 27538
rect 28724 27474 28776 27480
rect 28632 27328 28684 27334
rect 28632 27270 28684 27276
rect 28080 26444 28132 26450
rect 28080 26386 28132 26392
rect 28264 26444 28316 26450
rect 28264 26386 28316 26392
rect 28368 26438 28488 26466
rect 28540 26444 28592 26450
rect 27988 25900 28040 25906
rect 27988 25842 28040 25848
rect 27896 25832 27948 25838
rect 27896 25774 27948 25780
rect 27988 25696 28040 25702
rect 27988 25638 28040 25644
rect 28000 25430 28028 25638
rect 27988 25424 28040 25430
rect 27988 25366 28040 25372
rect 28000 25226 28028 25366
rect 28092 25294 28120 26386
rect 28172 25832 28224 25838
rect 28172 25774 28224 25780
rect 28080 25288 28132 25294
rect 28080 25230 28132 25236
rect 27988 25220 28040 25226
rect 27988 25162 28040 25168
rect 27896 25152 27948 25158
rect 27896 25094 27948 25100
rect 27908 24993 27936 25094
rect 27894 24984 27950 24993
rect 27894 24919 27950 24928
rect 27802 24848 27858 24857
rect 27908 24818 27936 24919
rect 27802 24783 27858 24792
rect 27896 24812 27948 24818
rect 27896 24754 27948 24760
rect 27988 24744 28040 24750
rect 27986 24712 27988 24721
rect 28040 24712 28042 24721
rect 27986 24647 28042 24656
rect 27896 24608 27948 24614
rect 27896 24550 27948 24556
rect 28078 24576 28134 24585
rect 27802 24304 27858 24313
rect 27802 24239 27804 24248
rect 27856 24239 27858 24248
rect 27804 24210 27856 24216
rect 27816 24018 27844 24210
rect 27908 24206 27936 24550
rect 28078 24511 28134 24520
rect 27896 24200 27948 24206
rect 27896 24142 27948 24148
rect 27988 24200 28040 24206
rect 27988 24142 28040 24148
rect 27816 23990 27936 24018
rect 27804 23860 27856 23866
rect 27804 23802 27856 23808
rect 27712 23520 27764 23526
rect 27712 23462 27764 23468
rect 27436 23044 27488 23050
rect 27436 22986 27488 22992
rect 27344 22772 27396 22778
rect 27344 22714 27396 22720
rect 27344 22228 27396 22234
rect 27344 22170 27396 22176
rect 27356 20874 27384 22170
rect 27344 20868 27396 20874
rect 27344 20810 27396 20816
rect 27342 20632 27398 20641
rect 27342 20567 27398 20576
rect 27356 19990 27384 20567
rect 27448 20398 27476 22986
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 27540 22030 27568 22714
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 27528 22024 27580 22030
rect 27528 21966 27580 21972
rect 27528 21344 27580 21350
rect 27632 21332 27660 22578
rect 27816 22098 27844 23802
rect 27908 22234 27936 23990
rect 28000 23322 28028 24142
rect 27988 23316 28040 23322
rect 27988 23258 28040 23264
rect 27988 23044 28040 23050
rect 27988 22986 28040 22992
rect 28000 22234 28028 22986
rect 27896 22228 27948 22234
rect 27896 22170 27948 22176
rect 27988 22228 28040 22234
rect 27988 22170 28040 22176
rect 27804 22092 27856 22098
rect 28092 22094 28120 24511
rect 27804 22034 27856 22040
rect 28000 22066 28120 22094
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 27580 21304 27660 21332
rect 27528 21286 27580 21292
rect 27632 21078 27660 21304
rect 27620 21072 27672 21078
rect 27620 21014 27672 21020
rect 27816 21010 27844 21422
rect 27804 21004 27856 21010
rect 27804 20946 27856 20952
rect 27712 20800 27764 20806
rect 27712 20742 27764 20748
rect 27436 20392 27488 20398
rect 27436 20334 27488 20340
rect 27528 20256 27580 20262
rect 27448 20216 27528 20244
rect 27344 19984 27396 19990
rect 27344 19926 27396 19932
rect 27252 19916 27304 19922
rect 27252 19858 27304 19864
rect 27448 19854 27476 20216
rect 27528 20198 27580 20204
rect 27436 19848 27488 19854
rect 27356 19796 27436 19802
rect 27356 19790 27488 19796
rect 27252 19780 27304 19786
rect 27252 19722 27304 19728
rect 27356 19774 27476 19790
rect 27160 19508 27212 19514
rect 27160 19450 27212 19456
rect 27068 19304 27120 19310
rect 27068 19246 27120 19252
rect 26976 18896 27028 18902
rect 26976 18838 27028 18844
rect 27080 18766 27108 19246
rect 26792 18760 26844 18766
rect 26792 18702 26844 18708
rect 27068 18760 27120 18766
rect 27068 18702 27120 18708
rect 27172 18170 27200 19450
rect 27264 19378 27292 19722
rect 27356 19514 27384 19774
rect 27434 19680 27490 19689
rect 27434 19615 27490 19624
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 27264 18290 27292 19314
rect 27448 19009 27476 19615
rect 27620 19304 27672 19310
rect 27620 19246 27672 19252
rect 27434 19000 27490 19009
rect 27434 18935 27490 18944
rect 27344 18896 27396 18902
rect 27344 18838 27396 18844
rect 27356 18737 27384 18838
rect 27528 18760 27580 18766
rect 27342 18728 27398 18737
rect 27398 18686 27476 18714
rect 27632 18748 27660 19246
rect 27724 18850 27752 20742
rect 28000 20398 28028 22066
rect 28080 22024 28132 22030
rect 28080 21966 28132 21972
rect 28092 21690 28120 21966
rect 28080 21684 28132 21690
rect 28080 21626 28132 21632
rect 27988 20392 28040 20398
rect 27988 20334 28040 20340
rect 27896 20324 27948 20330
rect 27896 20266 27948 20272
rect 27908 19378 27936 20266
rect 27896 19372 27948 19378
rect 28184 19334 28212 25774
rect 28276 23662 28304 26386
rect 28368 25702 28396 26438
rect 28540 26386 28592 26392
rect 28448 26376 28500 26382
rect 28448 26318 28500 26324
rect 28356 25696 28408 25702
rect 28356 25638 28408 25644
rect 28354 25528 28410 25537
rect 28354 25463 28410 25472
rect 28368 25226 28396 25463
rect 28356 25220 28408 25226
rect 28356 25162 28408 25168
rect 28368 24954 28396 25162
rect 28356 24948 28408 24954
rect 28356 24890 28408 24896
rect 28356 24336 28408 24342
rect 28356 24278 28408 24284
rect 28264 23656 28316 23662
rect 28264 23598 28316 23604
rect 28262 23352 28318 23361
rect 28262 23287 28318 23296
rect 28276 22642 28304 23287
rect 28368 23050 28396 24278
rect 28460 23730 28488 26318
rect 28552 25673 28580 26386
rect 28538 25664 28594 25673
rect 28538 25599 28594 25608
rect 28644 24993 28672 27270
rect 28736 25838 28764 27474
rect 28828 26450 28856 28358
rect 28920 27470 28948 28426
rect 29012 28082 29040 30359
rect 29104 30190 29132 31198
rect 29276 31136 29328 31142
rect 29276 31078 29328 31084
rect 29288 30938 29316 31078
rect 29276 30932 29328 30938
rect 29276 30874 29328 30880
rect 29380 30569 29408 32914
rect 29472 32434 29500 33798
rect 29564 32978 29592 33895
rect 29656 33590 29684 37159
rect 29920 36576 29972 36582
rect 29920 36518 29972 36524
rect 29828 36372 29880 36378
rect 29828 36314 29880 36320
rect 29840 35873 29868 36314
rect 29932 36310 29960 36518
rect 29920 36304 29972 36310
rect 29920 36246 29972 36252
rect 29826 35864 29882 35873
rect 29826 35799 29882 35808
rect 29840 35698 29868 35799
rect 29932 35698 29960 36246
rect 29828 35692 29880 35698
rect 29748 35652 29828 35680
rect 29644 33584 29696 33590
rect 29644 33526 29696 33532
rect 29644 33312 29696 33318
rect 29644 33254 29696 33260
rect 29552 32972 29604 32978
rect 29552 32914 29604 32920
rect 29460 32428 29512 32434
rect 29512 32388 29592 32416
rect 29460 32370 29512 32376
rect 29458 32056 29514 32065
rect 29458 31991 29514 32000
rect 29366 30560 29422 30569
rect 29366 30495 29422 30504
rect 29092 30184 29144 30190
rect 29092 30126 29144 30132
rect 29104 28082 29132 30126
rect 29274 29880 29330 29889
rect 29274 29815 29330 29824
rect 29184 29572 29236 29578
rect 29184 29514 29236 29520
rect 29196 29238 29224 29514
rect 29288 29306 29316 29815
rect 29380 29646 29408 30495
rect 29368 29640 29420 29646
rect 29368 29582 29420 29588
rect 29276 29300 29328 29306
rect 29276 29242 29328 29248
rect 29184 29232 29236 29238
rect 29184 29174 29236 29180
rect 29380 29170 29408 29582
rect 29368 29164 29420 29170
rect 29368 29106 29420 29112
rect 29276 28960 29328 28966
rect 29182 28928 29238 28937
rect 29276 28902 29328 28908
rect 29368 28960 29420 28966
rect 29368 28902 29420 28908
rect 29182 28863 29238 28872
rect 29196 28626 29224 28863
rect 29288 28626 29316 28902
rect 29184 28620 29236 28626
rect 29184 28562 29236 28568
rect 29276 28620 29328 28626
rect 29276 28562 29328 28568
rect 29000 28076 29052 28082
rect 29000 28018 29052 28024
rect 29092 28076 29144 28082
rect 29092 28018 29144 28024
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 28920 26489 28948 27406
rect 29000 27056 29052 27062
rect 28998 27024 29000 27033
rect 29052 27024 29054 27033
rect 29104 26994 29132 28018
rect 29196 27538 29224 28562
rect 29184 27532 29236 27538
rect 29184 27474 29236 27480
rect 29276 27464 29328 27470
rect 29276 27406 29328 27412
rect 29288 27033 29316 27406
rect 29274 27024 29330 27033
rect 28998 26959 29054 26968
rect 29092 26988 29144 26994
rect 29274 26959 29330 26968
rect 29092 26930 29144 26936
rect 29000 26920 29052 26926
rect 29000 26862 29052 26868
rect 28906 26480 28962 26489
rect 28816 26444 28868 26450
rect 28906 26415 28962 26424
rect 28816 26386 28868 26392
rect 28828 25945 28856 26386
rect 29012 26330 29040 26862
rect 29184 26376 29236 26382
rect 28920 26302 29040 26330
rect 29104 26336 29184 26364
rect 28920 26246 28948 26302
rect 28908 26240 28960 26246
rect 28908 26182 28960 26188
rect 28998 26208 29054 26217
rect 28998 26143 29054 26152
rect 28814 25936 28870 25945
rect 28814 25871 28870 25880
rect 28908 25900 28960 25906
rect 28724 25832 28776 25838
rect 28724 25774 28776 25780
rect 28722 25664 28778 25673
rect 28722 25599 28778 25608
rect 28630 24984 28686 24993
rect 28630 24919 28686 24928
rect 28630 24848 28686 24857
rect 28630 24783 28686 24792
rect 28540 24744 28592 24750
rect 28540 24686 28592 24692
rect 28552 23730 28580 24686
rect 28448 23724 28500 23730
rect 28448 23666 28500 23672
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28446 23488 28502 23497
rect 28446 23423 28502 23432
rect 28460 23254 28488 23423
rect 28644 23338 28672 24783
rect 28736 23508 28764 25599
rect 28828 23746 28856 25871
rect 28908 25842 28960 25848
rect 28920 25537 28948 25842
rect 28906 25528 28962 25537
rect 28906 25463 28908 25472
rect 28960 25463 28962 25472
rect 28908 25434 28960 25440
rect 28908 25356 28960 25362
rect 28908 25298 28960 25304
rect 28920 25158 28948 25298
rect 29012 25158 29040 26143
rect 28908 25152 28960 25158
rect 28908 25094 28960 25100
rect 29000 25152 29052 25158
rect 29000 25094 29052 25100
rect 29104 24970 29132 26336
rect 29184 26318 29236 26324
rect 29276 26376 29328 26382
rect 29276 26318 29328 26324
rect 29184 25900 29236 25906
rect 29184 25842 29236 25848
rect 29196 25226 29224 25842
rect 29184 25220 29236 25226
rect 29184 25162 29236 25168
rect 28920 24942 29132 24970
rect 29182 24984 29238 24993
rect 28920 23866 28948 24942
rect 29182 24919 29184 24928
rect 29236 24919 29238 24928
rect 29184 24890 29236 24896
rect 29092 24880 29144 24886
rect 29090 24848 29092 24857
rect 29144 24848 29146 24857
rect 29090 24783 29146 24792
rect 29184 24812 29236 24818
rect 29288 24800 29316 26318
rect 29236 24772 29316 24800
rect 29184 24754 29236 24760
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 29012 23905 29040 24550
rect 29092 24064 29144 24070
rect 29090 24032 29092 24041
rect 29144 24032 29146 24041
rect 29090 23967 29146 23976
rect 28998 23896 29054 23905
rect 28908 23860 28960 23866
rect 28998 23831 29054 23840
rect 28908 23802 28960 23808
rect 28828 23718 28948 23746
rect 28816 23520 28868 23526
rect 28736 23480 28816 23508
rect 28816 23462 28868 23468
rect 28644 23310 28856 23338
rect 28448 23248 28500 23254
rect 28448 23190 28500 23196
rect 28540 23248 28592 23254
rect 28540 23190 28592 23196
rect 28356 23044 28408 23050
rect 28356 22986 28408 22992
rect 28446 22808 28502 22817
rect 28446 22743 28502 22752
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 28460 22506 28488 22743
rect 28448 22500 28500 22506
rect 28448 22442 28500 22448
rect 28552 22098 28580 23190
rect 28724 23044 28776 23050
rect 28724 22986 28776 22992
rect 28632 22976 28684 22982
rect 28632 22918 28684 22924
rect 28644 22778 28672 22918
rect 28632 22772 28684 22778
rect 28632 22714 28684 22720
rect 28644 22166 28672 22714
rect 28736 22642 28764 22986
rect 28724 22636 28776 22642
rect 28724 22578 28776 22584
rect 28632 22160 28684 22166
rect 28632 22102 28684 22108
rect 28540 22092 28592 22098
rect 28540 22034 28592 22040
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 28540 21956 28592 21962
rect 28540 21898 28592 21904
rect 28264 21888 28316 21894
rect 28264 21830 28316 21836
rect 28356 21888 28408 21894
rect 28356 21830 28408 21836
rect 28276 21486 28304 21830
rect 28264 21480 28316 21486
rect 28264 21422 28316 21428
rect 28368 20754 28396 21830
rect 28460 21554 28488 21898
rect 28552 21554 28580 21898
rect 28644 21622 28672 22102
rect 28828 22094 28856 23310
rect 28736 22066 28856 22094
rect 28632 21616 28684 21622
rect 28632 21558 28684 21564
rect 28448 21548 28500 21554
rect 28448 21490 28500 21496
rect 28540 21548 28592 21554
rect 28540 21490 28592 21496
rect 28460 21350 28488 21490
rect 28448 21344 28500 21350
rect 28448 21286 28500 21292
rect 28538 20904 28594 20913
rect 28538 20839 28594 20848
rect 28368 20726 28488 20754
rect 28354 20632 28410 20641
rect 28354 20567 28410 20576
rect 28368 20534 28396 20567
rect 28356 20528 28408 20534
rect 28356 20470 28408 20476
rect 28354 20360 28410 20369
rect 28354 20295 28356 20304
rect 28408 20295 28410 20304
rect 28356 20266 28408 20272
rect 28262 19816 28318 19825
rect 28262 19751 28318 19760
rect 28276 19718 28304 19751
rect 28264 19712 28316 19718
rect 28264 19654 28316 19660
rect 27896 19314 27948 19320
rect 27724 18834 27844 18850
rect 27712 18828 27844 18834
rect 27764 18822 27844 18828
rect 27712 18770 27764 18776
rect 27580 18720 27660 18748
rect 27528 18702 27580 18708
rect 27342 18663 27398 18672
rect 27344 18624 27396 18630
rect 27344 18566 27396 18572
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 26896 18142 27200 18170
rect 26896 17354 26924 18142
rect 27160 17808 27212 17814
rect 27160 17750 27212 17756
rect 26976 17536 27028 17542
rect 26976 17478 27028 17484
rect 26700 17332 26752 17338
rect 26700 17274 26752 17280
rect 26804 17326 26924 17354
rect 26608 17264 26660 17270
rect 26608 17206 26660 17212
rect 26424 16176 26476 16182
rect 26424 16118 26476 16124
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 26516 16108 26568 16114
rect 26516 16050 26568 16056
rect 25964 16040 26016 16046
rect 25964 15982 26016 15988
rect 25976 12986 26004 15982
rect 26068 14822 26096 16050
rect 26528 15570 26556 16050
rect 26620 15570 26648 17206
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26056 14816 26108 14822
rect 26056 14758 26108 14764
rect 26068 14482 26096 14758
rect 26056 14476 26108 14482
rect 26056 14418 26108 14424
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 26528 14226 26556 15506
rect 26620 14346 26648 15506
rect 26608 14340 26660 14346
rect 26608 14282 26660 14288
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 26160 13818 26188 14010
rect 26160 13790 26280 13818
rect 26148 13728 26200 13734
rect 26148 13670 26200 13676
rect 26160 13326 26188 13670
rect 26148 13320 26200 13326
rect 26148 13262 26200 13268
rect 26252 13190 26280 13790
rect 26344 13410 26372 14214
rect 26528 14198 26648 14226
rect 26344 13382 26556 13410
rect 26332 13320 26384 13326
rect 26332 13262 26384 13268
rect 26240 13184 26292 13190
rect 26240 13126 26292 13132
rect 25964 12980 26016 12986
rect 25964 12922 26016 12928
rect 26056 12912 26108 12918
rect 26056 12854 26108 12860
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 26068 11830 26096 12854
rect 26344 12850 26372 13262
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26332 12640 26384 12646
rect 26332 12582 26384 12588
rect 26344 12306 26372 12582
rect 26332 12300 26384 12306
rect 26332 12242 26384 12248
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 26056 11824 26108 11830
rect 26056 11766 26108 11772
rect 24860 11756 24912 11762
rect 24860 11698 24912 11704
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 24308 11688 24360 11694
rect 24308 11630 24360 11636
rect 24320 11218 24348 11630
rect 26436 11218 26464 12106
rect 26528 11898 26556 13382
rect 26620 12850 26648 14198
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 26804 12646 26832 17326
rect 26884 13184 26936 13190
rect 26884 13126 26936 13132
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 26608 12436 26660 12442
rect 26608 12378 26660 12384
rect 26620 12322 26648 12378
rect 26620 12294 26740 12322
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26620 11898 26648 12174
rect 26712 12084 26740 12294
rect 26896 12238 26924 13126
rect 26988 12374 27016 17478
rect 27068 12844 27120 12850
rect 27068 12786 27120 12792
rect 26976 12368 27028 12374
rect 26976 12310 27028 12316
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26976 12232 27028 12238
rect 26976 12174 27028 12180
rect 26988 12084 27016 12174
rect 26712 12056 27016 12084
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26608 11892 26660 11898
rect 26608 11834 26660 11840
rect 26792 11688 26844 11694
rect 26792 11630 26844 11636
rect 26804 11354 26832 11630
rect 27080 11558 27108 12786
rect 27068 11552 27120 11558
rect 27068 11494 27120 11500
rect 27080 11354 27108 11494
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 27068 11348 27120 11354
rect 27068 11290 27120 11296
rect 24216 11212 24268 11218
rect 24216 11154 24268 11160
rect 24308 11212 24360 11218
rect 24308 11154 24360 11160
rect 26424 11212 26476 11218
rect 26424 11154 26476 11160
rect 26804 11150 26832 11290
rect 27080 11218 27108 11290
rect 27068 11212 27120 11218
rect 27068 11154 27120 11160
rect 27172 11150 27200 17750
rect 27356 17610 27384 18566
rect 27344 17604 27396 17610
rect 27344 17546 27396 17552
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 27252 16584 27304 16590
rect 27252 16526 27304 16532
rect 27264 15706 27292 16526
rect 27356 16454 27384 17138
rect 27344 16448 27396 16454
rect 27344 16390 27396 16396
rect 27344 15904 27396 15910
rect 27344 15846 27396 15852
rect 27252 15700 27304 15706
rect 27252 15642 27304 15648
rect 27356 15502 27384 15846
rect 27344 15496 27396 15502
rect 27344 15438 27396 15444
rect 27448 15434 27476 18686
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27540 17882 27568 18566
rect 27632 18358 27660 18720
rect 27712 18692 27764 18698
rect 27712 18634 27764 18640
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 27528 17876 27580 17882
rect 27528 17818 27580 17824
rect 27540 17134 27568 17818
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 27632 17134 27660 17614
rect 27724 17202 27752 18634
rect 27712 17196 27764 17202
rect 27712 17138 27764 17144
rect 27528 17128 27580 17134
rect 27528 17070 27580 17076
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27724 16794 27752 17138
rect 27712 16788 27764 16794
rect 27712 16730 27764 16736
rect 27816 16658 27844 18822
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27804 16652 27856 16658
rect 27804 16594 27856 16600
rect 27436 15428 27488 15434
rect 27436 15370 27488 15376
rect 27344 15020 27396 15026
rect 27344 14962 27396 14968
rect 27436 15020 27488 15026
rect 27436 14962 27488 14968
rect 27356 14618 27384 14962
rect 27344 14612 27396 14618
rect 27344 14554 27396 14560
rect 27448 14074 27476 14962
rect 27436 14068 27488 14074
rect 27436 14010 27488 14016
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27356 13258 27384 13466
rect 27344 13252 27396 13258
rect 27344 13194 27396 13200
rect 27356 12628 27384 13194
rect 27448 12782 27476 14010
rect 27540 14006 27568 16594
rect 27712 16244 27764 16250
rect 27712 16186 27764 16192
rect 27724 14482 27752 16186
rect 27712 14476 27764 14482
rect 27712 14418 27764 14424
rect 27528 14000 27580 14006
rect 27528 13942 27580 13948
rect 27540 13394 27568 13942
rect 27620 13864 27672 13870
rect 27620 13806 27672 13812
rect 27528 13388 27580 13394
rect 27528 13330 27580 13336
rect 27632 13190 27660 13806
rect 27908 13802 27936 19314
rect 28092 19306 28212 19334
rect 27986 17776 28042 17785
rect 27986 17711 28042 17720
rect 28000 17610 28028 17711
rect 27988 17604 28040 17610
rect 27988 17546 28040 17552
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 28000 14414 28028 14962
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 27896 13796 27948 13802
rect 27896 13738 27948 13744
rect 27804 13388 27856 13394
rect 27804 13330 27856 13336
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27632 12850 27660 13126
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27436 12776 27488 12782
rect 27436 12718 27488 12724
rect 27436 12640 27488 12646
rect 27356 12600 27436 12628
rect 27436 12582 27488 12588
rect 27252 12164 27304 12170
rect 27252 12106 27304 12112
rect 27264 11898 27292 12106
rect 27252 11892 27304 11898
rect 27252 11834 27304 11840
rect 26792 11144 26844 11150
rect 26792 11086 26844 11092
rect 27160 11144 27212 11150
rect 27212 11104 27292 11132
rect 27160 11086 27212 11092
rect 27264 10130 27292 11104
rect 27252 10124 27304 10130
rect 27252 10066 27304 10072
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23848 10056 23900 10062
rect 23848 9998 23900 10004
rect 27160 9988 27212 9994
rect 27160 9930 27212 9936
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 27172 9722 27200 9930
rect 27160 9716 27212 9722
rect 27160 9658 27212 9664
rect 27264 9654 27292 10066
rect 27252 9648 27304 9654
rect 27252 9590 27304 9596
rect 27448 9586 27476 12582
rect 27528 11620 27580 11626
rect 27528 11562 27580 11568
rect 27540 10266 27568 11562
rect 27816 11218 27844 13330
rect 27896 13320 27948 13326
rect 28092 13308 28120 19306
rect 28172 18760 28224 18766
rect 28170 18728 28172 18737
rect 28356 18760 28408 18766
rect 28224 18728 28226 18737
rect 28356 18702 28408 18708
rect 28170 18663 28226 18672
rect 28368 18329 28396 18702
rect 28354 18320 28410 18329
rect 28354 18255 28410 18264
rect 28264 18080 28316 18086
rect 28264 18022 28316 18028
rect 28172 17808 28224 17814
rect 28172 17750 28224 17756
rect 27948 13280 28120 13308
rect 27896 13262 27948 13268
rect 27896 12980 27948 12986
rect 27896 12922 27948 12928
rect 27908 12646 27936 12922
rect 28092 12850 28120 13280
rect 28080 12844 28132 12850
rect 28080 12786 28132 12792
rect 27896 12640 27948 12646
rect 27896 12582 27948 12588
rect 28184 11558 28212 17750
rect 28276 17241 28304 18022
rect 28368 17542 28396 18255
rect 28356 17536 28408 17542
rect 28356 17478 28408 17484
rect 28354 17368 28410 17377
rect 28354 17303 28410 17312
rect 28262 17232 28318 17241
rect 28262 17167 28318 17176
rect 28276 16590 28304 17167
rect 28264 16584 28316 16590
rect 28264 16526 28316 16532
rect 28368 16522 28396 17303
rect 28356 16516 28408 16522
rect 28356 16458 28408 16464
rect 28460 16232 28488 20726
rect 28552 20602 28580 20839
rect 28540 20596 28592 20602
rect 28540 20538 28592 20544
rect 28736 20466 28764 22066
rect 28920 21962 28948 23718
rect 29012 22681 29040 23831
rect 29092 23724 29144 23730
rect 29092 23666 29144 23672
rect 29104 23497 29132 23666
rect 29090 23488 29146 23497
rect 29090 23423 29146 23432
rect 29092 22772 29144 22778
rect 29092 22714 29144 22720
rect 28998 22672 29054 22681
rect 28998 22607 29054 22616
rect 28998 22536 29054 22545
rect 28998 22471 29054 22480
rect 29012 22030 29040 22471
rect 29000 22024 29052 22030
rect 28998 21992 29000 22001
rect 29052 21992 29054 22001
rect 28908 21956 28960 21962
rect 28998 21927 29054 21936
rect 28908 21898 28960 21904
rect 29000 21888 29052 21894
rect 29000 21830 29052 21836
rect 29012 21690 29040 21830
rect 29000 21684 29052 21690
rect 29000 21626 29052 21632
rect 28906 21584 28962 21593
rect 28906 21519 28962 21528
rect 29000 21548 29052 21554
rect 28816 21480 28868 21486
rect 28816 21422 28868 21428
rect 28828 20942 28856 21422
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28816 20800 28868 20806
rect 28816 20742 28868 20748
rect 28724 20460 28776 20466
rect 28724 20402 28776 20408
rect 28540 20392 28592 20398
rect 28540 20334 28592 20340
rect 28552 18834 28580 20334
rect 28724 19984 28776 19990
rect 28724 19926 28776 19932
rect 28736 19446 28764 19926
rect 28724 19440 28776 19446
rect 28724 19382 28776 19388
rect 28724 19168 28776 19174
rect 28724 19110 28776 19116
rect 28632 18964 28684 18970
rect 28632 18906 28684 18912
rect 28644 18873 28672 18906
rect 28630 18864 28686 18873
rect 28540 18828 28592 18834
rect 28630 18799 28686 18808
rect 28540 18770 28592 18776
rect 28538 18184 28594 18193
rect 28538 18119 28594 18128
rect 28552 17542 28580 18119
rect 28632 17604 28684 17610
rect 28632 17546 28684 17552
rect 28540 17536 28592 17542
rect 28540 17478 28592 17484
rect 28540 17196 28592 17202
rect 28540 17138 28592 17144
rect 28276 16204 28488 16232
rect 28276 12782 28304 16204
rect 28552 16114 28580 17138
rect 28644 16794 28672 17546
rect 28632 16788 28684 16794
rect 28632 16730 28684 16736
rect 28448 16108 28500 16114
rect 28448 16050 28500 16056
rect 28540 16108 28592 16114
rect 28540 16050 28592 16056
rect 28460 15706 28488 16050
rect 28448 15700 28500 15706
rect 28448 15642 28500 15648
rect 28460 15026 28488 15642
rect 28552 15570 28580 16050
rect 28540 15564 28592 15570
rect 28540 15506 28592 15512
rect 28448 15020 28500 15026
rect 28448 14962 28500 14968
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 28368 14550 28396 14894
rect 28356 14544 28408 14550
rect 28356 14486 28408 14492
rect 28368 14414 28396 14486
rect 28540 14476 28592 14482
rect 28540 14418 28592 14424
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 28356 13932 28408 13938
rect 28356 13874 28408 13880
rect 28368 12918 28396 13874
rect 28356 12912 28408 12918
rect 28356 12854 28408 12860
rect 28264 12776 28316 12782
rect 28264 12718 28316 12724
rect 28552 12238 28580 14418
rect 28632 13252 28684 13258
rect 28632 13194 28684 13200
rect 28644 12986 28672 13194
rect 28632 12980 28684 12986
rect 28632 12922 28684 12928
rect 28736 12434 28764 19110
rect 28828 16289 28856 20742
rect 28920 20534 28948 21519
rect 29000 21490 29052 21496
rect 29012 21418 29040 21490
rect 29000 21412 29052 21418
rect 29000 21354 29052 21360
rect 28998 20632 29054 20641
rect 28998 20567 29054 20576
rect 28908 20528 28960 20534
rect 28908 20470 28960 20476
rect 29012 19990 29040 20567
rect 29000 19984 29052 19990
rect 28998 19952 29000 19961
rect 29052 19952 29054 19961
rect 28998 19887 29054 19896
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 28814 16280 28870 16289
rect 28814 16215 28870 16224
rect 28816 16108 28868 16114
rect 28816 16050 28868 16056
rect 28828 15162 28856 16050
rect 28816 15156 28868 15162
rect 28816 15098 28868 15104
rect 28920 14074 28948 19790
rect 28998 19544 29054 19553
rect 28998 19479 29054 19488
rect 29012 19446 29040 19479
rect 29000 19440 29052 19446
rect 29000 19382 29052 19388
rect 29000 18624 29052 18630
rect 29000 18566 29052 18572
rect 29012 16998 29040 18566
rect 29104 18290 29132 22714
rect 29196 21554 29224 24754
rect 29276 24200 29328 24206
rect 29276 24142 29328 24148
rect 29288 23798 29316 24142
rect 29276 23792 29328 23798
rect 29276 23734 29328 23740
rect 29276 23656 29328 23662
rect 29276 23598 29328 23604
rect 29288 23254 29316 23598
rect 29276 23248 29328 23254
rect 29276 23190 29328 23196
rect 29276 23112 29328 23118
rect 29276 23054 29328 23060
rect 29288 22438 29316 23054
rect 29276 22432 29328 22438
rect 29276 22374 29328 22380
rect 29288 21622 29316 22374
rect 29276 21616 29328 21622
rect 29276 21558 29328 21564
rect 29184 21548 29236 21554
rect 29184 21490 29236 21496
rect 29276 21072 29328 21078
rect 29276 21014 29328 21020
rect 29288 20466 29316 21014
rect 29276 20460 29328 20466
rect 29276 20402 29328 20408
rect 29182 20360 29238 20369
rect 29182 20295 29238 20304
rect 29092 18284 29144 18290
rect 29092 18226 29144 18232
rect 29090 18184 29146 18193
rect 29090 18119 29146 18128
rect 29104 18086 29132 18119
rect 29092 18080 29144 18086
rect 29092 18022 29144 18028
rect 29196 17270 29224 20295
rect 29288 17610 29316 20402
rect 29380 20398 29408 28902
rect 29472 24886 29500 31991
rect 29564 31822 29592 32388
rect 29552 31816 29604 31822
rect 29552 31758 29604 31764
rect 29552 31680 29604 31686
rect 29552 31622 29604 31628
rect 29564 30977 29592 31622
rect 29550 30968 29606 30977
rect 29550 30903 29606 30912
rect 29552 30796 29604 30802
rect 29552 30738 29604 30744
rect 29564 30190 29592 30738
rect 29552 30184 29604 30190
rect 29552 30126 29604 30132
rect 29550 30016 29606 30025
rect 29550 29951 29606 29960
rect 29564 26761 29592 29951
rect 29656 29209 29684 33254
rect 29748 32978 29776 35652
rect 29828 35634 29880 35640
rect 29920 35692 29972 35698
rect 29920 35634 29972 35640
rect 29932 35154 29960 35634
rect 29920 35148 29972 35154
rect 29920 35090 29972 35096
rect 29826 34368 29882 34377
rect 29826 34303 29882 34312
rect 29840 33590 29868 34303
rect 29828 33584 29880 33590
rect 29828 33526 29880 33532
rect 29736 32972 29788 32978
rect 29788 32932 29868 32960
rect 29736 32914 29788 32920
rect 29736 32836 29788 32842
rect 29736 32778 29788 32784
rect 29748 32473 29776 32778
rect 29840 32502 29868 32932
rect 29828 32496 29880 32502
rect 29734 32464 29790 32473
rect 29828 32438 29880 32444
rect 29734 32399 29790 32408
rect 29828 32224 29880 32230
rect 29828 32166 29880 32172
rect 29840 32042 29868 32166
rect 29748 32014 29868 32042
rect 29748 31793 29776 32014
rect 29828 31884 29880 31890
rect 29828 31826 29880 31832
rect 29734 31784 29790 31793
rect 29734 31719 29790 31728
rect 29736 31408 29788 31414
rect 29734 31376 29736 31385
rect 29788 31376 29790 31385
rect 29734 31311 29790 31320
rect 29736 31136 29788 31142
rect 29736 31078 29788 31084
rect 29748 29753 29776 31078
rect 29840 30734 29868 31826
rect 29828 30728 29880 30734
rect 29828 30670 29880 30676
rect 29828 30592 29880 30598
rect 29828 30534 29880 30540
rect 29840 30394 29868 30534
rect 29828 30388 29880 30394
rect 29828 30330 29880 30336
rect 29828 30184 29880 30190
rect 29932 30172 29960 35090
rect 30024 33930 30052 38791
rect 34244 38752 34296 38758
rect 34244 38694 34296 38700
rect 31944 38616 31996 38622
rect 31944 38558 31996 38564
rect 31760 38344 31812 38350
rect 31760 38286 31812 38292
rect 30564 38072 30616 38078
rect 30194 38040 30250 38049
rect 30564 38014 30616 38020
rect 30656 38072 30708 38078
rect 30656 38014 30708 38020
rect 30194 37975 30250 37984
rect 30102 37904 30158 37913
rect 30102 37839 30158 37848
rect 30116 36825 30144 37839
rect 30102 36816 30158 36825
rect 30102 36751 30158 36760
rect 30116 36242 30144 36751
rect 30104 36236 30156 36242
rect 30104 36178 30156 36184
rect 30104 36100 30156 36106
rect 30104 36042 30156 36048
rect 30116 35018 30144 36042
rect 30104 35012 30156 35018
rect 30104 34954 30156 34960
rect 30104 34604 30156 34610
rect 30104 34546 30156 34552
rect 30012 33924 30064 33930
rect 30012 33866 30064 33872
rect 30024 33522 30052 33866
rect 30012 33516 30064 33522
rect 30012 33458 30064 33464
rect 30024 32473 30052 33458
rect 30010 32464 30066 32473
rect 30116 32434 30144 34546
rect 30208 33658 30236 37975
rect 30288 37256 30340 37262
rect 30288 37198 30340 37204
rect 30300 35601 30328 37198
rect 30380 36236 30432 36242
rect 30380 36178 30432 36184
rect 30392 35630 30420 36178
rect 30380 35624 30432 35630
rect 30286 35592 30342 35601
rect 30380 35566 30432 35572
rect 30286 35527 30342 35536
rect 30288 35488 30340 35494
rect 30286 35456 30288 35465
rect 30340 35456 30342 35465
rect 30286 35391 30342 35400
rect 30300 35193 30328 35391
rect 30286 35184 30342 35193
rect 30286 35119 30342 35128
rect 30392 34728 30420 35566
rect 30472 35488 30524 35494
rect 30472 35430 30524 35436
rect 30300 34700 30420 34728
rect 30300 33998 30328 34700
rect 30380 34604 30432 34610
rect 30380 34546 30432 34552
rect 30288 33992 30340 33998
rect 30288 33934 30340 33940
rect 30196 33652 30248 33658
rect 30196 33594 30248 33600
rect 30208 33454 30236 33594
rect 30196 33448 30248 33454
rect 30196 33390 30248 33396
rect 30194 33280 30250 33289
rect 30194 33215 30250 33224
rect 30208 32910 30236 33215
rect 30196 32904 30248 32910
rect 30196 32846 30248 32852
rect 30010 32399 30066 32408
rect 30104 32428 30156 32434
rect 30024 31958 30052 32399
rect 30104 32370 30156 32376
rect 30012 31952 30064 31958
rect 30012 31894 30064 31900
rect 30104 31884 30156 31890
rect 30104 31826 30156 31832
rect 30012 31816 30064 31822
rect 30012 31758 30064 31764
rect 30024 30802 30052 31758
rect 30116 30802 30144 31826
rect 30208 31822 30236 32846
rect 30300 32586 30328 33934
rect 30392 33522 30420 34546
rect 30484 34241 30512 35430
rect 30470 34232 30526 34241
rect 30470 34167 30526 34176
rect 30472 33856 30524 33862
rect 30472 33798 30524 33804
rect 30380 33516 30432 33522
rect 30380 33458 30432 33464
rect 30378 33416 30434 33425
rect 30378 33351 30434 33360
rect 30392 32978 30420 33351
rect 30484 33114 30512 33798
rect 30576 33658 30604 38014
rect 30668 37738 30696 38014
rect 31392 37800 31444 37806
rect 31392 37742 31444 37748
rect 30656 37732 30708 37738
rect 30656 37674 30708 37680
rect 31116 37188 31168 37194
rect 31116 37130 31168 37136
rect 30840 36168 30892 36174
rect 30840 36110 30892 36116
rect 30656 35624 30708 35630
rect 30656 35566 30708 35572
rect 30668 34610 30696 35566
rect 30748 34944 30800 34950
rect 30746 34912 30748 34921
rect 30800 34912 30802 34921
rect 30746 34847 30802 34856
rect 30746 34776 30802 34785
rect 30746 34711 30802 34720
rect 30760 34610 30788 34711
rect 30656 34604 30708 34610
rect 30656 34546 30708 34552
rect 30748 34604 30800 34610
rect 30748 34546 30800 34552
rect 30668 34513 30696 34546
rect 30654 34504 30710 34513
rect 30654 34439 30710 34448
rect 30852 34406 30880 36110
rect 31024 34536 31076 34542
rect 31024 34478 31076 34484
rect 30840 34400 30892 34406
rect 30840 34342 30892 34348
rect 30654 34232 30710 34241
rect 30654 34167 30710 34176
rect 30668 33697 30696 34167
rect 30748 33924 30800 33930
rect 30748 33866 30800 33872
rect 30654 33688 30710 33697
rect 30564 33652 30616 33658
rect 30654 33623 30710 33632
rect 30564 33594 30616 33600
rect 30656 33312 30708 33318
rect 30576 33272 30656 33300
rect 30472 33108 30524 33114
rect 30472 33050 30524 33056
rect 30380 32972 30432 32978
rect 30380 32914 30432 32920
rect 30300 32558 30420 32586
rect 30288 32496 30340 32502
rect 30288 32438 30340 32444
rect 30300 31890 30328 32438
rect 30288 31884 30340 31890
rect 30288 31826 30340 31832
rect 30196 31816 30248 31822
rect 30196 31758 30248 31764
rect 30196 31680 30248 31686
rect 30196 31622 30248 31628
rect 30208 31414 30236 31622
rect 30196 31408 30248 31414
rect 30196 31350 30248 31356
rect 30196 31136 30248 31142
rect 30196 31078 30248 31084
rect 30012 30796 30064 30802
rect 30012 30738 30064 30744
rect 30104 30796 30156 30802
rect 30104 30738 30156 30744
rect 30116 30394 30144 30738
rect 30208 30394 30236 31078
rect 30392 30920 30420 32558
rect 30470 32464 30526 32473
rect 30470 32399 30526 32408
rect 30484 31929 30512 32399
rect 30470 31920 30526 31929
rect 30470 31855 30472 31864
rect 30524 31855 30526 31864
rect 30472 31826 30524 31832
rect 30576 31754 30604 33272
rect 30656 33254 30708 33260
rect 30656 33108 30708 33114
rect 30656 33050 30708 33056
rect 30668 32434 30696 33050
rect 30656 32428 30708 32434
rect 30656 32370 30708 32376
rect 30668 32201 30696 32370
rect 30654 32192 30710 32201
rect 30654 32127 30710 32136
rect 30484 31726 30604 31754
rect 30484 31249 30512 31726
rect 30668 31521 30696 32127
rect 30654 31512 30710 31521
rect 30654 31447 30710 31456
rect 30668 31346 30696 31447
rect 30656 31340 30708 31346
rect 30656 31282 30708 31288
rect 30470 31240 30526 31249
rect 30760 31226 30788 33866
rect 30470 31175 30526 31184
rect 30576 31198 30788 31226
rect 30852 31210 30880 34342
rect 31036 34218 31064 34478
rect 30944 34190 31064 34218
rect 30944 33114 30972 34190
rect 31024 34128 31076 34134
rect 31024 34070 31076 34076
rect 31036 33522 31064 34070
rect 31024 33516 31076 33522
rect 31024 33458 31076 33464
rect 30932 33108 30984 33114
rect 30932 33050 30984 33056
rect 31024 32972 31076 32978
rect 31024 32914 31076 32920
rect 31036 32434 31064 32914
rect 31024 32428 31076 32434
rect 31024 32370 31076 32376
rect 30932 32360 30984 32366
rect 30932 32302 30984 32308
rect 30944 31890 30972 32302
rect 30932 31884 30984 31890
rect 30932 31826 30984 31832
rect 30930 31648 30986 31657
rect 30930 31583 30986 31592
rect 30840 31204 30892 31210
rect 30484 31142 30512 31175
rect 30472 31136 30524 31142
rect 30472 31078 30524 31084
rect 30300 30892 30420 30920
rect 30104 30388 30156 30394
rect 30104 30330 30156 30336
rect 30196 30388 30248 30394
rect 30196 30330 30248 30336
rect 29880 30144 29960 30172
rect 29828 30126 29880 30132
rect 29840 29850 29868 30126
rect 30116 30122 30144 30330
rect 30300 30258 30328 30892
rect 30380 30796 30432 30802
rect 30380 30738 30432 30744
rect 30392 30666 30420 30738
rect 30380 30660 30432 30666
rect 30380 30602 30432 30608
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30104 30116 30156 30122
rect 30104 30058 30156 30064
rect 30196 30048 30248 30054
rect 30196 29990 30248 29996
rect 29918 29880 29974 29889
rect 29828 29844 29880 29850
rect 29918 29815 29974 29824
rect 29828 29786 29880 29792
rect 29734 29744 29790 29753
rect 29734 29679 29790 29688
rect 29828 29572 29880 29578
rect 29828 29514 29880 29520
rect 29736 29504 29788 29510
rect 29734 29472 29736 29481
rect 29788 29472 29790 29481
rect 29734 29407 29790 29416
rect 29840 29238 29868 29514
rect 29828 29232 29880 29238
rect 29642 29200 29698 29209
rect 29828 29174 29880 29180
rect 29642 29135 29698 29144
rect 29644 27872 29696 27878
rect 29644 27814 29696 27820
rect 29736 27872 29788 27878
rect 29736 27814 29788 27820
rect 29656 27577 29684 27814
rect 29642 27568 29698 27577
rect 29642 27503 29698 27512
rect 29642 27024 29698 27033
rect 29642 26959 29698 26968
rect 29550 26752 29606 26761
rect 29550 26687 29606 26696
rect 29550 26344 29606 26353
rect 29550 26279 29606 26288
rect 29564 25650 29592 26279
rect 29656 25974 29684 26959
rect 29748 26858 29776 27814
rect 29932 27577 29960 29815
rect 30010 29744 30066 29753
rect 30208 29714 30236 29990
rect 30288 29844 30340 29850
rect 30288 29786 30340 29792
rect 30472 29844 30524 29850
rect 30472 29786 30524 29792
rect 30010 29679 30066 29688
rect 30196 29708 30248 29714
rect 30024 27985 30052 29679
rect 30196 29650 30248 29656
rect 30104 29572 30156 29578
rect 30104 29514 30156 29520
rect 30010 27976 30066 27985
rect 30010 27911 30066 27920
rect 30012 27600 30064 27606
rect 29918 27568 29974 27577
rect 30012 27542 30064 27548
rect 29918 27503 29974 27512
rect 29736 26852 29788 26858
rect 29736 26794 29788 26800
rect 29748 26314 29776 26794
rect 29736 26308 29788 26314
rect 29736 26250 29788 26256
rect 29644 25968 29696 25974
rect 29644 25910 29696 25916
rect 29656 25809 29684 25910
rect 29642 25800 29698 25809
rect 29642 25735 29698 25744
rect 29564 25622 29684 25650
rect 29552 25492 29604 25498
rect 29552 25434 29604 25440
rect 29564 25226 29592 25434
rect 29552 25220 29604 25226
rect 29552 25162 29604 25168
rect 29460 24880 29512 24886
rect 29460 24822 29512 24828
rect 29472 24313 29500 24822
rect 29564 24818 29592 25162
rect 29656 24818 29684 25622
rect 29748 25537 29776 26250
rect 29734 25528 29790 25537
rect 29734 25463 29790 25472
rect 29932 25362 29960 27503
rect 30024 27470 30052 27542
rect 30012 27464 30064 27470
rect 30012 27406 30064 27412
rect 30116 27169 30144 29514
rect 30300 29481 30328 29786
rect 30380 29708 30432 29714
rect 30380 29650 30432 29656
rect 30286 29472 30342 29481
rect 30286 29407 30342 29416
rect 30286 28792 30342 28801
rect 30392 28762 30420 29650
rect 30484 29628 30512 29786
rect 30576 29782 30604 31198
rect 30840 31146 30892 31152
rect 30840 30932 30892 30938
rect 30840 30874 30892 30880
rect 30746 30288 30802 30297
rect 30746 30223 30802 30232
rect 30656 30048 30708 30054
rect 30654 30016 30656 30025
rect 30708 30016 30710 30025
rect 30654 29951 30710 29960
rect 30564 29776 30616 29782
rect 30760 29753 30788 30223
rect 30564 29718 30616 29724
rect 30746 29744 30802 29753
rect 30746 29679 30802 29688
rect 30564 29640 30616 29646
rect 30484 29600 30564 29628
rect 30564 29582 30616 29588
rect 30656 29572 30708 29578
rect 30656 29514 30708 29520
rect 30748 29572 30800 29578
rect 30748 29514 30800 29520
rect 30472 29504 30524 29510
rect 30472 29446 30524 29452
rect 30484 29170 30512 29446
rect 30562 29200 30618 29209
rect 30472 29164 30524 29170
rect 30668 29170 30696 29514
rect 30562 29135 30564 29144
rect 30472 29106 30524 29112
rect 30616 29135 30618 29144
rect 30656 29164 30708 29170
rect 30564 29106 30616 29112
rect 30656 29106 30708 29112
rect 30564 29028 30616 29034
rect 30564 28970 30616 28976
rect 30472 28960 30524 28966
rect 30472 28902 30524 28908
rect 30286 28727 30342 28736
rect 30380 28756 30432 28762
rect 30102 27160 30158 27169
rect 30102 27095 30158 27104
rect 30012 26852 30064 26858
rect 30012 26794 30064 26800
rect 30024 25537 30052 26794
rect 30300 26353 30328 28727
rect 30380 28698 30432 28704
rect 30484 28642 30512 28902
rect 30392 28614 30512 28642
rect 30392 28558 30420 28614
rect 30380 28552 30432 28558
rect 30380 28494 30432 28500
rect 30392 27985 30420 28494
rect 30576 28218 30604 28970
rect 30654 28656 30710 28665
rect 30654 28591 30710 28600
rect 30668 28558 30696 28591
rect 30656 28552 30708 28558
rect 30656 28494 30708 28500
rect 30564 28212 30616 28218
rect 30564 28154 30616 28160
rect 30668 28082 30696 28494
rect 30656 28076 30708 28082
rect 30656 28018 30708 28024
rect 30472 28008 30524 28014
rect 30378 27976 30434 27985
rect 30472 27950 30524 27956
rect 30378 27911 30434 27920
rect 30378 27568 30434 27577
rect 30378 27503 30434 27512
rect 30392 27470 30420 27503
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 30392 26790 30420 27406
rect 30380 26784 30432 26790
rect 30380 26726 30432 26732
rect 30484 26586 30512 27950
rect 30564 27668 30616 27674
rect 30564 27610 30616 27616
rect 30576 27470 30604 27610
rect 30656 27600 30708 27606
rect 30656 27542 30708 27548
rect 30564 27464 30616 27470
rect 30564 27406 30616 27412
rect 30576 27033 30604 27406
rect 30562 27024 30618 27033
rect 30562 26959 30618 26968
rect 30472 26580 30524 26586
rect 30472 26522 30524 26528
rect 30668 26518 30696 27542
rect 30760 26926 30788 29514
rect 30852 29209 30880 30874
rect 30944 30433 30972 31583
rect 31022 31240 31078 31249
rect 31022 31175 31078 31184
rect 30930 30424 30986 30433
rect 30930 30359 30986 30368
rect 31036 30025 31064 31175
rect 31022 30016 31078 30025
rect 31022 29951 31078 29960
rect 30932 29232 30984 29238
rect 30838 29200 30894 29209
rect 30932 29174 30984 29180
rect 30838 29135 30894 29144
rect 30944 29050 30972 29174
rect 30852 29022 30972 29050
rect 31024 29096 31076 29102
rect 31024 29038 31076 29044
rect 30852 28014 30880 29022
rect 30930 28928 30986 28937
rect 30930 28863 30986 28872
rect 30840 28008 30892 28014
rect 30838 27976 30840 27985
rect 30892 27976 30894 27985
rect 30838 27911 30894 27920
rect 30748 26920 30800 26926
rect 30748 26862 30800 26868
rect 30748 26580 30800 26586
rect 30748 26522 30800 26528
rect 30656 26512 30708 26518
rect 30656 26454 30708 26460
rect 30286 26344 30342 26353
rect 30286 26279 30342 26288
rect 30472 26240 30524 26246
rect 30472 26182 30524 26188
rect 30102 26072 30158 26081
rect 30102 26007 30158 26016
rect 30010 25528 30066 25537
rect 30010 25463 30066 25472
rect 29920 25356 29972 25362
rect 29920 25298 29972 25304
rect 29932 25140 29960 25298
rect 30024 25265 30052 25463
rect 30010 25256 30066 25265
rect 30010 25191 30066 25200
rect 29932 25112 30052 25140
rect 29552 24812 29604 24818
rect 29552 24754 29604 24760
rect 29644 24812 29696 24818
rect 29644 24754 29696 24760
rect 29458 24304 29514 24313
rect 29458 24239 29514 24248
rect 29564 24206 29592 24754
rect 29656 24614 29684 24754
rect 29644 24608 29696 24614
rect 29644 24550 29696 24556
rect 29644 24336 29696 24342
rect 29696 24284 29868 24290
rect 29644 24278 29868 24284
rect 29656 24262 29868 24278
rect 29552 24200 29604 24206
rect 29840 24188 29868 24262
rect 29840 24160 29960 24188
rect 29552 24142 29604 24148
rect 29564 23866 29592 24142
rect 29826 24032 29882 24041
rect 29826 23967 29882 23976
rect 29460 23860 29512 23866
rect 29460 23802 29512 23808
rect 29552 23860 29604 23866
rect 29552 23802 29604 23808
rect 29472 23633 29500 23802
rect 29734 23760 29790 23769
rect 29734 23695 29790 23704
rect 29458 23624 29514 23633
rect 29748 23594 29776 23695
rect 29458 23559 29514 23568
rect 29736 23588 29788 23594
rect 29736 23530 29788 23536
rect 29644 23520 29696 23526
rect 29644 23462 29696 23468
rect 29458 23216 29514 23225
rect 29458 23151 29514 23160
rect 29472 22642 29500 23151
rect 29656 22642 29684 23462
rect 29736 23112 29788 23118
rect 29736 23054 29788 23060
rect 29748 22817 29776 23054
rect 29734 22808 29790 22817
rect 29734 22743 29790 22752
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 29644 22636 29696 22642
rect 29644 22578 29696 22584
rect 29550 22536 29606 22545
rect 29550 22471 29552 22480
rect 29604 22471 29606 22480
rect 29552 22442 29604 22448
rect 29550 22128 29606 22137
rect 29840 22094 29868 23967
rect 29550 22063 29552 22072
rect 29604 22063 29606 22072
rect 29748 22066 29868 22094
rect 29552 22034 29604 22040
rect 29460 21480 29512 21486
rect 29460 21422 29512 21428
rect 29472 20942 29500 21422
rect 29552 21344 29604 21350
rect 29552 21286 29604 21292
rect 29564 21010 29592 21286
rect 29552 21004 29604 21010
rect 29552 20946 29604 20952
rect 29460 20936 29512 20942
rect 29460 20878 29512 20884
rect 29368 20392 29420 20398
rect 29368 20334 29420 20340
rect 29472 20244 29500 20878
rect 29748 20641 29776 22066
rect 29828 21684 29880 21690
rect 29828 21626 29880 21632
rect 29734 20632 29790 20641
rect 29734 20567 29790 20576
rect 29550 20496 29606 20505
rect 29550 20431 29606 20440
rect 29380 20216 29500 20244
rect 29380 19310 29408 20216
rect 29458 19816 29514 19825
rect 29458 19751 29460 19760
rect 29512 19751 29514 19760
rect 29460 19722 29512 19728
rect 29460 19440 29512 19446
rect 29460 19382 29512 19388
rect 29368 19304 29420 19310
rect 29368 19246 29420 19252
rect 29368 18896 29420 18902
rect 29366 18864 29368 18873
rect 29420 18864 29422 18873
rect 29472 18834 29500 19382
rect 29366 18799 29422 18808
rect 29460 18828 29512 18834
rect 29460 18770 29512 18776
rect 29368 18692 29420 18698
rect 29368 18634 29420 18640
rect 29276 17604 29328 17610
rect 29276 17546 29328 17552
rect 29184 17264 29236 17270
rect 29184 17206 29236 17212
rect 29006 16992 29058 16998
rect 29006 16934 29058 16940
rect 29092 16788 29144 16794
rect 29092 16730 29144 16736
rect 28998 16688 29054 16697
rect 29104 16674 29132 16730
rect 29182 16688 29238 16697
rect 29104 16646 29182 16674
rect 28998 16623 29054 16632
rect 29182 16623 29238 16632
rect 29012 15706 29040 16623
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 28908 14068 28960 14074
rect 28908 14010 28960 14016
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 28816 13796 28868 13802
rect 28816 13738 28868 13744
rect 28828 13326 28856 13738
rect 28816 13320 28868 13326
rect 28816 13262 28868 13268
rect 28736 12406 28856 12434
rect 28632 12300 28684 12306
rect 28632 12242 28684 12248
rect 28540 12232 28592 12238
rect 28540 12174 28592 12180
rect 28552 11898 28580 12174
rect 28540 11892 28592 11898
rect 28540 11834 28592 11840
rect 28644 11830 28672 12242
rect 28632 11824 28684 11830
rect 28632 11766 28684 11772
rect 28724 11756 28776 11762
rect 28724 11698 28776 11704
rect 28172 11552 28224 11558
rect 28172 11494 28224 11500
rect 27804 11212 27856 11218
rect 27804 11154 27856 11160
rect 27816 10674 27844 11154
rect 28736 10810 28764 11698
rect 28724 10804 28776 10810
rect 28724 10746 28776 10752
rect 27712 10668 27764 10674
rect 27712 10610 27764 10616
rect 27804 10668 27856 10674
rect 27804 10610 27856 10616
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 27724 10266 27752 10610
rect 27528 10260 27580 10266
rect 27528 10202 27580 10208
rect 27712 10260 27764 10266
rect 27712 10202 27764 10208
rect 27540 9722 27568 10202
rect 27816 10062 27844 10610
rect 27804 10056 27856 10062
rect 27804 9998 27856 10004
rect 28368 9722 28396 10610
rect 28736 10062 28764 10746
rect 28724 10056 28776 10062
rect 28724 9998 28776 10004
rect 28828 9722 28856 12406
rect 29012 12374 29040 13806
rect 29276 13184 29328 13190
rect 29276 13126 29328 13132
rect 29092 12980 29144 12986
rect 29092 12922 29144 12928
rect 29104 12782 29132 12922
rect 29288 12850 29316 13126
rect 29380 12918 29408 18634
rect 29472 18290 29500 18770
rect 29460 18284 29512 18290
rect 29460 18226 29512 18232
rect 29472 14822 29500 18226
rect 29564 16522 29592 20431
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29644 20256 29696 20262
rect 29644 20198 29696 20204
rect 29656 19786 29684 20198
rect 29644 19780 29696 19786
rect 29644 19722 29696 19728
rect 29644 19304 29696 19310
rect 29644 19246 29696 19252
rect 29656 17542 29684 19246
rect 29748 17678 29776 20334
rect 29840 18850 29868 21626
rect 29932 19378 29960 24160
rect 30024 23644 30052 25112
rect 30116 23798 30144 26007
rect 30196 25968 30248 25974
rect 30196 25910 30248 25916
rect 30208 25770 30236 25910
rect 30286 25800 30342 25809
rect 30196 25764 30248 25770
rect 30286 25735 30342 25744
rect 30196 25706 30248 25712
rect 30194 25664 30250 25673
rect 30194 25599 30250 25608
rect 30208 25378 30236 25599
rect 30300 25498 30328 25735
rect 30484 25702 30512 26182
rect 30562 25936 30618 25945
rect 30562 25871 30618 25880
rect 30576 25770 30604 25871
rect 30564 25764 30616 25770
rect 30564 25706 30616 25712
rect 30380 25696 30432 25702
rect 30380 25638 30432 25644
rect 30472 25696 30524 25702
rect 30472 25638 30524 25644
rect 30288 25492 30340 25498
rect 30288 25434 30340 25440
rect 30208 25350 30328 25378
rect 30300 25294 30328 25350
rect 30196 25288 30248 25294
rect 30196 25230 30248 25236
rect 30288 25288 30340 25294
rect 30288 25230 30340 25236
rect 30208 25158 30236 25230
rect 30196 25152 30248 25158
rect 30196 25094 30248 25100
rect 30208 24818 30236 25094
rect 30288 24880 30340 24886
rect 30288 24822 30340 24828
rect 30196 24812 30248 24818
rect 30196 24754 30248 24760
rect 30208 24206 30236 24754
rect 30300 24698 30328 24822
rect 30392 24818 30420 25638
rect 30472 25492 30524 25498
rect 30472 25434 30524 25440
rect 30484 25226 30512 25434
rect 30576 25226 30604 25706
rect 30472 25220 30524 25226
rect 30472 25162 30524 25168
rect 30564 25220 30616 25226
rect 30564 25162 30616 25168
rect 30470 24984 30526 24993
rect 30470 24919 30526 24928
rect 30484 24886 30512 24919
rect 30472 24880 30524 24886
rect 30472 24822 30524 24828
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 30300 24670 30512 24698
rect 30484 24614 30512 24670
rect 30288 24608 30340 24614
rect 30380 24608 30432 24614
rect 30288 24550 30340 24556
rect 30378 24576 30380 24585
rect 30472 24608 30524 24614
rect 30432 24576 30434 24585
rect 30300 24206 30328 24550
rect 30472 24550 30524 24556
rect 30378 24511 30434 24520
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30196 24200 30248 24206
rect 30196 24142 30248 24148
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30104 23792 30156 23798
rect 30104 23734 30156 23740
rect 30392 23730 30420 24346
rect 30472 24336 30524 24342
rect 30472 24278 30524 24284
rect 30196 23724 30248 23730
rect 30196 23666 30248 23672
rect 30380 23724 30432 23730
rect 30380 23666 30432 23672
rect 30024 23616 30144 23644
rect 30010 23216 30066 23225
rect 30010 23151 30066 23160
rect 30024 23118 30052 23151
rect 30012 23112 30064 23118
rect 30012 23054 30064 23060
rect 30012 22976 30064 22982
rect 30012 22918 30064 22924
rect 30024 22234 30052 22918
rect 30012 22228 30064 22234
rect 30012 22170 30064 22176
rect 30116 22114 30144 23616
rect 30208 23118 30236 23666
rect 30380 23520 30432 23526
rect 30380 23462 30432 23468
rect 30392 23186 30420 23462
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 30196 23112 30248 23118
rect 30196 23054 30248 23060
rect 30288 22976 30340 22982
rect 30286 22944 30288 22953
rect 30380 22976 30432 22982
rect 30340 22944 30342 22953
rect 30380 22918 30432 22924
rect 30286 22879 30342 22888
rect 30392 22710 30420 22918
rect 30484 22778 30512 24278
rect 30576 22982 30604 25162
rect 30668 24818 30696 26454
rect 30760 26382 30788 26522
rect 30944 26489 30972 28863
rect 31036 28762 31064 29038
rect 31024 28756 31076 28762
rect 31024 28698 31076 28704
rect 31036 28422 31064 28698
rect 31024 28416 31076 28422
rect 31024 28358 31076 28364
rect 31024 27396 31076 27402
rect 31024 27338 31076 27344
rect 31036 26994 31064 27338
rect 31024 26988 31076 26994
rect 31024 26930 31076 26936
rect 31036 26518 31064 26930
rect 31128 26926 31156 37130
rect 31300 36712 31352 36718
rect 31206 36680 31262 36689
rect 31300 36654 31352 36660
rect 31206 36615 31262 36624
rect 31220 35698 31248 36615
rect 31208 35692 31260 35698
rect 31208 35634 31260 35640
rect 31220 34134 31248 35634
rect 31312 35018 31340 36654
rect 31300 35012 31352 35018
rect 31300 34954 31352 34960
rect 31312 34542 31340 34954
rect 31300 34536 31352 34542
rect 31300 34478 31352 34484
rect 31208 34128 31260 34134
rect 31208 34070 31260 34076
rect 31220 33998 31248 34070
rect 31404 33998 31432 37742
rect 31668 36712 31720 36718
rect 31668 36654 31720 36660
rect 31484 35080 31536 35086
rect 31484 35022 31536 35028
rect 31208 33992 31260 33998
rect 31208 33934 31260 33940
rect 31392 33992 31444 33998
rect 31392 33934 31444 33940
rect 31496 32978 31524 35022
rect 31574 34912 31630 34921
rect 31574 34847 31630 34856
rect 31588 34202 31616 34847
rect 31576 34196 31628 34202
rect 31576 34138 31628 34144
rect 31484 32972 31536 32978
rect 31484 32914 31536 32920
rect 31206 32736 31262 32745
rect 31206 32671 31262 32680
rect 31220 32502 31248 32671
rect 31208 32496 31260 32502
rect 31208 32438 31260 32444
rect 31208 31884 31260 31890
rect 31208 31826 31260 31832
rect 31220 31278 31248 31826
rect 31496 31822 31524 32914
rect 31576 32428 31628 32434
rect 31576 32370 31628 32376
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 31392 31340 31444 31346
rect 31392 31282 31444 31288
rect 31208 31272 31260 31278
rect 31208 31214 31260 31220
rect 31208 31136 31260 31142
rect 31208 31078 31260 31084
rect 31220 30938 31248 31078
rect 31208 30932 31260 30938
rect 31208 30874 31260 30880
rect 31404 30598 31432 31282
rect 31496 30870 31524 31758
rect 31588 31686 31616 32370
rect 31576 31680 31628 31686
rect 31576 31622 31628 31628
rect 31680 31498 31708 36654
rect 31772 35766 31800 38286
rect 31850 36952 31906 36961
rect 31850 36887 31852 36896
rect 31904 36887 31906 36896
rect 31852 36858 31904 36864
rect 31864 36242 31892 36858
rect 31852 36236 31904 36242
rect 31852 36178 31904 36184
rect 31956 36106 31984 38558
rect 32496 38480 32548 38486
rect 32496 38422 32548 38428
rect 32404 37324 32456 37330
rect 32404 37266 32456 37272
rect 32036 37256 32088 37262
rect 32312 37256 32364 37262
rect 32036 37198 32088 37204
rect 32310 37224 32312 37233
rect 32364 37224 32366 37233
rect 32048 36378 32076 37198
rect 32310 37159 32366 37168
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 32232 36786 32260 37062
rect 32220 36780 32272 36786
rect 32220 36722 32272 36728
rect 32036 36372 32088 36378
rect 32036 36314 32088 36320
rect 32324 36281 32352 37159
rect 32310 36272 32366 36281
rect 32310 36207 32366 36216
rect 31944 36100 31996 36106
rect 31944 36042 31996 36048
rect 32310 35864 32366 35873
rect 32310 35799 32312 35808
rect 32364 35799 32366 35808
rect 32312 35770 32364 35776
rect 31760 35760 31812 35766
rect 31760 35702 31812 35708
rect 32128 35624 32180 35630
rect 32128 35566 32180 35572
rect 32140 35290 32168 35566
rect 32310 35456 32366 35465
rect 32310 35391 32366 35400
rect 32128 35284 32180 35290
rect 32128 35226 32180 35232
rect 31852 35148 31904 35154
rect 31852 35090 31904 35096
rect 31758 35048 31814 35057
rect 31758 34983 31814 34992
rect 31772 34105 31800 34983
rect 31864 34746 31892 35090
rect 32034 34776 32090 34785
rect 31852 34740 31904 34746
rect 32034 34711 32090 34720
rect 31852 34682 31904 34688
rect 31942 34640 31998 34649
rect 31942 34575 31998 34584
rect 31852 34196 31904 34202
rect 31852 34138 31904 34144
rect 31758 34096 31814 34105
rect 31864 34066 31892 34138
rect 31758 34031 31814 34040
rect 31852 34060 31904 34066
rect 31852 34002 31904 34008
rect 31956 33697 31984 34575
rect 31942 33688 31998 33697
rect 31942 33623 31998 33632
rect 31760 33040 31812 33046
rect 31760 32982 31812 32988
rect 31772 32774 31800 32982
rect 31760 32768 31812 32774
rect 31760 32710 31812 32716
rect 31944 32428 31996 32434
rect 31944 32370 31996 32376
rect 31956 32026 31984 32370
rect 31760 32020 31812 32026
rect 31760 31962 31812 31968
rect 31944 32020 31996 32026
rect 31944 31962 31996 31968
rect 31588 31470 31708 31498
rect 31484 30864 31536 30870
rect 31484 30806 31536 30812
rect 31392 30592 31444 30598
rect 31298 30560 31354 30569
rect 31392 30534 31444 30540
rect 31298 30495 31354 30504
rect 31208 30048 31260 30054
rect 31208 29990 31260 29996
rect 31220 28966 31248 29990
rect 31312 29646 31340 30495
rect 31404 29646 31432 30534
rect 31300 29640 31352 29646
rect 31300 29582 31352 29588
rect 31392 29640 31444 29646
rect 31392 29582 31444 29588
rect 31312 29492 31340 29582
rect 31496 29510 31524 30806
rect 31484 29504 31536 29510
rect 31312 29464 31432 29492
rect 31300 29164 31352 29170
rect 31300 29106 31352 29112
rect 31208 28960 31260 28966
rect 31208 28902 31260 28908
rect 31312 28626 31340 29106
rect 31300 28620 31352 28626
rect 31300 28562 31352 28568
rect 31312 28098 31340 28562
rect 31220 28070 31340 28098
rect 31116 26920 31168 26926
rect 31116 26862 31168 26868
rect 31024 26512 31076 26518
rect 30930 26480 30986 26489
rect 31024 26454 31076 26460
rect 30930 26415 30986 26424
rect 31220 26382 31248 28070
rect 31300 27396 31352 27402
rect 31300 27338 31352 27344
rect 30748 26376 30800 26382
rect 30932 26376 30984 26382
rect 30748 26318 30800 26324
rect 30930 26344 30932 26353
rect 31208 26376 31260 26382
rect 30984 26344 30986 26353
rect 31208 26318 31260 26324
rect 30930 26279 30986 26288
rect 30748 26240 30800 26246
rect 30748 26182 30800 26188
rect 31208 26240 31260 26246
rect 31208 26182 31260 26188
rect 30760 25922 30788 26182
rect 31220 26024 31248 26182
rect 31129 25996 31248 26024
rect 31129 25922 31157 25996
rect 30760 25894 30972 25922
rect 30748 25832 30800 25838
rect 30748 25774 30800 25780
rect 30656 24812 30708 24818
rect 30656 24754 30708 24760
rect 30668 24138 30696 24754
rect 30760 24585 30788 25774
rect 30944 25673 30972 25894
rect 31036 25894 31157 25922
rect 31206 25936 31262 25945
rect 30930 25664 30986 25673
rect 30930 25599 30986 25608
rect 30932 25424 30984 25430
rect 30932 25366 30984 25372
rect 30944 24857 30972 25366
rect 30930 24848 30986 24857
rect 30930 24783 30986 24792
rect 30840 24608 30892 24614
rect 30746 24576 30802 24585
rect 30840 24550 30892 24556
rect 30746 24511 30802 24520
rect 30656 24132 30708 24138
rect 30656 24074 30708 24080
rect 30668 23594 30696 24074
rect 30852 24070 30880 24550
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 30838 23896 30894 23905
rect 30838 23831 30894 23840
rect 30746 23760 30802 23769
rect 30746 23695 30802 23704
rect 30656 23588 30708 23594
rect 30656 23530 30708 23536
rect 30668 23225 30696 23530
rect 30654 23216 30710 23225
rect 30654 23151 30710 23160
rect 30654 23080 30710 23089
rect 30654 23015 30710 23024
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30380 22704 30432 22710
rect 30380 22646 30432 22652
rect 30194 22536 30250 22545
rect 30194 22471 30250 22480
rect 30024 22086 30144 22114
rect 30024 21690 30052 22086
rect 30104 22024 30156 22030
rect 30104 21966 30156 21972
rect 30116 21865 30144 21966
rect 30102 21856 30158 21865
rect 30102 21791 30158 21800
rect 30012 21684 30064 21690
rect 30012 21626 30064 21632
rect 30208 21622 30236 22471
rect 30378 22128 30434 22137
rect 30378 22063 30434 22072
rect 30392 21962 30420 22063
rect 30470 21992 30526 22001
rect 30380 21956 30432 21962
rect 30470 21927 30526 21936
rect 30564 21956 30616 21962
rect 30380 21898 30432 21904
rect 30196 21616 30248 21622
rect 30288 21616 30340 21622
rect 30196 21558 30248 21564
rect 30286 21584 30288 21593
rect 30340 21584 30342 21593
rect 30286 21519 30342 21528
rect 30484 21418 30512 21927
rect 30564 21898 30616 21904
rect 30472 21412 30524 21418
rect 30472 21354 30524 21360
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 30012 21004 30064 21010
rect 30012 20946 30064 20952
rect 30024 19514 30052 20946
rect 30012 19508 30064 19514
rect 30012 19450 30064 19456
rect 30024 19394 30052 19450
rect 29920 19372 29972 19378
rect 30024 19366 30144 19394
rect 29920 19314 29972 19320
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 29918 19000 29974 19009
rect 29918 18935 29920 18944
rect 29972 18935 29974 18944
rect 29920 18906 29972 18912
rect 30024 18902 30052 19110
rect 30012 18896 30064 18902
rect 29840 18822 29960 18850
rect 30012 18838 30064 18844
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29840 17898 29868 18702
rect 29932 18426 29960 18822
rect 30012 18760 30064 18766
rect 30012 18702 30064 18708
rect 30024 18601 30052 18702
rect 30010 18592 30066 18601
rect 30010 18527 30066 18536
rect 29920 18420 29972 18426
rect 29920 18362 29972 18368
rect 30012 18148 30064 18154
rect 30012 18090 30064 18096
rect 30024 18057 30052 18090
rect 30010 18048 30066 18057
rect 30010 17983 30066 17992
rect 29840 17870 30052 17898
rect 29736 17672 29788 17678
rect 29736 17614 29788 17620
rect 29644 17536 29696 17542
rect 29644 17478 29696 17484
rect 30024 17354 30052 17870
rect 29932 17338 30052 17354
rect 30116 17338 30144 19366
rect 29920 17332 30052 17338
rect 29972 17326 30052 17332
rect 29920 17274 29972 17280
rect 29736 17264 29788 17270
rect 29736 17206 29788 17212
rect 29552 16516 29604 16522
rect 29552 16458 29604 16464
rect 29564 16046 29592 16458
rect 29552 16040 29604 16046
rect 29552 15982 29604 15988
rect 29564 15502 29592 15982
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 29552 15360 29604 15366
rect 29552 15302 29604 15308
rect 29460 14816 29512 14822
rect 29460 14758 29512 14764
rect 29460 13184 29512 13190
rect 29460 13126 29512 13132
rect 29472 12986 29500 13126
rect 29460 12980 29512 12986
rect 29460 12922 29512 12928
rect 29368 12912 29420 12918
rect 29368 12854 29420 12860
rect 29276 12844 29328 12850
rect 29276 12786 29328 12792
rect 29092 12776 29144 12782
rect 29092 12718 29144 12724
rect 29000 12368 29052 12374
rect 29000 12310 29052 12316
rect 29564 12306 29592 15302
rect 29748 15094 29776 17206
rect 29920 15904 29972 15910
rect 29920 15846 29972 15852
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29736 15088 29788 15094
rect 29736 15030 29788 15036
rect 29644 14000 29696 14006
rect 29644 13942 29696 13948
rect 29656 12434 29684 13942
rect 29840 13394 29868 15438
rect 29932 15162 29960 15846
rect 29920 15156 29972 15162
rect 29920 15098 29972 15104
rect 29932 14006 29960 15098
rect 29920 14000 29972 14006
rect 29920 13942 29972 13948
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 29656 12406 29776 12434
rect 29552 12300 29604 12306
rect 29552 12242 29604 12248
rect 29000 12232 29052 12238
rect 29000 12174 29052 12180
rect 29184 12232 29236 12238
rect 29184 12174 29236 12180
rect 27528 9716 27580 9722
rect 27528 9658 27580 9664
rect 28356 9716 28408 9722
rect 28356 9658 28408 9664
rect 28816 9716 28868 9722
rect 28816 9658 28868 9664
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 29012 9382 29040 12174
rect 29196 9518 29224 12174
rect 29748 12170 29776 12406
rect 29644 12164 29696 12170
rect 29644 12106 29696 12112
rect 29736 12164 29788 12170
rect 29736 12106 29788 12112
rect 29552 11552 29604 11558
rect 29552 11494 29604 11500
rect 29564 11150 29592 11494
rect 29552 11144 29604 11150
rect 29552 11086 29604 11092
rect 29656 10810 29684 12106
rect 29644 10804 29696 10810
rect 29644 10746 29696 10752
rect 29460 10464 29512 10470
rect 29460 10406 29512 10412
rect 29472 9654 29500 10406
rect 29748 9926 29776 12106
rect 29840 11218 29868 13330
rect 29920 12844 29972 12850
rect 29920 12786 29972 12792
rect 29932 12238 29960 12786
rect 29920 12232 29972 12238
rect 29920 12174 29972 12180
rect 30024 11898 30052 17326
rect 30104 17332 30156 17338
rect 30104 17274 30156 17280
rect 30104 16788 30156 16794
rect 30104 16730 30156 16736
rect 30116 16697 30144 16730
rect 30102 16688 30158 16697
rect 30102 16623 30158 16632
rect 30208 16425 30236 21286
rect 30576 21146 30604 21898
rect 30668 21554 30696 23015
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 30760 21418 30788 23695
rect 30852 23322 30880 23831
rect 30932 23724 30984 23730
rect 30932 23666 30984 23672
rect 30840 23316 30892 23322
rect 30840 23258 30892 23264
rect 30838 22672 30894 22681
rect 30838 22607 30840 22616
rect 30892 22607 30894 22616
rect 30840 22578 30892 22584
rect 30852 22166 30880 22578
rect 30944 22574 30972 23666
rect 31036 23118 31064 25894
rect 31206 25871 31262 25880
rect 31114 25664 31170 25673
rect 31114 25599 31170 25608
rect 31128 25158 31156 25599
rect 31116 25152 31168 25158
rect 31116 25094 31168 25100
rect 31128 24750 31156 25094
rect 31220 24954 31248 25871
rect 31312 25820 31340 27338
rect 31404 26382 31432 29464
rect 31484 29446 31536 29452
rect 31484 29096 31536 29102
rect 31482 29064 31484 29073
rect 31536 29064 31538 29073
rect 31482 28999 31538 29008
rect 31484 28756 31536 28762
rect 31484 28698 31536 28704
rect 31392 26376 31444 26382
rect 31392 26318 31444 26324
rect 31392 25832 31444 25838
rect 31312 25792 31392 25820
rect 31208 24948 31260 24954
rect 31208 24890 31260 24896
rect 31312 24886 31340 25792
rect 31392 25774 31444 25780
rect 31390 25664 31446 25673
rect 31390 25599 31446 25608
rect 31404 25498 31432 25599
rect 31392 25492 31444 25498
rect 31392 25434 31444 25440
rect 31392 25356 31444 25362
rect 31392 25298 31444 25304
rect 31300 24880 31352 24886
rect 31300 24822 31352 24828
rect 31404 24818 31432 25298
rect 31496 25294 31524 28698
rect 31588 28082 31616 31470
rect 31772 31278 31800 31962
rect 31852 31884 31904 31890
rect 31852 31826 31904 31832
rect 31760 31272 31812 31278
rect 31760 31214 31812 31220
rect 31760 30932 31812 30938
rect 31760 30874 31812 30880
rect 31668 30796 31720 30802
rect 31668 30738 31720 30744
rect 31680 30326 31708 30738
rect 31772 30734 31800 30874
rect 31864 30734 31892 31826
rect 31760 30728 31812 30734
rect 31760 30670 31812 30676
rect 31852 30728 31904 30734
rect 31852 30670 31904 30676
rect 31864 30433 31892 30670
rect 31850 30424 31906 30433
rect 31850 30359 31906 30368
rect 31668 30320 31720 30326
rect 31668 30262 31720 30268
rect 31850 30288 31906 30297
rect 31850 30223 31906 30232
rect 31760 30184 31812 30190
rect 31760 30126 31812 30132
rect 31668 30048 31720 30054
rect 31668 29990 31720 29996
rect 31680 28558 31708 29990
rect 31772 28994 31800 30126
rect 31864 29186 31892 30223
rect 31956 30190 31984 31962
rect 32048 31793 32076 34711
rect 32140 34377 32168 35226
rect 32126 34368 32182 34377
rect 32126 34303 32182 34312
rect 32128 34128 32180 34134
rect 32128 34070 32180 34076
rect 32140 33046 32168 34070
rect 32324 33425 32352 35391
rect 32416 35154 32444 37266
rect 32404 35148 32456 35154
rect 32404 35090 32456 35096
rect 32404 34468 32456 34474
rect 32404 34410 32456 34416
rect 32310 33416 32366 33425
rect 32310 33351 32366 33360
rect 32128 33040 32180 33046
rect 32128 32982 32180 32988
rect 32140 32910 32168 32982
rect 32324 32910 32352 33351
rect 32128 32904 32180 32910
rect 32128 32846 32180 32852
rect 32312 32904 32364 32910
rect 32312 32846 32364 32852
rect 32312 32428 32364 32434
rect 32312 32370 32364 32376
rect 32324 32337 32352 32370
rect 32310 32328 32366 32337
rect 32310 32263 32366 32272
rect 32416 32230 32444 34410
rect 32508 34406 32536 38422
rect 33692 38208 33744 38214
rect 33692 38150 33744 38156
rect 32772 38072 32824 38078
rect 32772 38014 32824 38020
rect 32588 37256 32640 37262
rect 32588 37198 32640 37204
rect 32600 36582 32628 37198
rect 32588 36576 32640 36582
rect 32588 36518 32640 36524
rect 32784 35834 32812 38014
rect 33324 37868 33376 37874
rect 33324 37810 33376 37816
rect 32956 37460 33008 37466
rect 32956 37402 33008 37408
rect 32968 36825 32996 37402
rect 33140 37256 33192 37262
rect 33140 37198 33192 37204
rect 32954 36816 33010 36825
rect 32954 36751 33010 36760
rect 33048 36780 33100 36786
rect 32864 36304 32916 36310
rect 32864 36246 32916 36252
rect 32772 35828 32824 35834
rect 32772 35770 32824 35776
rect 32588 35760 32640 35766
rect 32588 35702 32640 35708
rect 32496 34400 32548 34406
rect 32496 34342 32548 34348
rect 32496 34060 32548 34066
rect 32496 34002 32548 34008
rect 32508 33590 32536 34002
rect 32496 33584 32548 33590
rect 32496 33526 32548 33532
rect 32600 33386 32628 35702
rect 32680 35624 32732 35630
rect 32680 35566 32732 35572
rect 32692 35494 32720 35566
rect 32680 35488 32732 35494
rect 32680 35430 32732 35436
rect 32772 35080 32824 35086
rect 32772 35022 32824 35028
rect 32680 35012 32732 35018
rect 32680 34954 32732 34960
rect 32692 34649 32720 34954
rect 32678 34640 32734 34649
rect 32678 34575 32734 34584
rect 32680 34536 32732 34542
rect 32678 34504 32680 34513
rect 32732 34504 32734 34513
rect 32678 34439 32734 34448
rect 32588 33380 32640 33386
rect 32588 33322 32640 33328
rect 32692 33266 32720 34439
rect 32784 33318 32812 35022
rect 32876 34610 32904 36246
rect 32968 36242 32996 36751
rect 33048 36722 33100 36728
rect 32956 36236 33008 36242
rect 32956 36178 33008 36184
rect 32956 35828 33008 35834
rect 32956 35770 33008 35776
rect 32968 35290 32996 35770
rect 33060 35698 33088 36722
rect 33048 35692 33100 35698
rect 33048 35634 33100 35640
rect 32956 35284 33008 35290
rect 32956 35226 33008 35232
rect 33152 35034 33180 37198
rect 33232 36576 33284 36582
rect 33232 36518 33284 36524
rect 33244 35630 33272 36518
rect 33336 36038 33364 37810
rect 33704 37330 33732 38150
rect 34152 37664 34204 37670
rect 34152 37606 34204 37612
rect 33692 37324 33744 37330
rect 33692 37266 33744 37272
rect 33784 37256 33836 37262
rect 33784 37198 33836 37204
rect 33324 36032 33376 36038
rect 33324 35974 33376 35980
rect 33416 36032 33468 36038
rect 33416 35974 33468 35980
rect 33336 35834 33364 35974
rect 33324 35828 33376 35834
rect 33324 35770 33376 35776
rect 33324 35692 33376 35698
rect 33324 35634 33376 35640
rect 33232 35624 33284 35630
rect 33232 35566 33284 35572
rect 33336 35193 33364 35634
rect 33428 35465 33456 35974
rect 33796 35816 33824 37198
rect 34164 36768 34192 37606
rect 34256 37262 34284 38694
rect 34900 37754 34928 39200
rect 35622 38992 35678 39001
rect 35622 38927 35678 38936
rect 35530 38448 35586 38457
rect 35530 38383 35586 38392
rect 35438 38312 35494 38321
rect 35438 38247 35494 38256
rect 35348 38140 35400 38146
rect 35348 38082 35400 38088
rect 34808 37726 34928 37754
rect 34520 37392 34572 37398
rect 34520 37334 34572 37340
rect 34702 37360 34758 37369
rect 34244 37256 34296 37262
rect 34244 37198 34296 37204
rect 34532 36786 34560 37334
rect 34702 37295 34758 37304
rect 34520 36780 34572 36786
rect 34164 36740 34284 36768
rect 34152 36644 34204 36650
rect 34152 36586 34204 36592
rect 33874 36408 33930 36417
rect 33874 36343 33930 36352
rect 33704 35788 33824 35816
rect 33600 35488 33652 35494
rect 33414 35456 33470 35465
rect 33600 35430 33652 35436
rect 33414 35391 33470 35400
rect 33414 35320 33470 35329
rect 33414 35255 33470 35264
rect 33322 35184 33378 35193
rect 33322 35119 33378 35128
rect 32968 35006 33180 35034
rect 32864 34604 32916 34610
rect 32864 34546 32916 34552
rect 32864 34468 32916 34474
rect 32864 34410 32916 34416
rect 32876 34241 32904 34410
rect 32862 34232 32918 34241
rect 32862 34167 32918 34176
rect 32968 34184 32996 35006
rect 33048 34944 33100 34950
rect 33048 34886 33100 34892
rect 33060 34241 33088 34886
rect 33428 34542 33456 35255
rect 33612 34610 33640 35430
rect 33704 34678 33732 35788
rect 33784 35692 33836 35698
rect 33784 35634 33836 35640
rect 33692 34672 33744 34678
rect 33692 34614 33744 34620
rect 33508 34604 33560 34610
rect 33508 34546 33560 34552
rect 33600 34604 33652 34610
rect 33600 34546 33652 34552
rect 33416 34536 33468 34542
rect 33230 34504 33286 34513
rect 33140 34468 33192 34474
rect 33230 34439 33286 34448
rect 33336 34496 33416 34524
rect 33140 34410 33192 34416
rect 33046 34232 33102 34241
rect 32968 34156 32997 34184
rect 33152 34202 33180 34410
rect 33046 34167 33102 34176
rect 33140 34196 33192 34202
rect 32969 34116 32997 34156
rect 33140 34138 33192 34144
rect 32876 34088 32997 34116
rect 32876 33998 32904 34088
rect 33244 33998 33272 34439
rect 32864 33992 32916 33998
rect 32864 33934 32916 33940
rect 33232 33992 33284 33998
rect 33232 33934 33284 33940
rect 33336 33946 33364 34496
rect 33416 34478 33468 34484
rect 33416 33992 33468 33998
rect 32876 33810 32904 33934
rect 33336 33918 33369 33946
rect 33416 33934 33468 33940
rect 33428 33918 33461 33934
rect 33341 33810 33369 33918
rect 33433 33844 33461 33918
rect 32876 33782 32997 33810
rect 32969 33674 32997 33782
rect 32864 33652 32916 33658
rect 32864 33594 32916 33600
rect 32968 33646 32997 33674
rect 33244 33782 33369 33810
rect 33428 33816 33461 33844
rect 32876 33522 32904 33594
rect 32864 33516 32916 33522
rect 32864 33458 32916 33464
rect 32600 33238 32720 33266
rect 32772 33312 32824 33318
rect 32772 33254 32824 33260
rect 32496 33108 32548 33114
rect 32496 33050 32548 33056
rect 32508 32416 32536 33050
rect 32600 32910 32628 33238
rect 32678 33144 32734 33153
rect 32678 33079 32734 33088
rect 32692 32910 32720 33079
rect 32876 32910 32904 33458
rect 32968 33436 32996 33646
rect 33140 33584 33192 33590
rect 33140 33526 33192 33532
rect 32968 33408 33088 33436
rect 32588 32904 32640 32910
rect 32588 32846 32640 32852
rect 32680 32904 32732 32910
rect 32864 32904 32916 32910
rect 32680 32846 32732 32852
rect 32784 32864 32864 32892
rect 32588 32428 32640 32434
rect 32508 32388 32588 32416
rect 32404 32224 32456 32230
rect 32404 32166 32456 32172
rect 32508 32042 32536 32388
rect 32588 32370 32640 32376
rect 32586 32192 32642 32201
rect 32586 32127 32642 32136
rect 32416 32014 32536 32042
rect 32034 31784 32090 31793
rect 32034 31719 32090 31728
rect 32220 31748 32272 31754
rect 32220 31690 32272 31696
rect 32034 31648 32090 31657
rect 32034 31583 32090 31592
rect 32048 31482 32076 31583
rect 32126 31512 32182 31521
rect 32036 31476 32088 31482
rect 32126 31447 32182 31456
rect 32036 31418 32088 31424
rect 32140 31210 32168 31447
rect 32128 31204 32180 31210
rect 32128 31146 32180 31152
rect 32034 31104 32090 31113
rect 32034 31039 32090 31048
rect 31944 30184 31996 30190
rect 31944 30126 31996 30132
rect 31942 29744 31998 29753
rect 31942 29679 31998 29688
rect 31956 29306 31984 29679
rect 31944 29300 31996 29306
rect 31944 29242 31996 29248
rect 31864 29158 31984 29186
rect 31772 28966 31892 28994
rect 31668 28552 31720 28558
rect 31668 28494 31720 28500
rect 31864 28150 31892 28966
rect 31668 28144 31720 28150
rect 31666 28112 31668 28121
rect 31852 28144 31904 28150
rect 31720 28112 31722 28121
rect 31576 28076 31628 28082
rect 31852 28086 31904 28092
rect 31666 28047 31722 28056
rect 31576 28018 31628 28024
rect 31666 27840 31722 27849
rect 31666 27775 31722 27784
rect 31574 27568 31630 27577
rect 31574 27503 31630 27512
rect 31588 26314 31616 27503
rect 31680 27441 31708 27775
rect 31666 27432 31722 27441
rect 31666 27367 31722 27376
rect 31758 27024 31814 27033
rect 31680 26982 31758 27010
rect 31576 26308 31628 26314
rect 31576 26250 31628 26256
rect 31484 25288 31536 25294
rect 31484 25230 31536 25236
rect 31496 24954 31524 25230
rect 31576 25220 31628 25226
rect 31576 25162 31628 25168
rect 31484 24948 31536 24954
rect 31484 24890 31536 24896
rect 31392 24812 31444 24818
rect 31392 24754 31444 24760
rect 31116 24744 31168 24750
rect 31116 24686 31168 24692
rect 31208 24608 31260 24614
rect 31208 24550 31260 24556
rect 31116 24064 31168 24070
rect 31116 24006 31168 24012
rect 31024 23112 31076 23118
rect 31024 23054 31076 23060
rect 30932 22568 30984 22574
rect 30932 22510 30984 22516
rect 30840 22160 30892 22166
rect 30840 22102 30892 22108
rect 31128 22030 31156 24006
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31116 22024 31168 22030
rect 31116 21966 31168 21972
rect 31036 21690 31064 21966
rect 31128 21865 31156 21966
rect 31114 21856 31170 21865
rect 31114 21791 31170 21800
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 31116 21548 31168 21554
rect 31116 21490 31168 21496
rect 30748 21412 30800 21418
rect 30748 21354 30800 21360
rect 30564 21140 30616 21146
rect 30564 21082 30616 21088
rect 30380 21004 30432 21010
rect 30380 20946 30432 20952
rect 30392 20534 30420 20946
rect 30564 20936 30616 20942
rect 30564 20878 30616 20884
rect 30380 20528 30432 20534
rect 30380 20470 30432 20476
rect 30378 20224 30434 20233
rect 30378 20159 30434 20168
rect 30288 19304 30340 19310
rect 30288 19246 30340 19252
rect 30300 19145 30328 19246
rect 30286 19136 30342 19145
rect 30286 19071 30342 19080
rect 30300 18290 30328 19071
rect 30392 18290 30420 20159
rect 30472 19780 30524 19786
rect 30472 19722 30524 19728
rect 30484 19242 30512 19722
rect 30472 19236 30524 19242
rect 30472 19178 30524 19184
rect 30470 19000 30526 19009
rect 30470 18935 30526 18944
rect 30484 18698 30512 18935
rect 30472 18692 30524 18698
rect 30472 18634 30524 18640
rect 30576 18630 30604 20878
rect 30760 20874 30788 21354
rect 31128 21298 31156 21490
rect 31220 21457 31248 24550
rect 31404 23798 31432 24754
rect 31392 23792 31444 23798
rect 31298 23760 31354 23769
rect 31444 23752 31524 23780
rect 31392 23734 31444 23740
rect 31298 23695 31300 23704
rect 31352 23695 31354 23704
rect 31300 23666 31352 23672
rect 31392 23520 31444 23526
rect 31392 23462 31444 23468
rect 31298 23216 31354 23225
rect 31298 23151 31354 23160
rect 31312 22710 31340 23151
rect 31300 22704 31352 22710
rect 31300 22646 31352 22652
rect 31404 22574 31432 23462
rect 31300 22568 31352 22574
rect 31300 22510 31352 22516
rect 31392 22568 31444 22574
rect 31392 22510 31444 22516
rect 31206 21448 31262 21457
rect 31206 21383 31262 21392
rect 30944 21270 31156 21298
rect 31208 21344 31260 21350
rect 31208 21286 31260 21292
rect 30748 20868 30800 20874
rect 30668 20828 30748 20856
rect 30668 20466 30696 20828
rect 30748 20810 30800 20816
rect 30748 20596 30800 20602
rect 30800 20556 30880 20584
rect 30748 20538 30800 20544
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30748 20392 30800 20398
rect 30748 20334 30800 20340
rect 30760 19174 30788 20334
rect 30852 20262 30880 20556
rect 30840 20256 30892 20262
rect 30840 20198 30892 20204
rect 30852 19378 30880 20198
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 30748 19168 30800 19174
rect 30748 19110 30800 19116
rect 30564 18624 30616 18630
rect 30562 18592 30564 18601
rect 30616 18592 30618 18601
rect 30562 18527 30618 18536
rect 30288 18284 30340 18290
rect 30288 18226 30340 18232
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 30564 18284 30616 18290
rect 30564 18226 30616 18232
rect 30576 17678 30604 18226
rect 30760 18154 30788 19110
rect 30840 18896 30892 18902
rect 30944 18873 30972 21270
rect 31116 20868 31168 20874
rect 31116 20810 31168 20816
rect 31024 19984 31076 19990
rect 31024 19926 31076 19932
rect 31036 19514 31064 19926
rect 31128 19514 31156 20810
rect 31024 19508 31076 19514
rect 31024 19450 31076 19456
rect 31116 19508 31168 19514
rect 31116 19450 31168 19456
rect 31220 19394 31248 21286
rect 31312 20942 31340 22510
rect 31496 22030 31524 23752
rect 31588 23254 31616 25162
rect 31680 24070 31708 26982
rect 31864 26994 31892 28086
rect 31758 26959 31814 26968
rect 31852 26988 31904 26994
rect 31852 26930 31904 26936
rect 31852 26784 31904 26790
rect 31852 26726 31904 26732
rect 31864 26353 31892 26726
rect 31850 26344 31906 26353
rect 31850 26279 31906 26288
rect 31956 26234 31984 29158
rect 31864 26206 31984 26234
rect 31760 25968 31812 25974
rect 31760 25910 31812 25916
rect 31772 24682 31800 25910
rect 31760 24676 31812 24682
rect 31760 24618 31812 24624
rect 31758 24440 31814 24449
rect 31758 24375 31760 24384
rect 31812 24375 31814 24384
rect 31760 24346 31812 24352
rect 31864 24290 31892 26206
rect 31942 25528 31998 25537
rect 31942 25463 31998 25472
rect 31772 24262 31892 24290
rect 31668 24064 31720 24070
rect 31772 24041 31800 24262
rect 31852 24200 31904 24206
rect 31852 24142 31904 24148
rect 31668 24006 31720 24012
rect 31758 24032 31814 24041
rect 31758 23967 31814 23976
rect 31758 23488 31814 23497
rect 31758 23423 31814 23432
rect 31576 23248 31628 23254
rect 31576 23190 31628 23196
rect 31588 23118 31616 23190
rect 31576 23112 31628 23118
rect 31576 23054 31628 23060
rect 31576 22704 31628 22710
rect 31628 22664 31708 22692
rect 31576 22646 31628 22652
rect 31484 22024 31536 22030
rect 31484 21966 31536 21972
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 31300 20936 31352 20942
rect 31300 20878 31352 20884
rect 31300 20800 31352 20806
rect 31404 20788 31432 21490
rect 31496 21010 31524 21966
rect 31576 21888 31628 21894
rect 31576 21830 31628 21836
rect 31588 21350 31616 21830
rect 31576 21344 31628 21350
rect 31576 21286 31628 21292
rect 31484 21004 31536 21010
rect 31484 20946 31536 20952
rect 31352 20760 31432 20788
rect 31300 20742 31352 20748
rect 31312 20058 31340 20742
rect 31392 20392 31444 20398
rect 31392 20334 31444 20340
rect 31300 20052 31352 20058
rect 31300 19994 31352 20000
rect 31300 19712 31352 19718
rect 31300 19654 31352 19660
rect 31024 19372 31076 19378
rect 31024 19314 31076 19320
rect 31128 19366 31248 19394
rect 31036 19174 31064 19314
rect 31024 19168 31076 19174
rect 31024 19110 31076 19116
rect 30840 18838 30892 18844
rect 30930 18864 30986 18873
rect 30852 18578 30880 18838
rect 30930 18799 30986 18808
rect 30852 18550 30972 18578
rect 30840 18420 30892 18426
rect 30840 18362 30892 18368
rect 30852 18154 30880 18362
rect 30748 18148 30800 18154
rect 30748 18090 30800 18096
rect 30840 18148 30892 18154
rect 30840 18090 30892 18096
rect 30654 17912 30710 17921
rect 30654 17847 30710 17856
rect 30564 17672 30616 17678
rect 30562 17640 30564 17649
rect 30616 17640 30618 17649
rect 30562 17575 30618 17584
rect 30564 17536 30616 17542
rect 30564 17478 30616 17484
rect 30286 16552 30342 16561
rect 30286 16487 30342 16496
rect 30300 16454 30328 16487
rect 30288 16448 30340 16454
rect 30194 16416 30250 16425
rect 30288 16390 30340 16396
rect 30194 16351 30250 16360
rect 30102 16280 30158 16289
rect 30102 16215 30158 16224
rect 30116 15162 30144 16215
rect 30380 15904 30432 15910
rect 30380 15846 30432 15852
rect 30392 15434 30420 15846
rect 30380 15428 30432 15434
rect 30380 15370 30432 15376
rect 30104 15156 30156 15162
rect 30104 15098 30156 15104
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 30196 14952 30248 14958
rect 30196 14894 30248 14900
rect 30208 12782 30236 14894
rect 30484 13802 30512 14962
rect 30472 13796 30524 13802
rect 30472 13738 30524 13744
rect 30288 13252 30340 13258
rect 30288 13194 30340 13200
rect 30300 12986 30328 13194
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 30576 12850 30604 17478
rect 30668 17202 30696 17847
rect 30760 17814 30788 18090
rect 30748 17808 30800 17814
rect 30748 17750 30800 17756
rect 30944 17746 30972 18550
rect 30840 17740 30892 17746
rect 30840 17682 30892 17688
rect 30932 17740 30984 17746
rect 30932 17682 30984 17688
rect 30746 17368 30802 17377
rect 30746 17303 30802 17312
rect 30760 17202 30788 17303
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30748 17196 30800 17202
rect 30748 17138 30800 17144
rect 30746 16280 30802 16289
rect 30746 16215 30748 16224
rect 30800 16215 30802 16224
rect 30748 16186 30800 16192
rect 30748 16108 30800 16114
rect 30748 16050 30800 16056
rect 30760 15366 30788 16050
rect 30748 15360 30800 15366
rect 30748 15302 30800 15308
rect 30656 14476 30708 14482
rect 30656 14418 30708 14424
rect 30668 13938 30696 14418
rect 30760 13938 30788 15302
rect 30656 13932 30708 13938
rect 30656 13874 30708 13880
rect 30748 13932 30800 13938
rect 30748 13874 30800 13880
rect 30748 13252 30800 13258
rect 30748 13194 30800 13200
rect 30656 13184 30708 13190
rect 30656 13126 30708 13132
rect 30668 12986 30696 13126
rect 30760 12986 30788 13194
rect 30852 12986 30880 17682
rect 30932 17196 30984 17202
rect 31036 17184 31064 19110
rect 30984 17156 31064 17184
rect 30932 17138 30984 17144
rect 31128 16182 31156 19366
rect 31206 19272 31262 19281
rect 31206 19207 31262 19216
rect 31220 18766 31248 19207
rect 31312 18834 31340 19654
rect 31300 18828 31352 18834
rect 31300 18770 31352 18776
rect 31208 18760 31260 18766
rect 31208 18702 31260 18708
rect 31208 18624 31260 18630
rect 31208 18566 31260 18572
rect 31300 18624 31352 18630
rect 31300 18566 31352 18572
rect 31220 17202 31248 18566
rect 31312 18086 31340 18566
rect 31300 18080 31352 18086
rect 31300 18022 31352 18028
rect 31404 17882 31432 20334
rect 31484 20324 31536 20330
rect 31484 20266 31536 20272
rect 31392 17876 31444 17882
rect 31392 17818 31444 17824
rect 31496 17678 31524 20266
rect 31680 19718 31708 22664
rect 31668 19712 31720 19718
rect 31668 19654 31720 19660
rect 31680 19378 31708 19654
rect 31772 19417 31800 23423
rect 31864 23118 31892 24142
rect 31956 23905 31984 25463
rect 31942 23896 31998 23905
rect 31942 23831 31998 23840
rect 32048 23662 32076 31039
rect 32128 30932 32180 30938
rect 32128 30874 32180 30880
rect 32140 30433 32168 30874
rect 32126 30424 32182 30433
rect 32126 30359 32182 30368
rect 32128 30048 32180 30054
rect 32128 29990 32180 29996
rect 32140 29209 32168 29990
rect 32126 29200 32182 29209
rect 32126 29135 32182 29144
rect 32232 28994 32260 31690
rect 32312 31340 32364 31346
rect 32312 31282 32364 31288
rect 32324 30870 32352 31282
rect 32312 30864 32364 30870
rect 32312 30806 32364 30812
rect 32312 30728 32364 30734
rect 32312 30670 32364 30676
rect 32324 30122 32352 30670
rect 32312 30116 32364 30122
rect 32312 30058 32364 30064
rect 32324 29646 32352 30058
rect 32312 29640 32364 29646
rect 32312 29582 32364 29588
rect 32140 28966 32260 28994
rect 32140 24274 32168 28966
rect 32324 28540 32352 29582
rect 32416 28642 32444 32014
rect 32496 31952 32548 31958
rect 32600 31929 32628 32127
rect 32496 31894 32548 31900
rect 32586 31920 32642 31929
rect 32508 31482 32536 31894
rect 32586 31855 32642 31864
rect 32496 31476 32548 31482
rect 32496 31418 32548 31424
rect 32496 31340 32548 31346
rect 32496 31282 32548 31288
rect 32508 30938 32536 31282
rect 32496 30932 32548 30938
rect 32496 30874 32548 30880
rect 32508 28801 32536 30874
rect 32588 30592 32640 30598
rect 32588 30534 32640 30540
rect 32600 29889 32628 30534
rect 32586 29880 32642 29889
rect 32586 29815 32642 29824
rect 32588 29708 32640 29714
rect 32588 29650 32640 29656
rect 32494 28792 32550 28801
rect 32494 28727 32550 28736
rect 32416 28614 32536 28642
rect 32324 28512 32444 28540
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 32218 27568 32274 27577
rect 32218 27503 32220 27512
rect 32272 27503 32274 27512
rect 32220 27474 32272 27480
rect 32232 27305 32260 27474
rect 32218 27296 32274 27305
rect 32218 27231 32274 27240
rect 32220 26920 32272 26926
rect 32220 26862 32272 26868
rect 32232 25974 32260 26862
rect 32220 25968 32272 25974
rect 32220 25910 32272 25916
rect 32220 25696 32272 25702
rect 32220 25638 32272 25644
rect 32232 25294 32260 25638
rect 32220 25288 32272 25294
rect 32220 25230 32272 25236
rect 32220 24676 32272 24682
rect 32220 24618 32272 24624
rect 32128 24268 32180 24274
rect 32128 24210 32180 24216
rect 32232 24138 32260 24618
rect 32220 24132 32272 24138
rect 32220 24074 32272 24080
rect 32128 24064 32180 24070
rect 32128 24006 32180 24012
rect 32140 23730 32168 24006
rect 32128 23724 32180 23730
rect 32128 23666 32180 23672
rect 32036 23656 32088 23662
rect 32036 23598 32088 23604
rect 32232 23118 32260 24074
rect 32324 23730 32352 28018
rect 32416 27305 32444 28512
rect 32402 27296 32458 27305
rect 32402 27231 32458 27240
rect 32508 26994 32536 28614
rect 32404 26988 32456 26994
rect 32404 26930 32456 26936
rect 32496 26988 32548 26994
rect 32496 26930 32548 26936
rect 32416 26625 32444 26930
rect 32508 26790 32536 26930
rect 32496 26784 32548 26790
rect 32496 26726 32548 26732
rect 32402 26616 32458 26625
rect 32402 26551 32458 26560
rect 32404 26308 32456 26314
rect 32404 26250 32456 26256
rect 32416 25974 32444 26250
rect 32404 25968 32456 25974
rect 32404 25910 32456 25916
rect 32496 25900 32548 25906
rect 32496 25842 32548 25848
rect 32404 25764 32456 25770
rect 32404 25706 32456 25712
rect 32416 25294 32444 25706
rect 32404 25288 32456 25294
rect 32404 25230 32456 25236
rect 32404 24744 32456 24750
rect 32404 24686 32456 24692
rect 32416 24449 32444 24686
rect 32402 24440 32458 24449
rect 32402 24375 32458 24384
rect 32508 24138 32536 25842
rect 32600 24138 32628 29650
rect 32692 29306 32720 32846
rect 32680 29300 32732 29306
rect 32680 29242 32732 29248
rect 32784 29170 32812 32864
rect 32864 32846 32916 32852
rect 33060 32552 33088 33408
rect 33152 32910 33180 33526
rect 33140 32904 33192 32910
rect 33140 32846 33192 32852
rect 32968 32524 33088 32552
rect 32862 32328 32918 32337
rect 32862 32263 32918 32272
rect 32876 31958 32904 32263
rect 32968 32230 32996 32524
rect 33048 32428 33100 32434
rect 33048 32370 33100 32376
rect 32956 32224 33008 32230
rect 32956 32166 33008 32172
rect 32864 31952 32916 31958
rect 32864 31894 32916 31900
rect 32968 31822 32996 32166
rect 32956 31816 33008 31822
rect 32876 31776 32956 31804
rect 32876 31346 32904 31776
rect 32956 31758 33008 31764
rect 32956 31680 33008 31686
rect 32956 31622 33008 31628
rect 32864 31340 32916 31346
rect 32864 31282 32916 31288
rect 32876 30870 32904 31282
rect 32864 30864 32916 30870
rect 32864 30806 32916 30812
rect 32968 30802 32996 31622
rect 32956 30796 33008 30802
rect 32956 30738 33008 30744
rect 32968 30297 32996 30738
rect 32954 30288 33010 30297
rect 32954 30223 33010 30232
rect 32956 30184 33008 30190
rect 32956 30126 33008 30132
rect 32864 30048 32916 30054
rect 32864 29990 32916 29996
rect 32772 29164 32824 29170
rect 32772 29106 32824 29112
rect 32772 28960 32824 28966
rect 32772 28902 32824 28908
rect 32680 28484 32732 28490
rect 32680 28426 32732 28432
rect 32692 25208 32720 28426
rect 32784 28014 32812 28902
rect 32772 28008 32824 28014
rect 32772 27950 32824 27956
rect 32772 27328 32824 27334
rect 32772 27270 32824 27276
rect 32784 25906 32812 27270
rect 32876 26382 32904 29990
rect 32968 28694 32996 30126
rect 33060 29238 33088 32370
rect 33152 31736 33180 32846
rect 33244 32502 33272 33782
rect 33322 33688 33378 33697
rect 33322 33623 33378 33632
rect 33336 33114 33364 33623
rect 33428 33425 33456 33816
rect 33414 33416 33470 33425
rect 33414 33351 33470 33360
rect 33324 33108 33376 33114
rect 33324 33050 33376 33056
rect 33324 32904 33376 32910
rect 33324 32846 33376 32852
rect 33416 32904 33468 32910
rect 33416 32846 33468 32852
rect 33336 32745 33364 32846
rect 33322 32736 33378 32745
rect 33322 32671 33378 32680
rect 33232 32496 33284 32502
rect 33232 32438 33284 32444
rect 33324 32428 33376 32434
rect 33324 32370 33376 32376
rect 33336 31754 33364 32370
rect 33428 31822 33456 32846
rect 33520 32026 33548 34546
rect 33692 34060 33744 34066
rect 33612 34020 33692 34048
rect 33612 33862 33640 34020
rect 33692 34002 33744 34008
rect 33692 33924 33744 33930
rect 33692 33866 33744 33872
rect 33600 33856 33652 33862
rect 33600 33798 33652 33804
rect 33598 33688 33654 33697
rect 33598 33623 33654 33632
rect 33612 33318 33640 33623
rect 33704 33590 33732 33866
rect 33692 33584 33744 33590
rect 33692 33526 33744 33532
rect 33692 33448 33744 33454
rect 33692 33390 33744 33396
rect 33600 33312 33652 33318
rect 33600 33254 33652 33260
rect 33508 32020 33560 32026
rect 33508 31962 33560 31968
rect 33598 31920 33654 31929
rect 33598 31855 33654 31864
rect 33612 31822 33640 31855
rect 33416 31816 33468 31822
rect 33416 31758 33468 31764
rect 33600 31816 33652 31822
rect 33600 31758 33652 31764
rect 33232 31748 33284 31754
rect 33152 31708 33232 31736
rect 33232 31690 33284 31696
rect 33324 31748 33376 31754
rect 33324 31690 33376 31696
rect 33244 31464 33272 31690
rect 33324 31476 33376 31482
rect 33244 31436 33324 31464
rect 33324 31418 33376 31424
rect 33140 31272 33192 31278
rect 33140 31214 33192 31220
rect 33232 31272 33284 31278
rect 33232 31214 33284 31220
rect 33152 30870 33180 31214
rect 33140 30864 33192 30870
rect 33140 30806 33192 30812
rect 33244 30734 33272 31214
rect 33232 30728 33284 30734
rect 33232 30670 33284 30676
rect 33140 30660 33192 30666
rect 33140 30602 33192 30608
rect 33152 30569 33180 30602
rect 33138 30560 33194 30569
rect 33138 30495 33194 30504
rect 33244 30258 33272 30670
rect 33336 30598 33364 31418
rect 33428 31278 33456 31758
rect 33508 31680 33560 31686
rect 33704 31668 33732 33390
rect 33508 31622 33560 31628
rect 33612 31640 33732 31668
rect 33520 31414 33548 31622
rect 33508 31408 33560 31414
rect 33508 31350 33560 31356
rect 33416 31272 33468 31278
rect 33416 31214 33468 31220
rect 33520 31113 33548 31350
rect 33506 31104 33562 31113
rect 33506 31039 33562 31048
rect 33612 30954 33640 31640
rect 33796 30954 33824 35634
rect 33888 35154 33916 36343
rect 33966 35864 34022 35873
rect 33966 35799 34022 35808
rect 33980 35766 34008 35799
rect 33968 35760 34020 35766
rect 33968 35702 34020 35708
rect 34164 35630 34192 36586
rect 34152 35624 34204 35630
rect 34150 35592 34152 35601
rect 34204 35592 34206 35601
rect 34150 35527 34206 35536
rect 34060 35216 34112 35222
rect 34060 35158 34112 35164
rect 33876 35148 33928 35154
rect 33876 35090 33928 35096
rect 33888 34746 33916 35090
rect 33876 34740 33928 34746
rect 33876 34682 33928 34688
rect 33876 34400 33928 34406
rect 33876 34342 33928 34348
rect 33888 33522 33916 34342
rect 34072 34241 34100 35158
rect 34256 35057 34284 36740
rect 34520 36722 34572 36728
rect 34612 36712 34664 36718
rect 34612 36654 34664 36660
rect 34426 36544 34482 36553
rect 34426 36479 34482 36488
rect 34440 36378 34468 36479
rect 34428 36372 34480 36378
rect 34428 36314 34480 36320
rect 34520 35284 34572 35290
rect 34520 35226 34572 35232
rect 34428 35080 34480 35086
rect 34242 35048 34298 35057
rect 34428 35022 34480 35028
rect 34242 34983 34298 34992
rect 34152 34604 34204 34610
rect 34152 34546 34204 34552
rect 34058 34232 34114 34241
rect 34164 34202 34192 34546
rect 34256 34202 34284 34983
rect 34336 34672 34388 34678
rect 34336 34614 34388 34620
rect 34058 34167 34114 34176
rect 34152 34196 34204 34202
rect 34152 34138 34204 34144
rect 34244 34196 34296 34202
rect 34244 34138 34296 34144
rect 34060 33992 34112 33998
rect 34060 33934 34112 33940
rect 33876 33516 33928 33522
rect 33876 33458 33928 33464
rect 34072 33402 34100 33934
rect 34348 33862 34376 34614
rect 34440 34474 34468 35022
rect 34428 34468 34480 34474
rect 34428 34410 34480 34416
rect 34428 34196 34480 34202
rect 34428 34138 34480 34144
rect 34336 33856 34388 33862
rect 34256 33816 34336 33844
rect 34256 33522 34284 33816
rect 34336 33798 34388 33804
rect 34244 33516 34296 33522
rect 34244 33458 34296 33464
rect 34336 33516 34388 33522
rect 34440 33504 34468 34138
rect 34532 34082 34560 35226
rect 34624 34746 34652 36654
rect 34716 35154 34744 37295
rect 34808 35290 34836 37726
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35164 37256 35216 37262
rect 35164 37198 35216 37204
rect 35176 36961 35204 37198
rect 35360 36961 35388 38082
rect 35452 38010 35480 38247
rect 35440 38004 35492 38010
rect 35440 37946 35492 37952
rect 35544 37346 35572 38383
rect 35452 37318 35572 37346
rect 35162 36952 35218 36961
rect 35162 36887 35218 36896
rect 35346 36952 35402 36961
rect 35346 36887 35402 36896
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35348 35488 35400 35494
rect 35348 35430 35400 35436
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34796 35284 34848 35290
rect 34796 35226 34848 35232
rect 34704 35148 34756 35154
rect 34704 35090 34756 35096
rect 35256 35080 35308 35086
rect 35256 35022 35308 35028
rect 34980 34944 35032 34950
rect 34980 34886 35032 34892
rect 35072 34944 35124 34950
rect 35268 34898 35296 35022
rect 35124 34892 35296 34898
rect 35072 34886 35296 34892
rect 34612 34740 34664 34746
rect 34612 34682 34664 34688
rect 34992 34626 35020 34886
rect 35084 34870 35296 34886
rect 34808 34610 35112 34626
rect 34808 34604 35124 34610
rect 34808 34598 35072 34604
rect 34704 34468 34756 34474
rect 34704 34410 34756 34416
rect 34610 34368 34666 34377
rect 34610 34303 34666 34312
rect 34624 34202 34652 34303
rect 34716 34202 34744 34410
rect 34612 34196 34664 34202
rect 34612 34138 34664 34144
rect 34704 34196 34756 34202
rect 34704 34138 34756 34144
rect 34532 34054 34744 34082
rect 34520 33992 34572 33998
rect 34520 33934 34572 33940
rect 34388 33476 34468 33504
rect 34336 33458 34388 33464
rect 33888 33374 34100 33402
rect 33888 32473 33916 33374
rect 34060 33312 34112 33318
rect 34060 33254 34112 33260
rect 34150 33280 34206 33289
rect 34072 32892 34100 33254
rect 34150 33215 34206 33224
rect 34164 33046 34192 33215
rect 34152 33040 34204 33046
rect 34152 32982 34204 32988
rect 34072 32864 34192 32892
rect 33874 32464 33930 32473
rect 33874 32399 33930 32408
rect 33876 32292 33928 32298
rect 33876 32234 33928 32240
rect 33888 31657 33916 32234
rect 34060 31952 34112 31958
rect 34060 31894 34112 31900
rect 33968 31816 34020 31822
rect 33966 31784 33968 31793
rect 34020 31784 34022 31793
rect 33966 31719 34022 31728
rect 33874 31648 33930 31657
rect 33874 31583 33930 31592
rect 34072 31482 34100 31894
rect 34060 31476 34112 31482
rect 34060 31418 34112 31424
rect 34164 31142 34192 32864
rect 34256 31414 34284 33458
rect 34428 33380 34480 33386
rect 34428 33322 34480 33328
rect 34336 32972 34388 32978
rect 34336 32914 34388 32920
rect 34348 32881 34376 32914
rect 34334 32872 34390 32881
rect 34334 32807 34390 32816
rect 34440 32722 34468 33322
rect 34532 33114 34560 33934
rect 34612 33856 34664 33862
rect 34612 33798 34664 33804
rect 34520 33108 34572 33114
rect 34520 33050 34572 33056
rect 34624 33017 34652 33798
rect 34610 33008 34666 33017
rect 34610 32943 34666 32952
rect 34520 32904 34572 32910
rect 34520 32846 34572 32852
rect 34716 32858 34744 34054
rect 34808 33590 34836 34598
rect 35072 34546 35124 34552
rect 35164 34604 35216 34610
rect 35164 34546 35216 34552
rect 35176 34474 35204 34546
rect 35164 34468 35216 34474
rect 35164 34410 35216 34416
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34888 34128 34940 34134
rect 35360 34082 35388 35430
rect 35452 35086 35480 37318
rect 35532 37256 35584 37262
rect 35532 37198 35584 37204
rect 35440 35080 35492 35086
rect 35440 35022 35492 35028
rect 35452 34921 35480 35022
rect 35438 34912 35494 34921
rect 35438 34847 35494 34856
rect 35440 34536 35492 34542
rect 35440 34478 35492 34484
rect 34888 34070 34940 34076
rect 34796 33584 34848 33590
rect 34796 33526 34848 33532
rect 34900 33454 34928 34070
rect 35268 34066 35388 34082
rect 35256 34060 35388 34066
rect 35308 34054 35388 34060
rect 35256 34002 35308 34008
rect 35254 33552 35310 33561
rect 35072 33516 35124 33522
rect 35254 33487 35256 33496
rect 35072 33458 35124 33464
rect 35308 33487 35310 33496
rect 35256 33458 35308 33464
rect 34888 33448 34940 33454
rect 35084 33425 35112 33458
rect 34888 33390 34940 33396
rect 35070 33416 35126 33425
rect 35070 33351 35126 33360
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35072 32904 35124 32910
rect 34978 32872 35034 32881
rect 34348 32694 34468 32722
rect 34244 31408 34296 31414
rect 34244 31350 34296 31356
rect 34152 31136 34204 31142
rect 34152 31078 34204 31084
rect 33428 30926 33640 30954
rect 33704 30926 33824 30954
rect 33324 30592 33376 30598
rect 33324 30534 33376 30540
rect 33232 30252 33284 30258
rect 33232 30194 33284 30200
rect 33140 30048 33192 30054
rect 33140 29990 33192 29996
rect 33152 29782 33180 29990
rect 33140 29776 33192 29782
rect 33140 29718 33192 29724
rect 33048 29232 33100 29238
rect 33048 29174 33100 29180
rect 33060 28762 33088 29174
rect 33048 28756 33100 28762
rect 33048 28698 33100 28704
rect 32956 28688 33008 28694
rect 32956 28630 33008 28636
rect 33152 28540 33180 29718
rect 33244 29510 33272 30194
rect 33336 29782 33364 30534
rect 33324 29776 33376 29782
rect 33324 29718 33376 29724
rect 33232 29504 33284 29510
rect 33232 29446 33284 29452
rect 33232 29300 33284 29306
rect 33232 29242 33284 29248
rect 32968 28512 33180 28540
rect 32968 26586 32996 28512
rect 33046 28112 33102 28121
rect 33046 28047 33102 28056
rect 33060 26761 33088 28047
rect 33140 27396 33192 27402
rect 33140 27338 33192 27344
rect 33046 26752 33102 26761
rect 33046 26687 33102 26696
rect 32956 26580 33008 26586
rect 32956 26522 33008 26528
rect 32864 26376 32916 26382
rect 32864 26318 32916 26324
rect 32864 26240 32916 26246
rect 32968 26217 32996 26522
rect 33048 26308 33100 26314
rect 33048 26250 33100 26256
rect 32864 26182 32916 26188
rect 32954 26208 33010 26217
rect 32876 26042 32904 26182
rect 32954 26143 33010 26152
rect 32864 26036 32916 26042
rect 32864 25978 32916 25984
rect 32956 26036 33008 26042
rect 32956 25978 33008 25984
rect 32772 25900 32824 25906
rect 32772 25842 32824 25848
rect 32784 25378 32812 25842
rect 32784 25350 32904 25378
rect 32968 25362 32996 25978
rect 33060 25974 33088 26250
rect 33048 25968 33100 25974
rect 33048 25910 33100 25916
rect 33152 25786 33180 27338
rect 33244 26081 33272 29242
rect 33322 28792 33378 28801
rect 33322 28727 33378 28736
rect 33336 27946 33364 28727
rect 33324 27940 33376 27946
rect 33324 27882 33376 27888
rect 33428 27470 33456 30926
rect 33508 30592 33560 30598
rect 33508 30534 33560 30540
rect 33600 30592 33652 30598
rect 33600 30534 33652 30540
rect 33520 30258 33548 30534
rect 33508 30252 33560 30258
rect 33508 30194 33560 30200
rect 33508 30116 33560 30122
rect 33508 30058 33560 30064
rect 33520 29345 33548 30058
rect 33612 30002 33640 30534
rect 33704 30297 33732 30926
rect 33968 30796 34020 30802
rect 33968 30738 34020 30744
rect 33784 30660 33836 30666
rect 33784 30602 33836 30608
rect 33690 30288 33746 30297
rect 33690 30223 33746 30232
rect 33692 30116 33744 30122
rect 33692 30058 33744 30064
rect 33612 29974 33641 30002
rect 33613 29764 33641 29974
rect 33612 29736 33641 29764
rect 33506 29336 33562 29345
rect 33506 29271 33562 29280
rect 33508 29232 33560 29238
rect 33508 29174 33560 29180
rect 33520 28762 33548 29174
rect 33508 28756 33560 28762
rect 33508 28698 33560 28704
rect 33508 27872 33560 27878
rect 33508 27814 33560 27820
rect 33416 27464 33468 27470
rect 33416 27406 33468 27412
rect 33324 27328 33376 27334
rect 33324 27270 33376 27276
rect 33230 26072 33286 26081
rect 33230 26007 33286 26016
rect 33060 25758 33180 25786
rect 32876 25294 32904 25350
rect 32956 25356 33008 25362
rect 32956 25298 33008 25304
rect 32864 25288 32916 25294
rect 32864 25230 32916 25236
rect 32692 25180 32812 25208
rect 32678 25120 32734 25129
rect 32678 25055 32734 25064
rect 32692 24410 32720 25055
rect 32680 24404 32732 24410
rect 32680 24346 32732 24352
rect 32496 24132 32548 24138
rect 32496 24074 32548 24080
rect 32588 24132 32640 24138
rect 32588 24074 32640 24080
rect 32784 23848 32812 25180
rect 32862 24984 32918 24993
rect 32862 24919 32918 24928
rect 32876 24886 32904 24919
rect 32864 24880 32916 24886
rect 32864 24822 32916 24828
rect 32876 24177 32904 24822
rect 32956 24744 33008 24750
rect 32956 24686 33008 24692
rect 32968 24585 32996 24686
rect 32954 24576 33010 24585
rect 32954 24511 33010 24520
rect 32862 24168 32918 24177
rect 32862 24103 32918 24112
rect 32864 24064 32916 24070
rect 32862 24032 32864 24041
rect 32916 24032 32918 24041
rect 32862 23967 32918 23976
rect 32416 23820 32812 23848
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32416 23610 32444 23820
rect 32968 23798 32996 24511
rect 32956 23792 33008 23798
rect 32494 23760 32550 23769
rect 32956 23734 33008 23740
rect 32494 23695 32550 23704
rect 32588 23724 32640 23730
rect 32324 23582 32444 23610
rect 31852 23112 31904 23118
rect 31852 23054 31904 23060
rect 32220 23112 32272 23118
rect 32220 23054 32272 23060
rect 32220 22432 32272 22438
rect 32220 22374 32272 22380
rect 32036 21888 32088 21894
rect 32036 21830 32088 21836
rect 32128 21888 32180 21894
rect 32128 21830 32180 21836
rect 32048 21010 32076 21830
rect 32140 21622 32168 21830
rect 32128 21616 32180 21622
rect 32128 21558 32180 21564
rect 32232 21298 32260 22374
rect 32324 22030 32352 23582
rect 32508 23168 32536 23695
rect 32588 23666 32640 23672
rect 32772 23724 32824 23730
rect 32772 23666 32824 23672
rect 32416 23140 32536 23168
rect 32416 23050 32444 23140
rect 32494 23080 32550 23089
rect 32404 23044 32456 23050
rect 32494 23015 32550 23024
rect 32404 22986 32456 22992
rect 32402 22944 32458 22953
rect 32402 22879 32458 22888
rect 32416 22545 32444 22879
rect 32508 22681 32536 23015
rect 32494 22672 32550 22681
rect 32494 22607 32550 22616
rect 32402 22536 32458 22545
rect 32402 22471 32458 22480
rect 32496 22160 32548 22166
rect 32496 22102 32548 22108
rect 32312 22024 32364 22030
rect 32312 21966 32364 21972
rect 32310 21856 32366 21865
rect 32310 21791 32366 21800
rect 32324 21554 32352 21791
rect 32508 21622 32536 22102
rect 32496 21616 32548 21622
rect 32496 21558 32548 21564
rect 32312 21548 32364 21554
rect 32364 21508 32444 21536
rect 32312 21490 32364 21496
rect 32140 21270 32260 21298
rect 32312 21344 32364 21350
rect 32312 21286 32364 21292
rect 32036 21004 32088 21010
rect 32036 20946 32088 20952
rect 31944 20800 31996 20806
rect 31944 20742 31996 20748
rect 31850 20496 31906 20505
rect 31850 20431 31906 20440
rect 31864 20398 31892 20431
rect 31852 20392 31904 20398
rect 31852 20334 31904 20340
rect 31852 20256 31904 20262
rect 31852 20198 31904 20204
rect 31758 19408 31814 19417
rect 31668 19372 31720 19378
rect 31758 19343 31814 19352
rect 31668 19314 31720 19320
rect 31760 19236 31812 19242
rect 31760 19178 31812 19184
rect 31668 19168 31720 19174
rect 31668 19110 31720 19116
rect 31576 18896 31628 18902
rect 31574 18864 31576 18873
rect 31628 18864 31630 18873
rect 31574 18799 31630 18808
rect 31680 18766 31708 19110
rect 31668 18760 31720 18766
rect 31668 18702 31720 18708
rect 31772 18290 31800 19178
rect 31760 18284 31812 18290
rect 31760 18226 31812 18232
rect 31576 18216 31628 18222
rect 31576 18158 31628 18164
rect 31392 17672 31444 17678
rect 31392 17614 31444 17620
rect 31484 17672 31536 17678
rect 31484 17614 31536 17620
rect 31300 17604 31352 17610
rect 31300 17546 31352 17552
rect 31312 17270 31340 17546
rect 31300 17264 31352 17270
rect 31300 17206 31352 17212
rect 31208 17196 31260 17202
rect 31208 17138 31260 17144
rect 31116 16176 31168 16182
rect 31116 16118 31168 16124
rect 31116 16040 31168 16046
rect 31116 15982 31168 15988
rect 31024 14408 31076 14414
rect 31024 14350 31076 14356
rect 30932 14340 30984 14346
rect 30932 14282 30984 14288
rect 30656 12980 30708 12986
rect 30656 12922 30708 12928
rect 30748 12980 30800 12986
rect 30748 12922 30800 12928
rect 30840 12980 30892 12986
rect 30840 12922 30892 12928
rect 30564 12844 30616 12850
rect 30564 12786 30616 12792
rect 30196 12776 30248 12782
rect 30196 12718 30248 12724
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 30208 11694 30236 12718
rect 30668 12238 30696 12922
rect 30944 12238 30972 14282
rect 31036 13938 31064 14350
rect 31024 13932 31076 13938
rect 31024 13874 31076 13880
rect 31036 12238 31064 13874
rect 31128 12782 31156 15982
rect 31404 15502 31432 17614
rect 31496 16998 31524 17614
rect 31484 16992 31536 16998
rect 31484 16934 31536 16940
rect 31496 15570 31524 16934
rect 31588 16794 31616 18158
rect 31668 17740 31720 17746
rect 31668 17682 31720 17688
rect 31680 17134 31708 17682
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 31668 16992 31720 16998
rect 31668 16934 31720 16940
rect 31576 16788 31628 16794
rect 31576 16730 31628 16736
rect 31680 16590 31708 16934
rect 31668 16584 31720 16590
rect 31668 16526 31720 16532
rect 31772 16250 31800 18226
rect 31864 17202 31892 20198
rect 31956 19553 31984 20742
rect 32036 20052 32088 20058
rect 32036 19994 32088 20000
rect 32048 19786 32076 19994
rect 32036 19780 32088 19786
rect 32036 19722 32088 19728
rect 31942 19544 31998 19553
rect 31942 19479 31998 19488
rect 31944 17876 31996 17882
rect 31944 17818 31996 17824
rect 31852 17196 31904 17202
rect 31852 17138 31904 17144
rect 31852 17060 31904 17066
rect 31852 17002 31904 17008
rect 31760 16244 31812 16250
rect 31760 16186 31812 16192
rect 31484 15564 31536 15570
rect 31484 15506 31536 15512
rect 31392 15496 31444 15502
rect 31392 15438 31444 15444
rect 31484 14952 31536 14958
rect 31484 14894 31536 14900
rect 31668 14952 31720 14958
rect 31668 14894 31720 14900
rect 31496 13462 31524 14894
rect 31576 14816 31628 14822
rect 31576 14758 31628 14764
rect 31588 13938 31616 14758
rect 31680 14056 31708 14894
rect 31680 14028 31800 14056
rect 31576 13932 31628 13938
rect 31576 13874 31628 13880
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 31484 13456 31536 13462
rect 31484 13398 31536 13404
rect 31116 12776 31168 12782
rect 31116 12718 31168 12724
rect 31128 12434 31156 12718
rect 31128 12406 31340 12434
rect 30656 12232 30708 12238
rect 30656 12174 30708 12180
rect 30932 12232 30984 12238
rect 30932 12174 30984 12180
rect 31024 12232 31076 12238
rect 31024 12174 31076 12180
rect 30472 12164 30524 12170
rect 30472 12106 30524 12112
rect 30380 11756 30432 11762
rect 30380 11698 30432 11704
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 30392 11354 30420 11698
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 29828 11212 29880 11218
rect 29828 11154 29880 11160
rect 29840 10674 29868 11154
rect 30288 10804 30340 10810
rect 30288 10746 30340 10752
rect 29828 10668 29880 10674
rect 29828 10610 29880 10616
rect 30196 10668 30248 10674
rect 30196 10610 30248 10616
rect 30208 10266 30236 10610
rect 30196 10260 30248 10266
rect 30196 10202 30248 10208
rect 30300 10198 30328 10746
rect 30392 10266 30420 11290
rect 30484 11082 30512 12106
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 30656 11552 30708 11558
rect 30656 11494 30708 11500
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 30668 11082 30696 11494
rect 30472 11076 30524 11082
rect 30472 11018 30524 11024
rect 30656 11076 30708 11082
rect 30656 11018 30708 11024
rect 30484 10282 30512 11018
rect 30380 10260 30432 10266
rect 30484 10254 30788 10282
rect 30380 10202 30432 10208
rect 30288 10192 30340 10198
rect 30288 10134 30340 10140
rect 30484 10130 30696 10146
rect 30472 10124 30708 10130
rect 30524 10118 30656 10124
rect 30472 10066 30524 10072
rect 30656 10066 30708 10072
rect 29736 9920 29788 9926
rect 29736 9862 29788 9868
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 29460 9648 29512 9654
rect 29460 9590 29512 9596
rect 29748 9586 29776 9862
rect 30668 9722 30696 9862
rect 30656 9716 30708 9722
rect 30656 9658 30708 9664
rect 29736 9580 29788 9586
rect 29736 9522 29788 9528
rect 30760 9518 30788 10254
rect 30852 9654 30880 11494
rect 31036 11354 31064 11698
rect 31312 11694 31340 12406
rect 31680 12374 31708 13874
rect 31668 12368 31720 12374
rect 31668 12310 31720 12316
rect 31772 12306 31800 14028
rect 31760 12300 31812 12306
rect 31760 12242 31812 12248
rect 31392 12164 31444 12170
rect 31392 12106 31444 12112
rect 31300 11688 31352 11694
rect 31300 11630 31352 11636
rect 31024 11348 31076 11354
rect 31024 11290 31076 11296
rect 30840 9648 30892 9654
rect 30840 9590 30892 9596
rect 31036 9586 31064 11290
rect 31312 10130 31340 11630
rect 31404 11558 31432 12106
rect 31760 12096 31812 12102
rect 31760 12038 31812 12044
rect 31772 11898 31800 12038
rect 31864 11898 31892 17002
rect 31956 15638 31984 17818
rect 32036 17672 32088 17678
rect 32036 17614 32088 17620
rect 31944 15632 31996 15638
rect 31944 15574 31996 15580
rect 32048 15484 32076 17614
rect 32140 16454 32168 21270
rect 32218 21176 32274 21185
rect 32218 21111 32274 21120
rect 32232 20942 32260 21111
rect 32324 20942 32352 21286
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 32312 20936 32364 20942
rect 32312 20878 32364 20884
rect 32310 20768 32366 20777
rect 32310 20703 32366 20712
rect 32218 19680 32274 19689
rect 32218 19615 32274 19624
rect 32232 19242 32260 19615
rect 32220 19236 32272 19242
rect 32220 19178 32272 19184
rect 32220 18964 32272 18970
rect 32220 18906 32272 18912
rect 32232 18426 32260 18906
rect 32324 18698 32352 20703
rect 32416 20330 32444 21508
rect 32600 21418 32628 23666
rect 32784 23474 32812 23666
rect 32862 23624 32918 23633
rect 32862 23559 32864 23568
rect 32916 23559 32918 23568
rect 32864 23530 32916 23536
rect 32692 23446 32812 23474
rect 32692 22710 32720 23446
rect 32772 23316 32824 23322
rect 32772 23258 32824 23264
rect 32784 23118 32812 23258
rect 32772 23112 32824 23118
rect 32772 23054 32824 23060
rect 32862 23080 32918 23089
rect 32680 22704 32732 22710
rect 32680 22646 32732 22652
rect 32784 22642 32812 23054
rect 32862 23015 32918 23024
rect 32772 22636 32824 22642
rect 32772 22578 32824 22584
rect 32784 22030 32812 22578
rect 32680 22024 32732 22030
rect 32680 21966 32732 21972
rect 32772 22024 32824 22030
rect 32772 21966 32824 21972
rect 32692 21554 32720 21966
rect 32772 21888 32824 21894
rect 32772 21830 32824 21836
rect 32784 21554 32812 21830
rect 32680 21548 32732 21554
rect 32680 21490 32732 21496
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 32588 21412 32640 21418
rect 32588 21354 32640 21360
rect 32588 20936 32640 20942
rect 32588 20878 32640 20884
rect 32404 20324 32456 20330
rect 32404 20266 32456 20272
rect 32416 19718 32444 20266
rect 32494 19952 32550 19961
rect 32494 19887 32550 19896
rect 32404 19712 32456 19718
rect 32404 19654 32456 19660
rect 32508 19417 32536 19887
rect 32494 19408 32550 19417
rect 32494 19343 32550 19352
rect 32508 19242 32536 19343
rect 32496 19236 32548 19242
rect 32496 19178 32548 19184
rect 32404 18760 32456 18766
rect 32600 18737 32628 20878
rect 32680 20868 32732 20874
rect 32680 20810 32732 20816
rect 32692 20466 32720 20810
rect 32876 20482 32904 23015
rect 32968 22982 32996 23734
rect 32956 22976 33008 22982
rect 32956 22918 33008 22924
rect 32968 22166 32996 22918
rect 32956 22160 33008 22166
rect 32956 22102 33008 22108
rect 32956 20800 33008 20806
rect 32954 20768 32956 20777
rect 33008 20768 33010 20777
rect 32954 20703 33010 20712
rect 32680 20460 32732 20466
rect 32680 20402 32732 20408
rect 32784 20454 32904 20482
rect 32954 20496 33010 20505
rect 32784 20369 32812 20454
rect 32954 20431 33010 20440
rect 32968 20398 32996 20431
rect 32956 20392 33008 20398
rect 32770 20360 32826 20369
rect 32956 20334 33008 20340
rect 32770 20295 32826 20304
rect 32864 20324 32916 20330
rect 32864 20266 32916 20272
rect 32770 19680 32826 19689
rect 32770 19615 32826 19624
rect 32404 18702 32456 18708
rect 32586 18728 32642 18737
rect 32312 18692 32364 18698
rect 32312 18634 32364 18640
rect 32220 18420 32272 18426
rect 32220 18362 32272 18368
rect 32218 18320 32274 18329
rect 32218 18255 32274 18264
rect 32232 18222 32260 18255
rect 32220 18216 32272 18222
rect 32220 18158 32272 18164
rect 32220 17672 32272 17678
rect 32324 17660 32352 18634
rect 32416 18358 32444 18702
rect 32586 18663 32642 18672
rect 32496 18624 32548 18630
rect 32588 18624 32640 18630
rect 32496 18566 32548 18572
rect 32586 18592 32588 18601
rect 32640 18592 32642 18601
rect 32404 18352 32456 18358
rect 32404 18294 32456 18300
rect 32508 18306 32536 18566
rect 32586 18527 32642 18536
rect 32678 18456 32734 18465
rect 32678 18391 32734 18400
rect 32272 17632 32352 17660
rect 32220 17614 32272 17620
rect 32312 17196 32364 17202
rect 32312 17138 32364 17144
rect 32128 16448 32180 16454
rect 32128 16390 32180 16396
rect 31956 15456 32076 15484
rect 31956 12238 31984 15456
rect 32220 15428 32272 15434
rect 32220 15370 32272 15376
rect 32232 15162 32260 15370
rect 32220 15156 32272 15162
rect 32220 15098 32272 15104
rect 32324 14618 32352 17138
rect 32416 16114 32444 18294
rect 32508 18278 32628 18306
rect 32600 18222 32628 18278
rect 32496 18216 32548 18222
rect 32496 18158 32548 18164
rect 32588 18216 32640 18222
rect 32588 18158 32640 18164
rect 32508 17882 32536 18158
rect 32496 17876 32548 17882
rect 32496 17818 32548 17824
rect 32588 17808 32640 17814
rect 32588 17750 32640 17756
rect 32600 17134 32628 17750
rect 32692 17270 32720 18391
rect 32680 17264 32732 17270
rect 32680 17206 32732 17212
rect 32588 17128 32640 17134
rect 32588 17070 32640 17076
rect 32600 16726 32628 17070
rect 32588 16720 32640 16726
rect 32588 16662 32640 16668
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 32680 16108 32732 16114
rect 32680 16050 32732 16056
rect 32588 16040 32640 16046
rect 32588 15982 32640 15988
rect 32496 15020 32548 15026
rect 32496 14962 32548 14968
rect 32312 14612 32364 14618
rect 32312 14554 32364 14560
rect 32036 14340 32088 14346
rect 32036 14282 32088 14288
rect 32048 13530 32076 14282
rect 32508 14278 32536 14962
rect 32496 14272 32548 14278
rect 32496 14214 32548 14220
rect 32036 13524 32088 13530
rect 32036 13466 32088 13472
rect 32496 13388 32548 13394
rect 32496 13330 32548 13336
rect 32128 13320 32180 13326
rect 32128 13262 32180 13268
rect 32140 12918 32168 13262
rect 32128 12912 32180 12918
rect 32128 12854 32180 12860
rect 32312 12844 32364 12850
rect 32312 12786 32364 12792
rect 32324 12442 32352 12786
rect 32312 12436 32364 12442
rect 32312 12378 32364 12384
rect 31944 12232 31996 12238
rect 31944 12174 31996 12180
rect 32312 12096 32364 12102
rect 32312 12038 32364 12044
rect 31760 11892 31812 11898
rect 31760 11834 31812 11840
rect 31852 11892 31904 11898
rect 31852 11834 31904 11840
rect 32324 11762 32352 12038
rect 32508 11830 32536 13330
rect 32496 11824 32548 11830
rect 32496 11766 32548 11772
rect 32312 11756 32364 11762
rect 32312 11698 32364 11704
rect 31392 11552 31444 11558
rect 31392 11494 31444 11500
rect 32404 11552 32456 11558
rect 32404 11494 32456 11500
rect 32496 11552 32548 11558
rect 32496 11494 32548 11500
rect 32416 11082 32444 11494
rect 32508 11354 32536 11494
rect 32496 11348 32548 11354
rect 32496 11290 32548 11296
rect 32404 11076 32456 11082
rect 32404 11018 32456 11024
rect 32404 10668 32456 10674
rect 32404 10610 32456 10616
rect 32416 10266 32444 10610
rect 32404 10260 32456 10266
rect 32404 10202 32456 10208
rect 31300 10124 31352 10130
rect 31300 10066 31352 10072
rect 31760 9920 31812 9926
rect 31760 9862 31812 9868
rect 31772 9586 31800 9862
rect 31024 9580 31076 9586
rect 31024 9522 31076 9528
rect 31760 9580 31812 9586
rect 31760 9522 31812 9528
rect 29184 9512 29236 9518
rect 29184 9454 29236 9460
rect 30748 9512 30800 9518
rect 30748 9454 30800 9460
rect 29000 9376 29052 9382
rect 29000 9318 29052 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 32600 9042 32628 15982
rect 32692 12374 32720 16050
rect 32784 14074 32812 19615
rect 32876 19514 32904 20266
rect 32956 20256 33008 20262
rect 32956 20198 33008 20204
rect 32864 19508 32916 19514
rect 32864 19450 32916 19456
rect 32864 19372 32916 19378
rect 32864 19314 32916 19320
rect 32876 18970 32904 19314
rect 32864 18964 32916 18970
rect 32864 18906 32916 18912
rect 32876 18766 32904 18906
rect 32864 18760 32916 18766
rect 32864 18702 32916 18708
rect 32864 18216 32916 18222
rect 32864 18158 32916 18164
rect 32876 17678 32904 18158
rect 32968 17746 32996 20198
rect 33060 19922 33088 25758
rect 33232 25288 33284 25294
rect 33232 25230 33284 25236
rect 33140 25152 33192 25158
rect 33140 25094 33192 25100
rect 33152 24886 33180 25094
rect 33140 24880 33192 24886
rect 33140 24822 33192 24828
rect 33140 24744 33192 24750
rect 33140 24686 33192 24692
rect 33152 23338 33180 24686
rect 33244 24410 33272 25230
rect 33232 24404 33284 24410
rect 33232 24346 33284 24352
rect 33244 23526 33272 24346
rect 33232 23520 33284 23526
rect 33232 23462 33284 23468
rect 33152 23310 33272 23338
rect 33244 23089 33272 23310
rect 33230 23080 33286 23089
rect 33140 23044 33192 23050
rect 33230 23015 33286 23024
rect 33140 22986 33192 22992
rect 33152 22953 33180 22986
rect 33232 22976 33284 22982
rect 33138 22944 33194 22953
rect 33232 22918 33284 22924
rect 33138 22879 33194 22888
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 33152 22234 33180 22578
rect 33140 22228 33192 22234
rect 33140 22170 33192 22176
rect 33244 22094 33272 22918
rect 33336 22438 33364 27270
rect 33520 27169 33548 27814
rect 33506 27160 33562 27169
rect 33506 27095 33562 27104
rect 33416 26988 33468 26994
rect 33416 26930 33468 26936
rect 33428 25430 33456 26930
rect 33612 26450 33640 29736
rect 33704 29714 33732 30058
rect 33692 29708 33744 29714
rect 33692 29650 33744 29656
rect 33692 29504 33744 29510
rect 33692 29446 33744 29452
rect 33704 29170 33732 29446
rect 33692 29164 33744 29170
rect 33692 29106 33744 29112
rect 33690 29064 33746 29073
rect 33690 28999 33692 29008
rect 33744 28999 33746 29008
rect 33692 28970 33744 28976
rect 33704 28694 33732 28970
rect 33692 28688 33744 28694
rect 33692 28630 33744 28636
rect 33692 28552 33744 28558
rect 33692 28494 33744 28500
rect 33704 28422 33732 28494
rect 33692 28416 33744 28422
rect 33692 28358 33744 28364
rect 33692 27464 33744 27470
rect 33692 27406 33744 27412
rect 33600 26444 33652 26450
rect 33600 26386 33652 26392
rect 33508 26376 33560 26382
rect 33508 26318 33560 26324
rect 33520 25498 33548 26318
rect 33508 25492 33560 25498
rect 33508 25434 33560 25440
rect 33416 25424 33468 25430
rect 33416 25366 33468 25372
rect 33520 24886 33548 25434
rect 33600 25220 33652 25226
rect 33600 25162 33652 25168
rect 33612 25129 33640 25162
rect 33598 25120 33654 25129
rect 33598 25055 33654 25064
rect 33508 24880 33560 24886
rect 33508 24822 33560 24828
rect 33416 24608 33468 24614
rect 33416 24550 33468 24556
rect 33428 24138 33456 24550
rect 33520 24449 33548 24822
rect 33506 24440 33562 24449
rect 33506 24375 33562 24384
rect 33520 24206 33548 24375
rect 33612 24342 33640 25055
rect 33600 24336 33652 24342
rect 33600 24278 33652 24284
rect 33508 24200 33560 24206
rect 33508 24142 33560 24148
rect 33598 24168 33654 24177
rect 33416 24132 33468 24138
rect 33598 24103 33654 24112
rect 33416 24074 33468 24080
rect 33506 24032 33562 24041
rect 33506 23967 33562 23976
rect 33416 23860 33468 23866
rect 33416 23802 33468 23808
rect 33428 23118 33456 23802
rect 33520 23662 33548 23967
rect 33612 23798 33640 24103
rect 33600 23792 33652 23798
rect 33600 23734 33652 23740
rect 33508 23656 33560 23662
rect 33508 23598 33560 23604
rect 33600 23656 33652 23662
rect 33600 23598 33652 23604
rect 33416 23112 33468 23118
rect 33416 23054 33468 23060
rect 33324 22432 33376 22438
rect 33324 22374 33376 22380
rect 33428 22166 33456 23054
rect 33508 22976 33560 22982
rect 33508 22918 33560 22924
rect 33416 22160 33468 22166
rect 33416 22102 33468 22108
rect 33152 22066 33272 22094
rect 33152 20466 33180 22066
rect 33232 22024 33284 22030
rect 33232 21966 33284 21972
rect 33416 22024 33468 22030
rect 33416 21966 33468 21972
rect 33244 20942 33272 21966
rect 33324 21684 33376 21690
rect 33324 21626 33376 21632
rect 33336 21078 33364 21626
rect 33324 21072 33376 21078
rect 33324 21014 33376 21020
rect 33232 20936 33284 20942
rect 33232 20878 33284 20884
rect 33324 20936 33376 20942
rect 33324 20878 33376 20884
rect 33244 20641 33272 20878
rect 33230 20632 33286 20641
rect 33336 20602 33364 20878
rect 33230 20567 33286 20576
rect 33324 20596 33376 20602
rect 33324 20538 33376 20544
rect 33140 20460 33192 20466
rect 33140 20402 33192 20408
rect 33324 20460 33376 20466
rect 33324 20402 33376 20408
rect 33232 20392 33284 20398
rect 33232 20334 33284 20340
rect 33140 20256 33192 20262
rect 33140 20198 33192 20204
rect 33048 19916 33100 19922
rect 33048 19858 33100 19864
rect 33048 19304 33100 19310
rect 33048 19246 33100 19252
rect 33060 19145 33088 19246
rect 33046 19136 33102 19145
rect 33046 19071 33102 19080
rect 32956 17740 33008 17746
rect 32956 17682 33008 17688
rect 32864 17672 32916 17678
rect 32864 17614 32916 17620
rect 33060 17354 33088 19071
rect 33152 18970 33180 20198
rect 33244 20058 33272 20334
rect 33232 20052 33284 20058
rect 33232 19994 33284 20000
rect 33230 19952 33286 19961
rect 33230 19887 33286 19896
rect 33244 19854 33272 19887
rect 33232 19848 33284 19854
rect 33232 19790 33284 19796
rect 33230 19544 33286 19553
rect 33336 19514 33364 20402
rect 33428 20262 33456 21966
rect 33520 21350 33548 22918
rect 33612 22574 33640 23598
rect 33704 23361 33732 27406
rect 33796 27112 33824 30602
rect 33876 30252 33928 30258
rect 33876 30194 33928 30200
rect 33888 30025 33916 30194
rect 33874 30016 33930 30025
rect 33874 29951 33930 29960
rect 33876 29640 33928 29646
rect 33876 29582 33928 29588
rect 33888 29306 33916 29582
rect 33876 29300 33928 29306
rect 33876 29242 33928 29248
rect 33980 29050 34008 30738
rect 34060 30592 34112 30598
rect 34060 30534 34112 30540
rect 34072 29481 34100 30534
rect 34256 30326 34284 31350
rect 34244 30320 34296 30326
rect 34244 30262 34296 30268
rect 34152 30252 34204 30258
rect 34152 30194 34204 30200
rect 34058 29472 34114 29481
rect 34058 29407 34114 29416
rect 34072 29238 34100 29407
rect 34060 29232 34112 29238
rect 34060 29174 34112 29180
rect 34164 29170 34192 30194
rect 34256 29306 34284 30262
rect 34244 29300 34296 29306
rect 34244 29242 34296 29248
rect 34242 29200 34298 29209
rect 34152 29164 34204 29170
rect 34242 29135 34298 29144
rect 34152 29106 34204 29112
rect 33980 29022 34100 29050
rect 34072 28994 34100 29022
rect 33980 28966 34100 28994
rect 33876 28756 33928 28762
rect 33876 28698 33928 28704
rect 33888 28082 33916 28698
rect 33876 28076 33928 28082
rect 33876 28018 33928 28024
rect 33980 27282 34008 28966
rect 34164 28914 34192 29106
rect 34256 29102 34284 29135
rect 34244 29096 34296 29102
rect 34244 29038 34296 29044
rect 34072 28886 34192 28914
rect 34072 28472 34100 28886
rect 34348 28778 34376 32694
rect 34428 32496 34480 32502
rect 34428 32438 34480 32444
rect 34440 31686 34468 32438
rect 34532 32065 34560 32846
rect 34716 32830 34928 32858
rect 34704 32768 34756 32774
rect 34704 32710 34756 32716
rect 34612 32428 34664 32434
rect 34612 32370 34664 32376
rect 34518 32056 34574 32065
rect 34624 32042 34652 32370
rect 34716 32201 34744 32710
rect 34900 32434 34928 32830
rect 35072 32846 35124 32852
rect 34978 32807 35034 32816
rect 34888 32428 34940 32434
rect 34888 32370 34940 32376
rect 34796 32360 34848 32366
rect 34900 32337 34928 32370
rect 34796 32302 34848 32308
rect 34886 32328 34942 32337
rect 34702 32192 34758 32201
rect 34702 32127 34758 32136
rect 34624 32026 34744 32042
rect 34518 31991 34574 32000
rect 34612 32020 34744 32026
rect 34664 32014 34744 32020
rect 34612 31962 34664 31968
rect 34518 31784 34574 31793
rect 34716 31754 34744 32014
rect 34518 31719 34520 31728
rect 34572 31719 34574 31728
rect 34704 31748 34756 31754
rect 34520 31690 34572 31696
rect 34704 31690 34756 31696
rect 34428 31680 34480 31686
rect 34612 31680 34664 31686
rect 34428 31622 34480 31628
rect 34610 31648 34612 31657
rect 34664 31648 34666 31657
rect 34610 31583 34666 31592
rect 34808 31498 34836 32302
rect 34886 32263 34942 32272
rect 34992 32230 35020 32807
rect 35084 32609 35112 32846
rect 35360 32774 35388 34054
rect 35348 32768 35400 32774
rect 35348 32710 35400 32716
rect 35070 32600 35126 32609
rect 35070 32535 35126 32544
rect 34980 32224 35032 32230
rect 34980 32166 35032 32172
rect 35348 32224 35400 32230
rect 35348 32166 35400 32172
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35162 31920 35218 31929
rect 35162 31855 35218 31864
rect 35176 31822 35204 31855
rect 35164 31816 35216 31822
rect 34978 31784 35034 31793
rect 34888 31748 34940 31754
rect 34940 31728 34978 31736
rect 35164 31758 35216 31764
rect 34940 31719 35034 31728
rect 34940 31708 35020 31719
rect 34888 31690 34940 31696
rect 35256 31680 35308 31686
rect 35256 31622 35308 31628
rect 34520 31476 34572 31482
rect 34520 31418 34572 31424
rect 34624 31470 34836 31498
rect 34428 31340 34480 31346
rect 34428 31282 34480 31288
rect 34440 31142 34468 31282
rect 34428 31136 34480 31142
rect 34428 31078 34480 31084
rect 34440 30258 34468 31078
rect 34428 30252 34480 30258
rect 34428 30194 34480 30200
rect 34532 29850 34560 31418
rect 34624 30394 34652 31470
rect 34704 31408 34756 31414
rect 34704 31350 34756 31356
rect 34794 31376 34850 31385
rect 34612 30388 34664 30394
rect 34612 30330 34664 30336
rect 34610 30288 34666 30297
rect 34610 30223 34666 30232
rect 34520 29844 34572 29850
rect 34520 29786 34572 29792
rect 34624 29782 34652 30223
rect 34716 30025 34744 31350
rect 35268 31346 35296 31622
rect 34794 31311 34796 31320
rect 34848 31311 34850 31320
rect 35256 31340 35308 31346
rect 34796 31282 34848 31288
rect 35256 31282 35308 31288
rect 34978 31240 35034 31249
rect 34978 31175 35034 31184
rect 34992 31142 35020 31175
rect 34980 31136 35032 31142
rect 34980 31078 35032 31084
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34888 30728 34940 30734
rect 34888 30670 34940 30676
rect 34900 30054 34928 30670
rect 35360 30258 35388 32166
rect 35452 31906 35480 34478
rect 35544 32026 35572 37198
rect 35636 35601 35664 38927
rect 35716 38276 35768 38282
rect 35716 38218 35768 38224
rect 35728 36854 35756 38218
rect 35820 37210 35848 39335
rect 38198 39200 38254 40000
rect 38014 38176 38070 38185
rect 38014 38111 38070 38120
rect 35820 37182 35940 37210
rect 38028 37194 38056 38111
rect 38212 37346 38240 39200
rect 38476 37460 38528 37466
rect 38476 37402 38528 37408
rect 38120 37318 38240 37346
rect 38120 37262 38148 37318
rect 38108 37256 38160 37262
rect 38108 37198 38160 37204
rect 35808 37120 35860 37126
rect 35808 37062 35860 37068
rect 35820 36854 35848 37062
rect 35716 36848 35768 36854
rect 35716 36790 35768 36796
rect 35808 36848 35860 36854
rect 35808 36790 35860 36796
rect 35912 36700 35940 37182
rect 37556 37188 37608 37194
rect 37556 37130 37608 37136
rect 38016 37188 38068 37194
rect 38016 37130 38068 37136
rect 37372 37120 37424 37126
rect 37372 37062 37424 37068
rect 37462 37088 37518 37097
rect 36084 36780 36136 36786
rect 36084 36722 36136 36728
rect 35820 36672 35940 36700
rect 35714 35728 35770 35737
rect 35714 35663 35770 35672
rect 35622 35592 35678 35601
rect 35622 35527 35678 35536
rect 35624 34604 35676 34610
rect 35624 34546 35676 34552
rect 35636 33658 35664 34546
rect 35728 34241 35756 35663
rect 35714 34232 35770 34241
rect 35714 34167 35716 34176
rect 35768 34167 35770 34176
rect 35716 34138 35768 34144
rect 35728 34066 35756 34138
rect 35716 34060 35768 34066
rect 35716 34002 35768 34008
rect 35820 33946 35848 36672
rect 36096 36310 36124 36722
rect 36176 36576 36228 36582
rect 36176 36518 36228 36524
rect 36452 36576 36504 36582
rect 36452 36518 36504 36524
rect 36084 36304 36136 36310
rect 36084 36246 36136 36252
rect 36188 36174 36216 36518
rect 36084 36168 36136 36174
rect 36084 36110 36136 36116
rect 36176 36168 36228 36174
rect 36176 36110 36228 36116
rect 35898 35184 35954 35193
rect 35898 35119 35954 35128
rect 35912 34241 35940 35119
rect 36096 35086 36124 36110
rect 36360 35624 36412 35630
rect 36360 35566 36412 35572
rect 36084 35080 36136 35086
rect 36084 35022 36136 35028
rect 36176 35080 36228 35086
rect 36176 35022 36228 35028
rect 35898 34232 35954 34241
rect 35898 34167 35954 34176
rect 36096 34066 36124 35022
rect 36188 34542 36216 35022
rect 36176 34536 36228 34542
rect 36174 34504 36176 34513
rect 36228 34504 36230 34513
rect 36174 34439 36230 34448
rect 36084 34060 36136 34066
rect 36084 34002 36136 34008
rect 35992 33992 36044 33998
rect 35990 33960 35992 33969
rect 36044 33960 36046 33969
rect 35716 33924 35768 33930
rect 35820 33918 35940 33946
rect 35716 33866 35768 33872
rect 35728 33833 35756 33866
rect 35808 33856 35860 33862
rect 35714 33824 35770 33833
rect 35808 33798 35860 33804
rect 35714 33759 35770 33768
rect 35624 33652 35676 33658
rect 35624 33594 35676 33600
rect 35820 33590 35848 33798
rect 35808 33584 35860 33590
rect 35622 33552 35678 33561
rect 35808 33526 35860 33532
rect 35912 33538 35940 33918
rect 35990 33895 36046 33904
rect 36268 33924 36320 33930
rect 36268 33866 36320 33872
rect 36176 33856 36228 33862
rect 36176 33798 36228 33804
rect 35912 33510 36032 33538
rect 35622 33487 35678 33496
rect 35636 32366 35664 33487
rect 35716 33448 35768 33454
rect 35716 33390 35768 33396
rect 35900 33448 35952 33454
rect 35900 33390 35952 33396
rect 35728 33289 35756 33390
rect 35714 33280 35770 33289
rect 35714 33215 35770 33224
rect 35714 33008 35770 33017
rect 35714 32943 35716 32952
rect 35768 32943 35770 32952
rect 35716 32914 35768 32920
rect 35912 32858 35940 33390
rect 35820 32842 35940 32858
rect 35808 32836 35940 32842
rect 35860 32830 35940 32836
rect 35808 32778 35860 32784
rect 35716 32768 35768 32774
rect 35716 32710 35768 32716
rect 35624 32360 35676 32366
rect 35624 32302 35676 32308
rect 35532 32020 35584 32026
rect 35532 31962 35584 31968
rect 35452 31878 35664 31906
rect 35438 31784 35494 31793
rect 35438 31719 35494 31728
rect 35452 31346 35480 31719
rect 35440 31340 35492 31346
rect 35440 31282 35492 31288
rect 35452 30734 35480 31282
rect 35440 30728 35492 30734
rect 35440 30670 35492 30676
rect 35348 30252 35400 30258
rect 35348 30194 35400 30200
rect 34888 30048 34940 30054
rect 34702 30016 34758 30025
rect 35452 30025 35480 30670
rect 34888 29990 34940 29996
rect 35438 30016 35494 30025
rect 34702 29951 34758 29960
rect 34934 29948 35242 29957
rect 35438 29951 35494 29960
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34980 29844 35032 29850
rect 34980 29786 35032 29792
rect 34612 29776 34664 29782
rect 34612 29718 34664 29724
rect 34796 29708 34848 29714
rect 34848 29668 34928 29696
rect 34796 29650 34848 29656
rect 34428 29640 34480 29646
rect 34428 29582 34480 29588
rect 34256 28750 34376 28778
rect 34256 28744 34284 28750
rect 34164 28716 34284 28744
rect 34164 28540 34192 28716
rect 34164 28512 34376 28540
rect 34072 28444 34192 28472
rect 34164 28082 34192 28444
rect 34244 28416 34296 28422
rect 34244 28358 34296 28364
rect 34060 28076 34112 28082
rect 34060 28018 34112 28024
rect 34152 28076 34204 28082
rect 34152 28018 34204 28024
rect 34072 27878 34100 28018
rect 34060 27872 34112 27878
rect 34060 27814 34112 27820
rect 33980 27254 34100 27282
rect 33796 27084 34008 27112
rect 33784 26988 33836 26994
rect 33784 26930 33836 26936
rect 33796 26450 33824 26930
rect 33876 26852 33928 26858
rect 33876 26794 33928 26800
rect 33784 26444 33836 26450
rect 33784 26386 33836 26392
rect 33796 25673 33824 26386
rect 33888 26382 33916 26794
rect 33876 26376 33928 26382
rect 33876 26318 33928 26324
rect 33980 25906 34008 27084
rect 34072 26994 34100 27254
rect 34060 26988 34112 26994
rect 34060 26930 34112 26936
rect 34152 26784 34204 26790
rect 34152 26726 34204 26732
rect 33968 25900 34020 25906
rect 33968 25842 34020 25848
rect 33876 25764 33928 25770
rect 33876 25706 33928 25712
rect 33782 25664 33838 25673
rect 33782 25599 33838 25608
rect 33784 25356 33836 25362
rect 33784 25298 33836 25304
rect 33796 24410 33824 25298
rect 33888 25158 33916 25706
rect 33980 25702 34008 25842
rect 33968 25696 34020 25702
rect 33968 25638 34020 25644
rect 33876 25152 33928 25158
rect 33876 25094 33928 25100
rect 34058 24984 34114 24993
rect 34058 24919 34114 24928
rect 33876 24812 33928 24818
rect 33928 24772 34008 24800
rect 33876 24754 33928 24760
rect 33876 24608 33928 24614
rect 33876 24550 33928 24556
rect 33784 24404 33836 24410
rect 33784 24346 33836 24352
rect 33796 24206 33824 24346
rect 33784 24200 33836 24206
rect 33784 24142 33836 24148
rect 33888 23848 33916 24550
rect 33796 23820 33916 23848
rect 33796 23730 33824 23820
rect 33784 23724 33836 23730
rect 33784 23666 33836 23672
rect 33876 23724 33928 23730
rect 33876 23666 33928 23672
rect 33690 23352 33746 23361
rect 33888 23322 33916 23666
rect 33690 23287 33746 23296
rect 33876 23316 33928 23322
rect 33876 23258 33928 23264
rect 33782 22944 33838 22953
rect 33782 22879 33838 22888
rect 33600 22568 33652 22574
rect 33600 22510 33652 22516
rect 33796 22098 33824 22879
rect 33980 22642 34008 24772
rect 34072 24750 34100 24919
rect 34060 24744 34112 24750
rect 34060 24686 34112 24692
rect 34058 24032 34114 24041
rect 34058 23967 34114 23976
rect 33876 22636 33928 22642
rect 33876 22578 33928 22584
rect 33968 22636 34020 22642
rect 33968 22578 34020 22584
rect 33888 22409 33916 22578
rect 33874 22400 33930 22409
rect 33874 22335 33930 22344
rect 33784 22092 33836 22098
rect 33784 22034 33836 22040
rect 33876 22092 33928 22098
rect 33876 22034 33928 22040
rect 33692 22024 33744 22030
rect 33692 21966 33744 21972
rect 33600 21548 33652 21554
rect 33600 21490 33652 21496
rect 33508 21344 33560 21350
rect 33508 21286 33560 21292
rect 33416 20256 33468 20262
rect 33416 20198 33468 20204
rect 33612 20097 33640 21490
rect 33598 20088 33654 20097
rect 33598 20023 33654 20032
rect 33704 19922 33732 21966
rect 33796 21049 33824 22034
rect 33782 21040 33838 21049
rect 33782 20975 33838 20984
rect 33784 20596 33836 20602
rect 33784 20538 33836 20544
rect 33796 20466 33824 20538
rect 33784 20460 33836 20466
rect 33784 20402 33836 20408
rect 33692 19916 33744 19922
rect 33692 19858 33744 19864
rect 33508 19780 33560 19786
rect 33508 19722 33560 19728
rect 33600 19780 33652 19786
rect 33600 19722 33652 19728
rect 33230 19479 33286 19488
rect 33324 19508 33376 19514
rect 33244 19446 33272 19479
rect 33324 19450 33376 19456
rect 33232 19440 33284 19446
rect 33232 19382 33284 19388
rect 33140 18964 33192 18970
rect 33140 18906 33192 18912
rect 33244 18834 33272 19382
rect 33232 18828 33284 18834
rect 33232 18770 33284 18776
rect 33140 18692 33192 18698
rect 33140 18634 33192 18640
rect 33152 18193 33180 18634
rect 33244 18290 33272 18770
rect 33232 18284 33284 18290
rect 33232 18226 33284 18232
rect 33138 18184 33194 18193
rect 33138 18119 33194 18128
rect 33138 18048 33194 18057
rect 33138 17983 33194 17992
rect 32876 17326 33088 17354
rect 32772 14068 32824 14074
rect 32772 14010 32824 14016
rect 32876 12850 32904 17326
rect 32956 16652 33008 16658
rect 32956 16594 33008 16600
rect 32968 16538 32996 16594
rect 32968 16510 33088 16538
rect 32956 16108 33008 16114
rect 32956 16050 33008 16056
rect 32968 13734 32996 16050
rect 33060 14414 33088 16510
rect 33152 15706 33180 17983
rect 33244 17270 33272 18226
rect 33336 18057 33364 19450
rect 33520 19310 33548 19722
rect 33508 19304 33560 19310
rect 33508 19246 33560 19252
rect 33520 19122 33548 19246
rect 33428 19094 33548 19122
rect 33428 18290 33456 19094
rect 33612 18970 33640 19722
rect 33704 19378 33732 19858
rect 33692 19372 33744 19378
rect 33692 19314 33744 19320
rect 33508 18964 33560 18970
rect 33508 18906 33560 18912
rect 33600 18964 33652 18970
rect 33600 18906 33652 18912
rect 33416 18284 33468 18290
rect 33416 18226 33468 18232
rect 33322 18048 33378 18057
rect 33322 17983 33378 17992
rect 33428 17898 33456 18226
rect 33520 18057 33548 18906
rect 33612 18290 33640 18906
rect 33692 18624 33744 18630
rect 33692 18566 33744 18572
rect 33600 18284 33652 18290
rect 33600 18226 33652 18232
rect 33506 18048 33562 18057
rect 33506 17983 33562 17992
rect 33336 17870 33456 17898
rect 33336 17678 33364 17870
rect 33612 17864 33640 18226
rect 33704 18154 33732 18566
rect 33796 18272 33824 20402
rect 33888 19854 33916 22034
rect 33980 22030 34008 22578
rect 33968 22024 34020 22030
rect 33968 21966 34020 21972
rect 34072 21434 34100 23967
rect 34164 23662 34192 26726
rect 34256 24614 34284 28358
rect 34244 24608 34296 24614
rect 34244 24550 34296 24556
rect 34244 23724 34296 23730
rect 34348 23712 34376 28512
rect 34440 28257 34468 29582
rect 34704 29572 34756 29578
rect 34704 29514 34756 29520
rect 34612 29504 34664 29510
rect 34612 29446 34664 29452
rect 34520 29096 34572 29102
rect 34520 29038 34572 29044
rect 34426 28248 34482 28257
rect 34426 28183 34482 28192
rect 34428 28076 34480 28082
rect 34428 28018 34480 28024
rect 34440 27985 34468 28018
rect 34426 27976 34482 27985
rect 34426 27911 34482 27920
rect 34428 27872 34480 27878
rect 34426 27840 34428 27849
rect 34480 27840 34482 27849
rect 34426 27775 34482 27784
rect 34532 27577 34560 29038
rect 34624 28393 34652 29446
rect 34610 28384 34666 28393
rect 34610 28319 34666 28328
rect 34612 27872 34664 27878
rect 34612 27814 34664 27820
rect 34624 27713 34652 27814
rect 34610 27704 34666 27713
rect 34610 27639 34666 27648
rect 34518 27568 34574 27577
rect 34716 27554 34744 29514
rect 34900 29102 34928 29668
rect 34888 29096 34940 29102
rect 34888 29038 34940 29044
rect 34992 28994 35020 29786
rect 35530 29744 35586 29753
rect 35530 29679 35532 29688
rect 35584 29679 35586 29688
rect 35532 29650 35584 29656
rect 35532 29300 35584 29306
rect 35532 29242 35584 29248
rect 35072 29164 35124 29170
rect 35072 29106 35124 29112
rect 34808 28966 35020 28994
rect 35084 28994 35112 29106
rect 35440 29028 35492 29034
rect 35084 28966 35388 28994
rect 35440 28970 35492 28976
rect 34808 28801 34836 28966
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34794 28792 34850 28801
rect 34934 28795 35242 28804
rect 34794 28727 34850 28736
rect 34808 28257 34836 28727
rect 34886 28656 34942 28665
rect 34886 28591 34888 28600
rect 34940 28591 34942 28600
rect 34888 28562 34940 28568
rect 34794 28248 34850 28257
rect 34794 28183 34850 28192
rect 34796 28144 34848 28150
rect 34796 28086 34848 28092
rect 34808 27674 34836 28086
rect 34900 28064 34928 28562
rect 35360 28218 35388 28966
rect 35348 28212 35400 28218
rect 35348 28154 35400 28160
rect 35164 28076 35216 28082
rect 34900 28036 35164 28064
rect 35164 28018 35216 28024
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 27668 34848 27674
rect 34796 27610 34848 27616
rect 35162 27568 35218 27577
rect 34716 27526 35112 27554
rect 34518 27503 34574 27512
rect 35084 27470 35112 27526
rect 35162 27503 35218 27512
rect 34888 27464 34940 27470
rect 34888 27406 34940 27412
rect 35072 27464 35124 27470
rect 35072 27406 35124 27412
rect 34428 27396 34480 27402
rect 34428 27338 34480 27344
rect 34796 27396 34848 27402
rect 34796 27338 34848 27344
rect 34440 26790 34468 27338
rect 34520 27328 34572 27334
rect 34520 27270 34572 27276
rect 34428 26784 34480 26790
rect 34428 26726 34480 26732
rect 34532 25945 34560 27270
rect 34612 27056 34664 27062
rect 34612 26998 34664 27004
rect 34518 25936 34574 25945
rect 34518 25871 34574 25880
rect 34428 25832 34480 25838
rect 34428 25774 34480 25780
rect 34440 25362 34468 25774
rect 34428 25356 34480 25362
rect 34428 25298 34480 25304
rect 34624 24936 34652 26998
rect 34704 26784 34756 26790
rect 34704 26726 34756 26732
rect 34532 24908 34652 24936
rect 34428 24336 34480 24342
rect 34428 24278 34480 24284
rect 34296 23684 34376 23712
rect 34244 23666 34296 23672
rect 34152 23656 34204 23662
rect 34152 23598 34204 23604
rect 34336 23520 34388 23526
rect 34150 23488 34206 23497
rect 34336 23462 34388 23468
rect 34150 23423 34206 23432
rect 34164 22710 34192 23423
rect 34244 23112 34296 23118
rect 34244 23054 34296 23060
rect 34152 22704 34204 22710
rect 34152 22646 34204 22652
rect 34164 22098 34192 22646
rect 34152 22092 34204 22098
rect 34152 22034 34204 22040
rect 34256 21729 34284 23054
rect 34242 21720 34298 21729
rect 34242 21655 34298 21664
rect 34072 21406 34192 21434
rect 33968 21344 34020 21350
rect 33968 21286 34020 21292
rect 34060 21344 34112 21350
rect 34060 21286 34112 21292
rect 33980 20777 34008 21286
rect 34072 20942 34100 21286
rect 34164 20942 34192 21406
rect 34060 20936 34112 20942
rect 34060 20878 34112 20884
rect 34152 20936 34204 20942
rect 34152 20878 34204 20884
rect 33966 20768 34022 20777
rect 33966 20703 34022 20712
rect 34164 20618 34192 20878
rect 34036 20590 34192 20618
rect 34242 20632 34298 20641
rect 34036 20482 34064 20590
rect 34242 20567 34298 20576
rect 34036 20466 34100 20482
rect 34036 20460 34112 20466
rect 34036 20454 34060 20460
rect 34060 20402 34112 20408
rect 34152 20460 34204 20466
rect 34152 20402 34204 20408
rect 33966 20224 34022 20233
rect 33966 20159 34022 20168
rect 33876 19848 33928 19854
rect 33876 19790 33928 19796
rect 33888 19553 33916 19790
rect 33874 19544 33930 19553
rect 33874 19479 33930 19488
rect 33980 19394 34008 20159
rect 34072 19446 34100 20402
rect 34164 20058 34192 20402
rect 34152 20052 34204 20058
rect 34152 19994 34204 20000
rect 33888 19378 34008 19394
rect 34060 19440 34112 19446
rect 34060 19382 34112 19388
rect 33876 19372 34008 19378
rect 33928 19366 34008 19372
rect 34072 19334 34100 19382
rect 34256 19334 34284 20567
rect 33876 19314 33928 19320
rect 33980 19306 34100 19334
rect 34164 19306 34284 19334
rect 33980 18902 34008 19306
rect 34060 19236 34112 19242
rect 34060 19178 34112 19184
rect 33968 18896 34020 18902
rect 33968 18838 34020 18844
rect 33968 18624 34020 18630
rect 33968 18566 34020 18572
rect 33876 18284 33928 18290
rect 33796 18244 33876 18272
rect 33692 18148 33744 18154
rect 33692 18090 33744 18096
rect 33520 17836 33640 17864
rect 33414 17776 33470 17785
rect 33414 17711 33470 17720
rect 33428 17678 33456 17711
rect 33520 17678 33548 17836
rect 33704 17785 33732 18090
rect 33690 17776 33746 17785
rect 33600 17740 33652 17746
rect 33690 17711 33746 17720
rect 33600 17682 33652 17688
rect 33324 17672 33376 17678
rect 33324 17614 33376 17620
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 33508 17672 33560 17678
rect 33508 17614 33560 17620
rect 33416 17536 33468 17542
rect 33416 17478 33468 17484
rect 33232 17264 33284 17270
rect 33232 17206 33284 17212
rect 33428 16674 33456 17478
rect 33612 17270 33640 17682
rect 33796 17678 33824 18244
rect 33876 18226 33928 18232
rect 33874 18048 33930 18057
rect 33874 17983 33930 17992
rect 33784 17672 33836 17678
rect 33784 17614 33836 17620
rect 33692 17604 33744 17610
rect 33692 17546 33744 17552
rect 33704 17377 33732 17546
rect 33690 17368 33746 17377
rect 33690 17303 33746 17312
rect 33600 17264 33652 17270
rect 33600 17206 33652 17212
rect 33704 16794 33732 17303
rect 33692 16788 33744 16794
rect 33692 16730 33744 16736
rect 33428 16646 33548 16674
rect 33520 16590 33548 16646
rect 33508 16584 33560 16590
rect 33508 16526 33560 16532
rect 33600 16516 33652 16522
rect 33600 16458 33652 16464
rect 33612 16250 33640 16458
rect 33704 16250 33732 16730
rect 33600 16244 33652 16250
rect 33600 16186 33652 16192
rect 33692 16244 33744 16250
rect 33692 16186 33744 16192
rect 33140 15700 33192 15706
rect 33140 15642 33192 15648
rect 33888 15450 33916 17983
rect 33980 16658 34008 18566
rect 34072 17814 34100 19178
rect 34164 18193 34192 19306
rect 34348 19224 34376 23462
rect 34440 23322 34468 24278
rect 34532 24177 34560 24908
rect 34612 24812 34664 24818
rect 34612 24754 34664 24760
rect 34518 24168 34574 24177
rect 34518 24103 34574 24112
rect 34624 23730 34652 24754
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34428 23316 34480 23322
rect 34428 23258 34480 23264
rect 34428 23044 34480 23050
rect 34428 22986 34480 22992
rect 34440 22953 34468 22986
rect 34426 22944 34482 22953
rect 34426 22879 34482 22888
rect 34428 22568 34480 22574
rect 34428 22510 34480 22516
rect 34440 22234 34468 22510
rect 34532 22506 34560 23462
rect 34612 23044 34664 23050
rect 34612 22986 34664 22992
rect 34520 22500 34572 22506
rect 34520 22442 34572 22448
rect 34518 22400 34574 22409
rect 34518 22335 34574 22344
rect 34428 22228 34480 22234
rect 34428 22170 34480 22176
rect 34532 21554 34560 22335
rect 34624 22273 34652 22986
rect 34610 22264 34666 22273
rect 34610 22199 34666 22208
rect 34716 21842 34744 26726
rect 34808 26246 34836 27338
rect 34900 27305 34928 27406
rect 35176 27402 35204 27503
rect 35164 27396 35216 27402
rect 35164 27338 35216 27344
rect 34886 27296 34942 27305
rect 34886 27231 34942 27240
rect 34900 27130 34928 27231
rect 34888 27124 34940 27130
rect 34888 27066 34940 27072
rect 34978 27024 35034 27033
rect 34978 26959 34980 26968
rect 35032 26959 35034 26968
rect 34980 26930 35032 26936
rect 35360 26761 35388 28154
rect 35452 27577 35480 28970
rect 35438 27568 35494 27577
rect 35438 27503 35494 27512
rect 35440 26988 35492 26994
rect 35440 26930 35492 26936
rect 35346 26752 35402 26761
rect 34934 26684 35242 26693
rect 35346 26687 35402 26696
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34886 26480 34942 26489
rect 34886 26415 34942 26424
rect 35162 26480 35218 26489
rect 35162 26415 35218 26424
rect 34900 26382 34928 26415
rect 34888 26376 34940 26382
rect 34888 26318 34940 26324
rect 35176 26314 35204 26415
rect 35072 26308 35124 26314
rect 35072 26250 35124 26256
rect 35164 26308 35216 26314
rect 35164 26250 35216 26256
rect 35348 26308 35400 26314
rect 35452 26296 35480 26930
rect 35400 26268 35480 26296
rect 35348 26250 35400 26256
rect 34796 26240 34848 26246
rect 34796 26182 34848 26188
rect 35084 26042 35112 26250
rect 35072 26036 35124 26042
rect 35072 25978 35124 25984
rect 35164 26036 35216 26042
rect 35164 25978 35216 25984
rect 35072 25832 35124 25838
rect 35176 25820 35204 25978
rect 35124 25792 35204 25820
rect 35072 25774 35124 25780
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35256 25288 35308 25294
rect 35254 25256 35256 25265
rect 35308 25256 35310 25265
rect 34980 25220 35032 25226
rect 35254 25191 35310 25200
rect 34980 25162 35032 25168
rect 34796 25152 34848 25158
rect 34796 25094 34848 25100
rect 34808 23866 34836 25094
rect 34886 24984 34942 24993
rect 34992 24954 35020 25162
rect 35360 25158 35388 26250
rect 35544 25430 35572 29242
rect 35532 25424 35584 25430
rect 35532 25366 35584 25372
rect 35348 25152 35400 25158
rect 35348 25094 35400 25100
rect 35440 25152 35492 25158
rect 35440 25094 35492 25100
rect 34886 24919 34942 24928
rect 34980 24948 35032 24954
rect 34900 24818 34928 24919
rect 34980 24890 35032 24896
rect 34888 24812 34940 24818
rect 34888 24754 34940 24760
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 34900 24596 34928 24754
rect 34864 24568 34928 24596
rect 34864 24392 34892 24568
rect 35360 24562 35388 24754
rect 35452 24682 35480 25094
rect 35544 24818 35572 25366
rect 35636 25362 35664 31878
rect 35728 31249 35756 32710
rect 35806 32600 35862 32609
rect 36004 32586 36032 33510
rect 36188 33386 36216 33798
rect 36280 33697 36308 33866
rect 36266 33688 36322 33697
rect 36266 33623 36322 33632
rect 36280 33522 36308 33623
rect 36268 33516 36320 33522
rect 36268 33458 36320 33464
rect 36176 33380 36228 33386
rect 36176 33322 36228 33328
rect 36268 33380 36320 33386
rect 36268 33322 36320 33328
rect 36176 32768 36228 32774
rect 36176 32710 36228 32716
rect 36004 32558 36124 32586
rect 36188 32570 36216 32710
rect 35806 32535 35862 32544
rect 35820 32450 35848 32535
rect 36096 32473 36124 32558
rect 36176 32564 36228 32570
rect 36176 32506 36228 32512
rect 36082 32464 36138 32473
rect 35820 32422 36032 32450
rect 35808 32360 35860 32366
rect 35808 32302 35860 32308
rect 35820 31686 35848 32302
rect 35900 32224 35952 32230
rect 35900 32166 35952 32172
rect 35808 31680 35860 31686
rect 35808 31622 35860 31628
rect 35808 31272 35860 31278
rect 35714 31240 35770 31249
rect 35808 31214 35860 31220
rect 35714 31175 35770 31184
rect 35716 31136 35768 31142
rect 35716 31078 35768 31084
rect 35728 29646 35756 31078
rect 35820 30569 35848 31214
rect 35912 30734 35940 32166
rect 35900 30728 35952 30734
rect 35900 30670 35952 30676
rect 35806 30560 35862 30569
rect 35806 30495 35862 30504
rect 35808 30048 35860 30054
rect 35808 29990 35860 29996
rect 35716 29640 35768 29646
rect 35716 29582 35768 29588
rect 35716 29164 35768 29170
rect 35716 29106 35768 29112
rect 35728 28966 35756 29106
rect 35716 28960 35768 28966
rect 35716 28902 35768 28908
rect 35714 28656 35770 28665
rect 35714 28591 35770 28600
rect 35728 28422 35756 28591
rect 35716 28416 35768 28422
rect 35716 28358 35768 28364
rect 35820 27418 35848 29990
rect 36004 29170 36032 32422
rect 36082 32399 36138 32408
rect 36176 32428 36228 32434
rect 36176 32370 36228 32376
rect 36084 32292 36136 32298
rect 36084 32234 36136 32240
rect 36096 31346 36124 32234
rect 36188 32065 36216 32370
rect 36174 32056 36230 32065
rect 36174 31991 36230 32000
rect 36084 31340 36136 31346
rect 36084 31282 36136 31288
rect 36280 31226 36308 33322
rect 36372 31754 36400 35566
rect 36464 33862 36492 36518
rect 36542 36272 36598 36281
rect 36542 36207 36598 36216
rect 36556 36106 36584 36207
rect 36910 36136 36966 36145
rect 36544 36100 36596 36106
rect 36910 36071 36966 36080
rect 36544 36042 36596 36048
rect 36634 36000 36690 36009
rect 36634 35935 36690 35944
rect 36544 35760 36596 35766
rect 36544 35702 36596 35708
rect 36556 35154 36584 35702
rect 36648 35494 36676 35935
rect 36924 35766 36952 36071
rect 37188 36032 37240 36038
rect 37188 35974 37240 35980
rect 36912 35760 36964 35766
rect 36912 35702 36964 35708
rect 36728 35556 36780 35562
rect 36728 35498 36780 35504
rect 36636 35488 36688 35494
rect 36636 35430 36688 35436
rect 36740 35442 36768 35498
rect 36648 35222 36676 35430
rect 36740 35414 36860 35442
rect 36636 35216 36688 35222
rect 36636 35158 36688 35164
rect 36544 35148 36596 35154
rect 36544 35090 36596 35096
rect 36726 35048 36782 35057
rect 36726 34983 36728 34992
rect 36780 34983 36782 34992
rect 36728 34954 36780 34960
rect 36832 34950 36860 35414
rect 36820 34944 36872 34950
rect 36820 34886 36872 34892
rect 36648 34610 36768 34626
rect 36544 34604 36596 34610
rect 36544 34546 36596 34552
rect 36648 34604 36780 34610
rect 36648 34598 36728 34604
rect 36452 33856 36504 33862
rect 36452 33798 36504 33804
rect 36464 33522 36492 33798
rect 36452 33516 36504 33522
rect 36452 33458 36504 33464
rect 36556 33386 36584 34546
rect 36648 33522 36676 34598
rect 36728 34546 36780 34552
rect 36832 34474 36860 34886
rect 36924 34746 36952 35702
rect 37004 35692 37056 35698
rect 37004 35634 37056 35640
rect 36912 34740 36964 34746
rect 36912 34682 36964 34688
rect 36728 34468 36780 34474
rect 36728 34410 36780 34416
rect 36820 34468 36872 34474
rect 36820 34410 36872 34416
rect 36636 33516 36688 33522
rect 36636 33458 36688 33464
rect 36544 33380 36596 33386
rect 36544 33322 36596 33328
rect 36648 32910 36676 33458
rect 36740 33318 36768 34410
rect 36820 34060 36872 34066
rect 36820 34002 36872 34008
rect 36728 33312 36780 33318
rect 36728 33254 36780 33260
rect 36740 32978 36768 33254
rect 36728 32972 36780 32978
rect 36728 32914 36780 32920
rect 36636 32904 36688 32910
rect 36636 32846 36688 32852
rect 36544 32836 36596 32842
rect 36544 32778 36596 32784
rect 36450 32328 36506 32337
rect 36450 32263 36506 32272
rect 36464 31958 36492 32263
rect 36556 32026 36584 32778
rect 36544 32020 36596 32026
rect 36544 31962 36596 31968
rect 36452 31952 36504 31958
rect 36450 31920 36452 31929
rect 36504 31920 36506 31929
rect 36450 31855 36506 31864
rect 36372 31726 36492 31754
rect 36360 31680 36412 31686
rect 36360 31622 36412 31628
rect 36372 31346 36400 31622
rect 36360 31340 36412 31346
rect 36360 31282 36412 31288
rect 36188 31210 36308 31226
rect 36176 31204 36308 31210
rect 36228 31198 36308 31204
rect 36176 31146 36228 31152
rect 36084 30932 36136 30938
rect 36084 30874 36136 30880
rect 36096 30734 36124 30874
rect 36084 30728 36136 30734
rect 36084 30670 36136 30676
rect 36096 30394 36124 30670
rect 36188 30666 36216 31146
rect 36268 31136 36320 31142
rect 36268 31078 36320 31084
rect 36280 30666 36308 31078
rect 36176 30660 36228 30666
rect 36176 30602 36228 30608
rect 36268 30660 36320 30666
rect 36268 30602 36320 30608
rect 36084 30388 36136 30394
rect 36084 30330 36136 30336
rect 36084 29844 36136 29850
rect 36084 29786 36136 29792
rect 35992 29164 36044 29170
rect 35992 29106 36044 29112
rect 35900 29096 35952 29102
rect 35900 29038 35952 29044
rect 35728 27390 35848 27418
rect 35728 27062 35756 27390
rect 35808 27328 35860 27334
rect 35808 27270 35860 27276
rect 35820 27062 35848 27270
rect 35716 27056 35768 27062
rect 35716 26998 35768 27004
rect 35808 27056 35860 27062
rect 35808 26998 35860 27004
rect 35912 26994 35940 29038
rect 35992 28960 36044 28966
rect 35992 28902 36044 28908
rect 36004 28393 36032 28902
rect 36096 28762 36124 29786
rect 36188 29510 36216 30602
rect 36360 30048 36412 30054
rect 36266 30016 36322 30025
rect 36360 29990 36412 29996
rect 36266 29951 36322 29960
rect 36176 29504 36228 29510
rect 36176 29446 36228 29452
rect 36084 28756 36136 28762
rect 36084 28698 36136 28704
rect 35990 28384 36046 28393
rect 35990 28319 36046 28328
rect 35992 27600 36044 27606
rect 35992 27542 36044 27548
rect 35900 26988 35952 26994
rect 35900 26930 35952 26936
rect 35808 26920 35860 26926
rect 35714 26888 35770 26897
rect 35860 26868 35940 26874
rect 35808 26862 35940 26868
rect 35820 26846 35940 26862
rect 35714 26823 35770 26832
rect 35624 25356 35676 25362
rect 35624 25298 35676 25304
rect 35624 24948 35676 24954
rect 35624 24890 35676 24896
rect 35532 24812 35584 24818
rect 35532 24754 35584 24760
rect 35440 24676 35492 24682
rect 35440 24618 35492 24624
rect 35360 24534 35480 24562
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35348 24404 35400 24410
rect 34864 24364 35204 24392
rect 34888 24200 34940 24206
rect 34888 24142 34940 24148
rect 35072 24200 35124 24206
rect 35072 24142 35124 24148
rect 34900 23866 34928 24142
rect 35084 24041 35112 24142
rect 35070 24032 35126 24041
rect 35070 23967 35126 23976
rect 34796 23860 34848 23866
rect 34796 23802 34848 23808
rect 34888 23860 34940 23866
rect 34888 23802 34940 23808
rect 34796 23724 34848 23730
rect 35176 23712 35204 24364
rect 35348 24346 35400 24352
rect 35256 24132 35308 24138
rect 35256 24074 35308 24080
rect 35268 24041 35296 24074
rect 35254 24032 35310 24041
rect 35254 23967 35310 23976
rect 35256 23724 35308 23730
rect 35176 23684 35256 23712
rect 34796 23666 34848 23672
rect 35256 23666 35308 23672
rect 34808 23202 34836 23666
rect 35268 23526 35296 23666
rect 35256 23520 35308 23526
rect 35256 23462 35308 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35164 23316 35216 23322
rect 35164 23258 35216 23264
rect 34808 23174 34928 23202
rect 34796 23112 34848 23118
rect 34796 23054 34848 23060
rect 34808 22030 34836 23054
rect 34900 22545 34928 23174
rect 35176 23118 35204 23258
rect 35360 23118 35388 24346
rect 35452 23769 35480 24534
rect 35438 23760 35494 23769
rect 35438 23695 35440 23704
rect 35492 23695 35494 23704
rect 35440 23666 35492 23672
rect 35164 23112 35216 23118
rect 35164 23054 35216 23060
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 35176 22710 35204 23054
rect 35164 22704 35216 22710
rect 35164 22646 35216 22652
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 34886 22536 34942 22545
rect 34886 22471 34942 22480
rect 35360 22409 35388 22578
rect 35346 22400 35402 22409
rect 34934 22332 35242 22341
rect 35346 22335 35402 22344
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35452 22216 35480 23666
rect 35544 23186 35572 24754
rect 35636 24698 35664 24890
rect 35728 24857 35756 26823
rect 35808 26784 35860 26790
rect 35808 26726 35860 26732
rect 35820 26586 35848 26726
rect 35808 26580 35860 26586
rect 35808 26522 35860 26528
rect 35912 26518 35940 26846
rect 35900 26512 35952 26518
rect 35900 26454 35952 26460
rect 35808 26444 35860 26450
rect 35808 26386 35860 26392
rect 35820 25401 35848 26386
rect 35900 26376 35952 26382
rect 35900 26318 35952 26324
rect 35912 26246 35940 26318
rect 35900 26240 35952 26246
rect 35900 26182 35952 26188
rect 35806 25392 35862 25401
rect 35806 25327 35862 25336
rect 35808 25220 35860 25226
rect 35860 25180 35940 25208
rect 35808 25162 35860 25168
rect 35714 24848 35770 24857
rect 35714 24783 35770 24792
rect 35808 24812 35860 24818
rect 35808 24754 35860 24760
rect 35820 24721 35848 24754
rect 35806 24712 35862 24721
rect 35636 24670 35756 24698
rect 35728 24342 35756 24670
rect 35806 24647 35862 24656
rect 35808 24608 35860 24614
rect 35808 24550 35860 24556
rect 35624 24336 35676 24342
rect 35624 24278 35676 24284
rect 35716 24336 35768 24342
rect 35716 24278 35768 24284
rect 35532 23180 35584 23186
rect 35532 23122 35584 23128
rect 35532 22704 35584 22710
rect 35532 22646 35584 22652
rect 35360 22188 35480 22216
rect 34888 22160 34940 22166
rect 34888 22102 34940 22108
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 34624 21814 34744 21842
rect 34624 21690 34652 21814
rect 34612 21684 34664 21690
rect 34612 21626 34664 21632
rect 34520 21548 34572 21554
rect 34520 21490 34572 21496
rect 34428 21480 34480 21486
rect 34428 21422 34480 21428
rect 34440 21010 34468 21422
rect 34428 21004 34480 21010
rect 34428 20946 34480 20952
rect 34426 20496 34482 20505
rect 34426 20431 34428 20440
rect 34480 20431 34482 20440
rect 34428 20402 34480 20408
rect 34428 20256 34480 20262
rect 34428 20198 34480 20204
rect 34256 19196 34376 19224
rect 34150 18184 34206 18193
rect 34150 18119 34206 18128
rect 34152 17876 34204 17882
rect 34152 17818 34204 17824
rect 34060 17808 34112 17814
rect 34060 17750 34112 17756
rect 34164 17082 34192 17818
rect 34256 17202 34284 19196
rect 34244 17196 34296 17202
rect 34244 17138 34296 17144
rect 34164 17054 34284 17082
rect 33968 16652 34020 16658
rect 33968 16594 34020 16600
rect 33796 15422 33916 15450
rect 33600 15360 33652 15366
rect 33600 15302 33652 15308
rect 33508 15020 33560 15026
rect 33508 14962 33560 14968
rect 33324 14952 33376 14958
rect 33324 14894 33376 14900
rect 33048 14408 33100 14414
rect 33048 14350 33100 14356
rect 32956 13728 33008 13734
rect 32956 13670 33008 13676
rect 32864 12844 32916 12850
rect 32864 12786 32916 12792
rect 32680 12368 32732 12374
rect 32680 12310 32732 12316
rect 32956 12300 33008 12306
rect 32956 12242 33008 12248
rect 32864 11688 32916 11694
rect 32864 11630 32916 11636
rect 32876 10130 32904 11630
rect 32968 11082 32996 12242
rect 33060 12170 33088 14350
rect 33336 14278 33364 14894
rect 33232 14272 33284 14278
rect 33232 14214 33284 14220
rect 33324 14272 33376 14278
rect 33324 14214 33376 14220
rect 33244 13938 33272 14214
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 33244 13002 33272 13874
rect 33336 13190 33364 14214
rect 33520 13938 33548 14962
rect 33508 13932 33560 13938
rect 33508 13874 33560 13880
rect 33324 13184 33376 13190
rect 33324 13126 33376 13132
rect 33244 12974 33364 13002
rect 33336 12850 33364 12974
rect 33520 12850 33548 13874
rect 33324 12844 33376 12850
rect 33324 12786 33376 12792
rect 33508 12844 33560 12850
rect 33508 12786 33560 12792
rect 33140 12708 33192 12714
rect 33140 12650 33192 12656
rect 33048 12164 33100 12170
rect 33048 12106 33100 12112
rect 33060 11558 33088 12106
rect 33152 11762 33180 12650
rect 33336 12238 33364 12786
rect 33520 12306 33548 12786
rect 33508 12300 33560 12306
rect 33508 12242 33560 12248
rect 33324 12232 33376 12238
rect 33324 12174 33376 12180
rect 33612 11762 33640 15302
rect 33796 15162 33824 15422
rect 33876 15360 33928 15366
rect 33876 15302 33928 15308
rect 33784 15156 33836 15162
rect 33784 15098 33836 15104
rect 33888 15094 33916 15302
rect 33876 15088 33928 15094
rect 33876 15030 33928 15036
rect 33784 14612 33836 14618
rect 33784 14554 33836 14560
rect 33692 12844 33744 12850
rect 33692 12786 33744 12792
rect 33140 11756 33192 11762
rect 33140 11698 33192 11704
rect 33600 11756 33652 11762
rect 33600 11698 33652 11704
rect 33048 11552 33100 11558
rect 33048 11494 33100 11500
rect 33152 11354 33180 11698
rect 33140 11348 33192 11354
rect 33140 11290 33192 11296
rect 32956 11076 33008 11082
rect 32956 11018 33008 11024
rect 32968 10130 32996 11018
rect 33704 10810 33732 12786
rect 33796 11762 33824 14554
rect 33980 14346 34008 16594
rect 34152 16584 34204 16590
rect 34152 16526 34204 16532
rect 34164 14346 34192 16526
rect 33968 14340 34020 14346
rect 33968 14282 34020 14288
rect 34152 14340 34204 14346
rect 34152 14282 34204 14288
rect 33968 14068 34020 14074
rect 33968 14010 34020 14016
rect 33980 13802 34008 14010
rect 33968 13796 34020 13802
rect 33968 13738 34020 13744
rect 33980 13190 34008 13738
rect 34256 13462 34284 17054
rect 34440 16572 34468 20198
rect 34532 19378 34560 21490
rect 34704 21480 34756 21486
rect 34704 21422 34756 21428
rect 34612 21004 34664 21010
rect 34612 20946 34664 20952
rect 34624 19802 34652 20946
rect 34716 20058 34744 21422
rect 34704 20052 34756 20058
rect 34704 19994 34756 20000
rect 34808 19854 34836 21966
rect 34900 21554 34928 22102
rect 35072 22024 35124 22030
rect 35070 21992 35072 22001
rect 35124 21992 35126 22001
rect 35070 21927 35126 21936
rect 35256 21956 35308 21962
rect 35256 21898 35308 21904
rect 35268 21622 35296 21898
rect 35256 21616 35308 21622
rect 35256 21558 35308 21564
rect 35360 21554 35388 22188
rect 35438 22128 35494 22137
rect 35544 22098 35572 22646
rect 35636 22574 35664 24278
rect 35820 24206 35848 24550
rect 35808 24200 35860 24206
rect 35912 24188 35940 25180
rect 36004 24954 36032 27542
rect 36084 27396 36136 27402
rect 36084 27338 36136 27344
rect 36096 25809 36124 27338
rect 36174 27160 36230 27169
rect 36174 27095 36230 27104
rect 36188 26382 36216 27095
rect 36280 26382 36308 29951
rect 36372 29714 36400 29990
rect 36464 29850 36492 31726
rect 36648 31346 36676 32846
rect 36728 32292 36780 32298
rect 36728 32234 36780 32240
rect 36740 32065 36768 32234
rect 36726 32056 36782 32065
rect 36726 31991 36782 32000
rect 36832 31906 36860 34002
rect 37016 33810 37044 35634
rect 37096 34740 37148 34746
rect 37096 34682 37148 34688
rect 37108 33998 37136 34682
rect 37200 34678 37228 35974
rect 37384 35698 37412 37062
rect 37462 37023 37518 37032
rect 37476 35714 37504 37023
rect 37568 35834 37596 37130
rect 38028 36718 38056 37130
rect 38016 36712 38068 36718
rect 38016 36654 38068 36660
rect 38106 36680 38162 36689
rect 38106 36615 38162 36624
rect 38120 36310 38148 36615
rect 38108 36304 38160 36310
rect 38108 36246 38160 36252
rect 37556 35828 37608 35834
rect 37556 35770 37608 35776
rect 37372 35692 37424 35698
rect 37476 35686 37596 35714
rect 37372 35634 37424 35640
rect 37280 35284 37332 35290
rect 37280 35226 37332 35232
rect 37188 34672 37240 34678
rect 37188 34614 37240 34620
rect 37188 34468 37240 34474
rect 37188 34410 37240 34416
rect 37096 33992 37148 33998
rect 37096 33934 37148 33940
rect 37016 33782 37136 33810
rect 36912 33448 36964 33454
rect 36912 33390 36964 33396
rect 36924 32745 36952 33390
rect 36910 32736 36966 32745
rect 36910 32671 36966 32680
rect 37004 32020 37056 32026
rect 36740 31890 36860 31906
rect 36924 31980 37004 32008
rect 36740 31884 36872 31890
rect 36740 31878 36820 31884
rect 36636 31340 36688 31346
rect 36556 31300 36636 31328
rect 36556 30734 36584 31300
rect 36636 31282 36688 31288
rect 36636 31204 36688 31210
rect 36636 31146 36688 31152
rect 36648 30734 36676 31146
rect 36544 30728 36596 30734
rect 36544 30670 36596 30676
rect 36636 30728 36688 30734
rect 36636 30670 36688 30676
rect 36452 29844 36504 29850
rect 36452 29786 36504 29792
rect 36360 29708 36412 29714
rect 36360 29650 36412 29656
rect 36556 29646 36584 30670
rect 36740 30326 36768 31878
rect 36820 31826 36872 31832
rect 36820 31680 36872 31686
rect 36820 31622 36872 31628
rect 36832 31346 36860 31622
rect 36820 31340 36872 31346
rect 36820 31282 36872 31288
rect 36820 31136 36872 31142
rect 36820 31078 36872 31084
rect 36832 30870 36860 31078
rect 36820 30864 36872 30870
rect 36820 30806 36872 30812
rect 36820 30728 36872 30734
rect 36820 30670 36872 30676
rect 36728 30320 36780 30326
rect 36728 30262 36780 30268
rect 36544 29640 36596 29646
rect 36358 29608 36414 29617
rect 36544 29582 36596 29588
rect 36636 29640 36688 29646
rect 36636 29582 36688 29588
rect 36358 29543 36414 29552
rect 36372 29510 36400 29543
rect 36360 29504 36412 29510
rect 36360 29446 36412 29452
rect 36544 29504 36596 29510
rect 36544 29446 36596 29452
rect 36372 29306 36400 29446
rect 36360 29300 36412 29306
rect 36360 29242 36412 29248
rect 36452 29232 36504 29238
rect 36452 29174 36504 29180
rect 36358 27160 36414 27169
rect 36358 27095 36414 27104
rect 36372 27062 36400 27095
rect 36360 27056 36412 27062
rect 36360 26998 36412 27004
rect 36360 26920 36412 26926
rect 36360 26862 36412 26868
rect 36176 26376 36228 26382
rect 36176 26318 36228 26324
rect 36268 26376 36320 26382
rect 36268 26318 36320 26324
rect 36372 26042 36400 26862
rect 36464 26586 36492 29174
rect 36452 26580 36504 26586
rect 36452 26522 36504 26528
rect 36556 26450 36584 29446
rect 36648 27470 36676 29582
rect 36740 27470 36768 30262
rect 36636 27464 36688 27470
rect 36636 27406 36688 27412
rect 36728 27464 36780 27470
rect 36728 27406 36780 27412
rect 36636 27328 36688 27334
rect 36636 27270 36688 27276
rect 36648 27033 36676 27270
rect 36634 27024 36690 27033
rect 36634 26959 36690 26968
rect 36636 26852 36688 26858
rect 36636 26794 36688 26800
rect 36544 26444 36596 26450
rect 36544 26386 36596 26392
rect 36360 26036 36412 26042
rect 36360 25978 36412 25984
rect 36082 25800 36138 25809
rect 36082 25735 36138 25744
rect 36648 25498 36676 26794
rect 36740 25702 36768 27406
rect 36832 26314 36860 30670
rect 36924 29646 36952 31980
rect 37004 31962 37056 31968
rect 37108 31754 37136 33782
rect 37016 31726 37136 31754
rect 36912 29640 36964 29646
rect 36912 29582 36964 29588
rect 36912 26376 36964 26382
rect 36912 26318 36964 26324
rect 36820 26308 36872 26314
rect 36820 26250 36872 26256
rect 36924 25974 36952 26318
rect 36912 25968 36964 25974
rect 36912 25910 36964 25916
rect 36728 25696 36780 25702
rect 36728 25638 36780 25644
rect 36820 25696 36872 25702
rect 36820 25638 36872 25644
rect 36084 25492 36136 25498
rect 36084 25434 36136 25440
rect 36636 25492 36688 25498
rect 36636 25434 36688 25440
rect 36728 25492 36780 25498
rect 36728 25434 36780 25440
rect 36096 25294 36124 25434
rect 36084 25288 36136 25294
rect 36084 25230 36136 25236
rect 36176 25288 36228 25294
rect 36176 25230 36228 25236
rect 36082 25120 36138 25129
rect 36082 25055 36138 25064
rect 35992 24948 36044 24954
rect 35992 24890 36044 24896
rect 35992 24812 36044 24818
rect 36096 24800 36124 25055
rect 36044 24772 36124 24800
rect 35992 24754 36044 24760
rect 35992 24200 36044 24206
rect 35912 24160 35992 24188
rect 35808 24142 35860 24148
rect 35992 24142 36044 24148
rect 36188 23905 36216 25230
rect 36268 24812 36320 24818
rect 36268 24754 36320 24760
rect 36280 24410 36308 24754
rect 36452 24744 36504 24750
rect 36452 24686 36504 24692
rect 36268 24404 36320 24410
rect 36268 24346 36320 24352
rect 36268 24200 36320 24206
rect 36268 24142 36320 24148
rect 36174 23896 36230 23905
rect 36174 23831 36230 23840
rect 35716 23792 35768 23798
rect 35716 23734 35768 23740
rect 35728 23050 35756 23734
rect 35900 23724 35952 23730
rect 35900 23666 35952 23672
rect 35912 23322 35940 23666
rect 35992 23656 36044 23662
rect 35992 23598 36044 23604
rect 35900 23316 35952 23322
rect 35900 23258 35952 23264
rect 35808 23112 35860 23118
rect 35808 23054 35860 23060
rect 35716 23044 35768 23050
rect 35716 22986 35768 22992
rect 35716 22636 35768 22642
rect 35716 22578 35768 22584
rect 35624 22568 35676 22574
rect 35624 22510 35676 22516
rect 35622 22400 35678 22409
rect 35622 22335 35678 22344
rect 35636 22234 35664 22335
rect 35624 22228 35676 22234
rect 35624 22170 35676 22176
rect 35438 22063 35494 22072
rect 35532 22092 35584 22098
rect 35452 21622 35480 22063
rect 35584 22052 35664 22080
rect 35532 22034 35584 22040
rect 35440 21616 35492 21622
rect 35440 21558 35492 21564
rect 34888 21548 34940 21554
rect 34888 21490 34940 21496
rect 35348 21548 35400 21554
rect 35348 21490 35400 21496
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35256 20936 35308 20942
rect 35256 20878 35308 20884
rect 34978 20496 35034 20505
rect 34978 20431 34980 20440
rect 35032 20431 35034 20440
rect 34980 20402 35032 20408
rect 35268 20398 35296 20878
rect 35256 20392 35308 20398
rect 35256 20334 35308 20340
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34980 20052 35032 20058
rect 34980 19994 35032 20000
rect 35256 20052 35308 20058
rect 35256 19994 35308 20000
rect 34796 19848 34848 19854
rect 34624 19774 34744 19802
rect 34796 19790 34848 19796
rect 34610 19544 34666 19553
rect 34610 19479 34666 19488
rect 34624 19446 34652 19479
rect 34612 19440 34664 19446
rect 34612 19382 34664 19388
rect 34520 19372 34572 19378
rect 34520 19314 34572 19320
rect 34532 18766 34560 19314
rect 34520 18760 34572 18766
rect 34520 18702 34572 18708
rect 34716 18170 34744 19774
rect 34808 19242 34836 19790
rect 34888 19712 34940 19718
rect 34888 19654 34940 19660
rect 34900 19378 34928 19654
rect 34992 19417 35020 19994
rect 35268 19854 35296 19994
rect 35072 19848 35124 19854
rect 35070 19816 35072 19825
rect 35256 19848 35308 19854
rect 35124 19816 35126 19825
rect 35256 19790 35308 19796
rect 35070 19751 35126 19760
rect 35268 19530 35296 19790
rect 35084 19502 35296 19530
rect 34978 19408 35034 19417
rect 34888 19372 34940 19378
rect 34978 19343 34981 19352
rect 34888 19314 34940 19320
rect 35033 19343 35034 19352
rect 34981 19314 35033 19320
rect 35084 19334 35112 19502
rect 35254 19408 35310 19417
rect 35360 19378 35388 21490
rect 35532 21004 35584 21010
rect 35452 20964 35532 20992
rect 35254 19343 35310 19352
rect 35348 19372 35400 19378
rect 34796 19236 34848 19242
rect 34796 19178 34848 19184
rect 34808 18290 34836 19178
rect 34992 19174 35020 19314
rect 35084 19306 35204 19334
rect 35176 19174 35204 19306
rect 34980 19168 35032 19174
rect 34980 19110 35032 19116
rect 35164 19168 35216 19174
rect 35164 19110 35216 19116
rect 35268 19122 35296 19343
rect 35348 19314 35400 19320
rect 35268 19094 35301 19122
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35273 18986 35301 19094
rect 35072 18964 35124 18970
rect 35072 18906 35124 18912
rect 35268 18958 35301 18986
rect 34980 18760 35032 18766
rect 34980 18702 35032 18708
rect 34992 18358 35020 18702
rect 34980 18352 35032 18358
rect 34980 18294 35032 18300
rect 35084 18290 35112 18906
rect 35164 18760 35216 18766
rect 35268 18748 35296 18958
rect 35360 18766 35388 19314
rect 35216 18720 35296 18748
rect 35348 18760 35400 18766
rect 35164 18702 35216 18708
rect 35348 18702 35400 18708
rect 35348 18624 35400 18630
rect 35348 18566 35400 18572
rect 35256 18420 35308 18426
rect 35256 18362 35308 18368
rect 35268 18290 35296 18362
rect 35360 18358 35388 18566
rect 35348 18352 35400 18358
rect 35348 18294 35400 18300
rect 34796 18284 34848 18290
rect 34796 18226 34848 18232
rect 35072 18284 35124 18290
rect 35072 18226 35124 18232
rect 35256 18284 35308 18290
rect 35256 18226 35308 18232
rect 35254 18184 35310 18193
rect 34612 18148 34664 18154
rect 34716 18142 34836 18170
rect 34612 18090 34664 18096
rect 34520 18080 34572 18086
rect 34520 18022 34572 18028
rect 34532 17202 34560 18022
rect 34624 17202 34652 18090
rect 34704 17740 34756 17746
rect 34704 17682 34756 17688
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34612 17196 34664 17202
rect 34612 17138 34664 17144
rect 34610 16960 34666 16969
rect 34610 16895 34666 16904
rect 34440 16544 34560 16572
rect 34336 16448 34388 16454
rect 34336 16390 34388 16396
rect 34244 13456 34296 13462
rect 34244 13398 34296 13404
rect 33968 13184 34020 13190
rect 33968 13126 34020 13132
rect 33784 11756 33836 11762
rect 33784 11698 33836 11704
rect 33692 10804 33744 10810
rect 33692 10746 33744 10752
rect 32864 10124 32916 10130
rect 32864 10066 32916 10072
rect 32956 10124 33008 10130
rect 32956 10066 33008 10072
rect 33704 10062 33732 10746
rect 34348 10062 34376 16390
rect 34532 16250 34560 16544
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 34624 15162 34652 16895
rect 34716 16114 34744 17682
rect 34808 16794 34836 18142
rect 35254 18119 35310 18128
rect 35268 18034 35296 18119
rect 35348 18080 35400 18086
rect 35268 18006 35301 18034
rect 35348 18022 35400 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35273 17898 35301 18006
rect 35268 17870 35301 17898
rect 35360 17882 35388 18022
rect 35348 17876 35400 17882
rect 35164 17672 35216 17678
rect 35164 17614 35216 17620
rect 35176 17338 35204 17614
rect 35164 17332 35216 17338
rect 35164 17274 35216 17280
rect 35268 16946 35296 17870
rect 35348 17818 35400 17824
rect 35360 17066 35388 17818
rect 35348 17060 35400 17066
rect 35348 17002 35400 17008
rect 35268 16918 35388 16946
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 35256 16652 35308 16658
rect 35256 16594 35308 16600
rect 34796 16516 34848 16522
rect 34796 16458 34848 16464
rect 34704 16108 34756 16114
rect 34704 16050 34756 16056
rect 34808 16046 34836 16458
rect 35268 16182 35296 16594
rect 35256 16176 35308 16182
rect 35256 16118 35308 16124
rect 34796 16040 34848 16046
rect 34796 15982 34848 15988
rect 34704 15496 34756 15502
rect 34704 15438 34756 15444
rect 34612 15156 34664 15162
rect 34612 15098 34664 15104
rect 34520 14000 34572 14006
rect 34520 13942 34572 13948
rect 34532 13530 34560 13942
rect 34716 13938 34744 15438
rect 34808 14414 34836 15982
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34796 14408 34848 14414
rect 34796 14350 34848 14356
rect 35360 14362 35388 16918
rect 35452 15366 35480 20964
rect 35532 20946 35584 20952
rect 35636 20584 35664 22052
rect 35728 20874 35756 22578
rect 35820 22030 35848 23054
rect 35900 22568 35952 22574
rect 35900 22510 35952 22516
rect 35808 22024 35860 22030
rect 35808 21966 35860 21972
rect 35716 20868 35768 20874
rect 35716 20810 35768 20816
rect 35820 20602 35848 21966
rect 35544 20556 35664 20584
rect 35808 20596 35860 20602
rect 35544 20058 35572 20556
rect 35808 20538 35860 20544
rect 35624 20460 35676 20466
rect 35624 20402 35676 20408
rect 35532 20052 35584 20058
rect 35532 19994 35584 20000
rect 35636 19990 35664 20402
rect 35716 20392 35768 20398
rect 35716 20334 35768 20340
rect 35624 19984 35676 19990
rect 35624 19926 35676 19932
rect 35532 19848 35584 19854
rect 35532 19790 35584 19796
rect 35544 18426 35572 19790
rect 35624 19168 35676 19174
rect 35624 19110 35676 19116
rect 35636 18970 35664 19110
rect 35624 18964 35676 18970
rect 35624 18906 35676 18912
rect 35622 18728 35678 18737
rect 35622 18663 35678 18672
rect 35532 18420 35584 18426
rect 35532 18362 35584 18368
rect 35530 15464 35586 15473
rect 35530 15399 35586 15408
rect 35440 15360 35492 15366
rect 35440 15302 35492 15308
rect 35360 14334 35480 14362
rect 34796 14272 34848 14278
rect 34796 14214 34848 14220
rect 35348 14272 35400 14278
rect 35348 14214 35400 14220
rect 34704 13932 34756 13938
rect 34704 13874 34756 13880
rect 34808 13530 34836 14214
rect 35360 13938 35388 14214
rect 35348 13932 35400 13938
rect 35348 13874 35400 13880
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34520 13524 34572 13530
rect 34520 13466 34572 13472
rect 34796 13524 34848 13530
rect 34796 13466 34848 13472
rect 35164 13388 35216 13394
rect 35164 13330 35216 13336
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 34520 12776 34572 12782
rect 34520 12718 34572 12724
rect 34532 12102 34560 12718
rect 34612 12640 34664 12646
rect 34612 12582 34664 12588
rect 34624 12306 34652 12582
rect 34808 12442 34836 12786
rect 35176 12782 35204 13330
rect 35360 13190 35388 13874
rect 35452 13512 35480 14334
rect 35544 13938 35572 15399
rect 35532 13932 35584 13938
rect 35532 13874 35584 13880
rect 35452 13484 35572 13512
rect 35440 13388 35492 13394
rect 35440 13330 35492 13336
rect 35348 13184 35400 13190
rect 35348 13126 35400 13132
rect 35164 12776 35216 12782
rect 35164 12718 35216 12724
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34796 12436 34848 12442
rect 34796 12378 34848 12384
rect 34612 12300 34664 12306
rect 34612 12242 34664 12248
rect 34796 12232 34848 12238
rect 34796 12174 34848 12180
rect 34520 12096 34572 12102
rect 34520 12038 34572 12044
rect 34532 11082 34560 12038
rect 34808 11898 34836 12174
rect 34796 11892 34848 11898
rect 34796 11834 34848 11840
rect 35348 11892 35400 11898
rect 35348 11834 35400 11840
rect 34796 11756 34848 11762
rect 34796 11698 34848 11704
rect 34808 11354 34836 11698
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11348 34848 11354
rect 34796 11290 34848 11296
rect 35360 11150 35388 11834
rect 35452 11218 35480 13330
rect 35544 12782 35572 13484
rect 35636 12986 35664 18663
rect 35728 15434 35756 20334
rect 35820 19854 35848 20538
rect 35808 19848 35860 19854
rect 35808 19790 35860 19796
rect 35806 19408 35862 19417
rect 35806 19343 35808 19352
rect 35860 19343 35862 19352
rect 35808 19314 35860 19320
rect 35806 18592 35862 18601
rect 35806 18527 35862 18536
rect 35820 18358 35848 18527
rect 35808 18352 35860 18358
rect 35808 18294 35860 18300
rect 35806 16824 35862 16833
rect 35806 16759 35862 16768
rect 35820 16590 35848 16759
rect 35808 16584 35860 16590
rect 35808 16526 35860 16532
rect 35716 15428 35768 15434
rect 35716 15370 35768 15376
rect 35728 14634 35756 15370
rect 35912 15094 35940 22510
rect 36004 22030 36032 23598
rect 36280 23594 36308 24142
rect 36464 24138 36492 24686
rect 36740 24342 36768 25434
rect 36832 25158 36860 25638
rect 36924 25362 36952 25910
rect 36912 25356 36964 25362
rect 36912 25298 36964 25304
rect 36820 25152 36872 25158
rect 36820 25094 36872 25100
rect 36728 24336 36780 24342
rect 36728 24278 36780 24284
rect 36452 24132 36504 24138
rect 36452 24074 36504 24080
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 36268 23588 36320 23594
rect 36268 23530 36320 23536
rect 36084 23520 36136 23526
rect 36084 23462 36136 23468
rect 35992 22024 36044 22030
rect 35992 21966 36044 21972
rect 36096 21622 36124 23462
rect 36176 22432 36228 22438
rect 36176 22374 36228 22380
rect 36084 21616 36136 21622
rect 36084 21558 36136 21564
rect 35992 20460 36044 20466
rect 35992 20402 36044 20408
rect 36004 20369 36032 20402
rect 36084 20392 36136 20398
rect 35990 20360 36046 20369
rect 36188 20380 36216 22374
rect 36280 20602 36308 23530
rect 36372 22778 36400 23666
rect 36360 22772 36412 22778
rect 36360 22714 36412 22720
rect 36464 21554 36492 24074
rect 36636 24064 36688 24070
rect 36636 24006 36688 24012
rect 36648 23730 36676 24006
rect 36636 23724 36688 23730
rect 36636 23666 36688 23672
rect 36740 23594 36768 24278
rect 36924 24274 36952 25298
rect 37016 25226 37044 31726
rect 37200 31686 37228 34410
rect 37188 31680 37240 31686
rect 37188 31622 37240 31628
rect 37096 30796 37148 30802
rect 37096 30738 37148 30744
rect 37108 29481 37136 30738
rect 37188 30728 37240 30734
rect 37186 30696 37188 30705
rect 37240 30696 37242 30705
rect 37186 30631 37242 30640
rect 37186 29744 37242 29753
rect 37186 29679 37242 29688
rect 37094 29472 37150 29481
rect 37094 29407 37150 29416
rect 37200 29238 37228 29679
rect 37188 29232 37240 29238
rect 37188 29174 37240 29180
rect 37096 27124 37148 27130
rect 37096 27066 37148 27072
rect 37004 25220 37056 25226
rect 37004 25162 37056 25168
rect 36912 24268 36964 24274
rect 36912 24210 36964 24216
rect 36544 23588 36596 23594
rect 36544 23530 36596 23536
rect 36728 23588 36780 23594
rect 36728 23530 36780 23536
rect 36556 22438 36584 23530
rect 36924 23118 36952 24210
rect 36912 23112 36964 23118
rect 37004 23112 37056 23118
rect 36912 23054 36964 23060
rect 37002 23080 37004 23089
rect 37056 23080 37058 23089
rect 36728 23044 36780 23050
rect 36728 22986 36780 22992
rect 36740 22574 36768 22986
rect 36818 22808 36874 22817
rect 36818 22743 36874 22752
rect 36728 22568 36780 22574
rect 36728 22510 36780 22516
rect 36544 22432 36596 22438
rect 36544 22374 36596 22380
rect 36634 21584 36690 21593
rect 36452 21548 36504 21554
rect 36634 21519 36690 21528
rect 36452 21490 36504 21496
rect 36360 20936 36412 20942
rect 36412 20884 36584 20890
rect 36360 20878 36584 20884
rect 36372 20862 36584 20878
rect 36268 20596 36320 20602
rect 36268 20538 36320 20544
rect 36452 20460 36504 20466
rect 36452 20402 36504 20408
rect 36136 20352 36216 20380
rect 36084 20334 36136 20340
rect 35990 20295 36046 20304
rect 35992 19848 36044 19854
rect 35992 19790 36044 19796
rect 36004 15162 36032 19790
rect 36096 18086 36124 20334
rect 36176 20256 36228 20262
rect 36176 20198 36228 20204
rect 36188 19854 36216 20198
rect 36360 19916 36412 19922
rect 36360 19858 36412 19864
rect 36176 19848 36228 19854
rect 36176 19790 36228 19796
rect 36084 18080 36136 18086
rect 36084 18022 36136 18028
rect 36084 17672 36136 17678
rect 36084 17614 36136 17620
rect 35992 15156 36044 15162
rect 35992 15098 36044 15104
rect 35900 15088 35952 15094
rect 35900 15030 35952 15036
rect 35992 14952 36044 14958
rect 35992 14894 36044 14900
rect 35728 14618 35848 14634
rect 35728 14612 35860 14618
rect 35728 14606 35808 14612
rect 35808 14554 35860 14560
rect 36004 13326 36032 14894
rect 36096 14414 36124 17614
rect 36188 15026 36216 19790
rect 36372 19446 36400 19858
rect 36360 19440 36412 19446
rect 36360 19382 36412 19388
rect 36464 18970 36492 20402
rect 36556 19854 36584 20862
rect 36544 19848 36596 19854
rect 36544 19790 36596 19796
rect 36452 18964 36504 18970
rect 36452 18906 36504 18912
rect 36268 18828 36320 18834
rect 36268 18770 36320 18776
rect 36280 18290 36308 18770
rect 36556 18766 36584 19790
rect 36648 19718 36676 21519
rect 36636 19712 36688 19718
rect 36636 19654 36688 19660
rect 36726 19680 36782 19689
rect 36544 18760 36596 18766
rect 36544 18702 36596 18708
rect 36452 18692 36504 18698
rect 36452 18634 36504 18640
rect 36268 18284 36320 18290
rect 36268 18226 36320 18232
rect 36280 17082 36308 18226
rect 36360 18216 36412 18222
rect 36360 18158 36412 18164
rect 36372 17202 36400 18158
rect 36464 17882 36492 18634
rect 36452 17876 36504 17882
rect 36452 17818 36504 17824
rect 36556 17678 36584 18702
rect 36544 17672 36596 17678
rect 36544 17614 36596 17620
rect 36360 17196 36412 17202
rect 36360 17138 36412 17144
rect 36280 17054 36400 17082
rect 36266 16688 36322 16697
rect 36266 16623 36322 16632
rect 36280 16454 36308 16623
rect 36268 16448 36320 16454
rect 36268 16390 36320 16396
rect 36372 16250 36400 17054
rect 36360 16244 36412 16250
rect 36360 16186 36412 16192
rect 36360 16108 36412 16114
rect 36360 16050 36412 16056
rect 36268 15360 36320 15366
rect 36268 15302 36320 15308
rect 36280 15094 36308 15302
rect 36268 15088 36320 15094
rect 36268 15030 36320 15036
rect 36372 15026 36400 16050
rect 36176 15020 36228 15026
rect 36176 14962 36228 14968
rect 36360 15020 36412 15026
rect 36360 14962 36412 14968
rect 36360 14816 36412 14822
rect 36360 14758 36412 14764
rect 36084 14408 36136 14414
rect 36084 14350 36136 14356
rect 36268 13728 36320 13734
rect 36268 13670 36320 13676
rect 36084 13456 36136 13462
rect 36082 13424 36084 13433
rect 36136 13424 36138 13433
rect 36082 13359 36138 13368
rect 36280 13326 36308 13670
rect 35992 13320 36044 13326
rect 35992 13262 36044 13268
rect 36268 13320 36320 13326
rect 36268 13262 36320 13268
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 36372 12850 36400 14758
rect 36648 12850 36676 19654
rect 36726 19615 36782 19624
rect 36740 19378 36768 19615
rect 36728 19372 36780 19378
rect 36728 19314 36780 19320
rect 36832 19310 36860 22743
rect 36924 22098 36952 23054
rect 37002 23015 37058 23024
rect 37004 22636 37056 22642
rect 37004 22578 37056 22584
rect 36912 22092 36964 22098
rect 36912 22034 36964 22040
rect 36820 19304 36872 19310
rect 36820 19246 36872 19252
rect 36728 17740 36780 17746
rect 36728 17682 36780 17688
rect 36740 14346 36768 17682
rect 36820 17672 36872 17678
rect 36820 17614 36872 17620
rect 36832 16658 36860 17614
rect 37016 17218 37044 22578
rect 36924 17190 37044 17218
rect 36820 16652 36872 16658
rect 36820 16594 36872 16600
rect 36818 15328 36874 15337
rect 36818 15263 36874 15272
rect 36728 14340 36780 14346
rect 36728 14282 36780 14288
rect 36832 14074 36860 15263
rect 36924 15094 36952 17190
rect 37108 17116 37136 27066
rect 37188 25220 37240 25226
rect 37188 25162 37240 25168
rect 37200 24682 37228 25162
rect 37188 24676 37240 24682
rect 37188 24618 37240 24624
rect 37292 23633 37320 35226
rect 37384 35086 37412 35634
rect 37372 35080 37424 35086
rect 37372 35022 37424 35028
rect 37464 35080 37516 35086
rect 37464 35022 37516 35028
rect 37372 34944 37424 34950
rect 37372 34886 37424 34892
rect 37384 33590 37412 34886
rect 37476 34406 37504 35022
rect 37464 34400 37516 34406
rect 37464 34342 37516 34348
rect 37372 33584 37424 33590
rect 37372 33526 37424 33532
rect 37372 33312 37424 33318
rect 37372 33254 37424 33260
rect 37384 31142 37412 33254
rect 37464 32836 37516 32842
rect 37464 32778 37516 32784
rect 37476 32570 37504 32778
rect 37464 32564 37516 32570
rect 37464 32506 37516 32512
rect 37464 31816 37516 31822
rect 37464 31758 37516 31764
rect 37476 31482 37504 31758
rect 37464 31476 37516 31482
rect 37464 31418 37516 31424
rect 37372 31136 37424 31142
rect 37372 31078 37424 31084
rect 37568 30938 37596 35686
rect 38108 35624 38160 35630
rect 38108 35566 38160 35572
rect 37740 35216 37792 35222
rect 37740 35158 37792 35164
rect 37648 35012 37700 35018
rect 37648 34954 37700 34960
rect 37660 33561 37688 34954
rect 37646 33552 37702 33561
rect 37646 33487 37648 33496
rect 37700 33487 37702 33496
rect 37648 33458 37700 33464
rect 37556 30932 37608 30938
rect 37556 30874 37608 30880
rect 37372 30796 37424 30802
rect 37372 30738 37424 30744
rect 37384 28150 37412 30738
rect 37568 30326 37596 30874
rect 37648 30592 37700 30598
rect 37648 30534 37700 30540
rect 37556 30320 37608 30326
rect 37556 30262 37608 30268
rect 37464 30048 37516 30054
rect 37464 29990 37516 29996
rect 37476 29646 37504 29990
rect 37464 29640 37516 29646
rect 37464 29582 37516 29588
rect 37556 29572 37608 29578
rect 37556 29514 37608 29520
rect 37464 28960 37516 28966
rect 37464 28902 37516 28908
rect 37476 28558 37504 28902
rect 37464 28552 37516 28558
rect 37464 28494 37516 28500
rect 37372 28144 37424 28150
rect 37372 28086 37424 28092
rect 37462 28112 37518 28121
rect 37462 28047 37464 28056
rect 37516 28047 37518 28056
rect 37464 28018 37516 28024
rect 37464 27396 37516 27402
rect 37464 27338 37516 27344
rect 37476 27130 37504 27338
rect 37464 27124 37516 27130
rect 37464 27066 37516 27072
rect 37464 26308 37516 26314
rect 37464 26250 37516 26256
rect 37370 26072 37426 26081
rect 37476 26042 37504 26250
rect 37370 26007 37426 26016
rect 37464 26036 37516 26042
rect 37384 25974 37412 26007
rect 37464 25978 37516 25984
rect 37372 25968 37424 25974
rect 37372 25910 37424 25916
rect 37568 25106 37596 29514
rect 37660 25294 37688 30534
rect 37752 27130 37780 35158
rect 37924 35080 37976 35086
rect 37924 35022 37976 35028
rect 37832 34604 37884 34610
rect 37832 34546 37884 34552
rect 37844 33930 37872 34546
rect 37832 33924 37884 33930
rect 37832 33866 37884 33872
rect 37936 33522 37964 35022
rect 38120 34542 38148 35566
rect 38384 35148 38436 35154
rect 38384 35090 38436 35096
rect 38108 34536 38160 34542
rect 38108 34478 38160 34484
rect 37924 33516 37976 33522
rect 37924 33458 37976 33464
rect 37936 33289 37964 33458
rect 38016 33312 38068 33318
rect 37922 33280 37978 33289
rect 38016 33254 38068 33260
rect 37922 33215 37978 33224
rect 37830 33008 37886 33017
rect 37830 32943 37886 32952
rect 37844 32774 37872 32943
rect 37832 32768 37884 32774
rect 37832 32710 37884 32716
rect 37844 32570 37872 32710
rect 37832 32564 37884 32570
rect 37832 32506 37884 32512
rect 37936 32298 37964 33215
rect 38028 33114 38056 33254
rect 38016 33108 38068 33114
rect 38016 33050 38068 33056
rect 38014 32600 38070 32609
rect 38014 32535 38070 32544
rect 38028 32366 38056 32535
rect 38016 32360 38068 32366
rect 38120 32348 38148 34478
rect 38292 34196 38344 34202
rect 38292 34138 38344 34144
rect 38198 34096 38254 34105
rect 38198 34031 38254 34040
rect 38068 32320 38148 32348
rect 38016 32302 38068 32308
rect 37924 32292 37976 32298
rect 37924 32234 37976 32240
rect 38016 31748 38068 31754
rect 38016 31690 38068 31696
rect 37832 31680 37884 31686
rect 37832 31622 37884 31628
rect 37844 31414 37872 31622
rect 37832 31408 37884 31414
rect 37832 31350 37884 31356
rect 37924 31136 37976 31142
rect 37924 31078 37976 31084
rect 37936 29186 37964 31078
rect 38028 30598 38056 31690
rect 38120 31278 38148 32320
rect 38108 31272 38160 31278
rect 38108 31214 38160 31220
rect 38016 30592 38068 30598
rect 38016 30534 38068 30540
rect 37844 29158 37964 29186
rect 37844 28937 37872 29158
rect 37924 29096 37976 29102
rect 37924 29038 37976 29044
rect 37830 28928 37886 28937
rect 37830 28863 37886 28872
rect 37740 27124 37792 27130
rect 37740 27066 37792 27072
rect 37740 26240 37792 26246
rect 37740 26182 37792 26188
rect 37752 25974 37780 26182
rect 37740 25968 37792 25974
rect 37740 25910 37792 25916
rect 37648 25288 37700 25294
rect 37648 25230 37700 25236
rect 37832 25152 37884 25158
rect 37568 25078 37780 25106
rect 37832 25094 37884 25100
rect 37556 24948 37608 24954
rect 37556 24890 37608 24896
rect 37372 24608 37424 24614
rect 37372 24550 37424 24556
rect 37278 23624 37334 23633
rect 37278 23559 37334 23568
rect 37188 21956 37240 21962
rect 37188 21898 37240 21904
rect 37200 21690 37228 21898
rect 37188 21684 37240 21690
rect 37188 21626 37240 21632
rect 37280 21140 37332 21146
rect 37280 21082 37332 21088
rect 37016 17088 37136 17116
rect 37016 16794 37044 17088
rect 37096 16992 37148 16998
rect 37096 16934 37148 16940
rect 37004 16788 37056 16794
rect 37004 16730 37056 16736
rect 37108 16590 37136 16934
rect 37096 16584 37148 16590
rect 37096 16526 37148 16532
rect 36912 15088 36964 15094
rect 36912 15030 36964 15036
rect 36820 14068 36872 14074
rect 36820 14010 36872 14016
rect 36832 13802 36860 14010
rect 36820 13796 36872 13802
rect 36820 13738 36872 13744
rect 37292 13530 37320 21082
rect 37384 20534 37412 24550
rect 37464 24132 37516 24138
rect 37464 24074 37516 24080
rect 37476 23866 37504 24074
rect 37464 23860 37516 23866
rect 37464 23802 37516 23808
rect 37464 23724 37516 23730
rect 37464 23666 37516 23672
rect 37476 23322 37504 23666
rect 37464 23316 37516 23322
rect 37464 23258 37516 23264
rect 37462 23216 37518 23225
rect 37462 23151 37518 23160
rect 37476 22642 37504 23151
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37568 22094 37596 24890
rect 37648 24608 37700 24614
rect 37648 24550 37700 24556
rect 37476 22066 37596 22094
rect 37372 20528 37424 20534
rect 37372 20470 37424 20476
rect 37476 20380 37504 22066
rect 37556 22024 37608 22030
rect 37556 21966 37608 21972
rect 37384 20352 37504 20380
rect 37384 18873 37412 20352
rect 37464 20256 37516 20262
rect 37464 20198 37516 20204
rect 37476 19854 37504 20198
rect 37464 19848 37516 19854
rect 37464 19790 37516 19796
rect 37568 19378 37596 21966
rect 37660 21554 37688 24550
rect 37648 21548 37700 21554
rect 37648 21490 37700 21496
rect 37646 20904 37702 20913
rect 37646 20839 37702 20848
rect 37556 19372 37608 19378
rect 37556 19314 37608 19320
rect 37660 19258 37688 20839
rect 37568 19230 37688 19258
rect 37370 18864 37426 18873
rect 37370 18799 37426 18808
rect 37464 18080 37516 18086
rect 37464 18022 37516 18028
rect 37476 17678 37504 18022
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37568 17218 37596 19230
rect 37568 17190 37688 17218
rect 37370 16416 37426 16425
rect 37370 16351 37426 16360
rect 37280 13524 37332 13530
rect 37280 13466 37332 13472
rect 37384 13326 37412 16351
rect 37464 15904 37516 15910
rect 37464 15846 37516 15852
rect 37476 15502 37504 15846
rect 37464 15496 37516 15502
rect 37464 15438 37516 15444
rect 37554 14376 37610 14385
rect 37554 14311 37556 14320
rect 37608 14311 37610 14320
rect 37556 14282 37608 14288
rect 37568 14074 37596 14282
rect 37556 14068 37608 14074
rect 37556 14010 37608 14016
rect 37660 13326 37688 17190
rect 37752 14006 37780 25078
rect 37844 24954 37872 25094
rect 37832 24948 37884 24954
rect 37832 24890 37884 24896
rect 37936 24614 37964 29038
rect 38028 28642 38056 30534
rect 38120 30190 38148 31214
rect 38212 30938 38240 34031
rect 38304 33658 38332 34138
rect 38292 33652 38344 33658
rect 38292 33594 38344 33600
rect 38200 30932 38252 30938
rect 38200 30874 38252 30880
rect 38290 30832 38346 30841
rect 38290 30767 38292 30776
rect 38344 30767 38346 30776
rect 38292 30738 38344 30744
rect 38396 30734 38424 35090
rect 38384 30728 38436 30734
rect 38384 30670 38436 30676
rect 38292 30592 38344 30598
rect 38292 30534 38344 30540
rect 38200 30388 38252 30394
rect 38200 30330 38252 30336
rect 38108 30184 38160 30190
rect 38108 30126 38160 30132
rect 38120 29102 38148 30126
rect 38212 29850 38240 30330
rect 38200 29844 38252 29850
rect 38200 29786 38252 29792
rect 38304 29782 38332 30534
rect 38292 29776 38344 29782
rect 38292 29718 38344 29724
rect 38200 29232 38252 29238
rect 38200 29174 38252 29180
rect 38108 29096 38160 29102
rect 38108 29038 38160 29044
rect 38212 28762 38240 29174
rect 38200 28756 38252 28762
rect 38200 28698 38252 28704
rect 38028 28614 38240 28642
rect 38016 28008 38068 28014
rect 38016 27950 38068 27956
rect 38028 26926 38056 27950
rect 38108 27328 38160 27334
rect 38108 27270 38160 27276
rect 38120 26994 38148 27270
rect 38108 26988 38160 26994
rect 38108 26930 38160 26936
rect 38016 26920 38068 26926
rect 38016 26862 38068 26868
rect 38028 25838 38056 26862
rect 38016 25832 38068 25838
rect 38016 25774 38068 25780
rect 38028 24750 38056 25774
rect 38016 24744 38068 24750
rect 38016 24686 38068 24692
rect 37924 24608 37976 24614
rect 37924 24550 37976 24556
rect 37832 24064 37884 24070
rect 37832 24006 37884 24012
rect 37844 23866 37872 24006
rect 37832 23860 37884 23866
rect 37832 23802 37884 23808
rect 38028 23662 38056 24686
rect 38016 23656 38068 23662
rect 38016 23598 38068 23604
rect 37924 22500 37976 22506
rect 37924 22442 37976 22448
rect 37936 21486 37964 22442
rect 37924 21480 37976 21486
rect 38028 21468 38056 23598
rect 38212 21894 38240 28614
rect 38384 28484 38436 28490
rect 38384 28426 38436 28432
rect 38396 26194 38424 28426
rect 38488 26926 38516 37402
rect 38936 35488 38988 35494
rect 38936 35430 38988 35436
rect 38566 34776 38622 34785
rect 38566 34711 38622 34720
rect 38580 31754 38608 34711
rect 38948 31754 38976 35430
rect 39396 33448 39448 33454
rect 39396 33390 39448 33396
rect 39578 33416 39634 33425
rect 38580 31726 38884 31754
rect 38948 31726 39068 31754
rect 38750 30424 38806 30433
rect 38750 30359 38806 30368
rect 38476 26920 38528 26926
rect 38476 26862 38528 26868
rect 38396 26166 38700 26194
rect 38474 26072 38530 26081
rect 38474 26007 38530 26016
rect 38292 23112 38344 23118
rect 38292 23054 38344 23060
rect 38304 22030 38332 23054
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38200 21888 38252 21894
rect 38200 21830 38252 21836
rect 38292 21888 38344 21894
rect 38292 21830 38344 21836
rect 38304 21690 38332 21830
rect 38292 21684 38344 21690
rect 38292 21626 38344 21632
rect 38108 21480 38160 21486
rect 38028 21440 38108 21468
rect 37924 21422 37976 21428
rect 38108 21422 38160 21428
rect 37832 20460 37884 20466
rect 37832 20402 37884 20408
rect 37844 19786 37872 20402
rect 37832 19780 37884 19786
rect 37832 19722 37884 19728
rect 37936 19378 37964 21422
rect 38016 20528 38068 20534
rect 38016 20470 38068 20476
rect 37924 19372 37976 19378
rect 37924 19314 37976 19320
rect 37832 18624 37884 18630
rect 37832 18566 37884 18572
rect 37844 18290 37872 18566
rect 37832 18284 37884 18290
rect 37832 18226 37884 18232
rect 37844 17882 37872 18226
rect 37832 17876 37884 17882
rect 37832 17818 37884 17824
rect 37830 17776 37886 17785
rect 37830 17711 37886 17720
rect 37844 17338 37872 17711
rect 37832 17332 37884 17338
rect 37832 17274 37884 17280
rect 37844 16794 37872 17274
rect 37832 16788 37884 16794
rect 37832 16730 37884 16736
rect 37924 16176 37976 16182
rect 37924 16118 37976 16124
rect 37832 16108 37884 16114
rect 37832 16050 37884 16056
rect 37844 15706 37872 16050
rect 37832 15700 37884 15706
rect 37832 15642 37884 15648
rect 37936 14414 37964 16118
rect 38028 15502 38056 20470
rect 38120 20398 38148 21422
rect 38290 20768 38346 20777
rect 38290 20703 38346 20712
rect 38108 20392 38160 20398
rect 38108 20334 38160 20340
rect 38120 18222 38148 20334
rect 38108 18216 38160 18222
rect 38108 18158 38160 18164
rect 38120 17134 38148 18158
rect 38108 17128 38160 17134
rect 38108 17070 38160 17076
rect 38120 16046 38148 17070
rect 38304 16674 38332 20703
rect 38488 20505 38516 26007
rect 38568 25764 38620 25770
rect 38568 25706 38620 25712
rect 38474 20496 38530 20505
rect 38474 20431 38530 20440
rect 38212 16646 38332 16674
rect 38108 16040 38160 16046
rect 38108 15982 38160 15988
rect 38016 15496 38068 15502
rect 38016 15438 38068 15444
rect 38106 15192 38162 15201
rect 38106 15127 38162 15136
rect 38120 14482 38148 15127
rect 38108 14476 38160 14482
rect 38108 14418 38160 14424
rect 37924 14408 37976 14414
rect 37924 14350 37976 14356
rect 37740 14000 37792 14006
rect 37740 13942 37792 13948
rect 36912 13320 36964 13326
rect 36912 13262 36964 13268
rect 37372 13320 37424 13326
rect 37372 13262 37424 13268
rect 37648 13320 37700 13326
rect 37648 13262 37700 13268
rect 36360 12844 36412 12850
rect 36360 12786 36412 12792
rect 36636 12844 36688 12850
rect 36636 12786 36688 12792
rect 36924 12782 36952 13262
rect 35532 12776 35584 12782
rect 35532 12718 35584 12724
rect 36912 12776 36964 12782
rect 36912 12718 36964 12724
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 35348 11144 35400 11150
rect 35348 11086 35400 11092
rect 38106 11112 38162 11121
rect 34520 11076 34572 11082
rect 38106 11047 38108 11056
rect 34520 11018 34572 11024
rect 38160 11047 38162 11056
rect 38108 11018 38160 11024
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 33692 10056 33744 10062
rect 33692 9998 33744 10004
rect 34336 10056 34388 10062
rect 34336 9998 34388 10004
rect 38108 9988 38160 9994
rect 38108 9930 38160 9936
rect 38120 9761 38148 9930
rect 38106 9752 38162 9761
rect 38106 9687 38162 9696
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 32588 9036 32640 9042
rect 32588 8978 32640 8984
rect 37280 9036 37332 9042
rect 37280 8978 37332 8984
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 37292 5710 37320 8978
rect 37830 8528 37886 8537
rect 38212 8498 38240 16646
rect 38580 12986 38608 25706
rect 38672 13394 38700 26166
rect 38764 15609 38792 30359
rect 38856 27010 38884 31726
rect 39040 27146 39068 31726
rect 39040 27118 39344 27146
rect 38856 26982 39252 27010
rect 39120 26920 39172 26926
rect 39120 26862 39172 26868
rect 38934 24712 38990 24721
rect 38934 24647 38990 24656
rect 38842 23352 38898 23361
rect 38842 23287 38898 23296
rect 38856 22234 38884 23287
rect 38844 22228 38896 22234
rect 38844 22170 38896 22176
rect 38948 21554 38976 24647
rect 39026 21992 39082 22001
rect 39026 21927 39082 21936
rect 38936 21548 38988 21554
rect 38936 21490 38988 21496
rect 38934 20632 38990 20641
rect 38934 20567 38990 20576
rect 38842 19272 38898 19281
rect 38842 19207 38898 19216
rect 38856 17202 38884 19207
rect 38844 17196 38896 17202
rect 38844 17138 38896 17144
rect 38750 15600 38806 15609
rect 38948 15570 38976 20567
rect 39040 19446 39068 21927
rect 39028 19440 39080 19446
rect 39028 19382 39080 19388
rect 39026 19136 39082 19145
rect 39132 19122 39160 26862
rect 39224 22094 39252 26982
rect 39316 25498 39344 27118
rect 39304 25492 39356 25498
rect 39304 25434 39356 25440
rect 39408 24392 39436 33390
rect 39578 33351 39634 33360
rect 39486 29200 39542 29209
rect 39486 29135 39542 29144
rect 39316 24364 39436 24392
rect 39316 23254 39344 24364
rect 39394 24304 39450 24313
rect 39394 24239 39450 24248
rect 39304 23248 39356 23254
rect 39304 23190 39356 23196
rect 39224 22066 39344 22094
rect 39210 21448 39266 21457
rect 39210 21383 39266 21392
rect 39082 19094 39160 19122
rect 39026 19071 39082 19080
rect 39026 17912 39082 17921
rect 39026 17847 39082 17856
rect 39040 17066 39068 17847
rect 39028 17060 39080 17066
rect 39028 17002 39080 17008
rect 39026 16552 39082 16561
rect 39026 16487 39082 16496
rect 38750 15535 38806 15544
rect 38936 15564 38988 15570
rect 38936 15506 38988 15512
rect 39040 15094 39068 16487
rect 39028 15088 39080 15094
rect 39028 15030 39080 15036
rect 39026 13832 39082 13841
rect 39026 13767 39082 13776
rect 39040 13530 39068 13767
rect 39028 13524 39080 13530
rect 39028 13466 39080 13472
rect 38660 13388 38712 13394
rect 38660 13330 38712 13336
rect 38568 12980 38620 12986
rect 38568 12922 38620 12928
rect 38292 12640 38344 12646
rect 38292 12582 38344 12588
rect 38304 12481 38332 12582
rect 38290 12472 38346 12481
rect 38290 12407 38346 12416
rect 39224 11150 39252 21383
rect 39316 17105 39344 22066
rect 39302 17096 39358 17105
rect 39302 17031 39358 17040
rect 39408 14006 39436 24239
rect 39500 14074 39528 29135
rect 39592 24818 39620 33351
rect 39580 24812 39632 24818
rect 39580 24754 39632 24760
rect 39488 14068 39540 14074
rect 39488 14010 39540 14016
rect 39396 14000 39448 14006
rect 39396 13942 39448 13948
rect 39212 11144 39264 11150
rect 39212 11086 39264 11092
rect 37830 8463 37886 8472
rect 38200 8492 38252 8498
rect 37844 7410 37872 8463
rect 38200 8434 38252 8440
rect 38108 8424 38160 8430
rect 38106 8392 38108 8401
rect 38160 8392 38162 8401
rect 38106 8327 38162 8336
rect 37832 7404 37884 7410
rect 37832 7346 37884 7352
rect 38108 7336 38160 7342
rect 38108 7278 38160 7284
rect 38120 7041 38148 7278
rect 38106 7032 38162 7041
rect 38106 6967 38162 6976
rect 37830 6896 37886 6905
rect 37830 6831 37886 6840
rect 37370 6760 37426 6769
rect 37370 6695 37426 6704
rect 37280 5704 37332 5710
rect 37280 5646 37332 5652
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 37384 3058 37412 6695
rect 37844 4622 37872 6831
rect 38106 5672 38162 5681
rect 38106 5607 38108 5616
rect 38160 5607 38162 5616
rect 38108 5578 38160 5584
rect 37832 4616 37884 4622
rect 37832 4558 37884 4564
rect 38108 4548 38160 4554
rect 38108 4490 38160 4496
rect 38120 4321 38148 4490
rect 38106 4312 38162 4321
rect 38106 4247 38162 4256
rect 37372 3052 37424 3058
rect 37372 2994 37424 3000
rect 38108 2984 38160 2990
rect 38106 2952 38108 2961
rect 38160 2952 38162 2961
rect 38106 2887 38162 2896
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 37830 2544 37886 2553
rect 37830 2479 37886 2488
rect 37844 2446 37872 2479
rect 37832 2440 37884 2446
rect 37832 2382 37884 2388
rect 38108 2372 38160 2378
rect 38108 2314 38160 2320
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 38120 1601 38148 2314
rect 38106 1592 38162 1601
rect 38106 1527 38162 1536
<< via2 >>
rect 1674 36216 1730 36272
rect 1766 27920 1822 27976
rect 3606 38256 3662 38312
rect 4894 38664 4950 38720
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4342 35692 4398 35728
rect 4342 35672 4344 35692
rect 4344 35672 4396 35692
rect 4396 35672 4398 35692
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4342 34584 4398 34640
rect 4618 34312 4674 34368
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 3790 25064 3846 25120
rect 3698 22616 3754 22672
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4526 32544 4582 32600
rect 6826 39208 6882 39264
rect 35806 39344 35862 39400
rect 5354 38936 5410 38992
rect 5170 37712 5226 37768
rect 5078 36896 5134 36952
rect 4894 36352 4950 36408
rect 4802 34720 4858 34776
rect 5354 37304 5410 37360
rect 4986 35808 5042 35864
rect 5170 35808 5226 35864
rect 5446 36624 5502 36680
rect 5170 34856 5226 34912
rect 5078 34720 5134 34776
rect 5078 34584 5134 34640
rect 4710 32272 4766 32328
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4434 31884 4490 31920
rect 4434 31864 4436 31884
rect 4436 31864 4488 31884
rect 4488 31864 4490 31884
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4986 32852 4988 32872
rect 4988 32852 5040 32872
rect 5040 32852 5042 32872
rect 4986 32816 5042 32852
rect 4894 31456 4950 31512
rect 4894 26696 4950 26752
rect 4986 26152 5042 26208
rect 4802 25336 4858 25392
rect 4066 24792 4122 24848
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 5078 21936 5134 21992
rect 5722 36780 5778 36816
rect 5722 36760 5724 36780
rect 5724 36760 5776 36780
rect 5776 36760 5778 36780
rect 5446 33768 5502 33824
rect 6090 35944 6146 36000
rect 6458 38528 6514 38584
rect 5814 34040 5870 34096
rect 5814 33260 5816 33280
rect 5816 33260 5868 33280
rect 5868 33260 5870 33280
rect 5814 33224 5870 33260
rect 5262 31048 5318 31104
rect 5354 30676 5356 30696
rect 5356 30676 5408 30696
rect 5408 30676 5410 30696
rect 5354 30640 5410 30676
rect 5630 31320 5686 31376
rect 5814 32272 5870 32328
rect 5998 32272 6054 32328
rect 5722 30504 5778 30560
rect 5538 29416 5594 29472
rect 5906 31220 5908 31240
rect 5908 31220 5960 31240
rect 5960 31220 5962 31240
rect 5906 31184 5962 31220
rect 6090 31728 6146 31784
rect 6550 35808 6606 35864
rect 7102 37304 7158 37360
rect 7010 36488 7066 36544
rect 6826 35128 6882 35184
rect 7378 37848 7434 37904
rect 7010 34604 7066 34640
rect 7010 34584 7012 34604
rect 7012 34584 7064 34604
rect 7064 34584 7066 34604
rect 6550 33632 6606 33688
rect 6642 33496 6698 33552
rect 6642 33088 6698 33144
rect 6366 32544 6422 32600
rect 6274 32136 6330 32192
rect 6550 32544 6606 32600
rect 6274 31456 6330 31512
rect 6274 28600 6330 28656
rect 6642 29552 6698 29608
rect 6550 29144 6606 29200
rect 6918 32952 6974 33008
rect 7102 33516 7158 33552
rect 7102 33496 7104 33516
rect 7104 33496 7156 33516
rect 7156 33496 7158 33516
rect 7286 33940 7288 33960
rect 7288 33940 7340 33960
rect 7340 33940 7342 33960
rect 7286 33904 7342 33940
rect 8114 37576 8170 37632
rect 8758 38800 8814 38856
rect 8666 38392 8722 38448
rect 8390 36488 8446 36544
rect 7838 35400 7894 35456
rect 7746 34720 7802 34776
rect 7838 34604 7894 34640
rect 7838 34584 7840 34604
rect 7840 34584 7892 34604
rect 7892 34584 7894 34604
rect 7746 34176 7802 34232
rect 7562 33360 7618 33416
rect 7102 30912 7158 30968
rect 6918 29280 6974 29336
rect 7838 32136 7894 32192
rect 8206 34584 8262 34640
rect 8482 33632 8538 33688
rect 9402 35808 9458 35864
rect 11242 39072 11298 39128
rect 11058 38120 11114 38176
rect 9678 35980 9680 36000
rect 9680 35980 9732 36000
rect 9732 35980 9734 36000
rect 9678 35944 9734 35980
rect 10230 35808 10286 35864
rect 8114 32408 8170 32464
rect 8206 31864 8262 31920
rect 9034 32680 9090 32736
rect 8942 32544 8998 32600
rect 7562 30096 7618 30152
rect 6826 28872 6882 28928
rect 6734 27784 6790 27840
rect 6366 27240 6422 27296
rect 5446 26016 5502 26072
rect 7746 29824 7802 29880
rect 8390 31456 8446 31512
rect 8114 30776 8170 30832
rect 7930 29688 7986 29744
rect 8114 29300 8170 29336
rect 8114 29280 8116 29300
rect 8116 29280 8168 29300
rect 8168 29280 8170 29300
rect 7654 27648 7710 27704
rect 7010 23160 7066 23216
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 8758 29996 8760 30016
rect 8760 29996 8812 30016
rect 8812 29996 8814 30016
rect 8758 29960 8814 29996
rect 8758 29416 8814 29472
rect 9678 34584 9734 34640
rect 10322 35028 10324 35048
rect 10324 35028 10376 35048
rect 10376 35028 10378 35048
rect 10322 34992 10378 35028
rect 9954 33652 10010 33688
rect 9954 33632 9956 33652
rect 9956 33632 10008 33652
rect 10008 33632 10010 33652
rect 10782 34448 10838 34504
rect 9494 32680 9550 32736
rect 9402 32136 9458 32192
rect 9770 32816 9826 32872
rect 9770 32272 9826 32328
rect 9402 31456 9458 31512
rect 9034 29688 9090 29744
rect 9586 30912 9642 30968
rect 9494 30776 9550 30832
rect 9954 31320 10010 31376
rect 9770 30776 9826 30832
rect 9678 30232 9734 30288
rect 9402 29416 9458 29472
rect 9218 29044 9220 29064
rect 9220 29044 9272 29064
rect 9272 29044 9274 29064
rect 9218 29008 9274 29044
rect 8758 27512 8814 27568
rect 8666 27376 8722 27432
rect 10414 32952 10470 33008
rect 10690 32852 10692 32872
rect 10692 32852 10744 32872
rect 10744 32852 10746 32872
rect 10690 32816 10746 32852
rect 11058 34176 11114 34232
rect 11150 33224 11206 33280
rect 10874 32680 10930 32736
rect 10414 31864 10470 31920
rect 10322 31456 10378 31512
rect 10046 29688 10102 29744
rect 10322 29280 10378 29336
rect 9862 26988 9918 27024
rect 9862 26968 9864 26988
rect 9864 26968 9916 26988
rect 9916 26968 9918 26988
rect 10782 32000 10838 32056
rect 12254 37440 12310 37496
rect 11702 35536 11758 35592
rect 11886 34720 11942 34776
rect 11702 33904 11758 33960
rect 11702 33516 11758 33552
rect 12162 34720 12218 34776
rect 11978 33904 12034 33960
rect 11702 33496 11704 33516
rect 11704 33496 11756 33516
rect 11756 33496 11758 33516
rect 11518 32000 11574 32056
rect 11610 31864 11666 31920
rect 10874 30912 10930 30968
rect 10874 30504 10930 30560
rect 11058 31340 11114 31376
rect 11058 31320 11060 31340
rect 11060 31320 11112 31340
rect 11112 31320 11114 31340
rect 10966 30096 11022 30152
rect 10598 28736 10654 28792
rect 11150 30640 11206 30696
rect 11150 30268 11152 30288
rect 11152 30268 11204 30288
rect 11204 30268 11206 30288
rect 11150 30232 11206 30268
rect 11334 29824 11390 29880
rect 11518 30096 11574 30152
rect 11058 28464 11114 28520
rect 11242 28328 11298 28384
rect 11058 27104 11114 27160
rect 11518 29552 11574 29608
rect 11426 28736 11482 28792
rect 12070 33380 12126 33416
rect 12070 33360 12072 33380
rect 12072 33360 12124 33380
rect 12124 33360 12126 33380
rect 12070 33224 12126 33280
rect 11794 32952 11850 33008
rect 13358 37068 13360 37088
rect 13360 37068 13412 37088
rect 13412 37068 13414 37088
rect 13358 37032 13414 37068
rect 13266 36352 13322 36408
rect 12530 34992 12586 35048
rect 12346 32544 12402 32600
rect 11886 30232 11942 30288
rect 11702 29164 11758 29200
rect 11702 29144 11704 29164
rect 11704 29144 11756 29164
rect 11756 29144 11758 29164
rect 11886 29552 11942 29608
rect 12070 28736 12126 28792
rect 12438 30776 12494 30832
rect 12438 29572 12494 29608
rect 12438 29552 12440 29572
rect 12440 29552 12492 29572
rect 12492 29552 12494 29572
rect 13634 35980 13636 36000
rect 13636 35980 13688 36000
rect 13688 35980 13690 36000
rect 13634 35944 13690 35980
rect 14554 36352 14610 36408
rect 13542 35264 13598 35320
rect 13174 34856 13230 34912
rect 12898 32716 12900 32736
rect 12900 32716 12952 32736
rect 12952 32716 12954 32736
rect 12898 32680 12954 32716
rect 12990 32544 13046 32600
rect 14370 35400 14426 35456
rect 15382 37712 15438 37768
rect 16486 37712 16542 37768
rect 15106 36896 15162 36952
rect 15014 35400 15070 35456
rect 15198 35400 15254 35456
rect 13542 34040 13598 34096
rect 13818 34040 13874 34096
rect 13266 33108 13322 33144
rect 13266 33088 13268 33108
rect 13268 33088 13320 33108
rect 13320 33088 13322 33108
rect 13910 33904 13966 33960
rect 13358 32272 13414 32328
rect 13174 31592 13230 31648
rect 13082 30776 13138 30832
rect 13818 33088 13874 33144
rect 12806 30132 12808 30152
rect 12808 30132 12860 30152
rect 12860 30132 12862 30152
rect 12806 30096 12862 30132
rect 12990 29688 13046 29744
rect 11978 26968 12034 27024
rect 8390 19080 8446 19136
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 13450 30912 13506 30968
rect 13358 30776 13414 30832
rect 14370 33768 14426 33824
rect 14094 32680 14150 32736
rect 14002 32272 14058 32328
rect 14370 32544 14426 32600
rect 14738 34720 14794 34776
rect 15014 34720 15070 34776
rect 14922 34584 14978 34640
rect 14646 32544 14702 32600
rect 14646 32272 14702 32328
rect 14462 31592 14518 31648
rect 14094 31320 14150 31376
rect 13910 30504 13966 30560
rect 13542 28600 13598 28656
rect 13726 28736 13782 28792
rect 13450 26988 13506 27024
rect 13450 26968 13452 26988
rect 13452 26968 13504 26988
rect 13504 26968 13506 26988
rect 13266 26832 13322 26888
rect 12990 25744 13046 25800
rect 14094 28736 14150 28792
rect 14554 30912 14610 30968
rect 14554 26968 14610 27024
rect 14922 34040 14978 34096
rect 14830 32816 14886 32872
rect 15290 34448 15346 34504
rect 15934 37032 15990 37088
rect 15750 35536 15806 35592
rect 15750 34992 15806 35048
rect 15566 34176 15622 34232
rect 16486 36216 16542 36272
rect 16210 35264 16266 35320
rect 15934 34584 15990 34640
rect 15842 34448 15898 34504
rect 14922 31456 14978 31512
rect 14738 30776 14794 30832
rect 15842 33224 15898 33280
rect 15474 32544 15530 32600
rect 15382 32136 15438 32192
rect 15198 31204 15254 31240
rect 15198 31184 15200 31204
rect 15200 31184 15252 31204
rect 15252 31184 15254 31204
rect 15658 31320 15714 31376
rect 15934 32816 15990 32872
rect 16486 35808 16542 35864
rect 16394 34448 16450 34504
rect 16394 34176 16450 34232
rect 16302 33904 16358 33960
rect 16302 31592 16358 31648
rect 14462 25220 14518 25256
rect 14462 25200 14464 25220
rect 14464 25200 14516 25220
rect 14516 25200 14518 25220
rect 15106 27820 15108 27840
rect 15108 27820 15160 27840
rect 15160 27820 15162 27840
rect 15106 27784 15162 27820
rect 15750 29688 15806 29744
rect 15290 26968 15346 27024
rect 15750 27376 15806 27432
rect 16118 28872 16174 28928
rect 16118 28484 16174 28520
rect 16118 28464 16120 28484
rect 16120 28464 16172 28484
rect 16172 28464 16174 28484
rect 15842 27240 15898 27296
rect 15198 24928 15254 24984
rect 16578 32816 16634 32872
rect 16578 31900 16580 31920
rect 16580 31900 16632 31920
rect 16632 31900 16634 31920
rect 16578 31864 16634 31900
rect 17222 37168 17278 37224
rect 17038 36216 17094 36272
rect 17222 36624 17278 36680
rect 17406 36624 17462 36680
rect 17314 36080 17370 36136
rect 16854 33224 16910 33280
rect 16854 32680 16910 32736
rect 16486 30912 16542 30968
rect 16486 29960 16542 30016
rect 16670 30912 16726 30968
rect 16578 28600 16634 28656
rect 17406 34856 17462 34912
rect 17314 34720 17370 34776
rect 18050 35980 18052 36000
rect 18052 35980 18104 36000
rect 18104 35980 18106 36000
rect 18050 35944 18106 35980
rect 17958 35572 17960 35592
rect 17960 35572 18012 35592
rect 18012 35572 18014 35592
rect 17958 35536 18014 35572
rect 17866 34040 17922 34096
rect 17130 29688 17186 29744
rect 16762 28192 16818 28248
rect 17406 29144 17462 29200
rect 17866 32544 17922 32600
rect 19430 37304 19486 37360
rect 18234 34856 18290 34912
rect 18234 33088 18290 33144
rect 18418 33632 18474 33688
rect 18234 32544 18290 32600
rect 18418 32680 18474 32736
rect 17866 31456 17922 31512
rect 18050 30368 18106 30424
rect 18786 35536 18842 35592
rect 18602 32136 18658 32192
rect 18050 29416 18106 29472
rect 17406 26968 17462 27024
rect 17866 27512 17922 27568
rect 17682 27376 17738 27432
rect 12438 20596 12494 20632
rect 12438 20576 12440 20596
rect 12440 20576 12492 20596
rect 12492 20576 12494 20596
rect 14002 20576 14058 20632
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 3882 17040 3938 17096
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 17958 26968 18014 27024
rect 18050 26696 18106 26752
rect 17314 23432 17370 23488
rect 17958 26288 18014 26344
rect 18970 36524 18972 36544
rect 18972 36524 19024 36544
rect 19024 36524 19026 36544
rect 18970 36488 19026 36524
rect 18970 35944 19026 36000
rect 19338 36896 19394 36952
rect 19338 36216 19394 36272
rect 19246 35828 19302 35864
rect 19246 35808 19248 35828
rect 19248 35808 19300 35828
rect 19300 35808 19302 35828
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 20534 37304 20590 37360
rect 20166 36352 20222 36408
rect 19614 34448 19670 34504
rect 19430 34040 19486 34096
rect 19982 33904 20038 33960
rect 18786 31592 18842 31648
rect 18878 31456 18934 31512
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 20074 33632 20130 33688
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 18970 30504 19026 30560
rect 18786 30096 18842 30152
rect 18786 28328 18842 28384
rect 18786 26696 18842 26752
rect 18602 26288 18658 26344
rect 18602 26152 18658 26208
rect 18418 25608 18474 25664
rect 18418 25064 18474 25120
rect 18050 24656 18106 24712
rect 17774 24384 17830 24440
rect 17682 23704 17738 23760
rect 19338 31864 19394 31920
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 20994 37304 21050 37360
rect 20350 32272 20406 32328
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19062 26036 19118 26072
rect 19062 26016 19064 26036
rect 19064 26016 19116 26036
rect 19116 26016 19118 26036
rect 19062 24248 19118 24304
rect 18786 23568 18842 23624
rect 18970 23432 19026 23488
rect 20350 31592 20406 31648
rect 20074 29008 20130 29064
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19430 27784 19486 27840
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19430 25744 19486 25800
rect 21638 37032 21694 37088
rect 20718 33768 20774 33824
rect 20810 33224 20866 33280
rect 20810 32136 20866 32192
rect 20810 31884 20866 31920
rect 20810 31864 20812 31884
rect 20812 31864 20864 31884
rect 20864 31864 20866 31884
rect 21270 32272 21326 32328
rect 21178 31864 21234 31920
rect 21638 32544 21694 32600
rect 21638 32428 21694 32464
rect 21638 32408 21640 32428
rect 21640 32408 21692 32428
rect 21692 32408 21694 32428
rect 21546 30640 21602 30696
rect 20442 28056 20498 28112
rect 20166 25744 20222 25800
rect 19430 25336 19486 25392
rect 19430 25064 19486 25120
rect 19982 25064 20038 25120
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19246 23432 19302 23488
rect 19154 23296 19210 23352
rect 18050 22480 18106 22536
rect 17130 20868 17186 20904
rect 17130 20848 17132 20868
rect 17132 20848 17184 20868
rect 17184 20848 17186 20868
rect 18050 20440 18106 20496
rect 18234 20984 18290 21040
rect 18142 20304 18198 20360
rect 14738 15544 14794 15600
rect 19522 24112 19578 24168
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 20718 28212 20774 28248
rect 20718 28192 20720 28212
rect 20720 28192 20772 28212
rect 20772 28192 20774 28212
rect 20534 26324 20536 26344
rect 20536 26324 20588 26344
rect 20588 26324 20590 26344
rect 20534 26288 20590 26324
rect 20534 26152 20590 26208
rect 20626 25492 20682 25528
rect 20626 25472 20628 25492
rect 20628 25472 20680 25492
rect 20680 25472 20682 25492
rect 20350 24656 20406 24712
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19798 22480 19854 22536
rect 20994 26016 21050 26072
rect 20718 24556 20720 24576
rect 20720 24556 20772 24576
rect 20772 24556 20774 24576
rect 20718 24520 20774 24556
rect 20902 24656 20958 24712
rect 20718 23568 20774 23624
rect 20442 23296 20498 23352
rect 20258 22888 20314 22944
rect 20166 22344 20222 22400
rect 19890 21972 19892 21992
rect 19892 21972 19944 21992
rect 19944 21972 19946 21992
rect 19890 21936 19946 21972
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 20074 21664 20130 21720
rect 19890 21392 19946 21448
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 20718 23296 20774 23352
rect 20074 20032 20130 20088
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19798 18264 19854 18320
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 22374 38936 22430 38992
rect 22098 36080 22154 36136
rect 22006 35944 22062 36000
rect 22650 36624 22706 36680
rect 22098 33904 22154 33960
rect 22466 33904 22522 33960
rect 22282 33632 22338 33688
rect 23110 36488 23166 36544
rect 23018 36080 23074 36136
rect 22742 34312 22798 34368
rect 22190 32952 22246 33008
rect 21914 32680 21970 32736
rect 21822 32408 21878 32464
rect 22098 32136 22154 32192
rect 21638 29824 21694 29880
rect 21362 28872 21418 28928
rect 21454 28056 21510 28112
rect 21638 27920 21694 27976
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 20902 18128 20958 18184
rect 21730 24928 21786 24984
rect 21730 24248 21786 24304
rect 23110 35400 23166 35456
rect 22834 32680 22890 32736
rect 22926 32544 22982 32600
rect 22742 32408 22798 32464
rect 22742 32136 22798 32192
rect 22190 29144 22246 29200
rect 22098 28736 22154 28792
rect 22374 29008 22430 29064
rect 22190 24112 22246 24168
rect 22650 29552 22706 29608
rect 23386 36896 23442 36952
rect 24674 38120 24730 38176
rect 23386 34992 23442 35048
rect 23386 34620 23388 34640
rect 23388 34620 23440 34640
rect 23440 34620 23442 34640
rect 23386 34584 23442 34620
rect 23294 34448 23350 34504
rect 23110 32408 23166 32464
rect 22742 29144 22798 29200
rect 22650 27648 22706 27704
rect 23478 32952 23534 33008
rect 23386 32272 23442 32328
rect 23294 31864 23350 31920
rect 22926 27648 22982 27704
rect 23846 35672 23902 35728
rect 24490 37304 24546 37360
rect 24306 35264 24362 35320
rect 23754 32272 23810 32328
rect 23662 31592 23718 31648
rect 23754 31048 23810 31104
rect 24214 33360 24270 33416
rect 24030 32680 24086 32736
rect 24122 32000 24178 32056
rect 24122 31048 24178 31104
rect 23110 27240 23166 27296
rect 22466 26152 22522 26208
rect 22650 25472 22706 25528
rect 22466 25064 22522 25120
rect 22926 26832 22982 26888
rect 23294 26288 23350 26344
rect 22926 25200 22982 25256
rect 22742 24928 22798 24984
rect 22742 23024 22798 23080
rect 22282 22888 22338 22944
rect 22834 22888 22890 22944
rect 21638 21664 21694 21720
rect 22466 21120 22522 21176
rect 22190 19896 22246 19952
rect 22098 19760 22154 19816
rect 22466 19216 22522 19272
rect 22190 17212 22192 17232
rect 22192 17212 22244 17232
rect 22244 17212 22246 17232
rect 22190 17176 22246 17212
rect 22650 20576 22706 20632
rect 22834 20984 22890 21040
rect 22926 20440 22982 20496
rect 23846 28500 23848 28520
rect 23848 28500 23900 28520
rect 23900 28500 23902 28520
rect 30010 38800 30066 38856
rect 26422 38664 26478 38720
rect 25870 38120 25926 38176
rect 25502 36896 25558 36952
rect 25318 36488 25374 36544
rect 24582 35672 24638 35728
rect 24858 35808 24914 35864
rect 24582 33088 24638 33144
rect 24214 30096 24270 30152
rect 24214 29280 24270 29336
rect 23846 28464 23902 28500
rect 23754 28192 23810 28248
rect 23938 28192 23994 28248
rect 23846 27240 23902 27296
rect 23846 26288 23902 26344
rect 24030 27784 24086 27840
rect 23938 25608 23994 25664
rect 24214 26152 24270 26208
rect 23938 24812 23994 24848
rect 23938 24792 23940 24812
rect 23940 24792 23992 24812
rect 23992 24792 23994 24812
rect 23202 23568 23258 23624
rect 23202 22616 23258 22672
rect 23662 23044 23718 23080
rect 23662 23024 23664 23044
rect 23664 23024 23716 23044
rect 23716 23024 23718 23044
rect 23110 20576 23166 20632
rect 23202 19896 23258 19952
rect 24490 32816 24546 32872
rect 25226 35808 25282 35864
rect 25778 35672 25834 35728
rect 25134 34720 25190 34776
rect 24582 32544 24638 32600
rect 24674 31320 24730 31376
rect 24766 30912 24822 30968
rect 25502 34176 25558 34232
rect 26146 37168 26202 37224
rect 25410 33496 25466 33552
rect 25318 33088 25374 33144
rect 25042 32952 25098 33008
rect 24950 32852 24952 32872
rect 24952 32852 25004 32872
rect 25004 32852 25006 32872
rect 24950 32816 25006 32852
rect 24950 31728 25006 31784
rect 24490 28464 24546 28520
rect 24490 27920 24546 27976
rect 25318 32272 25374 32328
rect 25318 32136 25374 32192
rect 25410 31884 25466 31920
rect 25410 31864 25412 31884
rect 25412 31864 25464 31884
rect 25464 31864 25466 31884
rect 25686 32952 25742 33008
rect 25594 31456 25650 31512
rect 25226 30912 25282 30968
rect 25686 31184 25742 31240
rect 25686 30640 25742 30696
rect 25594 30132 25596 30152
rect 25596 30132 25648 30152
rect 25648 30132 25650 30152
rect 25594 30096 25650 30132
rect 25042 29552 25098 29608
rect 25042 29280 25098 29336
rect 24766 29008 24822 29064
rect 25042 29008 25098 29064
rect 24306 25744 24362 25800
rect 24306 23432 24362 23488
rect 24122 21936 24178 21992
rect 24582 26696 24638 26752
rect 24858 26424 24914 26480
rect 24950 25608 25006 25664
rect 25226 26696 25282 26752
rect 25134 26424 25190 26480
rect 24858 24928 24914 24984
rect 24582 23024 24638 23080
rect 24306 21256 24362 21312
rect 24030 20440 24086 20496
rect 24030 19896 24086 19952
rect 23754 19372 23810 19408
rect 23754 19352 23756 19372
rect 23756 19352 23808 19372
rect 23808 19352 23810 19372
rect 23110 17584 23166 17640
rect 23202 17312 23258 17368
rect 24030 19080 24086 19136
rect 25042 24248 25098 24304
rect 25226 24928 25282 24984
rect 24490 21120 24546 21176
rect 24122 18808 24178 18864
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 24306 18284 24362 18320
rect 24306 18264 24308 18284
rect 24308 18264 24360 18284
rect 24360 18264 24362 18284
rect 25042 21392 25098 21448
rect 24582 19080 24638 19136
rect 24766 17620 24768 17640
rect 24768 17620 24820 17640
rect 24820 17620 24822 17640
rect 24766 17584 24822 17620
rect 25410 25064 25466 25120
rect 25594 25880 25650 25936
rect 25594 25200 25650 25256
rect 25502 24676 25558 24712
rect 25502 24656 25504 24676
rect 25504 24656 25556 24676
rect 25556 24656 25558 24676
rect 26054 35400 26110 35456
rect 26146 34312 26202 34368
rect 26238 34176 26294 34232
rect 26698 35672 26754 35728
rect 26514 34720 26570 34776
rect 27894 38528 27950 38584
rect 26882 35264 26938 35320
rect 26330 34040 26386 34096
rect 26882 34040 26938 34096
rect 26422 33360 26478 33416
rect 26330 33260 26332 33280
rect 26332 33260 26384 33280
rect 26384 33260 26386 33280
rect 26330 33224 26386 33260
rect 26330 32136 26386 32192
rect 26146 31184 26202 31240
rect 26054 30368 26110 30424
rect 26330 31184 26386 31240
rect 26238 29144 26294 29200
rect 26054 28464 26110 28520
rect 26238 28464 26294 28520
rect 26422 29008 26478 29064
rect 26606 29300 26662 29336
rect 26606 29280 26608 29300
rect 26608 29280 26660 29300
rect 26660 29280 26662 29300
rect 26054 27532 26110 27568
rect 26054 27512 26056 27532
rect 26056 27512 26108 27532
rect 26108 27512 26110 27532
rect 25962 25744 26018 25800
rect 25962 25608 26018 25664
rect 26330 27648 26386 27704
rect 26146 26288 26202 26344
rect 26514 27648 26570 27704
rect 26514 25880 26570 25936
rect 26790 31456 26846 31512
rect 27066 35400 27122 35456
rect 27434 36488 27490 36544
rect 27342 35828 27398 35864
rect 27342 35808 27344 35828
rect 27344 35808 27396 35828
rect 27396 35808 27398 35828
rect 27342 35264 27398 35320
rect 27250 35012 27306 35048
rect 27250 34992 27252 35012
rect 27252 34992 27304 35012
rect 27304 34992 27306 35012
rect 27342 34856 27398 34912
rect 27618 36760 27674 36816
rect 27526 34992 27582 35048
rect 28998 37440 29054 37496
rect 27894 34856 27950 34912
rect 27894 34720 27950 34776
rect 27066 31592 27122 31648
rect 27342 33496 27398 33552
rect 27526 33632 27582 33688
rect 27526 32544 27582 32600
rect 27066 31048 27122 31104
rect 26974 29960 27030 30016
rect 27158 29688 27214 29744
rect 27894 32816 27950 32872
rect 27618 30776 27674 30832
rect 27526 30232 27582 30288
rect 27434 29824 27490 29880
rect 27158 29280 27214 29336
rect 27158 29144 27214 29200
rect 27158 28736 27214 28792
rect 27066 27512 27122 27568
rect 27158 27240 27214 27296
rect 27526 27512 27582 27568
rect 26790 26152 26846 26208
rect 25962 24656 26018 24712
rect 25410 23160 25466 23216
rect 25226 22480 25282 22536
rect 25686 22344 25742 22400
rect 25134 20032 25190 20088
rect 24950 19352 25006 19408
rect 24858 16768 24914 16824
rect 24582 16496 24638 16552
rect 25686 19080 25742 19136
rect 25686 18400 25742 18456
rect 26238 24656 26294 24712
rect 26146 24112 26202 24168
rect 25962 22480 26018 22536
rect 26054 20032 26110 20088
rect 26514 24012 26516 24032
rect 26516 24012 26568 24032
rect 26568 24012 26570 24032
rect 26514 23976 26570 24012
rect 26790 23160 26846 23216
rect 26606 20848 26662 20904
rect 25962 19488 26018 19544
rect 25870 19080 25926 19136
rect 26054 18400 26110 18456
rect 25778 17620 25780 17640
rect 25780 17620 25832 17640
rect 25832 17620 25834 17640
rect 25778 17584 25834 17620
rect 25778 16632 25834 16688
rect 26238 18672 26294 18728
rect 26238 18128 26294 18184
rect 26514 19216 26570 19272
rect 26422 18264 26478 18320
rect 26146 16632 26202 16688
rect 26514 18128 26570 18184
rect 27158 23704 27214 23760
rect 26882 19080 26938 19136
rect 27158 21120 27214 21176
rect 27894 31748 27950 31784
rect 27894 31728 27896 31748
rect 27896 31728 27948 31748
rect 27948 31728 27950 31748
rect 27894 30912 27950 30968
rect 27802 28328 27858 28384
rect 27802 27240 27858 27296
rect 27710 26188 27712 26208
rect 27712 26188 27764 26208
rect 27764 26188 27766 26208
rect 27710 26152 27766 26188
rect 27526 25336 27582 25392
rect 27434 23976 27490 24032
rect 27618 25236 27620 25256
rect 27620 25236 27672 25256
rect 27672 25236 27674 25256
rect 27618 25200 27674 25236
rect 27618 24112 27674 24168
rect 27526 23568 27582 23624
rect 28262 35808 28318 35864
rect 28722 36624 28778 36680
rect 29642 37168 29698 37224
rect 29182 36216 29238 36272
rect 28538 34856 28594 34912
rect 28354 34720 28410 34776
rect 28446 34040 28502 34096
rect 28906 34856 28962 34912
rect 28998 34620 29000 34640
rect 29000 34620 29052 34640
rect 29052 34620 29054 34640
rect 28998 34584 29054 34620
rect 28998 34040 29054 34096
rect 28538 33224 28594 33280
rect 28354 32952 28410 33008
rect 28078 30368 28134 30424
rect 28630 32952 28686 33008
rect 28538 32544 28594 32600
rect 28998 33768 29054 33824
rect 28906 33532 28908 33552
rect 28908 33532 28960 33552
rect 28960 33532 28962 33552
rect 28906 33496 28962 33532
rect 29090 33224 29146 33280
rect 28814 32680 28870 32736
rect 29090 32680 29146 32736
rect 29090 32408 29146 32464
rect 28814 32272 28870 32328
rect 29090 32272 29146 32328
rect 28630 32000 28686 32056
rect 28814 31864 28870 31920
rect 28722 31728 28778 31784
rect 28446 31320 28502 31376
rect 28170 29008 28226 29064
rect 28446 30368 28502 30424
rect 29458 34584 29514 34640
rect 29366 33904 29422 33960
rect 29550 33904 29606 33960
rect 28998 30368 29054 30424
rect 28446 29280 28502 29336
rect 27894 24928 27950 24984
rect 27802 24792 27858 24848
rect 27986 24692 27988 24712
rect 27988 24692 28040 24712
rect 28040 24692 28042 24712
rect 27986 24656 28042 24692
rect 27802 24268 27858 24304
rect 27802 24248 27804 24268
rect 27804 24248 27856 24268
rect 27856 24248 27858 24268
rect 28078 24520 28134 24576
rect 27342 20576 27398 20632
rect 27434 19624 27490 19680
rect 27434 18944 27490 19000
rect 27342 18672 27398 18728
rect 28354 25472 28410 25528
rect 28262 23296 28318 23352
rect 28538 25608 28594 25664
rect 29826 35808 29882 35864
rect 29458 32000 29514 32056
rect 29366 30504 29422 30560
rect 29274 29824 29330 29880
rect 29182 28872 29238 28928
rect 28998 27004 29000 27024
rect 29000 27004 29052 27024
rect 29052 27004 29054 27024
rect 28998 26968 29054 27004
rect 29274 26968 29330 27024
rect 28906 26424 28962 26480
rect 28998 26152 29054 26208
rect 28814 25880 28870 25936
rect 28722 25608 28778 25664
rect 28630 24928 28686 24984
rect 28630 24792 28686 24848
rect 28446 23432 28502 23488
rect 28906 25492 28962 25528
rect 28906 25472 28908 25492
rect 28908 25472 28960 25492
rect 28960 25472 28962 25492
rect 29182 24948 29238 24984
rect 29182 24928 29184 24948
rect 29184 24928 29236 24948
rect 29236 24928 29238 24948
rect 29090 24828 29092 24848
rect 29092 24828 29144 24848
rect 29144 24828 29146 24848
rect 29090 24792 29146 24828
rect 29090 24012 29092 24032
rect 29092 24012 29144 24032
rect 29144 24012 29146 24032
rect 29090 23976 29146 24012
rect 28998 23840 29054 23896
rect 28446 22752 28502 22808
rect 28538 20848 28594 20904
rect 28354 20576 28410 20632
rect 28354 20324 28410 20360
rect 28354 20304 28356 20324
rect 28356 20304 28408 20324
rect 28408 20304 28410 20324
rect 28262 19760 28318 19816
rect 27986 17720 28042 17776
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 28170 18708 28172 18728
rect 28172 18708 28224 18728
rect 28224 18708 28226 18728
rect 28170 18672 28226 18708
rect 28354 18264 28410 18320
rect 28354 17312 28410 17368
rect 28262 17176 28318 17232
rect 29090 23432 29146 23488
rect 28998 22616 29054 22672
rect 28998 22480 29054 22536
rect 28998 21972 29000 21992
rect 29000 21972 29052 21992
rect 29052 21972 29054 21992
rect 28998 21936 29054 21972
rect 28906 21528 28962 21584
rect 28630 18808 28686 18864
rect 28538 18128 28594 18184
rect 28998 20576 29054 20632
rect 28998 19932 29000 19952
rect 29000 19932 29052 19952
rect 29052 19932 29054 19952
rect 28998 19896 29054 19932
rect 28814 16224 28870 16280
rect 28998 19488 29054 19544
rect 29182 20304 29238 20360
rect 29090 18128 29146 18184
rect 29550 30912 29606 30968
rect 29550 29960 29606 30016
rect 29826 34312 29882 34368
rect 29734 32408 29790 32464
rect 29734 31728 29790 31784
rect 29734 31356 29736 31376
rect 29736 31356 29788 31376
rect 29788 31356 29790 31376
rect 29734 31320 29790 31356
rect 30194 37984 30250 38040
rect 30102 37848 30158 37904
rect 30102 36760 30158 36816
rect 30010 32408 30066 32464
rect 30286 35536 30342 35592
rect 30286 35436 30288 35456
rect 30288 35436 30340 35456
rect 30340 35436 30342 35456
rect 30286 35400 30342 35436
rect 30286 35128 30342 35184
rect 30194 33224 30250 33280
rect 30470 34176 30526 34232
rect 30378 33360 30434 33416
rect 30746 34892 30748 34912
rect 30748 34892 30800 34912
rect 30800 34892 30802 34912
rect 30746 34856 30802 34892
rect 30746 34720 30802 34776
rect 30654 34448 30710 34504
rect 30654 34176 30710 34232
rect 30654 33632 30710 33688
rect 30470 32408 30526 32464
rect 30470 31884 30526 31920
rect 30470 31864 30472 31884
rect 30472 31864 30524 31884
rect 30524 31864 30526 31884
rect 30654 32136 30710 32192
rect 30654 31456 30710 31512
rect 30470 31184 30526 31240
rect 30930 31592 30986 31648
rect 29918 29824 29974 29880
rect 29734 29688 29790 29744
rect 29734 29452 29736 29472
rect 29736 29452 29788 29472
rect 29788 29452 29790 29472
rect 29734 29416 29790 29452
rect 29642 29144 29698 29200
rect 29642 27512 29698 27568
rect 29642 26968 29698 27024
rect 29550 26696 29606 26752
rect 29550 26288 29606 26344
rect 30010 29688 30066 29744
rect 30010 27920 30066 27976
rect 29918 27512 29974 27568
rect 29642 25744 29698 25800
rect 29734 25472 29790 25528
rect 30286 29416 30342 29472
rect 30286 28736 30342 28792
rect 30746 30232 30802 30288
rect 30654 29996 30656 30016
rect 30656 29996 30708 30016
rect 30708 29996 30710 30016
rect 30654 29960 30710 29996
rect 30746 29688 30802 29744
rect 30562 29164 30618 29200
rect 30562 29144 30564 29164
rect 30564 29144 30616 29164
rect 30616 29144 30618 29164
rect 30102 27104 30158 27160
rect 30654 28600 30710 28656
rect 30378 27920 30434 27976
rect 30378 27512 30434 27568
rect 30562 26968 30618 27024
rect 31022 31184 31078 31240
rect 30930 30368 30986 30424
rect 31022 29960 31078 30016
rect 30838 29144 30894 29200
rect 30930 28872 30986 28928
rect 30838 27956 30840 27976
rect 30840 27956 30892 27976
rect 30892 27956 30894 27976
rect 30838 27920 30894 27956
rect 30286 26288 30342 26344
rect 30102 26016 30158 26072
rect 30010 25472 30066 25528
rect 30010 25200 30066 25256
rect 29458 24248 29514 24304
rect 29826 23976 29882 24032
rect 29734 23704 29790 23760
rect 29458 23568 29514 23624
rect 29458 23160 29514 23216
rect 29734 22752 29790 22808
rect 29550 22500 29606 22536
rect 29550 22480 29552 22500
rect 29552 22480 29604 22500
rect 29604 22480 29606 22500
rect 29550 22092 29606 22128
rect 29550 22072 29552 22092
rect 29552 22072 29604 22092
rect 29604 22072 29606 22092
rect 29734 20576 29790 20632
rect 29550 20440 29606 20496
rect 29458 19780 29514 19816
rect 29458 19760 29460 19780
rect 29460 19760 29512 19780
rect 29512 19760 29514 19780
rect 29366 18844 29368 18864
rect 29368 18844 29420 18864
rect 29420 18844 29422 18864
rect 29366 18808 29422 18844
rect 28998 16632 29054 16688
rect 29182 16632 29238 16688
rect 30286 25744 30342 25800
rect 30194 25608 30250 25664
rect 30562 25880 30618 25936
rect 30470 24928 30526 24984
rect 30378 24556 30380 24576
rect 30380 24556 30432 24576
rect 30432 24556 30434 24576
rect 30378 24520 30434 24556
rect 30010 23160 30066 23216
rect 30286 22924 30288 22944
rect 30288 22924 30340 22944
rect 30340 22924 30342 22944
rect 30286 22888 30342 22924
rect 31206 36624 31262 36680
rect 31574 34856 31630 34912
rect 31206 32680 31262 32736
rect 31850 36916 31906 36952
rect 31850 36896 31852 36916
rect 31852 36896 31904 36916
rect 31904 36896 31906 36916
rect 32310 37204 32312 37224
rect 32312 37204 32364 37224
rect 32364 37204 32366 37224
rect 32310 37168 32366 37204
rect 32310 36216 32366 36272
rect 32310 35828 32366 35864
rect 32310 35808 32312 35828
rect 32312 35808 32364 35828
rect 32364 35808 32366 35828
rect 32310 35400 32366 35456
rect 31758 34992 31814 35048
rect 32034 34720 32090 34776
rect 31942 34584 31998 34640
rect 31758 34040 31814 34096
rect 31942 33632 31998 33688
rect 31298 30504 31354 30560
rect 30930 26424 30986 26480
rect 30930 26324 30932 26344
rect 30932 26324 30984 26344
rect 30984 26324 30986 26344
rect 30930 26288 30986 26324
rect 30930 25608 30986 25664
rect 30930 24792 30986 24848
rect 30746 24520 30802 24576
rect 30838 23840 30894 23896
rect 30746 23704 30802 23760
rect 30654 23160 30710 23216
rect 30654 23024 30710 23080
rect 30194 22480 30250 22536
rect 30102 21800 30158 21856
rect 30378 22072 30434 22128
rect 30470 21936 30526 21992
rect 30286 21564 30288 21584
rect 30288 21564 30340 21584
rect 30340 21564 30342 21584
rect 30286 21528 30342 21564
rect 29918 18964 29974 19000
rect 29918 18944 29920 18964
rect 29920 18944 29972 18964
rect 29972 18944 29974 18964
rect 30010 18536 30066 18592
rect 30010 17992 30066 18048
rect 30102 16632 30158 16688
rect 30838 22636 30894 22672
rect 30838 22616 30840 22636
rect 30840 22616 30892 22636
rect 30892 22616 30894 22636
rect 31206 25880 31262 25936
rect 31114 25608 31170 25664
rect 31482 29044 31484 29064
rect 31484 29044 31536 29064
rect 31536 29044 31538 29064
rect 31482 29008 31538 29044
rect 31390 25608 31446 25664
rect 31850 30368 31906 30424
rect 31850 30232 31906 30288
rect 32126 34312 32182 34368
rect 32310 33360 32366 33416
rect 32310 32272 32366 32328
rect 32954 36760 33010 36816
rect 32678 34584 32734 34640
rect 32678 34484 32680 34504
rect 32680 34484 32732 34504
rect 32732 34484 32734 34504
rect 32678 34448 32734 34484
rect 35622 38936 35678 38992
rect 35530 38392 35586 38448
rect 35438 38256 35494 38312
rect 34702 37304 34758 37360
rect 33874 36352 33930 36408
rect 33414 35400 33470 35456
rect 33414 35264 33470 35320
rect 33322 35128 33378 35184
rect 32862 34176 32918 34232
rect 33230 34448 33286 34504
rect 33046 34176 33102 34232
rect 32678 33088 32734 33144
rect 32586 32136 32642 32192
rect 32034 31728 32090 31784
rect 32034 31592 32090 31648
rect 32126 31456 32182 31512
rect 32034 31048 32090 31104
rect 31942 29688 31998 29744
rect 31666 28092 31668 28112
rect 31668 28092 31720 28112
rect 31720 28092 31722 28112
rect 31666 28056 31722 28092
rect 31666 27784 31722 27840
rect 31574 27512 31630 27568
rect 31666 27376 31722 27432
rect 31114 21800 31170 21856
rect 30378 20168 30434 20224
rect 30286 19080 30342 19136
rect 30470 18944 30526 19000
rect 31298 23724 31354 23760
rect 31298 23704 31300 23724
rect 31300 23704 31352 23724
rect 31352 23704 31354 23724
rect 31298 23160 31354 23216
rect 31206 21392 31262 21448
rect 30562 18572 30564 18592
rect 30564 18572 30616 18592
rect 30616 18572 30618 18592
rect 30562 18536 30618 18572
rect 31758 26968 31814 27024
rect 31850 26288 31906 26344
rect 31758 24404 31814 24440
rect 31758 24384 31760 24404
rect 31760 24384 31812 24404
rect 31812 24384 31814 24404
rect 31942 25472 31998 25528
rect 31758 23976 31814 24032
rect 31758 23432 31814 23488
rect 30930 18808 30986 18864
rect 30654 17856 30710 17912
rect 30562 17620 30564 17640
rect 30564 17620 30616 17640
rect 30616 17620 30618 17640
rect 30562 17584 30618 17620
rect 30286 16496 30342 16552
rect 30194 16360 30250 16416
rect 30102 16224 30158 16280
rect 30746 17312 30802 17368
rect 30746 16244 30802 16280
rect 30746 16224 30748 16244
rect 30748 16224 30800 16244
rect 30800 16224 30802 16244
rect 31206 19216 31262 19272
rect 31942 23840 31998 23896
rect 32126 30368 32182 30424
rect 32126 29144 32182 29200
rect 32586 31864 32642 31920
rect 32586 29824 32642 29880
rect 32494 28736 32550 28792
rect 32218 27532 32274 27568
rect 32218 27512 32220 27532
rect 32220 27512 32272 27532
rect 32272 27512 32274 27532
rect 32218 27240 32274 27296
rect 32402 27240 32458 27296
rect 32402 26560 32458 26616
rect 32402 24384 32458 24440
rect 32862 32272 32918 32328
rect 32954 30232 33010 30288
rect 33322 33632 33378 33688
rect 33414 33360 33470 33416
rect 33322 32680 33378 32736
rect 33598 33632 33654 33688
rect 33598 31864 33654 31920
rect 33138 30504 33194 30560
rect 33506 31048 33562 31104
rect 33966 35808 34022 35864
rect 34150 35572 34152 35592
rect 34152 35572 34204 35592
rect 34204 35572 34206 35592
rect 34150 35536 34206 35572
rect 34426 36488 34482 36544
rect 34242 34992 34298 35048
rect 34058 34176 34114 34232
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35162 36896 35218 36952
rect 35346 36896 35402 36952
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34610 34312 34666 34368
rect 34150 33224 34206 33280
rect 33874 32408 33930 32464
rect 33966 31764 33968 31784
rect 33968 31764 34020 31784
rect 34020 31764 34022 31784
rect 33966 31728 34022 31764
rect 33874 31592 33930 31648
rect 34334 32816 34390 32872
rect 34610 32952 34666 33008
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35438 34856 35494 34912
rect 35254 33516 35310 33552
rect 35254 33496 35256 33516
rect 35256 33496 35308 33516
rect 35308 33496 35310 33516
rect 35070 33360 35126 33416
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 33046 28056 33102 28112
rect 33046 26696 33102 26752
rect 32954 26152 33010 26208
rect 33322 28736 33378 28792
rect 33690 30232 33746 30288
rect 33506 29280 33562 29336
rect 33230 26016 33286 26072
rect 32678 25064 32734 25120
rect 32862 24928 32918 24984
rect 32954 24520 33010 24576
rect 32862 24112 32918 24168
rect 32862 24012 32864 24032
rect 32864 24012 32916 24032
rect 32916 24012 32918 24032
rect 32862 23976 32918 24012
rect 32494 23704 32550 23760
rect 32494 23024 32550 23080
rect 32402 22888 32458 22944
rect 32494 22616 32550 22672
rect 32402 22480 32458 22536
rect 32310 21800 32366 21856
rect 31850 20440 31906 20496
rect 31758 19352 31814 19408
rect 31574 18844 31576 18864
rect 31576 18844 31628 18864
rect 31628 18844 31630 18864
rect 31574 18808 31630 18844
rect 31942 19488 31998 19544
rect 32218 21120 32274 21176
rect 32310 20712 32366 20768
rect 32218 19624 32274 19680
rect 32862 23588 32918 23624
rect 32862 23568 32864 23588
rect 32864 23568 32916 23588
rect 32916 23568 32918 23588
rect 32862 23024 32918 23080
rect 32494 19896 32550 19952
rect 32494 19352 32550 19408
rect 32954 20748 32956 20768
rect 32956 20748 33008 20768
rect 33008 20748 33010 20768
rect 32954 20712 33010 20748
rect 32954 20440 33010 20496
rect 32770 20304 32826 20360
rect 32770 19624 32826 19680
rect 32218 18264 32274 18320
rect 32586 18672 32642 18728
rect 32586 18572 32588 18592
rect 32588 18572 32640 18592
rect 32640 18572 32642 18592
rect 32586 18536 32642 18572
rect 32678 18400 32734 18456
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 33230 23024 33286 23080
rect 33138 22888 33194 22944
rect 33506 27104 33562 27160
rect 33690 29028 33746 29064
rect 33690 29008 33692 29028
rect 33692 29008 33744 29028
rect 33744 29008 33746 29028
rect 33598 25064 33654 25120
rect 33506 24384 33562 24440
rect 33598 24112 33654 24168
rect 33506 23976 33562 24032
rect 33230 20576 33286 20632
rect 33046 19080 33102 19136
rect 33230 19896 33286 19952
rect 33230 19488 33286 19544
rect 33874 29960 33930 30016
rect 34058 29416 34114 29472
rect 34242 29144 34298 29200
rect 34518 32000 34574 32056
rect 34978 32816 35034 32872
rect 34702 32136 34758 32192
rect 34518 31748 34574 31784
rect 34518 31728 34520 31748
rect 34520 31728 34572 31748
rect 34572 31728 34574 31748
rect 34610 31628 34612 31648
rect 34612 31628 34664 31648
rect 34664 31628 34666 31648
rect 34610 31592 34666 31628
rect 34886 32272 34942 32328
rect 35070 32544 35126 32600
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35162 31864 35218 31920
rect 34978 31728 35034 31784
rect 34610 30232 34666 30288
rect 34794 31340 34850 31376
rect 34794 31320 34796 31340
rect 34796 31320 34848 31340
rect 34848 31320 34850 31340
rect 34978 31184 35034 31240
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 38014 38120 38070 38176
rect 35714 35672 35770 35728
rect 35622 35536 35678 35592
rect 35714 34196 35770 34232
rect 35714 34176 35716 34196
rect 35716 34176 35768 34196
rect 35768 34176 35770 34196
rect 35898 35128 35954 35184
rect 35898 34176 35954 34232
rect 36174 34484 36176 34504
rect 36176 34484 36228 34504
rect 36228 34484 36230 34504
rect 36174 34448 36230 34484
rect 35714 33768 35770 33824
rect 35622 33496 35678 33552
rect 35990 33940 35992 33960
rect 35992 33940 36044 33960
rect 36044 33940 36046 33960
rect 35990 33904 36046 33940
rect 35714 33224 35770 33280
rect 35714 32972 35770 33008
rect 35714 32952 35716 32972
rect 35716 32952 35768 32972
rect 35768 32952 35770 32972
rect 35438 31728 35494 31784
rect 34702 29960 34758 30016
rect 35438 29960 35494 30016
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 33782 25608 33838 25664
rect 34058 24928 34114 24984
rect 33690 23296 33746 23352
rect 33782 22888 33838 22944
rect 34058 23976 34114 24032
rect 33874 22344 33930 22400
rect 33598 20032 33654 20088
rect 33782 20984 33838 21040
rect 33138 18128 33194 18184
rect 33138 17992 33194 18048
rect 33322 17992 33378 18048
rect 33506 17992 33562 18048
rect 34426 28192 34482 28248
rect 34426 27920 34482 27976
rect 34426 27820 34428 27840
rect 34428 27820 34480 27840
rect 34480 27820 34482 27840
rect 34426 27784 34482 27820
rect 34610 28328 34666 28384
rect 34610 27648 34666 27704
rect 34518 27512 34574 27568
rect 35530 29708 35586 29744
rect 35530 29688 35532 29708
rect 35532 29688 35584 29708
rect 35584 29688 35586 29708
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34794 28736 34850 28792
rect 34886 28620 34942 28656
rect 34886 28600 34888 28620
rect 34888 28600 34940 28620
rect 34940 28600 34942 28620
rect 34794 28192 34850 28248
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35162 27512 35218 27568
rect 34518 25880 34574 25936
rect 34150 23432 34206 23488
rect 34242 21664 34298 21720
rect 33966 20712 34022 20768
rect 34242 20576 34298 20632
rect 33966 20168 34022 20224
rect 33874 19488 33930 19544
rect 33414 17720 33470 17776
rect 33690 17720 33746 17776
rect 33874 17992 33930 18048
rect 33690 17312 33746 17368
rect 34518 24112 34574 24168
rect 34426 22888 34482 22944
rect 34518 22344 34574 22400
rect 34610 22208 34666 22264
rect 34886 27240 34942 27296
rect 34978 26988 35034 27024
rect 34978 26968 34980 26988
rect 34980 26968 35032 26988
rect 35032 26968 35034 26988
rect 35438 27512 35494 27568
rect 35346 26696 35402 26752
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34886 26424 34942 26480
rect 35162 26424 35218 26480
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35254 25236 35256 25256
rect 35256 25236 35308 25256
rect 35308 25236 35310 25256
rect 35254 25200 35310 25236
rect 34886 24928 34942 24984
rect 35806 32544 35862 32600
rect 36266 33632 36322 33688
rect 35714 31184 35770 31240
rect 35806 30504 35862 30560
rect 35714 28600 35770 28656
rect 36082 32408 36138 32464
rect 36174 32000 36230 32056
rect 36542 36216 36598 36272
rect 36910 36080 36966 36136
rect 36634 35944 36690 36000
rect 36726 35012 36782 35048
rect 36726 34992 36728 35012
rect 36728 34992 36780 35012
rect 36780 34992 36782 35012
rect 36450 32272 36506 32328
rect 36450 31900 36452 31920
rect 36452 31900 36504 31920
rect 36504 31900 36506 31920
rect 36450 31864 36506 31900
rect 36266 29960 36322 30016
rect 35990 28328 36046 28384
rect 35714 26832 35770 26888
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35070 23976 35126 24032
rect 35254 23976 35310 24032
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35438 23724 35494 23760
rect 35438 23704 35440 23724
rect 35440 23704 35492 23724
rect 35492 23704 35494 23724
rect 34886 22480 34942 22536
rect 35346 22344 35402 22400
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35806 25336 35862 25392
rect 35714 24792 35770 24848
rect 35806 24656 35862 24712
rect 34426 20460 34482 20496
rect 34426 20440 34428 20460
rect 34428 20440 34480 20460
rect 34480 20440 34482 20460
rect 34150 18128 34206 18184
rect 35070 21972 35072 21992
rect 35072 21972 35124 21992
rect 35124 21972 35126 21992
rect 35070 21936 35126 21972
rect 35438 22072 35494 22128
rect 36174 27104 36230 27160
rect 36726 32000 36782 32056
rect 37462 37032 37518 37088
rect 38106 36624 38162 36680
rect 36910 32680 36966 32736
rect 36358 29552 36414 29608
rect 36358 27104 36414 27160
rect 36634 26968 36690 27024
rect 36082 25744 36138 25800
rect 36082 25064 36138 25120
rect 36174 23840 36230 23896
rect 35622 22344 35678 22400
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34978 20460 35034 20496
rect 34978 20440 34980 20460
rect 34980 20440 35032 20460
rect 35032 20440 35034 20460
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34610 19488 34666 19544
rect 35070 19796 35072 19816
rect 35072 19796 35124 19816
rect 35124 19796 35126 19816
rect 35070 19760 35126 19796
rect 34978 19372 35034 19408
rect 34978 19352 34981 19372
rect 34981 19352 35033 19372
rect 35033 19352 35034 19372
rect 35254 19352 35310 19408
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34610 16904 34666 16960
rect 35254 18128 35310 18184
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35622 18672 35678 18728
rect 35530 15408 35586 15464
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35806 19372 35862 19408
rect 35806 19352 35808 19372
rect 35808 19352 35860 19372
rect 35860 19352 35862 19372
rect 35806 18536 35862 18592
rect 35806 16768 35862 16824
rect 35990 20304 36046 20360
rect 37186 30676 37188 30696
rect 37188 30676 37240 30696
rect 37240 30676 37242 30696
rect 37186 30640 37242 30676
rect 37186 29688 37242 29744
rect 37094 29416 37150 29472
rect 37002 23060 37004 23080
rect 37004 23060 37056 23080
rect 37056 23060 37058 23080
rect 36818 22752 36874 22808
rect 36634 21528 36690 21584
rect 36266 16632 36322 16688
rect 36082 13404 36084 13424
rect 36084 13404 36136 13424
rect 36136 13404 36138 13424
rect 36082 13368 36138 13404
rect 36726 19624 36782 19680
rect 37002 23024 37058 23060
rect 36818 15272 36874 15328
rect 37646 33516 37702 33552
rect 37646 33496 37648 33516
rect 37648 33496 37700 33516
rect 37700 33496 37702 33516
rect 37462 28076 37518 28112
rect 37462 28056 37464 28076
rect 37464 28056 37516 28076
rect 37516 28056 37518 28076
rect 37370 26016 37426 26072
rect 37922 33224 37978 33280
rect 37830 32952 37886 33008
rect 38014 32544 38070 32600
rect 38198 34040 38254 34096
rect 37830 28872 37886 28928
rect 37278 23568 37334 23624
rect 37462 23160 37518 23216
rect 37646 20848 37702 20904
rect 37370 18808 37426 18864
rect 37370 16360 37426 16416
rect 37554 14340 37610 14376
rect 37554 14320 37556 14340
rect 37556 14320 37608 14340
rect 37608 14320 37610 14340
rect 38290 30796 38346 30832
rect 38290 30776 38292 30796
rect 38292 30776 38344 30796
rect 38344 30776 38346 30796
rect 38566 34720 38622 34776
rect 38750 30368 38806 30424
rect 38474 26016 38530 26072
rect 37830 17720 37886 17776
rect 38290 20712 38346 20768
rect 38474 20440 38530 20496
rect 38106 15136 38162 15192
rect 38106 11076 38162 11112
rect 38106 11056 38108 11076
rect 38108 11056 38160 11076
rect 38160 11056 38162 11076
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 38106 9696 38162 9752
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 37830 8472 37886 8528
rect 38934 24656 38990 24712
rect 38842 23296 38898 23352
rect 39026 21936 39082 21992
rect 38934 20576 38990 20632
rect 38842 19216 38898 19272
rect 38750 15544 38806 15600
rect 39026 19080 39082 19136
rect 39578 33360 39634 33416
rect 39486 29144 39542 29200
rect 39394 24248 39450 24304
rect 39210 21392 39266 21448
rect 39026 17856 39082 17912
rect 39026 16496 39082 16552
rect 39026 13776 39082 13832
rect 38290 12416 38346 12472
rect 39302 17040 39358 17096
rect 38106 8372 38108 8392
rect 38108 8372 38160 8392
rect 38160 8372 38162 8392
rect 38106 8336 38162 8372
rect 38106 6976 38162 7032
rect 37830 6840 37886 6896
rect 37370 6704 37426 6760
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 38106 5636 38162 5672
rect 38106 5616 38108 5636
rect 38108 5616 38160 5636
rect 38160 5616 38162 5636
rect 38106 4256 38162 4312
rect 38106 2932 38108 2952
rect 38108 2932 38160 2952
rect 38160 2932 38162 2952
rect 38106 2896 38162 2932
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37830 2488 37886 2544
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 38106 1536 38162 1592
<< metal3 >>
rect 22134 39340 22140 39404
rect 22204 39402 22210 39404
rect 35801 39402 35867 39405
rect 22204 39400 35867 39402
rect 22204 39344 35806 39400
rect 35862 39344 35867 39400
rect 22204 39342 35867 39344
rect 22204 39340 22210 39342
rect 35801 39339 35867 39342
rect 6821 39266 6887 39269
rect 27470 39266 27476 39268
rect 6821 39264 27476 39266
rect 6821 39208 6826 39264
rect 6882 39208 27476 39264
rect 6821 39206 27476 39208
rect 6821 39203 6887 39206
rect 27470 39204 27476 39206
rect 27540 39204 27546 39268
rect 11237 39130 11303 39133
rect 27286 39130 27292 39132
rect 11237 39128 27292 39130
rect 11237 39072 11242 39128
rect 11298 39072 27292 39128
rect 11237 39070 27292 39072
rect 11237 39067 11303 39070
rect 27286 39068 27292 39070
rect 27356 39068 27362 39132
rect 5349 38994 5415 38997
rect 12566 38994 12572 38996
rect 5349 38992 12572 38994
rect 5349 38936 5354 38992
rect 5410 38936 12572 38992
rect 5349 38934 12572 38936
rect 5349 38931 5415 38934
rect 12566 38932 12572 38934
rect 12636 38932 12642 38996
rect 22369 38994 22435 38997
rect 35617 38994 35683 38997
rect 22369 38992 35683 38994
rect 22369 38936 22374 38992
rect 22430 38936 35622 38992
rect 35678 38936 35683 38992
rect 22369 38934 35683 38936
rect 22369 38931 22435 38934
rect 35617 38931 35683 38934
rect 8753 38858 8819 38861
rect 30005 38858 30071 38861
rect 8753 38856 30071 38858
rect 8753 38800 8758 38856
rect 8814 38800 30010 38856
rect 30066 38800 30071 38856
rect 8753 38798 30071 38800
rect 8753 38795 8819 38798
rect 30005 38795 30071 38798
rect 4889 38722 4955 38725
rect 26417 38722 26483 38725
rect 4889 38720 26483 38722
rect 4889 38664 4894 38720
rect 4950 38664 26422 38720
rect 26478 38664 26483 38720
rect 4889 38662 26483 38664
rect 4889 38659 4955 38662
rect 26417 38659 26483 38662
rect 6453 38586 6519 38589
rect 27889 38586 27955 38589
rect 6453 38584 27955 38586
rect 6453 38528 6458 38584
rect 6514 38528 27894 38584
rect 27950 38528 27955 38584
rect 6453 38526 27955 38528
rect 6453 38523 6519 38526
rect 27889 38523 27955 38526
rect 8661 38450 8727 38453
rect 35525 38450 35591 38453
rect 8661 38448 35591 38450
rect 8661 38392 8666 38448
rect 8722 38392 35530 38448
rect 35586 38392 35591 38448
rect 8661 38390 35591 38392
rect 8661 38387 8727 38390
rect 35525 38387 35591 38390
rect 3601 38314 3667 38317
rect 27838 38314 27844 38316
rect 3601 38312 27844 38314
rect 3601 38256 3606 38312
rect 3662 38256 27844 38312
rect 3601 38254 27844 38256
rect 3601 38251 3667 38254
rect 27838 38252 27844 38254
rect 27908 38252 27914 38316
rect 35433 38314 35499 38317
rect 39200 38314 40000 38344
rect 35433 38312 40000 38314
rect 35433 38256 35438 38312
rect 35494 38256 40000 38312
rect 35433 38254 40000 38256
rect 35433 38251 35499 38254
rect 39200 38224 40000 38254
rect 11053 38178 11119 38181
rect 24669 38178 24735 38181
rect 11053 38176 24735 38178
rect 11053 38120 11058 38176
rect 11114 38120 24674 38176
rect 24730 38120 24735 38176
rect 11053 38118 24735 38120
rect 11053 38115 11119 38118
rect 24669 38115 24735 38118
rect 25865 38178 25931 38181
rect 38009 38178 38075 38181
rect 25865 38176 38075 38178
rect 25865 38120 25870 38176
rect 25926 38120 38014 38176
rect 38070 38120 38075 38176
rect 25865 38118 38075 38120
rect 25865 38115 25931 38118
rect 38009 38115 38075 38118
rect 9622 37980 9628 38044
rect 9692 38042 9698 38044
rect 30189 38042 30255 38045
rect 9692 38040 30255 38042
rect 9692 37984 30194 38040
rect 30250 37984 30255 38040
rect 9692 37982 30255 37984
rect 9692 37980 9698 37982
rect 30189 37979 30255 37982
rect 7373 37906 7439 37909
rect 30097 37906 30163 37909
rect 7373 37904 30163 37906
rect 7373 37848 7378 37904
rect 7434 37848 30102 37904
rect 30158 37848 30163 37904
rect 7373 37846 30163 37848
rect 7373 37843 7439 37846
rect 30097 37843 30163 37846
rect 5165 37770 5231 37773
rect 15377 37770 15443 37773
rect 16481 37772 16547 37773
rect 16430 37770 16436 37772
rect 5165 37768 15443 37770
rect 5165 37712 5170 37768
rect 5226 37712 15382 37768
rect 15438 37712 15443 37768
rect 5165 37710 15443 37712
rect 16354 37710 16436 37770
rect 16500 37770 16547 37772
rect 29310 37770 29316 37772
rect 16500 37768 29316 37770
rect 16542 37712 29316 37768
rect 5165 37707 5231 37710
rect 15377 37707 15443 37710
rect 16430 37708 16436 37710
rect 16500 37710 29316 37712
rect 16500 37708 16547 37710
rect 29310 37708 29316 37710
rect 29380 37708 29386 37772
rect 16481 37707 16547 37708
rect 8109 37634 8175 37637
rect 23422 37634 23428 37636
rect 8109 37632 23428 37634
rect 8109 37576 8114 37632
rect 8170 37576 23428 37632
rect 8109 37574 23428 37576
rect 8109 37571 8175 37574
rect 23422 37572 23428 37574
rect 23492 37572 23498 37636
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 12249 37498 12315 37501
rect 12249 37496 23490 37498
rect 12249 37440 12254 37496
rect 12310 37440 23490 37496
rect 12249 37438 23490 37440
rect 12249 37435 12315 37438
rect 4838 37300 4844 37364
rect 4908 37362 4914 37364
rect 5349 37362 5415 37365
rect 4908 37360 5415 37362
rect 4908 37304 5354 37360
rect 5410 37304 5415 37360
rect 4908 37302 5415 37304
rect 4908 37300 4914 37302
rect 5349 37299 5415 37302
rect 7097 37362 7163 37365
rect 19425 37362 19491 37365
rect 7097 37360 19491 37362
rect 7097 37304 7102 37360
rect 7158 37304 19430 37360
rect 19486 37304 19491 37360
rect 7097 37302 19491 37304
rect 7097 37299 7163 37302
rect 19425 37299 19491 37302
rect 20529 37362 20595 37365
rect 20989 37362 21055 37365
rect 20529 37360 21055 37362
rect 20529 37304 20534 37360
rect 20590 37304 20994 37360
rect 21050 37304 21055 37360
rect 20529 37302 21055 37304
rect 23430 37362 23490 37438
rect 23606 37436 23612 37500
rect 23676 37498 23682 37500
rect 28993 37498 29059 37501
rect 23676 37496 29059 37498
rect 23676 37440 28998 37496
rect 29054 37440 29059 37496
rect 23676 37438 29059 37440
rect 23676 37436 23682 37438
rect 28993 37435 29059 37438
rect 24485 37362 24551 37365
rect 23430 37360 24551 37362
rect 23430 37304 24490 37360
rect 24546 37304 24551 37360
rect 23430 37302 24551 37304
rect 20529 37299 20595 37302
rect 20989 37299 21055 37302
rect 24485 37299 24551 37302
rect 26918 37300 26924 37364
rect 26988 37362 26994 37364
rect 34697 37362 34763 37365
rect 26988 37360 34763 37362
rect 26988 37304 34702 37360
rect 34758 37304 34763 37360
rect 26988 37302 34763 37304
rect 26988 37300 26994 37302
rect 34697 37299 34763 37302
rect 17217 37226 17283 37229
rect 26141 37226 26207 37229
rect 17217 37224 26207 37226
rect 17217 37168 17222 37224
rect 17278 37168 26146 37224
rect 26202 37168 26207 37224
rect 17217 37166 26207 37168
rect 17217 37163 17283 37166
rect 26141 37163 26207 37166
rect 29637 37226 29703 37229
rect 32305 37226 32371 37229
rect 29637 37224 32371 37226
rect 29637 37168 29642 37224
rect 29698 37168 32310 37224
rect 32366 37168 32371 37224
rect 29637 37166 32371 37168
rect 29637 37163 29703 37166
rect 32305 37163 32371 37166
rect 13353 37090 13419 37093
rect 15929 37090 15995 37093
rect 13353 37088 15995 37090
rect 13353 37032 13358 37088
rect 13414 37032 15934 37088
rect 15990 37032 15995 37088
rect 13353 37030 15995 37032
rect 13353 37027 13419 37030
rect 15929 37027 15995 37030
rect 21633 37090 21699 37093
rect 37457 37090 37523 37093
rect 21633 37088 37523 37090
rect 21633 37032 21638 37088
rect 21694 37032 37462 37088
rect 37518 37032 37523 37088
rect 21633 37030 37523 37032
rect 21633 37027 21699 37030
rect 37457 37027 37523 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 5073 36954 5139 36957
rect 15101 36954 15167 36957
rect 5073 36952 15167 36954
rect 5073 36896 5078 36952
rect 5134 36896 15106 36952
rect 15162 36896 15167 36952
rect 5073 36894 15167 36896
rect 5073 36891 5139 36894
rect 15101 36891 15167 36894
rect 15326 36892 15332 36956
rect 15396 36954 15402 36956
rect 19333 36954 19399 36957
rect 15396 36952 19399 36954
rect 15396 36896 19338 36952
rect 19394 36896 19399 36952
rect 15396 36894 19399 36896
rect 15396 36892 15402 36894
rect 19333 36891 19399 36894
rect 23381 36954 23447 36957
rect 25497 36954 25563 36957
rect 23381 36952 25563 36954
rect 23381 36896 23386 36952
rect 23442 36896 25502 36952
rect 25558 36896 25563 36952
rect 23381 36894 25563 36896
rect 23381 36891 23447 36894
rect 25497 36891 25563 36894
rect 31845 36954 31911 36957
rect 35157 36954 35223 36957
rect 31845 36952 35223 36954
rect 31845 36896 31850 36952
rect 31906 36896 35162 36952
rect 35218 36896 35223 36952
rect 31845 36894 35223 36896
rect 31845 36891 31911 36894
rect 35157 36891 35223 36894
rect 35341 36954 35407 36957
rect 39200 36954 40000 36984
rect 35341 36952 40000 36954
rect 35341 36896 35346 36952
rect 35402 36896 40000 36952
rect 35341 36894 40000 36896
rect 35341 36891 35407 36894
rect 39200 36864 40000 36894
rect 5717 36818 5783 36821
rect 27613 36818 27679 36821
rect 5717 36816 27679 36818
rect 5717 36760 5722 36816
rect 5778 36760 27618 36816
rect 27674 36760 27679 36816
rect 5717 36758 27679 36760
rect 5717 36755 5783 36758
rect 27613 36755 27679 36758
rect 30097 36818 30163 36821
rect 32949 36818 33015 36821
rect 30097 36816 33015 36818
rect 30097 36760 30102 36816
rect 30158 36760 32954 36816
rect 33010 36760 33015 36816
rect 30097 36758 33015 36760
rect 30097 36755 30163 36758
rect 32949 36755 33015 36758
rect 5441 36682 5507 36685
rect 17217 36682 17283 36685
rect 5441 36680 17283 36682
rect 5441 36624 5446 36680
rect 5502 36624 17222 36680
rect 17278 36624 17283 36680
rect 5441 36622 17283 36624
rect 5441 36619 5507 36622
rect 17217 36619 17283 36622
rect 17401 36682 17467 36685
rect 21950 36682 21956 36684
rect 17401 36680 21956 36682
rect 17401 36624 17406 36680
rect 17462 36624 21956 36680
rect 17401 36622 21956 36624
rect 17401 36619 17467 36622
rect 21950 36620 21956 36622
rect 22020 36682 22026 36684
rect 22645 36682 22711 36685
rect 28717 36682 28783 36685
rect 22020 36680 22711 36682
rect 22020 36624 22650 36680
rect 22706 36624 22711 36680
rect 22020 36622 22711 36624
rect 22020 36620 22026 36622
rect 22645 36619 22711 36622
rect 22832 36680 28783 36682
rect 22832 36624 28722 36680
rect 28778 36624 28783 36680
rect 22832 36622 28783 36624
rect 7005 36546 7071 36549
rect 7230 36546 7236 36548
rect 7005 36544 7236 36546
rect 7005 36488 7010 36544
rect 7066 36488 7236 36544
rect 7005 36486 7236 36488
rect 7005 36483 7071 36486
rect 7230 36484 7236 36486
rect 7300 36484 7306 36548
rect 8385 36546 8451 36549
rect 18965 36546 19031 36549
rect 8385 36544 19031 36546
rect 8385 36488 8390 36544
rect 8446 36488 18970 36544
rect 19026 36488 19031 36544
rect 8385 36486 19031 36488
rect 8385 36483 8451 36486
rect 18965 36483 19031 36486
rect 19374 36484 19380 36548
rect 19444 36546 19450 36548
rect 22832 36546 22892 36622
rect 28717 36619 28783 36622
rect 31201 36682 31267 36685
rect 38101 36682 38167 36685
rect 31201 36680 38167 36682
rect 31201 36624 31206 36680
rect 31262 36624 38106 36680
rect 38162 36624 38167 36680
rect 31201 36622 38167 36624
rect 31201 36619 31267 36622
rect 38101 36619 38167 36622
rect 19444 36486 22892 36546
rect 23105 36546 23171 36549
rect 24894 36546 24900 36548
rect 23105 36544 24900 36546
rect 23105 36488 23110 36544
rect 23166 36488 24900 36544
rect 23105 36486 24900 36488
rect 19444 36484 19450 36486
rect 23105 36483 23171 36486
rect 24894 36484 24900 36486
rect 24964 36546 24970 36548
rect 25313 36546 25379 36549
rect 24964 36544 25379 36546
rect 24964 36488 25318 36544
rect 25374 36488 25379 36544
rect 24964 36486 25379 36488
rect 24964 36484 24970 36486
rect 25313 36483 25379 36486
rect 27429 36546 27495 36549
rect 34421 36546 34487 36549
rect 27429 36544 34487 36546
rect 27429 36488 27434 36544
rect 27490 36488 34426 36544
rect 34482 36488 34487 36544
rect 27429 36486 34487 36488
rect 27429 36483 27495 36486
rect 34421 36483 34487 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 4889 36410 4955 36413
rect 13261 36410 13327 36413
rect 4889 36408 13327 36410
rect 4889 36352 4894 36408
rect 4950 36352 13266 36408
rect 13322 36352 13327 36408
rect 4889 36350 13327 36352
rect 4889 36347 4955 36350
rect 13261 36347 13327 36350
rect 14549 36410 14615 36413
rect 20161 36412 20227 36413
rect 18270 36410 18276 36412
rect 14549 36408 18276 36410
rect 14549 36352 14554 36408
rect 14610 36352 18276 36408
rect 14549 36350 18276 36352
rect 14549 36347 14615 36350
rect 18270 36348 18276 36350
rect 18340 36348 18346 36412
rect 20110 36410 20116 36412
rect 20070 36350 20116 36410
rect 20180 36408 20227 36412
rect 33869 36410 33935 36413
rect 20222 36352 20227 36408
rect 20110 36348 20116 36350
rect 20180 36348 20227 36352
rect 20161 36347 20227 36348
rect 22050 36408 33935 36410
rect 22050 36352 33874 36408
rect 33930 36352 33935 36408
rect 22050 36350 33935 36352
rect 1669 36274 1735 36277
rect 16481 36274 16547 36277
rect 1669 36272 16547 36274
rect 1669 36216 1674 36272
rect 1730 36216 16486 36272
rect 16542 36216 16547 36272
rect 1669 36214 16547 36216
rect 1669 36211 1735 36214
rect 16481 36211 16547 36214
rect 17033 36274 17099 36277
rect 17718 36274 17724 36276
rect 17033 36272 17724 36274
rect 17033 36216 17038 36272
rect 17094 36216 17724 36272
rect 17033 36214 17724 36216
rect 17033 36211 17099 36214
rect 17718 36212 17724 36214
rect 17788 36212 17794 36276
rect 19333 36274 19399 36277
rect 22050 36274 22110 36350
rect 33869 36347 33935 36350
rect 19333 36272 22110 36274
rect 19333 36216 19338 36272
rect 19394 36216 22110 36272
rect 19333 36214 22110 36216
rect 19333 36211 19399 36214
rect 25262 36212 25268 36276
rect 25332 36274 25338 36276
rect 29177 36274 29243 36277
rect 25332 36272 29243 36274
rect 25332 36216 29182 36272
rect 29238 36216 29243 36272
rect 25332 36214 29243 36216
rect 25332 36212 25338 36214
rect 29177 36211 29243 36214
rect 32305 36274 32371 36277
rect 36537 36274 36603 36277
rect 32305 36272 36603 36274
rect 32305 36216 32310 36272
rect 32366 36216 36542 36272
rect 36598 36216 36603 36272
rect 32305 36214 36603 36216
rect 32305 36211 32371 36214
rect 36537 36211 36603 36214
rect 17309 36140 17375 36141
rect 17309 36136 17356 36140
rect 17420 36138 17426 36140
rect 22093 36138 22159 36141
rect 17309 36080 17314 36136
rect 17309 36076 17356 36080
rect 17420 36078 17466 36138
rect 17910 36136 22159 36138
rect 17910 36080 22098 36136
rect 22154 36080 22159 36136
rect 17910 36078 22159 36080
rect 17420 36076 17426 36078
rect 17309 36075 17375 36076
rect 6085 36004 6151 36005
rect 6085 36000 6132 36004
rect 6196 36002 6202 36004
rect 9673 36002 9739 36005
rect 12750 36002 12756 36004
rect 6085 35944 6090 36000
rect 6085 35940 6132 35944
rect 6196 35942 6242 36002
rect 9673 36000 12756 36002
rect 9673 35944 9678 36000
rect 9734 35944 12756 36000
rect 9673 35942 12756 35944
rect 6196 35940 6202 35942
rect 6085 35939 6151 35940
rect 9673 35939 9739 35942
rect 12750 35940 12756 35942
rect 12820 35940 12826 36004
rect 13629 36002 13695 36005
rect 17910 36002 17970 36078
rect 22093 36075 22159 36078
rect 23013 36138 23079 36141
rect 26182 36138 26188 36140
rect 23013 36136 26188 36138
rect 23013 36080 23018 36136
rect 23074 36080 26188 36136
rect 23013 36078 26188 36080
rect 23013 36075 23079 36078
rect 26182 36076 26188 36078
rect 26252 36076 26258 36140
rect 36905 36138 36971 36141
rect 31710 36136 36971 36138
rect 31710 36080 36910 36136
rect 36966 36080 36971 36136
rect 31710 36078 36971 36080
rect 13629 36000 17970 36002
rect 13629 35944 13634 36000
rect 13690 35944 17970 36000
rect 13629 35942 17970 35944
rect 18045 36002 18111 36005
rect 18965 36002 19031 36005
rect 18045 36000 19031 36002
rect 18045 35944 18050 36000
rect 18106 35944 18970 36000
rect 19026 35944 19031 36000
rect 18045 35942 19031 35944
rect 13629 35939 13695 35942
rect 18045 35939 18111 35942
rect 18965 35939 19031 35942
rect 22001 36002 22067 36005
rect 31710 36002 31770 36078
rect 36905 36075 36971 36078
rect 22001 36000 31770 36002
rect 22001 35944 22006 36000
rect 22062 35944 31770 36000
rect 22001 35942 31770 35944
rect 22001 35939 22067 35942
rect 33174 35940 33180 36004
rect 33244 36002 33250 36004
rect 36629 36002 36695 36005
rect 33244 36000 36695 36002
rect 33244 35944 36634 36000
rect 36690 35944 36695 36000
rect 33244 35942 36695 35944
rect 33244 35940 33250 35942
rect 36629 35939 36695 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4981 35866 5047 35869
rect 5165 35866 5231 35869
rect 4981 35864 5231 35866
rect 4981 35808 4986 35864
rect 5042 35808 5170 35864
rect 5226 35808 5231 35864
rect 4981 35806 5231 35808
rect 4981 35803 5047 35806
rect 5165 35803 5231 35806
rect 6545 35866 6611 35869
rect 9397 35866 9463 35869
rect 10225 35866 10291 35869
rect 10358 35866 10364 35868
rect 6545 35864 10364 35866
rect 6545 35808 6550 35864
rect 6606 35808 9402 35864
rect 9458 35808 10230 35864
rect 10286 35808 10364 35864
rect 6545 35806 10364 35808
rect 6545 35803 6611 35806
rect 9397 35803 9463 35806
rect 10225 35803 10291 35806
rect 10358 35804 10364 35806
rect 10428 35804 10434 35868
rect 16481 35866 16547 35869
rect 18086 35866 18092 35868
rect 16481 35864 18092 35866
rect 16481 35808 16486 35864
rect 16542 35808 18092 35864
rect 16481 35806 18092 35808
rect 16481 35803 16547 35806
rect 18086 35804 18092 35806
rect 18156 35866 18162 35868
rect 19241 35866 19307 35869
rect 18156 35864 19307 35866
rect 18156 35808 19246 35864
rect 19302 35808 19307 35864
rect 18156 35806 19307 35808
rect 18156 35804 18162 35806
rect 19241 35803 19307 35806
rect 21030 35804 21036 35868
rect 21100 35866 21106 35868
rect 24853 35866 24919 35869
rect 21100 35864 24919 35866
rect 21100 35808 24858 35864
rect 24914 35808 24919 35864
rect 21100 35806 24919 35808
rect 21100 35804 21106 35806
rect 24853 35803 24919 35806
rect 25221 35866 25287 35869
rect 27337 35866 27403 35869
rect 25221 35864 27403 35866
rect 25221 35808 25226 35864
rect 25282 35808 27342 35864
rect 27398 35808 27403 35864
rect 25221 35806 27403 35808
rect 25221 35803 25287 35806
rect 27337 35803 27403 35806
rect 27470 35804 27476 35868
rect 27540 35866 27546 35868
rect 28257 35866 28323 35869
rect 29821 35866 29887 35869
rect 27540 35864 29887 35866
rect 27540 35808 28262 35864
rect 28318 35808 29826 35864
rect 29882 35808 29887 35864
rect 27540 35806 29887 35808
rect 27540 35804 27546 35806
rect 28257 35803 28323 35806
rect 29821 35803 29887 35806
rect 32305 35866 32371 35869
rect 33961 35866 34027 35869
rect 32305 35864 34027 35866
rect 32305 35808 32310 35864
rect 32366 35808 33966 35864
rect 34022 35808 34027 35864
rect 32305 35806 34027 35808
rect 32305 35803 32371 35806
rect 33961 35803 34027 35806
rect 4337 35730 4403 35733
rect 23841 35730 23907 35733
rect 4337 35728 23907 35730
rect 4337 35672 4342 35728
rect 4398 35672 23846 35728
rect 23902 35672 23907 35728
rect 4337 35670 23907 35672
rect 4337 35667 4403 35670
rect 23841 35667 23907 35670
rect 23974 35668 23980 35732
rect 24044 35730 24050 35732
rect 24577 35730 24643 35733
rect 24044 35728 24643 35730
rect 24044 35672 24582 35728
rect 24638 35672 24643 35728
rect 24044 35670 24643 35672
rect 24044 35668 24050 35670
rect 24577 35667 24643 35670
rect 25773 35730 25839 35733
rect 26693 35730 26759 35733
rect 35709 35730 35775 35733
rect 25773 35728 26759 35730
rect 25773 35672 25778 35728
rect 25834 35672 26698 35728
rect 26754 35672 26759 35728
rect 25773 35670 26759 35672
rect 25773 35667 25839 35670
rect 26693 35667 26759 35670
rect 26926 35728 35775 35730
rect 26926 35672 35714 35728
rect 35770 35672 35775 35728
rect 26926 35670 35775 35672
rect 11697 35594 11763 35597
rect 15745 35594 15811 35597
rect 11697 35592 15811 35594
rect 11697 35536 11702 35592
rect 11758 35536 15750 35592
rect 15806 35536 15811 35592
rect 11697 35534 15811 35536
rect 11697 35531 11763 35534
rect 15745 35531 15811 35534
rect 17953 35594 18019 35597
rect 18781 35594 18847 35597
rect 26926 35594 26986 35670
rect 35709 35667 35775 35670
rect 17953 35592 26986 35594
rect 17953 35536 17958 35592
rect 18014 35536 18786 35592
rect 18842 35536 26986 35592
rect 17953 35534 26986 35536
rect 30281 35594 30347 35597
rect 34145 35596 34211 35597
rect 34094 35594 34100 35596
rect 30281 35592 34100 35594
rect 34164 35592 34211 35596
rect 30281 35536 30286 35592
rect 30342 35536 34100 35592
rect 34206 35536 34211 35592
rect 30281 35534 34100 35536
rect 17953 35531 18019 35534
rect 18781 35531 18847 35534
rect 30281 35531 30347 35534
rect 34094 35532 34100 35534
rect 34164 35532 34211 35536
rect 34145 35531 34211 35532
rect 35617 35594 35683 35597
rect 39200 35594 40000 35624
rect 35617 35592 40000 35594
rect 35617 35536 35622 35592
rect 35678 35536 40000 35592
rect 35617 35534 40000 35536
rect 35617 35531 35683 35534
rect 39200 35504 40000 35534
rect 7833 35458 7899 35461
rect 14365 35458 14431 35461
rect 15009 35458 15075 35461
rect 7833 35456 15075 35458
rect 7833 35400 7838 35456
rect 7894 35400 14370 35456
rect 14426 35400 15014 35456
rect 15070 35400 15075 35456
rect 7833 35398 15075 35400
rect 7833 35395 7899 35398
rect 14365 35395 14431 35398
rect 15009 35395 15075 35398
rect 15193 35458 15259 35461
rect 23105 35458 23171 35461
rect 15193 35456 23171 35458
rect 15193 35400 15198 35456
rect 15254 35400 23110 35456
rect 23166 35400 23171 35456
rect 15193 35398 23171 35400
rect 15193 35395 15259 35398
rect 23105 35395 23171 35398
rect 26049 35458 26115 35461
rect 27061 35458 27127 35461
rect 26049 35456 27127 35458
rect 26049 35400 26054 35456
rect 26110 35400 27066 35456
rect 27122 35400 27127 35456
rect 26049 35398 27127 35400
rect 26049 35395 26115 35398
rect 27061 35395 27127 35398
rect 30281 35458 30347 35461
rect 32305 35458 32371 35461
rect 33409 35458 33475 35461
rect 30281 35456 33475 35458
rect 30281 35400 30286 35456
rect 30342 35400 32310 35456
rect 32366 35400 33414 35456
rect 33470 35400 33475 35456
rect 30281 35398 33475 35400
rect 30281 35395 30347 35398
rect 32305 35395 32371 35398
rect 33409 35395 33475 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 13537 35322 13603 35325
rect 16205 35322 16271 35325
rect 13537 35320 16271 35322
rect 13537 35264 13542 35320
rect 13598 35264 16210 35320
rect 16266 35264 16271 35320
rect 13537 35262 16271 35264
rect 13537 35259 13603 35262
rect 16205 35259 16271 35262
rect 18270 35260 18276 35324
rect 18340 35322 18346 35324
rect 24301 35322 24367 35325
rect 26877 35322 26943 35325
rect 18340 35320 26943 35322
rect 18340 35264 24306 35320
rect 24362 35264 26882 35320
rect 26938 35264 26943 35320
rect 18340 35262 26943 35264
rect 18340 35260 18346 35262
rect 24301 35259 24367 35262
rect 26877 35259 26943 35262
rect 27337 35322 27403 35325
rect 29494 35322 29500 35324
rect 27337 35320 29500 35322
rect 27337 35264 27342 35320
rect 27398 35264 29500 35320
rect 27337 35262 29500 35264
rect 27337 35259 27403 35262
rect 29494 35260 29500 35262
rect 29564 35322 29570 35324
rect 33409 35322 33475 35325
rect 29564 35320 33475 35322
rect 29564 35264 33414 35320
rect 33470 35264 33475 35320
rect 29564 35262 33475 35264
rect 29564 35260 29570 35262
rect 33409 35259 33475 35262
rect 6821 35186 6887 35189
rect 30281 35186 30347 35189
rect 6821 35184 30347 35186
rect 6821 35128 6826 35184
rect 6882 35128 30286 35184
rect 30342 35128 30347 35184
rect 6821 35126 30347 35128
rect 6821 35123 6887 35126
rect 30281 35123 30347 35126
rect 30414 35124 30420 35188
rect 30484 35186 30490 35188
rect 33317 35186 33383 35189
rect 35893 35186 35959 35189
rect 30484 35184 33383 35186
rect 30484 35128 33322 35184
rect 33378 35128 33383 35184
rect 30484 35126 33383 35128
rect 30484 35124 30490 35126
rect 33317 35123 33383 35126
rect 33504 35184 35959 35186
rect 33504 35128 35898 35184
rect 35954 35128 35959 35184
rect 33504 35126 35959 35128
rect 10317 35050 10383 35053
rect 12525 35050 12591 35053
rect 10317 35048 12591 35050
rect 10317 34992 10322 35048
rect 10378 34992 12530 35048
rect 12586 34992 12591 35048
rect 10317 34990 12591 34992
rect 10317 34987 10383 34990
rect 12525 34987 12591 34990
rect 15745 35050 15811 35053
rect 19190 35050 19196 35052
rect 15745 35048 19196 35050
rect 15745 34992 15750 35048
rect 15806 34992 19196 35048
rect 15745 34990 19196 34992
rect 15745 34987 15811 34990
rect 19190 34988 19196 34990
rect 19260 34988 19266 35052
rect 23381 35050 23447 35053
rect 19428 35048 23447 35050
rect 19428 34992 23386 35048
rect 23442 34992 23447 35048
rect 19428 34990 23447 34992
rect 5165 34914 5231 34917
rect 13169 34914 13235 34917
rect 17401 34914 17467 34917
rect 5165 34912 12450 34914
rect 5165 34856 5170 34912
rect 5226 34856 12450 34912
rect 5165 34854 12450 34856
rect 5165 34851 5231 34854
rect 4797 34780 4863 34781
rect 4797 34778 4844 34780
rect 4752 34776 4844 34778
rect 4752 34720 4802 34776
rect 4752 34718 4844 34720
rect 4797 34716 4844 34718
rect 4908 34716 4914 34780
rect 5073 34778 5139 34781
rect 5206 34778 5212 34780
rect 5073 34776 5212 34778
rect 5073 34720 5078 34776
rect 5134 34720 5212 34776
rect 5073 34718 5212 34720
rect 4797 34715 4863 34716
rect 5073 34715 5139 34718
rect 5206 34716 5212 34718
rect 5276 34716 5282 34780
rect 7741 34778 7807 34781
rect 11881 34778 11947 34781
rect 12157 34780 12223 34781
rect 12157 34778 12204 34780
rect 7741 34776 11947 34778
rect 7741 34720 7746 34776
rect 7802 34720 11886 34776
rect 11942 34720 11947 34776
rect 7741 34718 11947 34720
rect 12112 34776 12204 34778
rect 12112 34720 12162 34776
rect 12112 34718 12204 34720
rect 7741 34715 7807 34718
rect 11881 34715 11947 34718
rect 12157 34716 12204 34718
rect 12268 34716 12274 34780
rect 12390 34778 12450 34854
rect 13169 34912 17467 34914
rect 13169 34856 13174 34912
rect 13230 34856 17406 34912
rect 17462 34856 17467 34912
rect 13169 34854 17467 34856
rect 13169 34851 13235 34854
rect 17401 34851 17467 34854
rect 17902 34852 17908 34916
rect 17972 34914 17978 34916
rect 18229 34914 18295 34917
rect 19428 34914 19488 34990
rect 23381 34987 23447 34990
rect 24894 34988 24900 35052
rect 24964 35050 24970 35052
rect 27245 35050 27311 35053
rect 24964 35048 27311 35050
rect 24964 34992 27250 35048
rect 27306 34992 27311 35048
rect 24964 34990 27311 34992
rect 24964 34988 24970 34990
rect 27245 34987 27311 34990
rect 27521 35050 27587 35053
rect 31753 35050 31819 35053
rect 27521 35048 31819 35050
rect 27521 34992 27526 35048
rect 27582 34992 31758 35048
rect 31814 34992 31819 35048
rect 27521 34990 31819 34992
rect 27521 34987 27587 34990
rect 31753 34987 31819 34990
rect 27337 34914 27403 34917
rect 17972 34912 18295 34914
rect 17972 34856 18234 34912
rect 18290 34856 18295 34912
rect 17972 34854 18295 34856
rect 17972 34852 17978 34854
rect 18229 34851 18295 34854
rect 19290 34854 19488 34914
rect 22050 34912 27403 34914
rect 22050 34856 27342 34912
rect 27398 34856 27403 34912
rect 22050 34854 27403 34856
rect 14733 34778 14799 34781
rect 12390 34776 14799 34778
rect 12390 34720 14738 34776
rect 14794 34720 14799 34776
rect 12390 34718 14799 34720
rect 12157 34715 12223 34716
rect 14733 34715 14799 34718
rect 15009 34778 15075 34781
rect 17309 34778 17375 34781
rect 19290 34778 19350 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 15009 34776 19350 34778
rect 15009 34720 15014 34776
rect 15070 34720 17314 34776
rect 17370 34720 19350 34776
rect 15009 34718 19350 34720
rect 15009 34715 15075 34718
rect 17309 34715 17375 34718
rect 4337 34642 4403 34645
rect 5073 34642 5139 34645
rect 4337 34640 5139 34642
rect 4337 34584 4342 34640
rect 4398 34584 5078 34640
rect 5134 34584 5139 34640
rect 4337 34582 5139 34584
rect 4337 34579 4403 34582
rect 5073 34579 5139 34582
rect 7005 34642 7071 34645
rect 7833 34642 7899 34645
rect 8201 34644 8267 34645
rect 8150 34642 8156 34644
rect 7005 34640 7899 34642
rect 7005 34584 7010 34640
rect 7066 34584 7838 34640
rect 7894 34584 7899 34640
rect 7005 34582 7899 34584
rect 8110 34582 8156 34642
rect 8220 34640 8267 34644
rect 8262 34584 8267 34640
rect 7005 34579 7071 34582
rect 7833 34579 7899 34582
rect 8150 34580 8156 34582
rect 8220 34580 8267 34584
rect 8201 34579 8267 34580
rect 9673 34642 9739 34645
rect 11094 34642 11100 34644
rect 9673 34640 11100 34642
rect 9673 34584 9678 34640
rect 9734 34584 11100 34640
rect 9673 34582 11100 34584
rect 9673 34579 9739 34582
rect 11094 34580 11100 34582
rect 11164 34580 11170 34644
rect 11278 34580 11284 34644
rect 11348 34642 11354 34644
rect 14917 34642 14983 34645
rect 11348 34640 14983 34642
rect 11348 34584 14922 34640
rect 14978 34584 14983 34640
rect 11348 34582 14983 34584
rect 11348 34580 11354 34582
rect 14917 34579 14983 34582
rect 15929 34642 15995 34645
rect 22050 34642 22110 34854
rect 27337 34851 27403 34854
rect 27889 34914 27955 34917
rect 28533 34914 28599 34917
rect 27889 34912 28599 34914
rect 27889 34856 27894 34912
rect 27950 34856 28538 34912
rect 28594 34856 28599 34912
rect 27889 34854 28599 34856
rect 27889 34851 27955 34854
rect 28533 34851 28599 34854
rect 28901 34914 28967 34917
rect 30741 34914 30807 34917
rect 31569 34914 31635 34917
rect 33504 34914 33564 35126
rect 35893 35123 35959 35126
rect 34237 35050 34303 35053
rect 36721 35050 36787 35053
rect 34237 35048 36787 35050
rect 34237 34992 34242 35048
rect 34298 34992 36726 35048
rect 36782 34992 36787 35048
rect 34237 34990 36787 34992
rect 34237 34987 34303 34990
rect 36721 34987 36787 34990
rect 28901 34912 31402 34914
rect 28901 34856 28906 34912
rect 28962 34856 30746 34912
rect 30802 34856 31402 34912
rect 28901 34854 31402 34856
rect 28901 34851 28967 34854
rect 30741 34851 30807 34854
rect 25129 34778 25195 34781
rect 26509 34778 26575 34781
rect 27889 34780 27955 34781
rect 15929 34640 22110 34642
rect 15929 34584 15934 34640
rect 15990 34584 22110 34640
rect 15929 34582 22110 34584
rect 22188 34776 26575 34778
rect 22188 34720 25134 34776
rect 25190 34720 26514 34776
rect 26570 34720 26575 34776
rect 22188 34718 26575 34720
rect 15929 34579 15995 34582
rect 10777 34506 10843 34509
rect 15285 34506 15351 34509
rect 10777 34504 15351 34506
rect 10777 34448 10782 34504
rect 10838 34448 15290 34504
rect 15346 34448 15351 34504
rect 10777 34446 15351 34448
rect 10777 34443 10843 34446
rect 15285 34443 15351 34446
rect 15837 34506 15903 34509
rect 16389 34506 16455 34509
rect 15837 34504 16455 34506
rect 15837 34448 15842 34504
rect 15898 34448 16394 34504
rect 16450 34448 16455 34504
rect 15837 34446 16455 34448
rect 15837 34443 15903 34446
rect 16389 34443 16455 34446
rect 19609 34506 19675 34509
rect 22188 34506 22248 34718
rect 25129 34715 25195 34718
rect 26509 34715 26575 34718
rect 27838 34716 27844 34780
rect 27908 34778 27955 34780
rect 28349 34778 28415 34781
rect 30741 34778 30807 34781
rect 27908 34776 28000 34778
rect 27950 34720 28000 34776
rect 27908 34718 28000 34720
rect 28349 34776 30807 34778
rect 28349 34720 28354 34776
rect 28410 34720 30746 34776
rect 30802 34720 30807 34776
rect 28349 34718 30807 34720
rect 31342 34778 31402 34854
rect 31569 34912 33564 34914
rect 31569 34856 31574 34912
rect 31630 34856 33564 34912
rect 31569 34854 33564 34856
rect 35433 34914 35499 34917
rect 36118 34914 36124 34916
rect 35433 34912 36124 34914
rect 35433 34856 35438 34912
rect 35494 34856 36124 34912
rect 35433 34854 36124 34856
rect 31569 34851 31635 34854
rect 35433 34851 35499 34854
rect 36118 34852 36124 34854
rect 36188 34852 36194 34916
rect 32029 34778 32095 34781
rect 38561 34778 38627 34781
rect 31342 34776 32095 34778
rect 31342 34720 32034 34776
rect 32090 34720 32095 34776
rect 31342 34718 32095 34720
rect 27908 34716 27955 34718
rect 27889 34715 27955 34716
rect 28349 34715 28415 34718
rect 30741 34715 30807 34718
rect 32029 34715 32095 34718
rect 32446 34776 38627 34778
rect 32446 34720 38566 34776
rect 38622 34720 38627 34776
rect 32446 34718 38627 34720
rect 23238 34580 23244 34644
rect 23308 34642 23314 34644
rect 23381 34642 23447 34645
rect 28993 34642 29059 34645
rect 23308 34640 23447 34642
rect 23308 34584 23386 34640
rect 23442 34584 23447 34640
rect 23308 34582 23447 34584
rect 23308 34580 23314 34582
rect 23381 34579 23447 34582
rect 23614 34640 29059 34642
rect 23614 34584 28998 34640
rect 29054 34584 29059 34640
rect 23614 34582 29059 34584
rect 19609 34504 22248 34506
rect 19609 34448 19614 34504
rect 19670 34448 22248 34504
rect 19609 34446 22248 34448
rect 23289 34506 23355 34509
rect 23614 34506 23674 34582
rect 28993 34579 29059 34582
rect 29453 34642 29519 34645
rect 29678 34642 29684 34644
rect 29453 34640 29684 34642
rect 29453 34584 29458 34640
rect 29514 34584 29684 34640
rect 29453 34582 29684 34584
rect 29453 34579 29519 34582
rect 29678 34580 29684 34582
rect 29748 34642 29754 34644
rect 31937 34642 32003 34645
rect 29748 34640 32003 34642
rect 29748 34584 31942 34640
rect 31998 34584 32003 34640
rect 29748 34582 32003 34584
rect 29748 34580 29754 34582
rect 31937 34579 32003 34582
rect 23289 34504 23674 34506
rect 23289 34448 23294 34504
rect 23350 34448 23674 34504
rect 23289 34446 23674 34448
rect 30649 34506 30715 34509
rect 32446 34506 32506 34718
rect 38561 34715 38627 34718
rect 32673 34642 32739 34645
rect 37038 34642 37044 34644
rect 32673 34640 37044 34642
rect 32673 34584 32678 34640
rect 32734 34584 37044 34640
rect 32673 34582 37044 34584
rect 32673 34579 32739 34582
rect 37038 34580 37044 34582
rect 37108 34580 37114 34644
rect 32673 34506 32739 34509
rect 30649 34504 32368 34506
rect 30649 34448 30654 34504
rect 30710 34448 32368 34504
rect 30649 34446 32368 34448
rect 32446 34504 32739 34506
rect 32446 34448 32678 34504
rect 32734 34448 32739 34504
rect 32446 34446 32739 34448
rect 19609 34443 19675 34446
rect 23289 34443 23355 34446
rect 30649 34443 30715 34446
rect 4613 34370 4679 34373
rect 22737 34370 22803 34373
rect 4613 34368 22803 34370
rect 4613 34312 4618 34368
rect 4674 34312 22742 34368
rect 22798 34312 22803 34368
rect 4613 34310 22803 34312
rect 4613 34307 4679 34310
rect 22737 34307 22803 34310
rect 23422 34308 23428 34372
rect 23492 34370 23498 34372
rect 26141 34370 26207 34373
rect 29821 34370 29887 34373
rect 23492 34368 29887 34370
rect 23492 34312 26146 34368
rect 26202 34312 29826 34368
rect 29882 34312 29887 34368
rect 23492 34310 29887 34312
rect 23492 34308 23498 34310
rect 26141 34307 26207 34310
rect 29821 34307 29887 34310
rect 30782 34308 30788 34372
rect 30852 34370 30858 34372
rect 32121 34370 32187 34373
rect 30852 34368 32187 34370
rect 30852 34312 32126 34368
rect 32182 34312 32187 34368
rect 30852 34310 32187 34312
rect 32308 34370 32368 34446
rect 32673 34443 32739 34446
rect 33225 34506 33291 34509
rect 36169 34506 36235 34509
rect 33225 34504 36235 34506
rect 33225 34448 33230 34504
rect 33286 34448 36174 34504
rect 36230 34448 36235 34504
rect 33225 34446 36235 34448
rect 33225 34443 33291 34446
rect 36169 34443 36235 34446
rect 34605 34370 34671 34373
rect 32308 34368 34671 34370
rect 32308 34312 34610 34368
rect 34666 34312 34671 34368
rect 32308 34310 34671 34312
rect 30852 34308 30858 34310
rect 32121 34307 32187 34310
rect 34605 34307 34671 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 7741 34234 7807 34237
rect 9622 34234 9628 34236
rect 7741 34232 9628 34234
rect 7741 34176 7746 34232
rect 7802 34176 9628 34232
rect 7741 34174 9628 34176
rect 7741 34171 7807 34174
rect 9622 34172 9628 34174
rect 9692 34172 9698 34236
rect 11053 34234 11119 34237
rect 15561 34234 15627 34237
rect 11053 34232 15627 34234
rect 11053 34176 11058 34232
rect 11114 34176 15566 34232
rect 15622 34176 15627 34232
rect 11053 34174 15627 34176
rect 11053 34171 11119 34174
rect 15561 34171 15627 34174
rect 16389 34234 16455 34237
rect 25497 34234 25563 34237
rect 26233 34236 26299 34237
rect 16389 34232 25563 34234
rect 16389 34176 16394 34232
rect 16450 34176 25502 34232
rect 25558 34176 25563 34232
rect 16389 34174 25563 34176
rect 16389 34171 16455 34174
rect 25497 34171 25563 34174
rect 26182 34172 26188 34236
rect 26252 34234 26299 34236
rect 30465 34234 30531 34237
rect 30649 34234 30715 34237
rect 32857 34234 32923 34237
rect 26252 34232 30715 34234
rect 26294 34176 30470 34232
rect 30526 34176 30654 34232
rect 30710 34176 30715 34232
rect 26252 34174 30715 34176
rect 26252 34172 26299 34174
rect 26233 34171 26299 34172
rect 30465 34171 30531 34174
rect 30649 34171 30715 34174
rect 30790 34232 32923 34234
rect 30790 34176 32862 34232
rect 32918 34176 32923 34232
rect 30790 34174 32923 34176
rect 5809 34098 5875 34101
rect 13537 34098 13603 34101
rect 13813 34098 13879 34101
rect 5809 34096 13603 34098
rect 5809 34040 5814 34096
rect 5870 34040 13542 34096
rect 13598 34040 13603 34096
rect 5809 34038 13603 34040
rect 5809 34035 5875 34038
rect 13537 34035 13603 34038
rect 13678 34096 13879 34098
rect 13678 34040 13818 34096
rect 13874 34040 13879 34096
rect 13678 34038 13879 34040
rect 7281 33962 7347 33965
rect 11697 33962 11763 33965
rect 7281 33960 11763 33962
rect 7281 33904 7286 33960
rect 7342 33904 11702 33960
rect 11758 33904 11763 33960
rect 7281 33902 11763 33904
rect 7281 33899 7347 33902
rect 11697 33899 11763 33902
rect 11973 33962 12039 33965
rect 13678 33962 13738 34038
rect 13813 34035 13879 34038
rect 14917 34098 14983 34101
rect 17861 34098 17927 34101
rect 14917 34096 17927 34098
rect 14917 34040 14922 34096
rect 14978 34040 17866 34096
rect 17922 34040 17927 34096
rect 14917 34038 17927 34040
rect 14917 34035 14983 34038
rect 17861 34035 17927 34038
rect 19425 34098 19491 34101
rect 26325 34098 26391 34101
rect 19425 34096 26391 34098
rect 19425 34040 19430 34096
rect 19486 34040 26330 34096
rect 26386 34040 26391 34096
rect 19425 34038 26391 34040
rect 19425 34035 19491 34038
rect 26325 34035 26391 34038
rect 26877 34098 26943 34101
rect 28441 34098 28507 34101
rect 26877 34096 28507 34098
rect 26877 34040 26882 34096
rect 26938 34040 28446 34096
rect 28502 34040 28507 34096
rect 26877 34038 28507 34040
rect 26877 34035 26943 34038
rect 28441 34035 28507 34038
rect 28993 34098 29059 34101
rect 30790 34098 30850 34174
rect 32857 34171 32923 34174
rect 33041 34234 33107 34237
rect 33726 34234 33732 34236
rect 33041 34232 33732 34234
rect 33041 34176 33046 34232
rect 33102 34176 33732 34232
rect 33041 34174 33732 34176
rect 33041 34171 33107 34174
rect 33726 34172 33732 34174
rect 33796 34172 33802 34236
rect 34053 34234 34119 34237
rect 34278 34234 34284 34236
rect 34053 34232 34284 34234
rect 34053 34176 34058 34232
rect 34114 34176 34284 34232
rect 34053 34174 34284 34176
rect 34053 34171 34119 34174
rect 34278 34172 34284 34174
rect 34348 34172 34354 34236
rect 35566 34172 35572 34236
rect 35636 34234 35642 34236
rect 35709 34234 35775 34237
rect 35636 34232 35775 34234
rect 35636 34176 35714 34232
rect 35770 34176 35775 34232
rect 35636 34174 35775 34176
rect 35636 34172 35642 34174
rect 35709 34171 35775 34174
rect 35893 34234 35959 34237
rect 39200 34234 40000 34264
rect 35893 34232 40000 34234
rect 35893 34176 35898 34232
rect 35954 34176 40000 34232
rect 35893 34174 40000 34176
rect 35893 34171 35959 34174
rect 39200 34144 40000 34174
rect 28993 34096 30850 34098
rect 28993 34040 28998 34096
rect 29054 34040 30850 34096
rect 28993 34038 30850 34040
rect 31753 34098 31819 34101
rect 38193 34098 38259 34101
rect 31753 34096 38259 34098
rect 31753 34040 31758 34096
rect 31814 34040 38198 34096
rect 38254 34040 38259 34096
rect 31753 34038 38259 34040
rect 28993 34035 29059 34038
rect 31753 34035 31819 34038
rect 38193 34035 38259 34038
rect 11973 33960 13738 33962
rect 11973 33904 11978 33960
rect 12034 33904 13738 33960
rect 11973 33902 13738 33904
rect 13905 33962 13971 33965
rect 16297 33962 16363 33965
rect 13905 33960 16363 33962
rect 13905 33904 13910 33960
rect 13966 33904 16302 33960
rect 16358 33904 16363 33960
rect 13905 33902 16363 33904
rect 11973 33899 12039 33902
rect 13905 33899 13971 33902
rect 16297 33899 16363 33902
rect 19977 33962 20043 33965
rect 22093 33962 22159 33965
rect 19977 33960 22159 33962
rect 19977 33904 19982 33960
rect 20038 33904 22098 33960
rect 22154 33904 22159 33960
rect 19977 33902 22159 33904
rect 19977 33899 20043 33902
rect 22093 33899 22159 33902
rect 22461 33962 22527 33965
rect 29361 33962 29427 33965
rect 22461 33960 29427 33962
rect 22461 33904 22466 33960
rect 22522 33904 29366 33960
rect 29422 33904 29427 33960
rect 22461 33902 29427 33904
rect 22461 33899 22527 33902
rect 29361 33899 29427 33902
rect 29545 33962 29611 33965
rect 35985 33962 36051 33965
rect 29545 33960 36051 33962
rect 29545 33904 29550 33960
rect 29606 33904 35990 33960
rect 36046 33904 36051 33960
rect 29545 33902 36051 33904
rect 29545 33899 29611 33902
rect 35985 33899 36051 33902
rect 5441 33826 5507 33829
rect 14365 33826 14431 33829
rect 5441 33824 14431 33826
rect 5441 33768 5446 33824
rect 5502 33768 14370 33824
rect 14426 33768 14431 33824
rect 5441 33766 14431 33768
rect 5441 33763 5507 33766
rect 14365 33763 14431 33766
rect 20713 33826 20779 33829
rect 28993 33826 29059 33829
rect 35709 33826 35775 33829
rect 20713 33824 29059 33826
rect 20713 33768 20718 33824
rect 20774 33768 28998 33824
rect 29054 33768 29059 33824
rect 20713 33766 29059 33768
rect 20713 33763 20779 33766
rect 28993 33763 29059 33766
rect 31710 33824 35775 33826
rect 31710 33768 35714 33824
rect 35770 33768 35775 33824
rect 31710 33766 35775 33768
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 6545 33690 6611 33693
rect 8477 33690 8543 33693
rect 6545 33688 8543 33690
rect 6545 33632 6550 33688
rect 6606 33632 8482 33688
rect 8538 33632 8543 33688
rect 6545 33630 8543 33632
rect 6545 33627 6611 33630
rect 8477 33627 8543 33630
rect 9949 33690 10015 33693
rect 18413 33690 18479 33693
rect 9949 33688 18479 33690
rect 9949 33632 9954 33688
rect 10010 33632 18418 33688
rect 18474 33632 18479 33688
rect 9949 33630 18479 33632
rect 9949 33627 10015 33630
rect 18413 33627 18479 33630
rect 20069 33690 20135 33693
rect 22277 33690 22343 33693
rect 27521 33690 27587 33693
rect 20069 33688 22343 33690
rect 20069 33632 20074 33688
rect 20130 33632 22282 33688
rect 22338 33632 22343 33688
rect 20069 33630 22343 33632
rect 20069 33627 20135 33630
rect 22277 33627 22343 33630
rect 25270 33688 27587 33690
rect 25270 33632 27526 33688
rect 27582 33632 27587 33688
rect 25270 33630 27587 33632
rect 6637 33554 6703 33557
rect 7097 33554 7163 33557
rect 6637 33552 7163 33554
rect 6637 33496 6642 33552
rect 6698 33496 7102 33552
rect 7158 33496 7163 33552
rect 6637 33494 7163 33496
rect 6637 33491 6703 33494
rect 7097 33491 7163 33494
rect 11697 33554 11763 33557
rect 25270 33554 25330 33630
rect 27521 33627 27587 33630
rect 30649 33690 30715 33693
rect 31334 33690 31340 33692
rect 30649 33688 31340 33690
rect 30649 33632 30654 33688
rect 30710 33632 31340 33688
rect 30649 33630 31340 33632
rect 30649 33627 30715 33630
rect 31334 33628 31340 33630
rect 31404 33690 31410 33692
rect 31710 33690 31770 33766
rect 35709 33763 35775 33766
rect 31404 33630 31770 33690
rect 31937 33690 32003 33693
rect 33317 33690 33383 33693
rect 31937 33688 33383 33690
rect 31937 33632 31942 33688
rect 31998 33632 33322 33688
rect 33378 33632 33383 33688
rect 31937 33630 33383 33632
rect 31404 33628 31410 33630
rect 31937 33627 32003 33630
rect 33317 33627 33383 33630
rect 33593 33690 33659 33693
rect 35934 33690 35940 33692
rect 33593 33688 35940 33690
rect 33593 33632 33598 33688
rect 33654 33632 35940 33688
rect 33593 33630 35940 33632
rect 33593 33627 33659 33630
rect 35934 33628 35940 33630
rect 36004 33690 36010 33692
rect 36261 33690 36327 33693
rect 36004 33688 36327 33690
rect 36004 33632 36266 33688
rect 36322 33632 36327 33688
rect 36004 33630 36327 33632
rect 36004 33628 36010 33630
rect 36261 33627 36327 33630
rect 11697 33552 25330 33554
rect 11697 33496 11702 33552
rect 11758 33496 25330 33552
rect 11697 33494 25330 33496
rect 25405 33554 25471 33557
rect 27337 33556 27403 33557
rect 25405 33552 27216 33554
rect 25405 33496 25410 33552
rect 25466 33496 27216 33552
rect 25405 33494 27216 33496
rect 11697 33491 11763 33494
rect 25405 33491 25471 33494
rect 7557 33418 7623 33421
rect 12065 33418 12131 33421
rect 23974 33418 23980 33420
rect 7557 33416 23980 33418
rect 7557 33360 7562 33416
rect 7618 33360 12070 33416
rect 12126 33360 23980 33416
rect 7557 33358 23980 33360
rect 7557 33355 7623 33358
rect 12065 33355 12131 33358
rect 23974 33356 23980 33358
rect 24044 33356 24050 33420
rect 24209 33418 24275 33421
rect 26417 33418 26483 33421
rect 24209 33416 26483 33418
rect 24209 33360 24214 33416
rect 24270 33360 26422 33416
rect 26478 33360 26483 33416
rect 24209 33358 26483 33360
rect 24209 33355 24275 33358
rect 26417 33355 26483 33358
rect 5809 33282 5875 33285
rect 6310 33282 6316 33284
rect 5809 33280 6316 33282
rect 5809 33224 5814 33280
rect 5870 33224 6316 33280
rect 5809 33222 6316 33224
rect 5809 33219 5875 33222
rect 6310 33220 6316 33222
rect 6380 33220 6386 33284
rect 11145 33282 11211 33285
rect 12065 33282 12131 33285
rect 15837 33282 15903 33285
rect 11145 33280 12131 33282
rect 11145 33224 11150 33280
rect 11206 33224 12070 33280
rect 12126 33224 12131 33280
rect 11145 33222 12131 33224
rect 11145 33219 11211 33222
rect 12065 33219 12131 33222
rect 13310 33280 15903 33282
rect 13310 33224 15842 33280
rect 15898 33224 15903 33280
rect 13310 33222 15903 33224
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 13310 33149 13370 33222
rect 15837 33219 15903 33222
rect 16849 33282 16915 33285
rect 20805 33284 20871 33285
rect 26325 33284 26391 33285
rect 16849 33280 19350 33282
rect 16849 33224 16854 33280
rect 16910 33224 19350 33280
rect 16849 33222 19350 33224
rect 16849 33219 16915 33222
rect 6637 33146 6703 33149
rect 6637 33144 11714 33146
rect 6637 33088 6642 33144
rect 6698 33088 11714 33144
rect 6637 33086 11714 33088
rect 6637 33083 6703 33086
rect 6913 33010 6979 33013
rect 10409 33010 10475 33013
rect 6913 33008 10475 33010
rect 6913 32952 6918 33008
rect 6974 32952 10414 33008
rect 10470 32952 10475 33008
rect 6913 32950 10475 32952
rect 6913 32947 6979 32950
rect 10409 32947 10475 32950
rect 4981 32874 5047 32877
rect 9765 32874 9831 32877
rect 10685 32874 10751 32877
rect 4981 32872 10751 32874
rect 4981 32816 4986 32872
rect 5042 32816 9770 32872
rect 9826 32816 10690 32872
rect 10746 32816 10751 32872
rect 4981 32814 10751 32816
rect 11654 32874 11714 33086
rect 13261 33144 13370 33149
rect 13261 33088 13266 33144
rect 13322 33088 13370 33144
rect 13261 33086 13370 33088
rect 13813 33146 13879 33149
rect 18229 33146 18295 33149
rect 13813 33144 18295 33146
rect 13813 33088 13818 33144
rect 13874 33088 18234 33144
rect 18290 33088 18295 33144
rect 13813 33086 18295 33088
rect 19290 33146 19350 33222
rect 20805 33280 20852 33284
rect 20916 33282 20922 33284
rect 20805 33224 20810 33280
rect 20805 33220 20852 33224
rect 20916 33222 20962 33282
rect 21912 33222 24824 33282
rect 20916 33220 20922 33222
rect 20805 33219 20871 33220
rect 21912 33146 21972 33222
rect 24577 33146 24643 33149
rect 19290 33086 21972 33146
rect 22050 33144 24643 33146
rect 22050 33088 24582 33144
rect 24638 33088 24643 33144
rect 22050 33086 24643 33088
rect 24764 33146 24824 33222
rect 26325 33280 26372 33284
rect 26436 33282 26442 33284
rect 27156 33282 27216 33494
rect 27286 33492 27292 33556
rect 27356 33554 27403 33556
rect 28901 33554 28967 33557
rect 33910 33554 33916 33556
rect 27356 33552 27448 33554
rect 27398 33496 27448 33552
rect 27356 33494 27448 33496
rect 28901 33552 33916 33554
rect 28901 33496 28906 33552
rect 28962 33496 33916 33552
rect 28901 33494 33916 33496
rect 27356 33492 27403 33494
rect 27337 33491 27403 33492
rect 28901 33491 28967 33494
rect 33910 33492 33916 33494
rect 33980 33492 33986 33556
rect 35249 33554 35315 33557
rect 35617 33554 35683 33557
rect 37641 33554 37707 33557
rect 35249 33552 37707 33554
rect 35249 33496 35254 33552
rect 35310 33496 35622 33552
rect 35678 33496 37646 33552
rect 37702 33496 37707 33552
rect 35249 33494 37707 33496
rect 35249 33491 35315 33494
rect 35617 33491 35683 33494
rect 37641 33491 37707 33494
rect 27470 33356 27476 33420
rect 27540 33418 27546 33420
rect 30373 33418 30439 33421
rect 32305 33418 32371 33421
rect 27540 33416 30439 33418
rect 27540 33360 30378 33416
rect 30434 33360 30439 33416
rect 27540 33358 30439 33360
rect 27540 33356 27546 33358
rect 30373 33355 30439 33358
rect 30606 33416 32371 33418
rect 30606 33360 32310 33416
rect 32366 33360 32371 33416
rect 30606 33358 32371 33360
rect 28206 33282 28212 33284
rect 26325 33224 26330 33280
rect 26325 33220 26372 33224
rect 26436 33222 26482 33282
rect 27156 33222 28212 33282
rect 26436 33220 26442 33222
rect 28206 33220 28212 33222
rect 28276 33282 28282 33284
rect 28533 33282 28599 33285
rect 28276 33280 28599 33282
rect 28276 33224 28538 33280
rect 28594 33224 28599 33280
rect 28276 33222 28599 33224
rect 28276 33220 28282 33222
rect 26325 33219 26391 33220
rect 28533 33219 28599 33222
rect 28942 33220 28948 33284
rect 29012 33282 29018 33284
rect 29085 33282 29151 33285
rect 29012 33280 29151 33282
rect 29012 33224 29090 33280
rect 29146 33224 29151 33280
rect 29012 33222 29151 33224
rect 29012 33220 29018 33222
rect 29085 33219 29151 33222
rect 30189 33282 30255 33285
rect 30606 33282 30666 33358
rect 32305 33355 32371 33358
rect 33409 33418 33475 33421
rect 35065 33418 35131 33421
rect 39573 33418 39639 33421
rect 33409 33416 39639 33418
rect 33409 33360 33414 33416
rect 33470 33360 35070 33416
rect 35126 33360 39578 33416
rect 39634 33360 39639 33416
rect 33409 33358 39639 33360
rect 33409 33355 33475 33358
rect 35065 33355 35131 33358
rect 39573 33355 39639 33358
rect 33174 33282 33180 33284
rect 30189 33280 30666 33282
rect 30189 33224 30194 33280
rect 30250 33224 30666 33280
rect 30189 33222 30666 33224
rect 31710 33222 33180 33282
rect 30189 33219 30255 33222
rect 25313 33146 25379 33149
rect 31710 33146 31770 33222
rect 33174 33220 33180 33222
rect 33244 33220 33250 33284
rect 33542 33220 33548 33284
rect 33612 33282 33618 33284
rect 34145 33282 34211 33285
rect 33612 33280 34211 33282
rect 33612 33224 34150 33280
rect 34206 33224 34211 33280
rect 33612 33222 34211 33224
rect 33612 33220 33618 33222
rect 34145 33219 34211 33222
rect 35709 33282 35775 33285
rect 37917 33282 37983 33285
rect 35709 33280 37983 33282
rect 35709 33224 35714 33280
rect 35770 33224 37922 33280
rect 37978 33224 37983 33280
rect 35709 33222 37983 33224
rect 35709 33219 35775 33222
rect 37917 33219 37983 33222
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 24764 33144 25379 33146
rect 24764 33088 25318 33144
rect 25374 33088 25379 33144
rect 24764 33086 25379 33088
rect 13261 33083 13327 33086
rect 13813 33083 13879 33086
rect 18229 33083 18295 33086
rect 11789 33010 11855 33013
rect 22050 33010 22110 33086
rect 24577 33083 24643 33086
rect 25313 33083 25379 33086
rect 25500 33086 31770 33146
rect 32673 33146 32739 33149
rect 32673 33144 34852 33146
rect 32673 33088 32678 33144
rect 32734 33088 34852 33144
rect 32673 33086 34852 33088
rect 11789 33008 22110 33010
rect 11789 32952 11794 33008
rect 11850 32952 22110 33008
rect 11789 32950 22110 32952
rect 22185 33010 22251 33013
rect 23473 33010 23539 33013
rect 22185 33008 23539 33010
rect 22185 32952 22190 33008
rect 22246 32952 23478 33008
rect 23534 32952 23539 33008
rect 22185 32950 23539 32952
rect 11789 32947 11855 32950
rect 22185 32947 22251 32950
rect 23473 32947 23539 32950
rect 25037 33010 25103 33013
rect 25262 33010 25268 33012
rect 25037 33008 25268 33010
rect 25037 32952 25042 33008
rect 25098 32952 25268 33008
rect 25037 32950 25268 32952
rect 25037 32947 25103 32950
rect 25262 32948 25268 32950
rect 25332 32948 25338 33012
rect 14825 32874 14891 32877
rect 15929 32874 15995 32877
rect 11654 32872 15995 32874
rect 11654 32816 14830 32872
rect 14886 32816 15934 32872
rect 15990 32816 15995 32872
rect 11654 32814 15995 32816
rect 4981 32811 5047 32814
rect 9765 32811 9831 32814
rect 10685 32811 10751 32814
rect 14825 32811 14891 32814
rect 15929 32811 15995 32814
rect 16573 32874 16639 32877
rect 24485 32874 24551 32877
rect 24945 32874 25011 32877
rect 16573 32872 25011 32874
rect 16573 32816 16578 32872
rect 16634 32816 24490 32872
rect 24546 32816 24950 32872
rect 25006 32816 25011 32872
rect 16573 32814 25011 32816
rect 16573 32811 16639 32814
rect 24485 32811 24551 32814
rect 24945 32811 25011 32814
rect 9029 32738 9095 32741
rect 9489 32738 9555 32741
rect 9029 32736 9555 32738
rect 9029 32680 9034 32736
rect 9090 32680 9494 32736
rect 9550 32680 9555 32736
rect 9029 32678 9555 32680
rect 9029 32675 9095 32678
rect 9489 32675 9555 32678
rect 10869 32738 10935 32741
rect 12893 32738 12959 32741
rect 10869 32736 12959 32738
rect 10869 32680 10874 32736
rect 10930 32680 12898 32736
rect 12954 32680 12959 32736
rect 10869 32678 12959 32680
rect 10869 32675 10935 32678
rect 12893 32675 12959 32678
rect 14089 32738 14155 32741
rect 16849 32738 16915 32741
rect 18413 32738 18479 32741
rect 14089 32736 18479 32738
rect 14089 32680 14094 32736
rect 14150 32680 16854 32736
rect 16910 32680 18418 32736
rect 18474 32680 18479 32736
rect 14089 32678 18479 32680
rect 14089 32675 14155 32678
rect 16849 32675 16915 32678
rect 18413 32675 18479 32678
rect 21909 32738 21975 32741
rect 22829 32738 22895 32741
rect 21909 32736 22895 32738
rect 21909 32680 21914 32736
rect 21970 32680 22834 32736
rect 22890 32680 22895 32736
rect 21909 32678 22895 32680
rect 21909 32675 21975 32678
rect 22829 32675 22895 32678
rect 24025 32738 24091 32741
rect 25500 32738 25560 33086
rect 32673 33083 32739 33086
rect 25681 33010 25747 33013
rect 28349 33010 28415 33013
rect 28625 33012 28691 33013
rect 28574 33010 28580 33012
rect 25681 33008 28415 33010
rect 25681 32952 25686 33008
rect 25742 32952 28354 33008
rect 28410 32952 28415 33008
rect 25681 32950 28415 32952
rect 28534 32950 28580 33010
rect 28644 33008 28691 33012
rect 28686 32952 28691 33008
rect 25681 32947 25747 32950
rect 28349 32947 28415 32950
rect 28574 32948 28580 32950
rect 28644 32948 28691 32952
rect 29126 32948 29132 33012
rect 29196 33010 29202 33012
rect 34605 33010 34671 33013
rect 29196 33008 34671 33010
rect 29196 32952 34610 33008
rect 34666 32952 34671 33008
rect 29196 32950 34671 32952
rect 34792 33010 34852 33086
rect 35709 33010 35775 33013
rect 37825 33010 37891 33013
rect 34792 33008 37891 33010
rect 34792 32952 35714 33008
rect 35770 32952 37830 33008
rect 37886 32952 37891 33008
rect 34792 32950 37891 32952
rect 29196 32948 29202 32950
rect 28625 32947 28691 32948
rect 34605 32947 34671 32950
rect 35709 32947 35775 32950
rect 37825 32947 37891 32950
rect 27889 32874 27955 32877
rect 34329 32874 34395 32877
rect 27889 32872 34395 32874
rect 27889 32816 27894 32872
rect 27950 32816 34334 32872
rect 34390 32816 34395 32872
rect 27889 32814 34395 32816
rect 27889 32811 27955 32814
rect 34329 32811 34395 32814
rect 34973 32874 35039 32877
rect 39200 32874 40000 32904
rect 34973 32872 40000 32874
rect 34973 32816 34978 32872
rect 35034 32816 40000 32872
rect 34973 32814 40000 32816
rect 34973 32811 35039 32814
rect 39200 32784 40000 32814
rect 24025 32736 25560 32738
rect 24025 32680 24030 32736
rect 24086 32680 25560 32736
rect 24025 32678 25560 32680
rect 24025 32675 24091 32678
rect 28022 32676 28028 32740
rect 28092 32738 28098 32740
rect 28809 32738 28875 32741
rect 28092 32736 28875 32738
rect 28092 32680 28814 32736
rect 28870 32680 28875 32736
rect 28092 32678 28875 32680
rect 28092 32676 28098 32678
rect 28809 32675 28875 32678
rect 29085 32738 29151 32741
rect 31201 32738 31267 32741
rect 29085 32736 31267 32738
rect 29085 32680 29090 32736
rect 29146 32680 31206 32736
rect 31262 32680 31267 32736
rect 29085 32678 31267 32680
rect 29085 32675 29151 32678
rect 31201 32675 31267 32678
rect 33317 32738 33383 32741
rect 36905 32738 36971 32741
rect 33317 32736 36971 32738
rect 33317 32680 33322 32736
rect 33378 32680 36910 32736
rect 36966 32680 36971 32736
rect 33317 32678 36971 32680
rect 33317 32675 33383 32678
rect 36905 32675 36971 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4521 32602 4587 32605
rect 6361 32602 6427 32605
rect 4521 32600 6427 32602
rect 4521 32544 4526 32600
rect 4582 32544 6366 32600
rect 6422 32544 6427 32600
rect 4521 32542 6427 32544
rect 4521 32539 4587 32542
rect 6361 32539 6427 32542
rect 6545 32602 6611 32605
rect 8937 32602 9003 32605
rect 12341 32604 12407 32605
rect 11278 32602 11284 32604
rect 6545 32600 11284 32602
rect 6545 32544 6550 32600
rect 6606 32544 8942 32600
rect 8998 32544 11284 32600
rect 6545 32542 11284 32544
rect 6545 32539 6611 32542
rect 8937 32539 9003 32542
rect 11278 32540 11284 32542
rect 11348 32540 11354 32604
rect 12341 32602 12388 32604
rect 12300 32600 12388 32602
rect 12452 32602 12458 32604
rect 12985 32602 13051 32605
rect 12452 32600 13051 32602
rect 12300 32544 12346 32600
rect 12452 32544 12990 32600
rect 13046 32544 13051 32600
rect 12300 32542 12388 32544
rect 12341 32540 12388 32542
rect 12452 32542 13051 32544
rect 12452 32540 12458 32542
rect 12341 32539 12407 32540
rect 12985 32539 13051 32542
rect 14365 32602 14431 32605
rect 14641 32602 14707 32605
rect 14365 32600 14707 32602
rect 14365 32544 14370 32600
rect 14426 32544 14646 32600
rect 14702 32544 14707 32600
rect 14365 32542 14707 32544
rect 14365 32539 14431 32542
rect 14641 32539 14707 32542
rect 15469 32602 15535 32605
rect 17861 32602 17927 32605
rect 18229 32602 18295 32605
rect 15469 32600 18295 32602
rect 15469 32544 15474 32600
rect 15530 32544 17866 32600
rect 17922 32544 18234 32600
rect 18290 32544 18295 32600
rect 15469 32542 18295 32544
rect 15469 32539 15535 32542
rect 17861 32539 17927 32542
rect 18229 32539 18295 32542
rect 21633 32602 21699 32605
rect 22921 32602 22987 32605
rect 21633 32600 22987 32602
rect 21633 32544 21638 32600
rect 21694 32544 22926 32600
rect 22982 32544 22987 32600
rect 21633 32542 22987 32544
rect 21633 32539 21699 32542
rect 22921 32539 22987 32542
rect 24577 32602 24643 32605
rect 27521 32602 27587 32605
rect 28390 32602 28396 32604
rect 24577 32600 28396 32602
rect 24577 32544 24582 32600
rect 24638 32544 27526 32600
rect 27582 32544 28396 32600
rect 24577 32542 28396 32544
rect 24577 32539 24643 32542
rect 27521 32539 27587 32542
rect 28390 32540 28396 32542
rect 28460 32540 28466 32604
rect 28533 32602 28599 32605
rect 35065 32602 35131 32605
rect 35801 32602 35867 32605
rect 38009 32602 38075 32605
rect 28533 32600 35867 32602
rect 28533 32544 28538 32600
rect 28594 32544 35070 32600
rect 35126 32544 35806 32600
rect 35862 32544 35867 32600
rect 28533 32542 35867 32544
rect 28533 32539 28599 32542
rect 35065 32539 35131 32542
rect 35801 32539 35867 32542
rect 35942 32600 38075 32602
rect 35942 32544 38014 32600
rect 38070 32544 38075 32600
rect 35942 32542 38075 32544
rect 8109 32466 8175 32469
rect 21633 32466 21699 32469
rect 8109 32464 21699 32466
rect 8109 32408 8114 32464
rect 8170 32408 21638 32464
rect 21694 32408 21699 32464
rect 8109 32406 21699 32408
rect 8109 32403 8175 32406
rect 21633 32403 21699 32406
rect 21817 32466 21883 32469
rect 22737 32466 22803 32469
rect 21817 32464 22803 32466
rect 21817 32408 21822 32464
rect 21878 32408 22742 32464
rect 22798 32408 22803 32464
rect 21817 32406 22803 32408
rect 21817 32403 21883 32406
rect 22737 32403 22803 32406
rect 23105 32466 23171 32469
rect 29085 32466 29151 32469
rect 23105 32464 29151 32466
rect 23105 32408 23110 32464
rect 23166 32408 29090 32464
rect 29146 32408 29151 32464
rect 23105 32406 29151 32408
rect 23105 32403 23171 32406
rect 29085 32403 29151 32406
rect 29729 32466 29795 32469
rect 30005 32466 30071 32469
rect 29729 32464 30071 32466
rect 29729 32408 29734 32464
rect 29790 32408 30010 32464
rect 30066 32408 30071 32464
rect 29729 32406 30071 32408
rect 29729 32403 29795 32406
rect 30005 32403 30071 32406
rect 30465 32466 30531 32469
rect 31886 32466 31892 32468
rect 30465 32464 31892 32466
rect 30465 32408 30470 32464
rect 30526 32408 31892 32464
rect 30465 32406 31892 32408
rect 30465 32403 30531 32406
rect 31886 32404 31892 32406
rect 31956 32466 31962 32468
rect 33869 32466 33935 32469
rect 35942 32466 36002 32542
rect 38009 32539 38075 32542
rect 31956 32464 33935 32466
rect 31956 32408 33874 32464
rect 33930 32408 33935 32464
rect 31956 32406 33935 32408
rect 31956 32404 31962 32406
rect 33869 32403 33935 32406
rect 34516 32406 36002 32466
rect 36077 32466 36143 32469
rect 36077 32464 36370 32466
rect 36077 32408 36082 32464
rect 36138 32408 36370 32464
rect 36077 32406 36370 32408
rect 4705 32330 4771 32333
rect 4838 32330 4844 32332
rect 4705 32328 4844 32330
rect 4705 32272 4710 32328
rect 4766 32272 4844 32328
rect 4705 32270 4844 32272
rect 4705 32267 4771 32270
rect 4838 32268 4844 32270
rect 4908 32268 4914 32332
rect 5809 32328 5875 32333
rect 5809 32272 5814 32328
rect 5870 32272 5875 32328
rect 5809 32267 5875 32272
rect 5993 32330 6059 32333
rect 9765 32330 9831 32333
rect 13353 32330 13419 32333
rect 13997 32330 14063 32333
rect 5993 32328 9690 32330
rect 5993 32272 5998 32328
rect 6054 32272 9690 32328
rect 5993 32270 9690 32272
rect 5993 32267 6059 32270
rect 5812 32194 5872 32267
rect 6269 32194 6335 32197
rect 5812 32192 6335 32194
rect 5812 32136 6274 32192
rect 6330 32136 6335 32192
rect 5812 32134 6335 32136
rect 6269 32131 6335 32134
rect 7833 32194 7899 32197
rect 9397 32194 9463 32197
rect 7833 32192 9463 32194
rect 7833 32136 7838 32192
rect 7894 32136 9402 32192
rect 9458 32136 9463 32192
rect 7833 32134 9463 32136
rect 9630 32194 9690 32270
rect 9765 32328 14063 32330
rect 9765 32272 9770 32328
rect 9826 32272 13358 32328
rect 13414 32272 14002 32328
rect 14058 32272 14063 32328
rect 9765 32270 14063 32272
rect 9765 32267 9831 32270
rect 13353 32267 13419 32270
rect 13997 32267 14063 32270
rect 14641 32330 14707 32333
rect 20345 32330 20411 32333
rect 21265 32330 21331 32333
rect 23381 32330 23447 32333
rect 14641 32328 21098 32330
rect 14641 32272 14646 32328
rect 14702 32272 20350 32328
rect 20406 32272 21098 32328
rect 14641 32270 21098 32272
rect 14641 32267 14707 32270
rect 20345 32267 20411 32270
rect 13486 32194 13492 32196
rect 9630 32134 13492 32194
rect 7833 32131 7899 32134
rect 9397 32131 9463 32134
rect 13486 32132 13492 32134
rect 13556 32132 13562 32196
rect 13670 32132 13676 32196
rect 13740 32194 13746 32196
rect 15377 32194 15443 32197
rect 18597 32194 18663 32197
rect 13740 32192 18663 32194
rect 13740 32136 15382 32192
rect 15438 32136 18602 32192
rect 18658 32136 18663 32192
rect 13740 32134 18663 32136
rect 13740 32132 13746 32134
rect 15377 32131 15443 32134
rect 18597 32131 18663 32134
rect 20662 32132 20668 32196
rect 20732 32194 20738 32196
rect 20805 32194 20871 32197
rect 20732 32192 20871 32194
rect 20732 32136 20810 32192
rect 20866 32136 20871 32192
rect 20732 32134 20871 32136
rect 21038 32194 21098 32270
rect 21265 32328 23447 32330
rect 21265 32272 21270 32328
rect 21326 32272 23386 32328
rect 23442 32272 23447 32328
rect 21265 32270 23447 32272
rect 21265 32267 21331 32270
rect 23381 32267 23447 32270
rect 23749 32330 23815 32333
rect 25313 32330 25379 32333
rect 28809 32330 28875 32333
rect 23749 32328 25379 32330
rect 23749 32272 23754 32328
rect 23810 32272 25318 32328
rect 25374 32272 25379 32328
rect 23749 32270 25379 32272
rect 23749 32267 23815 32270
rect 25313 32267 25379 32270
rect 26190 32328 28875 32330
rect 26190 32272 28814 32328
rect 28870 32272 28875 32328
rect 26190 32270 28875 32272
rect 22093 32194 22159 32197
rect 22737 32194 22803 32197
rect 25313 32194 25379 32197
rect 26190 32194 26250 32270
rect 28809 32267 28875 32270
rect 29085 32330 29151 32333
rect 32305 32330 32371 32333
rect 29085 32328 32371 32330
rect 29085 32272 29090 32328
rect 29146 32272 32310 32328
rect 32366 32272 32371 32328
rect 29085 32270 32371 32272
rect 29085 32267 29151 32270
rect 32305 32267 32371 32270
rect 32857 32330 32923 32333
rect 34516 32330 34576 32406
rect 36077 32403 36143 32406
rect 32857 32328 34576 32330
rect 32857 32272 32862 32328
rect 32918 32272 34576 32328
rect 32857 32270 34576 32272
rect 32857 32267 32923 32270
rect 34646 32268 34652 32332
rect 34716 32330 34722 32332
rect 34881 32330 34947 32333
rect 34716 32328 34947 32330
rect 34716 32272 34886 32328
rect 34942 32272 34947 32328
rect 34716 32270 34947 32272
rect 36310 32330 36370 32406
rect 36445 32330 36511 32333
rect 36310 32328 36511 32330
rect 36310 32272 36450 32328
rect 36506 32272 36511 32328
rect 36310 32270 36511 32272
rect 34716 32268 34722 32270
rect 34881 32267 34947 32270
rect 36445 32267 36511 32270
rect 21038 32192 22803 32194
rect 21038 32136 22098 32192
rect 22154 32136 22742 32192
rect 22798 32136 22803 32192
rect 21038 32134 22803 32136
rect 20732 32132 20738 32134
rect 20805 32131 20871 32134
rect 22093 32131 22159 32134
rect 22737 32131 22803 32134
rect 23982 32192 26250 32194
rect 23982 32136 25318 32192
rect 25374 32136 26250 32192
rect 23982 32134 26250 32136
rect 26325 32194 26391 32197
rect 29678 32194 29684 32196
rect 26325 32192 29684 32194
rect 26325 32136 26330 32192
rect 26386 32136 29684 32192
rect 26325 32134 29684 32136
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 10777 32058 10843 32061
rect 7974 32056 10843 32058
rect 7974 32000 10782 32056
rect 10838 32000 10843 32056
rect 7974 31998 10843 32000
rect 4429 31922 4495 31925
rect 7974 31922 8034 31998
rect 10777 31995 10843 31998
rect 11513 32058 11579 32061
rect 23982 32058 24042 32134
rect 25313 32131 25379 32134
rect 26325 32131 26391 32134
rect 29678 32132 29684 32134
rect 29748 32132 29754 32196
rect 30649 32194 30715 32197
rect 32581 32194 32647 32197
rect 30649 32192 32647 32194
rect 30649 32136 30654 32192
rect 30710 32136 32586 32192
rect 32642 32136 32647 32192
rect 30649 32134 32647 32136
rect 30649 32131 30715 32134
rect 32581 32131 32647 32134
rect 33358 32132 33364 32196
rect 33428 32194 33434 32196
rect 34697 32194 34763 32197
rect 33428 32192 34763 32194
rect 33428 32136 34702 32192
rect 34758 32136 34763 32192
rect 33428 32134 34763 32136
rect 33428 32132 33434 32134
rect 34697 32131 34763 32134
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 11513 32056 24042 32058
rect 11513 32000 11518 32056
rect 11574 32000 24042 32056
rect 11513 31998 24042 32000
rect 24117 32058 24183 32061
rect 24710 32058 24716 32060
rect 24117 32056 24716 32058
rect 24117 32000 24122 32056
rect 24178 32000 24716 32056
rect 24117 31998 24716 32000
rect 11513 31995 11579 31998
rect 24117 31995 24183 31998
rect 24710 31996 24716 31998
rect 24780 31996 24786 32060
rect 28206 31996 28212 32060
rect 28276 32058 28282 32060
rect 28625 32058 28691 32061
rect 28276 32056 28691 32058
rect 28276 32000 28630 32056
rect 28686 32000 28691 32056
rect 28276 31998 28691 32000
rect 28276 31996 28282 31998
rect 28625 31995 28691 31998
rect 29453 32060 29519 32061
rect 29453 32056 29500 32060
rect 29564 32058 29570 32060
rect 34513 32058 34579 32061
rect 29453 32000 29458 32056
rect 29453 31996 29500 32000
rect 29564 31998 29610 32058
rect 31710 32056 34579 32058
rect 31710 32000 34518 32056
rect 34574 32000 34579 32056
rect 31710 31998 34579 32000
rect 29564 31996 29570 31998
rect 29453 31995 29519 31996
rect 4429 31920 8034 31922
rect 4429 31864 4434 31920
rect 4490 31864 8034 31920
rect 4429 31862 8034 31864
rect 8201 31922 8267 31925
rect 10409 31922 10475 31925
rect 8201 31920 10475 31922
rect 8201 31864 8206 31920
rect 8262 31864 10414 31920
rect 10470 31864 10475 31920
rect 8201 31862 10475 31864
rect 4429 31859 4495 31862
rect 8201 31859 8267 31862
rect 10409 31859 10475 31862
rect 11605 31922 11671 31925
rect 13302 31922 13308 31924
rect 11605 31920 13308 31922
rect 11605 31864 11610 31920
rect 11666 31864 13308 31920
rect 11605 31862 13308 31864
rect 11605 31859 11671 31862
rect 13302 31860 13308 31862
rect 13372 31860 13378 31924
rect 16573 31922 16639 31925
rect 19333 31922 19399 31925
rect 16573 31920 19399 31922
rect 16573 31864 16578 31920
rect 16634 31864 19338 31920
rect 19394 31864 19399 31920
rect 16573 31862 19399 31864
rect 16573 31859 16639 31862
rect 19333 31859 19399 31862
rect 20805 31922 20871 31925
rect 21030 31922 21036 31924
rect 20805 31920 21036 31922
rect 20805 31864 20810 31920
rect 20866 31864 21036 31920
rect 20805 31862 21036 31864
rect 20805 31859 20871 31862
rect 21030 31860 21036 31862
rect 21100 31860 21106 31924
rect 21173 31922 21239 31925
rect 23289 31922 23355 31925
rect 21173 31920 23355 31922
rect 21173 31864 21178 31920
rect 21234 31864 23294 31920
rect 23350 31864 23355 31920
rect 21173 31862 23355 31864
rect 21173 31859 21239 31862
rect 23289 31859 23355 31862
rect 23974 31860 23980 31924
rect 24044 31922 24050 31924
rect 25405 31922 25471 31925
rect 24044 31920 25471 31922
rect 24044 31864 25410 31920
rect 25466 31864 25471 31920
rect 24044 31862 25471 31864
rect 24044 31860 24050 31862
rect 25405 31859 25471 31862
rect 28809 31922 28875 31925
rect 30465 31922 30531 31925
rect 28809 31920 30531 31922
rect 28809 31864 28814 31920
rect 28870 31864 30470 31920
rect 30526 31864 30531 31920
rect 28809 31862 30531 31864
rect 28809 31859 28875 31862
rect 30465 31859 30531 31862
rect 6085 31786 6151 31789
rect 6085 31784 6332 31786
rect 6085 31728 6090 31784
rect 6146 31728 6332 31784
rect 6085 31726 6332 31728
rect 6085 31723 6151 31726
rect 6272 31517 6332 31726
rect 8710 31726 15394 31786
rect 4889 31516 4955 31517
rect 4838 31514 4844 31516
rect 4798 31454 4844 31514
rect 4908 31512 4955 31516
rect 4950 31456 4955 31512
rect 4838 31452 4844 31454
rect 4908 31452 4955 31456
rect 4889 31451 4955 31452
rect 6269 31512 6335 31517
rect 6269 31456 6274 31512
rect 6330 31456 6335 31512
rect 6269 31451 6335 31456
rect 8385 31514 8451 31517
rect 8710 31514 8770 31726
rect 12566 31588 12572 31652
rect 12636 31650 12642 31652
rect 13169 31650 13235 31653
rect 12636 31648 13235 31650
rect 12636 31592 13174 31648
rect 13230 31592 13235 31648
rect 12636 31590 13235 31592
rect 12636 31588 12642 31590
rect 13169 31587 13235 31590
rect 13486 31588 13492 31652
rect 13556 31650 13562 31652
rect 14457 31650 14523 31653
rect 13556 31648 14523 31650
rect 13556 31592 14462 31648
rect 14518 31592 14523 31648
rect 13556 31590 14523 31592
rect 13556 31588 13562 31590
rect 14457 31587 14523 31590
rect 8385 31512 8770 31514
rect 8385 31456 8390 31512
rect 8446 31456 8770 31512
rect 8385 31454 8770 31456
rect 9397 31516 9463 31517
rect 9397 31512 9444 31516
rect 9508 31514 9514 31516
rect 10317 31514 10383 31517
rect 14917 31514 14983 31517
rect 9397 31456 9402 31512
rect 8385 31451 8451 31454
rect 9397 31452 9444 31456
rect 9508 31454 9554 31514
rect 10317 31512 14983 31514
rect 10317 31456 10322 31512
rect 10378 31456 14922 31512
rect 14978 31456 14983 31512
rect 10317 31454 14983 31456
rect 9508 31452 9514 31454
rect 9397 31451 9463 31452
rect 10317 31451 10383 31454
rect 14917 31451 14983 31454
rect 5625 31378 5691 31381
rect 9949 31378 10015 31381
rect 5625 31376 10015 31378
rect 5625 31320 5630 31376
rect 5686 31320 9954 31376
rect 10010 31320 10015 31376
rect 5625 31318 10015 31320
rect 5625 31315 5691 31318
rect 9949 31315 10015 31318
rect 11053 31378 11119 31381
rect 12198 31378 12204 31380
rect 11053 31376 12204 31378
rect 11053 31320 11058 31376
rect 11114 31320 12204 31376
rect 11053 31318 12204 31320
rect 11053 31315 11119 31318
rect 12198 31316 12204 31318
rect 12268 31378 12274 31380
rect 14089 31378 14155 31381
rect 12268 31376 14155 31378
rect 12268 31320 14094 31376
rect 14150 31320 14155 31376
rect 12268 31318 14155 31320
rect 12268 31316 12274 31318
rect 14089 31315 14155 31318
rect 5901 31242 5967 31245
rect 15193 31242 15259 31245
rect 5901 31240 15259 31242
rect 5901 31184 5906 31240
rect 5962 31184 15198 31240
rect 15254 31184 15259 31240
rect 5901 31182 15259 31184
rect 5901 31179 5967 31182
rect 15193 31179 15259 31182
rect 5257 31106 5323 31109
rect 15142 31106 15148 31108
rect 5257 31104 15148 31106
rect 5257 31048 5262 31104
rect 5318 31048 15148 31104
rect 5257 31046 15148 31048
rect 5257 31043 5323 31046
rect 15142 31044 15148 31046
rect 15212 31044 15218 31108
rect 15334 31106 15394 31726
rect 18270 31724 18276 31788
rect 18340 31786 18346 31788
rect 24945 31786 25011 31789
rect 25078 31786 25084 31788
rect 18340 31784 25084 31786
rect 18340 31728 24950 31784
rect 25006 31728 25084 31784
rect 18340 31726 25084 31728
rect 18340 31724 18346 31726
rect 24945 31723 25011 31726
rect 25078 31724 25084 31726
rect 25148 31724 25154 31788
rect 26550 31724 26556 31788
rect 26620 31786 26626 31788
rect 27889 31786 27955 31789
rect 26620 31784 27955 31786
rect 26620 31728 27894 31784
rect 27950 31728 27955 31784
rect 26620 31726 27955 31728
rect 26620 31724 26626 31726
rect 27889 31723 27955 31726
rect 28390 31724 28396 31788
rect 28460 31786 28466 31788
rect 28717 31786 28783 31789
rect 28460 31784 28783 31786
rect 28460 31728 28722 31784
rect 28778 31728 28783 31784
rect 28460 31726 28783 31728
rect 28460 31724 28466 31726
rect 28717 31723 28783 31726
rect 29310 31724 29316 31788
rect 29380 31786 29386 31788
rect 29729 31786 29795 31789
rect 29380 31784 29795 31786
rect 29380 31728 29734 31784
rect 29790 31728 29795 31784
rect 29380 31726 29795 31728
rect 29380 31724 29386 31726
rect 16297 31650 16363 31653
rect 18781 31650 18847 31653
rect 16297 31648 18847 31650
rect 16297 31592 16302 31648
rect 16358 31592 18786 31648
rect 18842 31592 18847 31648
rect 16297 31590 18847 31592
rect 16297 31587 16363 31590
rect 18781 31587 18847 31590
rect 20110 31588 20116 31652
rect 20180 31650 20186 31652
rect 20345 31650 20411 31653
rect 20180 31648 20411 31650
rect 20180 31592 20350 31648
rect 20406 31592 20411 31648
rect 20180 31590 20411 31592
rect 20180 31588 20186 31590
rect 20345 31587 20411 31590
rect 23657 31650 23723 31653
rect 27061 31650 27127 31653
rect 23657 31648 27127 31650
rect 23657 31592 23662 31648
rect 23718 31592 27066 31648
rect 27122 31592 27127 31648
rect 23657 31590 27127 31592
rect 23657 31587 23723 31590
rect 27061 31587 27127 31590
rect 27286 31588 27292 31652
rect 27356 31650 27362 31652
rect 29502 31650 29562 31726
rect 29729 31723 29795 31726
rect 27356 31590 29562 31650
rect 30925 31650 30991 31653
rect 31710 31650 31770 31998
rect 34513 31995 34579 31998
rect 35382 31996 35388 32060
rect 35452 32058 35458 32060
rect 36169 32058 36235 32061
rect 35452 32056 36235 32058
rect 35452 32000 36174 32056
rect 36230 32000 36235 32056
rect 35452 31998 36235 32000
rect 35452 31996 35458 31998
rect 36169 31995 36235 31998
rect 36721 32056 36787 32061
rect 36721 32000 36726 32056
rect 36782 32000 36787 32056
rect 36721 31995 36787 32000
rect 32581 31922 32647 31925
rect 33593 31922 33659 31925
rect 32581 31920 33659 31922
rect 32581 31864 32586 31920
rect 32642 31864 33598 31920
rect 33654 31864 33659 31920
rect 32581 31862 33659 31864
rect 32581 31859 32647 31862
rect 33593 31859 33659 31862
rect 35157 31922 35223 31925
rect 36445 31922 36511 31925
rect 35157 31920 36511 31922
rect 35157 31864 35162 31920
rect 35218 31864 36450 31920
rect 36506 31864 36511 31920
rect 35157 31862 36511 31864
rect 35157 31859 35223 31862
rect 36445 31859 36511 31862
rect 32029 31786 32095 31789
rect 33961 31786 34027 31789
rect 34513 31788 34579 31789
rect 34462 31786 34468 31788
rect 32029 31784 34027 31786
rect 32029 31728 32034 31784
rect 32090 31728 33966 31784
rect 34022 31728 34027 31784
rect 32029 31726 34027 31728
rect 34422 31726 34468 31786
rect 34532 31784 34579 31788
rect 34574 31728 34579 31784
rect 32029 31723 32095 31726
rect 33961 31723 34027 31726
rect 34462 31724 34468 31726
rect 34532 31724 34579 31728
rect 34513 31723 34579 31724
rect 34973 31786 35039 31789
rect 35433 31786 35499 31789
rect 36724 31786 36784 31995
rect 34973 31784 36784 31786
rect 34973 31728 34978 31784
rect 35034 31728 35438 31784
rect 35494 31728 36784 31784
rect 34973 31726 36784 31728
rect 34973 31723 35039 31726
rect 35433 31723 35499 31726
rect 30925 31648 31770 31650
rect 30925 31592 30930 31648
rect 30986 31592 31770 31648
rect 30925 31590 31770 31592
rect 32029 31650 32095 31653
rect 33542 31650 33548 31652
rect 32029 31648 33548 31650
rect 32029 31592 32034 31648
rect 32090 31592 33548 31648
rect 32029 31590 33548 31592
rect 27356 31588 27362 31590
rect 30925 31587 30991 31590
rect 32029 31587 32095 31590
rect 33542 31588 33548 31590
rect 33612 31588 33618 31652
rect 33869 31650 33935 31653
rect 34605 31650 34671 31653
rect 33869 31648 34671 31650
rect 33869 31592 33874 31648
rect 33930 31592 34610 31648
rect 34666 31592 34671 31648
rect 33869 31590 34671 31592
rect 33869 31587 33935 31590
rect 34605 31587 34671 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 17861 31514 17927 31517
rect 18873 31514 18939 31517
rect 17861 31512 18939 31514
rect 17861 31456 17866 31512
rect 17922 31456 18878 31512
rect 18934 31456 18939 31512
rect 17861 31454 18939 31456
rect 17861 31451 17927 31454
rect 18873 31451 18939 31454
rect 20478 31452 20484 31516
rect 20548 31514 20554 31516
rect 25589 31514 25655 31517
rect 20548 31512 25655 31514
rect 20548 31456 25594 31512
rect 25650 31456 25655 31512
rect 20548 31454 25655 31456
rect 20548 31452 20554 31454
rect 25589 31451 25655 31454
rect 26785 31514 26851 31517
rect 30649 31514 30715 31517
rect 26785 31512 30715 31514
rect 26785 31456 26790 31512
rect 26846 31456 30654 31512
rect 30710 31456 30715 31512
rect 26785 31454 30715 31456
rect 26785 31451 26851 31454
rect 30649 31451 30715 31454
rect 32121 31514 32187 31517
rect 39200 31514 40000 31544
rect 32121 31512 40000 31514
rect 32121 31456 32126 31512
rect 32182 31456 40000 31512
rect 32121 31454 40000 31456
rect 32121 31451 32187 31454
rect 39200 31424 40000 31454
rect 15653 31378 15719 31381
rect 24669 31378 24735 31381
rect 15653 31376 24735 31378
rect 15653 31320 15658 31376
rect 15714 31320 24674 31376
rect 24730 31320 24735 31376
rect 15653 31318 24735 31320
rect 15653 31315 15719 31318
rect 24669 31315 24735 31318
rect 25446 31316 25452 31380
rect 25516 31378 25522 31380
rect 28441 31378 28507 31381
rect 25516 31376 28507 31378
rect 25516 31320 28446 31376
rect 28502 31320 28507 31376
rect 25516 31318 28507 31320
rect 25516 31316 25522 31318
rect 28441 31315 28507 31318
rect 29729 31378 29795 31381
rect 30046 31378 30052 31380
rect 29729 31376 30052 31378
rect 29729 31320 29734 31376
rect 29790 31320 30052 31376
rect 29729 31318 30052 31320
rect 29729 31315 29795 31318
rect 30046 31316 30052 31318
rect 30116 31378 30122 31380
rect 34646 31378 34652 31380
rect 30116 31318 34652 31378
rect 30116 31316 30122 31318
rect 34646 31316 34652 31318
rect 34716 31316 34722 31380
rect 34789 31378 34855 31381
rect 35382 31378 35388 31380
rect 34789 31376 35388 31378
rect 34789 31320 34794 31376
rect 34850 31320 35388 31376
rect 34789 31318 35388 31320
rect 34789 31315 34855 31318
rect 35382 31316 35388 31318
rect 35452 31316 35458 31380
rect 16246 31180 16252 31244
rect 16316 31242 16322 31244
rect 25681 31242 25747 31245
rect 16316 31240 25747 31242
rect 16316 31184 25686 31240
rect 25742 31184 25747 31240
rect 16316 31182 25747 31184
rect 16316 31180 16322 31182
rect 25681 31179 25747 31182
rect 26141 31242 26207 31245
rect 26325 31242 26391 31245
rect 30465 31242 30531 31245
rect 26141 31240 26391 31242
rect 26141 31184 26146 31240
rect 26202 31184 26330 31240
rect 26386 31184 26391 31240
rect 26141 31182 26391 31184
rect 26141 31179 26207 31182
rect 26325 31179 26391 31182
rect 26926 31240 30531 31242
rect 26926 31184 30470 31240
rect 30526 31184 30531 31240
rect 26926 31182 30531 31184
rect 23749 31106 23815 31109
rect 15334 31104 23815 31106
rect 15334 31048 23754 31104
rect 23810 31048 23815 31104
rect 15334 31046 23815 31048
rect 23749 31043 23815 31046
rect 24117 31106 24183 31109
rect 26926 31106 26986 31182
rect 30465 31179 30531 31182
rect 31017 31242 31083 31245
rect 34462 31242 34468 31244
rect 31017 31240 34468 31242
rect 31017 31184 31022 31240
rect 31078 31184 34468 31240
rect 31017 31182 34468 31184
rect 31017 31179 31083 31182
rect 34462 31180 34468 31182
rect 34532 31180 34538 31244
rect 34973 31242 35039 31245
rect 34654 31240 35039 31242
rect 34654 31184 34978 31240
rect 35034 31184 35039 31240
rect 34654 31182 35039 31184
rect 24117 31104 26986 31106
rect 24117 31048 24122 31104
rect 24178 31048 26986 31104
rect 24117 31046 26986 31048
rect 27061 31106 27127 31109
rect 32029 31106 32095 31109
rect 27061 31104 32095 31106
rect 27061 31048 27066 31104
rect 27122 31048 32034 31104
rect 32090 31048 32095 31104
rect 27061 31046 32095 31048
rect 24117 31043 24183 31046
rect 27061 31043 27127 31046
rect 32029 31043 32095 31046
rect 32990 31044 32996 31108
rect 33060 31106 33066 31108
rect 33501 31106 33567 31109
rect 33060 31104 33567 31106
rect 33060 31048 33506 31104
rect 33562 31048 33567 31104
rect 33060 31046 33567 31048
rect 33060 31044 33066 31046
rect 33501 31043 33567 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 7097 30970 7163 30973
rect 9581 30970 9647 30973
rect 7097 30968 9647 30970
rect 7097 30912 7102 30968
rect 7158 30912 9586 30968
rect 9642 30912 9647 30968
rect 7097 30910 9647 30912
rect 7097 30907 7163 30910
rect 9581 30907 9647 30910
rect 10869 30970 10935 30973
rect 13445 30970 13511 30973
rect 10869 30968 13511 30970
rect 10869 30912 10874 30968
rect 10930 30912 13450 30968
rect 13506 30912 13511 30968
rect 10869 30910 13511 30912
rect 10869 30907 10935 30910
rect 13445 30907 13511 30910
rect 14549 30970 14615 30973
rect 16481 30970 16547 30973
rect 14549 30968 16547 30970
rect 14549 30912 14554 30968
rect 14610 30912 16486 30968
rect 16542 30912 16547 30968
rect 14549 30910 16547 30912
rect 14549 30907 14615 30910
rect 16481 30907 16547 30910
rect 16665 30970 16731 30973
rect 24761 30970 24827 30973
rect 16665 30968 24827 30970
rect 16665 30912 16670 30968
rect 16726 30912 24766 30968
rect 24822 30912 24827 30968
rect 16665 30910 24827 30912
rect 16665 30907 16731 30910
rect 24761 30907 24827 30910
rect 25221 30970 25287 30973
rect 27889 30970 27955 30973
rect 25221 30968 28320 30970
rect 25221 30912 25226 30968
rect 25282 30912 27894 30968
rect 27950 30912 28320 30968
rect 25221 30910 28320 30912
rect 25221 30907 25287 30910
rect 27889 30907 27955 30910
rect 8109 30834 8175 30837
rect 9489 30834 9555 30837
rect 8109 30832 9555 30834
rect 8109 30776 8114 30832
rect 8170 30776 9494 30832
rect 9550 30776 9555 30832
rect 8109 30774 9555 30776
rect 8109 30771 8175 30774
rect 9489 30771 9555 30774
rect 9765 30834 9831 30837
rect 12433 30834 12499 30837
rect 9765 30832 12499 30834
rect 9765 30776 9770 30832
rect 9826 30776 12438 30832
rect 12494 30776 12499 30832
rect 9765 30774 12499 30776
rect 9765 30771 9831 30774
rect 12433 30771 12499 30774
rect 13077 30834 13143 30837
rect 13353 30834 13419 30837
rect 13077 30832 13419 30834
rect 13077 30776 13082 30832
rect 13138 30776 13358 30832
rect 13414 30776 13419 30832
rect 13077 30774 13419 30776
rect 13077 30771 13143 30774
rect 13353 30771 13419 30774
rect 14733 30834 14799 30837
rect 27613 30834 27679 30837
rect 14733 30832 27679 30834
rect 14733 30776 14738 30832
rect 14794 30776 27618 30832
rect 27674 30776 27679 30832
rect 14733 30774 27679 30776
rect 28260 30834 28320 30910
rect 28390 30908 28396 30972
rect 28460 30970 28466 30972
rect 29545 30970 29611 30973
rect 34654 30970 34714 31182
rect 34973 31179 35039 31182
rect 35709 31244 35775 31245
rect 35709 31240 35756 31244
rect 35820 31242 35826 31244
rect 35709 31184 35714 31240
rect 35709 31180 35756 31184
rect 35820 31182 35866 31242
rect 35820 31180 35826 31182
rect 35709 31179 35775 31180
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 28460 30968 34714 30970
rect 28460 30912 29550 30968
rect 29606 30912 34714 30968
rect 28460 30910 34714 30912
rect 28460 30908 28466 30910
rect 29545 30907 29611 30910
rect 38285 30834 38351 30837
rect 28260 30832 38351 30834
rect 28260 30776 38290 30832
rect 38346 30776 38351 30832
rect 28260 30774 38351 30776
rect 14733 30771 14799 30774
rect 27613 30771 27679 30774
rect 38285 30771 38351 30774
rect 5349 30698 5415 30701
rect 9622 30698 9628 30700
rect 5349 30696 9628 30698
rect 5349 30640 5354 30696
rect 5410 30640 9628 30696
rect 5349 30638 9628 30640
rect 5349 30635 5415 30638
rect 9622 30636 9628 30638
rect 9692 30636 9698 30700
rect 11145 30698 11211 30701
rect 21541 30698 21607 30701
rect 11145 30696 21607 30698
rect 11145 30640 11150 30696
rect 11206 30640 21546 30696
rect 21602 30640 21607 30696
rect 11145 30638 21607 30640
rect 11145 30635 11211 30638
rect 21541 30635 21607 30638
rect 25681 30698 25747 30701
rect 30414 30698 30420 30700
rect 25681 30696 30420 30698
rect 25681 30640 25686 30696
rect 25742 30640 30420 30696
rect 25681 30638 30420 30640
rect 25681 30635 25747 30638
rect 30414 30636 30420 30638
rect 30484 30636 30490 30700
rect 30598 30636 30604 30700
rect 30668 30698 30674 30700
rect 35382 30698 35388 30700
rect 30668 30638 35388 30698
rect 30668 30636 30674 30638
rect 35382 30636 35388 30638
rect 35452 30636 35458 30700
rect 37038 30636 37044 30700
rect 37108 30698 37114 30700
rect 37181 30698 37247 30701
rect 37108 30696 37247 30698
rect 37108 30640 37186 30696
rect 37242 30640 37247 30696
rect 37108 30638 37247 30640
rect 37108 30636 37114 30638
rect 37181 30635 37247 30638
rect 5717 30562 5783 30565
rect 10869 30562 10935 30565
rect 13905 30562 13971 30565
rect 5717 30560 9690 30562
rect 5717 30504 5722 30560
rect 5778 30504 9690 30560
rect 5717 30502 9690 30504
rect 5717 30499 5783 30502
rect 7230 30364 7236 30428
rect 7300 30426 7306 30428
rect 8886 30426 8892 30428
rect 7300 30366 8892 30426
rect 7300 30364 7306 30366
rect 8886 30364 8892 30366
rect 8956 30364 8962 30428
rect 9630 30426 9690 30502
rect 10869 30560 13971 30562
rect 10869 30504 10874 30560
rect 10930 30504 13910 30560
rect 13966 30504 13971 30560
rect 10869 30502 13971 30504
rect 10869 30499 10935 30502
rect 13905 30499 13971 30502
rect 15326 30500 15332 30564
rect 15396 30562 15402 30564
rect 18965 30562 19031 30565
rect 15396 30560 19031 30562
rect 15396 30504 18970 30560
rect 19026 30504 19031 30560
rect 15396 30502 19031 30504
rect 15396 30500 15402 30502
rect 18965 30499 19031 30502
rect 23606 30500 23612 30564
rect 23676 30562 23682 30564
rect 28942 30562 28948 30564
rect 23676 30502 28948 30562
rect 23676 30500 23682 30502
rect 28942 30500 28948 30502
rect 29012 30500 29018 30564
rect 29361 30562 29427 30565
rect 31293 30562 31359 30565
rect 29361 30560 31359 30562
rect 29361 30504 29366 30560
rect 29422 30504 31298 30560
rect 31354 30504 31359 30560
rect 29361 30502 31359 30504
rect 29361 30499 29427 30502
rect 31293 30499 31359 30502
rect 33133 30562 33199 30565
rect 34646 30562 34652 30564
rect 33133 30560 34652 30562
rect 33133 30504 33138 30560
rect 33194 30504 34652 30560
rect 33133 30502 34652 30504
rect 33133 30499 33199 30502
rect 34646 30500 34652 30502
rect 34716 30562 34722 30564
rect 35801 30562 35867 30565
rect 34716 30560 35867 30562
rect 34716 30504 35806 30560
rect 35862 30504 35867 30560
rect 34716 30502 35867 30504
rect 34716 30500 34722 30502
rect 35801 30499 35867 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 18045 30426 18111 30429
rect 26049 30428 26115 30429
rect 25998 30426 26004 30428
rect 9630 30424 18111 30426
rect 9630 30368 18050 30424
rect 18106 30368 18111 30424
rect 9630 30366 18111 30368
rect 25958 30366 26004 30426
rect 26068 30424 26115 30428
rect 28073 30426 28139 30429
rect 26110 30368 26115 30424
rect 18045 30363 18111 30366
rect 25998 30364 26004 30366
rect 26068 30364 26115 30368
rect 26049 30363 26115 30364
rect 27294 30424 28139 30426
rect 27294 30368 28078 30424
rect 28134 30368 28139 30424
rect 27294 30366 28139 30368
rect 9673 30290 9739 30293
rect 11145 30290 11211 30293
rect 9673 30288 11211 30290
rect 9673 30232 9678 30288
rect 9734 30232 11150 30288
rect 11206 30232 11211 30288
rect 9673 30230 11211 30232
rect 9673 30227 9739 30230
rect 11145 30227 11211 30230
rect 11881 30290 11947 30293
rect 11881 30288 24410 30290
rect 11881 30232 11886 30288
rect 11942 30232 24410 30288
rect 11881 30230 24410 30232
rect 11881 30227 11947 30230
rect 7557 30154 7623 30157
rect 10961 30154 11027 30157
rect 7557 30152 11027 30154
rect 7557 30096 7562 30152
rect 7618 30096 10966 30152
rect 11022 30096 11027 30152
rect 7557 30094 11027 30096
rect 7557 30091 7623 30094
rect 10961 30091 11027 30094
rect 11513 30154 11579 30157
rect 12801 30154 12867 30157
rect 11513 30152 12867 30154
rect 11513 30096 11518 30152
rect 11574 30096 12806 30152
rect 12862 30096 12867 30152
rect 11513 30094 12867 30096
rect 11513 30091 11579 30094
rect 12801 30091 12867 30094
rect 18781 30154 18847 30157
rect 24209 30154 24275 30157
rect 18781 30152 24275 30154
rect 18781 30096 18786 30152
rect 18842 30096 24214 30152
rect 24270 30096 24275 30152
rect 18781 30094 24275 30096
rect 24350 30154 24410 30230
rect 24526 30228 24532 30292
rect 24596 30290 24602 30292
rect 27294 30290 27354 30366
rect 28073 30363 28139 30366
rect 28441 30426 28507 30429
rect 28993 30426 29059 30429
rect 30925 30426 30991 30429
rect 31845 30426 31911 30429
rect 28441 30424 29059 30426
rect 28441 30368 28446 30424
rect 28502 30368 28998 30424
rect 29054 30368 29059 30424
rect 28441 30366 29059 30368
rect 28441 30363 28507 30366
rect 28993 30363 29059 30366
rect 30284 30424 30991 30426
rect 30284 30368 30930 30424
rect 30986 30368 30991 30424
rect 30284 30366 30991 30368
rect 24596 30230 27354 30290
rect 27521 30290 27587 30293
rect 28574 30290 28580 30292
rect 27521 30288 28580 30290
rect 27521 30232 27526 30288
rect 27582 30232 28580 30288
rect 27521 30230 28580 30232
rect 24596 30228 24602 30230
rect 27521 30227 27587 30230
rect 28574 30228 28580 30230
rect 28644 30228 28650 30292
rect 25589 30156 25655 30157
rect 25446 30154 25452 30156
rect 24350 30094 25452 30154
rect 18781 30091 18847 30094
rect 24209 30091 24275 30094
rect 25446 30092 25452 30094
rect 25516 30092 25522 30156
rect 25589 30152 25636 30156
rect 25700 30154 25706 30156
rect 30284 30154 30344 30366
rect 30925 30363 30991 30366
rect 31710 30424 31911 30426
rect 31710 30368 31850 30424
rect 31906 30368 31911 30424
rect 31710 30366 31911 30368
rect 30741 30290 30807 30293
rect 31710 30290 31770 30366
rect 31845 30363 31911 30366
rect 32121 30426 32187 30429
rect 32121 30424 35266 30426
rect 32121 30368 32126 30424
rect 32182 30368 35266 30424
rect 32121 30366 35266 30368
rect 32121 30363 32187 30366
rect 30741 30288 31770 30290
rect 30741 30232 30746 30288
rect 30802 30232 31770 30288
rect 30741 30230 31770 30232
rect 31845 30290 31911 30293
rect 32949 30290 33015 30293
rect 31845 30288 33015 30290
rect 31845 30232 31850 30288
rect 31906 30232 32954 30288
rect 33010 30232 33015 30288
rect 31845 30230 33015 30232
rect 30741 30227 30807 30230
rect 31845 30227 31911 30230
rect 32949 30227 33015 30230
rect 33174 30228 33180 30292
rect 33244 30290 33250 30292
rect 33685 30290 33751 30293
rect 33244 30288 33751 30290
rect 33244 30232 33690 30288
rect 33746 30232 33751 30288
rect 33244 30230 33751 30232
rect 33244 30228 33250 30230
rect 33685 30227 33751 30230
rect 33910 30228 33916 30292
rect 33980 30290 33986 30292
rect 34605 30290 34671 30293
rect 33980 30288 34671 30290
rect 33980 30232 34610 30288
rect 34666 30232 34671 30288
rect 33980 30230 34671 30232
rect 35206 30290 35266 30366
rect 35382 30364 35388 30428
rect 35452 30426 35458 30428
rect 35934 30426 35940 30428
rect 35452 30366 35940 30426
rect 35452 30364 35458 30366
rect 35934 30364 35940 30366
rect 36004 30364 36010 30428
rect 38745 30426 38811 30429
rect 36126 30424 38811 30426
rect 36126 30368 38750 30424
rect 38806 30368 38811 30424
rect 36126 30366 38811 30368
rect 36126 30290 36186 30366
rect 38745 30363 38811 30366
rect 35206 30230 36186 30290
rect 33980 30228 33986 30230
rect 34605 30227 34671 30230
rect 33358 30154 33364 30156
rect 25589 30096 25594 30152
rect 25589 30092 25636 30096
rect 25700 30094 30344 30154
rect 30422 30094 33364 30154
rect 25700 30092 25706 30094
rect 25589 30091 25655 30092
rect 8753 30018 8819 30021
rect 16481 30018 16547 30021
rect 8753 30016 16547 30018
rect 8753 29960 8758 30016
rect 8814 29960 16486 30016
rect 16542 29960 16547 30016
rect 8753 29958 16547 29960
rect 8753 29955 8819 29958
rect 16481 29955 16547 29958
rect 26969 30018 27035 30021
rect 29545 30018 29611 30021
rect 30422 30018 30482 30094
rect 33358 30092 33364 30094
rect 33428 30092 33434 30156
rect 33542 30092 33548 30156
rect 33612 30154 33618 30156
rect 39200 30154 40000 30184
rect 33612 30094 40000 30154
rect 33612 30092 33618 30094
rect 39200 30064 40000 30094
rect 26969 30016 29611 30018
rect 26969 29960 26974 30016
rect 27030 29960 29550 30016
rect 29606 29960 29611 30016
rect 26969 29958 29611 29960
rect 26969 29955 27035 29958
rect 29545 29955 29611 29958
rect 29686 29958 30482 30018
rect 30649 30018 30715 30021
rect 31017 30018 31083 30021
rect 31150 30018 31156 30020
rect 30649 30016 31156 30018
rect 30649 29960 30654 30016
rect 30710 29960 31022 30016
rect 31078 29960 31156 30016
rect 30649 29958 31156 29960
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 7741 29882 7807 29885
rect 11329 29882 11395 29885
rect 7741 29880 11395 29882
rect 7741 29824 7746 29880
rect 7802 29824 11334 29880
rect 11390 29824 11395 29880
rect 7741 29822 11395 29824
rect 7741 29819 7807 29822
rect 11329 29819 11395 29822
rect 21633 29882 21699 29885
rect 27429 29882 27495 29885
rect 21633 29880 27495 29882
rect 21633 29824 21638 29880
rect 21694 29824 27434 29880
rect 27490 29824 27495 29880
rect 21633 29822 27495 29824
rect 21633 29819 21699 29822
rect 27429 29819 27495 29822
rect 29269 29882 29335 29885
rect 29686 29882 29746 29958
rect 30649 29955 30715 29958
rect 31017 29955 31083 29958
rect 31150 29956 31156 29958
rect 31220 29956 31226 30020
rect 33869 30018 33935 30021
rect 34697 30018 34763 30021
rect 32308 30016 34763 30018
rect 32308 29960 33874 30016
rect 33930 29960 34702 30016
rect 34758 29960 34763 30016
rect 32308 29958 34763 29960
rect 29269 29880 29746 29882
rect 29269 29824 29274 29880
rect 29330 29824 29746 29880
rect 29269 29822 29746 29824
rect 29913 29882 29979 29885
rect 32308 29882 32368 29958
rect 33869 29955 33935 29958
rect 34697 29955 34763 29958
rect 35433 30018 35499 30021
rect 36261 30018 36327 30021
rect 35433 30016 36327 30018
rect 35433 29960 35438 30016
rect 35494 29960 36266 30016
rect 36322 29960 36327 30016
rect 35433 29958 36327 29960
rect 35433 29955 35499 29958
rect 36261 29955 36327 29958
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 29913 29880 32368 29882
rect 29913 29824 29918 29880
rect 29974 29824 32368 29880
rect 29913 29822 32368 29824
rect 29269 29819 29335 29822
rect 29913 29819 29979 29822
rect 32438 29820 32444 29884
rect 32508 29882 32514 29884
rect 32581 29882 32647 29885
rect 32508 29880 34852 29882
rect 32508 29824 32586 29880
rect 32642 29824 34852 29880
rect 32508 29822 34852 29824
rect 32508 29820 32514 29822
rect 32581 29819 32647 29822
rect 7925 29746 7991 29749
rect 9029 29746 9095 29749
rect 7925 29744 9095 29746
rect 7925 29688 7930 29744
rect 7986 29688 9034 29744
rect 9090 29688 9095 29744
rect 7925 29686 9095 29688
rect 7925 29683 7991 29686
rect 9029 29683 9095 29686
rect 10041 29746 10107 29749
rect 12985 29746 13051 29749
rect 10041 29744 13051 29746
rect 10041 29688 10046 29744
rect 10102 29688 12990 29744
rect 13046 29688 13051 29744
rect 10041 29686 13051 29688
rect 10041 29683 10107 29686
rect 12985 29683 13051 29686
rect 15745 29746 15811 29749
rect 17125 29746 17191 29749
rect 15745 29744 17191 29746
rect 15745 29688 15750 29744
rect 15806 29688 17130 29744
rect 17186 29688 17191 29744
rect 15745 29686 17191 29688
rect 15745 29683 15811 29686
rect 17125 29683 17191 29686
rect 19006 29684 19012 29748
rect 19076 29746 19082 29748
rect 26918 29746 26924 29748
rect 19076 29686 26924 29746
rect 19076 29684 19082 29686
rect 26918 29684 26924 29686
rect 26988 29746 26994 29748
rect 27153 29746 27219 29749
rect 26988 29744 27219 29746
rect 26988 29688 27158 29744
rect 27214 29688 27219 29744
rect 26988 29686 27219 29688
rect 26988 29684 26994 29686
rect 27153 29683 27219 29686
rect 28942 29684 28948 29748
rect 29012 29746 29018 29748
rect 29729 29746 29795 29749
rect 29012 29744 29795 29746
rect 29012 29688 29734 29744
rect 29790 29688 29795 29744
rect 29012 29686 29795 29688
rect 29012 29684 29018 29686
rect 29729 29683 29795 29686
rect 30005 29746 30071 29749
rect 30741 29746 30807 29749
rect 30005 29744 30807 29746
rect 30005 29688 30010 29744
rect 30066 29688 30746 29744
rect 30802 29688 30807 29744
rect 30005 29686 30807 29688
rect 30005 29683 30071 29686
rect 30741 29683 30807 29686
rect 31937 29746 32003 29749
rect 34462 29746 34468 29748
rect 31937 29744 34468 29746
rect 31937 29688 31942 29744
rect 31998 29688 34468 29744
rect 31937 29686 34468 29688
rect 31937 29683 32003 29686
rect 34462 29684 34468 29686
rect 34532 29684 34538 29748
rect 34792 29746 34852 29822
rect 35525 29746 35591 29749
rect 37181 29746 37247 29749
rect 34792 29744 37247 29746
rect 34792 29688 35530 29744
rect 35586 29688 37186 29744
rect 37242 29688 37247 29744
rect 34792 29686 37247 29688
rect 35525 29683 35591 29686
rect 37181 29683 37247 29686
rect 6637 29610 6703 29613
rect 11513 29610 11579 29613
rect 11881 29610 11947 29613
rect 12433 29612 12499 29613
rect 6637 29608 11947 29610
rect 6637 29552 6642 29608
rect 6698 29552 11518 29608
rect 11574 29552 11886 29608
rect 11942 29552 11947 29608
rect 6637 29550 11947 29552
rect 6637 29547 6703 29550
rect 11513 29547 11579 29550
rect 11881 29547 11947 29550
rect 12382 29548 12388 29612
rect 12452 29610 12499 29612
rect 12452 29608 12544 29610
rect 12494 29552 12544 29608
rect 12452 29550 12544 29552
rect 12452 29548 12499 29550
rect 13302 29548 13308 29612
rect 13372 29610 13378 29612
rect 22134 29610 22140 29612
rect 13372 29550 22140 29610
rect 13372 29548 13378 29550
rect 22134 29548 22140 29550
rect 22204 29548 22210 29612
rect 22645 29610 22711 29613
rect 25037 29610 25103 29613
rect 36353 29610 36419 29613
rect 22645 29608 25103 29610
rect 22645 29552 22650 29608
rect 22706 29552 25042 29608
rect 25098 29552 25103 29608
rect 22645 29550 25103 29552
rect 12433 29547 12499 29548
rect 22645 29547 22711 29550
rect 25037 29547 25103 29550
rect 26926 29608 36419 29610
rect 26926 29552 36358 29608
rect 36414 29552 36419 29608
rect 26926 29550 36419 29552
rect 5533 29474 5599 29477
rect 8753 29474 8819 29477
rect 9397 29476 9463 29477
rect 9397 29474 9444 29476
rect 5533 29472 8819 29474
rect 5533 29416 5538 29472
rect 5594 29416 8758 29472
rect 8814 29416 8819 29472
rect 5533 29414 8819 29416
rect 9352 29472 9444 29474
rect 9352 29416 9402 29472
rect 9352 29414 9444 29416
rect 5533 29411 5599 29414
rect 8753 29411 8819 29414
rect 9397 29412 9444 29414
rect 9508 29412 9514 29476
rect 12750 29412 12756 29476
rect 12820 29474 12826 29476
rect 18045 29474 18111 29477
rect 26926 29474 26986 29550
rect 36353 29547 36419 29550
rect 12820 29472 18111 29474
rect 12820 29416 18050 29472
rect 18106 29416 18111 29472
rect 12820 29414 18111 29416
rect 12820 29412 12826 29414
rect 9397 29411 9463 29412
rect 18045 29411 18111 29414
rect 20072 29414 26986 29474
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 6913 29338 6979 29341
rect 8109 29338 8175 29341
rect 10317 29338 10383 29341
rect 6913 29336 10383 29338
rect 6913 29280 6918 29336
rect 6974 29280 8114 29336
rect 8170 29280 10322 29336
rect 10378 29280 10383 29336
rect 6913 29278 10383 29280
rect 6913 29275 6979 29278
rect 8109 29275 8175 29278
rect 10317 29275 10383 29278
rect 11094 29276 11100 29340
rect 11164 29338 11170 29340
rect 19374 29338 19380 29340
rect 11164 29278 19380 29338
rect 11164 29276 11170 29278
rect 19374 29276 19380 29278
rect 19444 29276 19450 29340
rect 6545 29202 6611 29205
rect 11697 29202 11763 29205
rect 17401 29202 17467 29205
rect 6545 29200 17467 29202
rect 6545 29144 6550 29200
rect 6606 29144 11702 29200
rect 11758 29144 17406 29200
rect 17462 29144 17467 29200
rect 6545 29142 17467 29144
rect 6545 29139 6611 29142
rect 11697 29139 11763 29142
rect 17401 29139 17467 29142
rect 17718 29140 17724 29204
rect 17788 29202 17794 29204
rect 20072 29202 20132 29414
rect 28758 29412 28764 29476
rect 28828 29474 28834 29476
rect 29729 29474 29795 29477
rect 30281 29474 30347 29477
rect 34053 29474 34119 29477
rect 28828 29472 30347 29474
rect 28828 29416 29734 29472
rect 29790 29416 30286 29472
rect 30342 29416 30347 29472
rect 28828 29414 30347 29416
rect 28828 29412 28834 29414
rect 29729 29411 29795 29414
rect 30281 29411 30347 29414
rect 31710 29472 34119 29474
rect 31710 29416 34058 29472
rect 34114 29416 34119 29472
rect 31710 29414 34119 29416
rect 24209 29338 24275 29341
rect 25037 29338 25103 29341
rect 24209 29336 25103 29338
rect 24209 29280 24214 29336
rect 24270 29280 25042 29336
rect 25098 29280 25103 29336
rect 24209 29278 25103 29280
rect 24209 29275 24275 29278
rect 25037 29275 25103 29278
rect 26601 29338 26667 29341
rect 27153 29338 27219 29341
rect 26601 29336 27219 29338
rect 26601 29280 26606 29336
rect 26662 29280 27158 29336
rect 27214 29280 27219 29336
rect 26601 29278 27219 29280
rect 26601 29275 26667 29278
rect 27153 29275 27219 29278
rect 28441 29338 28507 29341
rect 31710 29338 31770 29414
rect 34053 29411 34119 29414
rect 34278 29412 34284 29476
rect 34348 29474 34354 29476
rect 37089 29474 37155 29477
rect 34348 29472 37155 29474
rect 34348 29416 37094 29472
rect 37150 29416 37155 29472
rect 34348 29414 37155 29416
rect 34348 29412 34354 29414
rect 37089 29411 37155 29414
rect 33358 29338 33364 29340
rect 28441 29336 31770 29338
rect 28441 29280 28446 29336
rect 28502 29280 31770 29336
rect 28441 29278 31770 29280
rect 31848 29278 33364 29338
rect 28441 29275 28507 29278
rect 17788 29142 20132 29202
rect 22185 29202 22251 29205
rect 22737 29202 22803 29205
rect 26233 29202 26299 29205
rect 22185 29200 26299 29202
rect 22185 29144 22190 29200
rect 22246 29144 22742 29200
rect 22798 29144 26238 29200
rect 26294 29144 26299 29200
rect 22185 29142 26299 29144
rect 17788 29140 17794 29142
rect 22185 29139 22251 29142
rect 22737 29139 22803 29142
rect 26233 29139 26299 29142
rect 27153 29202 27219 29205
rect 29637 29202 29703 29205
rect 30557 29202 30623 29205
rect 27153 29200 30623 29202
rect 27153 29144 27158 29200
rect 27214 29144 29642 29200
rect 29698 29144 30562 29200
rect 30618 29144 30623 29200
rect 27153 29142 30623 29144
rect 27153 29139 27219 29142
rect 29637 29139 29703 29142
rect 30557 29139 30623 29142
rect 30833 29202 30899 29205
rect 31848 29202 31908 29278
rect 33358 29276 33364 29278
rect 33428 29276 33434 29340
rect 33501 29338 33567 29341
rect 36302 29338 36308 29340
rect 33501 29336 36308 29338
rect 33501 29280 33506 29336
rect 33562 29280 36308 29336
rect 33501 29278 36308 29280
rect 33501 29275 33567 29278
rect 36302 29276 36308 29278
rect 36372 29276 36378 29340
rect 32121 29204 32187 29205
rect 32070 29202 32076 29204
rect 30833 29200 31908 29202
rect 30833 29144 30838 29200
rect 30894 29144 31908 29200
rect 30833 29142 31908 29144
rect 32030 29142 32076 29202
rect 32140 29200 32187 29204
rect 32182 29144 32187 29200
rect 30833 29139 30899 29142
rect 32070 29140 32076 29142
rect 32140 29140 32187 29144
rect 32254 29140 32260 29204
rect 32324 29202 32330 29204
rect 33726 29202 33732 29204
rect 32324 29142 33732 29202
rect 32324 29140 32330 29142
rect 33726 29140 33732 29142
rect 33796 29202 33802 29204
rect 34237 29202 34303 29205
rect 33796 29200 34303 29202
rect 33796 29144 34242 29200
rect 34298 29144 34303 29200
rect 33796 29142 34303 29144
rect 33796 29140 33802 29142
rect 32121 29139 32187 29140
rect 34237 29139 34303 29142
rect 34462 29140 34468 29204
rect 34532 29202 34538 29204
rect 39481 29202 39547 29205
rect 34532 29200 39547 29202
rect 34532 29144 39486 29200
rect 39542 29144 39547 29200
rect 34532 29142 39547 29144
rect 34532 29140 34538 29142
rect 39481 29139 39547 29142
rect 9213 29066 9279 29069
rect 20069 29066 20135 29069
rect 9213 29064 20135 29066
rect 9213 29008 9218 29064
rect 9274 29008 20074 29064
rect 20130 29008 20135 29064
rect 9213 29006 20135 29008
rect 9213 29003 9279 29006
rect 20069 29003 20135 29006
rect 22369 29066 22435 29069
rect 22502 29066 22508 29068
rect 22369 29064 22508 29066
rect 22369 29008 22374 29064
rect 22430 29008 22508 29064
rect 22369 29006 22508 29008
rect 22369 29003 22435 29006
rect 22502 29004 22508 29006
rect 22572 29004 22578 29068
rect 24761 29066 24827 29069
rect 24894 29066 24900 29068
rect 24761 29064 24900 29066
rect 24761 29008 24766 29064
rect 24822 29008 24900 29064
rect 24761 29006 24900 29008
rect 24761 29003 24827 29006
rect 24894 29004 24900 29006
rect 24964 29004 24970 29068
rect 25037 29066 25103 29069
rect 25630 29066 25636 29068
rect 25037 29064 25636 29066
rect 25037 29008 25042 29064
rect 25098 29008 25636 29064
rect 25037 29006 25636 29008
rect 25037 29003 25103 29006
rect 25630 29004 25636 29006
rect 25700 29004 25706 29068
rect 26417 29066 26483 29069
rect 28165 29066 28231 29069
rect 26417 29064 28231 29066
rect 26417 29008 26422 29064
rect 26478 29008 28170 29064
rect 28226 29008 28231 29064
rect 26417 29006 28231 29008
rect 26417 29003 26483 29006
rect 28165 29003 28231 29006
rect 29310 29004 29316 29068
rect 29380 29066 29386 29068
rect 31477 29066 31543 29069
rect 29380 29064 31543 29066
rect 29380 29008 31482 29064
rect 31538 29008 31543 29064
rect 29380 29006 31543 29008
rect 29380 29004 29386 29006
rect 31477 29003 31543 29006
rect 33358 29004 33364 29068
rect 33428 29066 33434 29068
rect 33685 29066 33751 29069
rect 33428 29064 33751 29066
rect 33428 29008 33690 29064
rect 33746 29008 33751 29064
rect 33428 29006 33751 29008
rect 33428 29004 33434 29006
rect 33685 29003 33751 29006
rect 34654 29006 35450 29066
rect 6821 28930 6887 28933
rect 16113 28930 16179 28933
rect 6821 28928 16179 28930
rect 6821 28872 6826 28928
rect 6882 28872 16118 28928
rect 16174 28872 16179 28928
rect 6821 28870 16179 28872
rect 6821 28867 6887 28870
rect 16113 28867 16179 28870
rect 19190 28868 19196 28932
rect 19260 28930 19266 28932
rect 21357 28930 21423 28933
rect 19260 28928 21423 28930
rect 19260 28872 21362 28928
rect 21418 28872 21423 28928
rect 19260 28870 21423 28872
rect 19260 28868 19266 28870
rect 21357 28867 21423 28870
rect 23790 28868 23796 28932
rect 23860 28930 23866 28932
rect 28022 28930 28028 28932
rect 23860 28870 28028 28930
rect 23860 28868 23866 28870
rect 28022 28868 28028 28870
rect 28092 28868 28098 28932
rect 29177 28930 29243 28933
rect 30782 28930 30788 28932
rect 29177 28928 30788 28930
rect 29177 28872 29182 28928
rect 29238 28872 30788 28928
rect 29177 28870 30788 28872
rect 29177 28867 29243 28870
rect 30782 28868 30788 28870
rect 30852 28868 30858 28932
rect 30925 28930 30991 28933
rect 34654 28930 34714 29006
rect 30925 28928 34714 28930
rect 30925 28872 30930 28928
rect 30986 28872 34714 28928
rect 30925 28870 34714 28872
rect 35390 28930 35450 29006
rect 37825 28930 37891 28933
rect 35390 28928 37891 28930
rect 35390 28872 37830 28928
rect 37886 28872 37891 28928
rect 35390 28870 37891 28872
rect 30925 28867 30991 28870
rect 37825 28867 37891 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 10593 28794 10659 28797
rect 11421 28794 11487 28797
rect 10593 28792 11487 28794
rect 10593 28736 10598 28792
rect 10654 28736 11426 28792
rect 11482 28736 11487 28792
rect 10593 28734 11487 28736
rect 10593 28731 10659 28734
rect 11421 28731 11487 28734
rect 12065 28794 12131 28797
rect 13721 28794 13787 28797
rect 12065 28792 13787 28794
rect 12065 28736 12070 28792
rect 12126 28736 13726 28792
rect 13782 28736 13787 28792
rect 12065 28734 13787 28736
rect 12065 28731 12131 28734
rect 13721 28731 13787 28734
rect 14089 28794 14155 28797
rect 22093 28794 22159 28797
rect 27153 28794 27219 28797
rect 14089 28792 18522 28794
rect 14089 28736 14094 28792
rect 14150 28736 18522 28792
rect 14089 28734 18522 28736
rect 14089 28731 14155 28734
rect 6269 28658 6335 28661
rect 13537 28658 13603 28661
rect 6269 28656 13603 28658
rect 6269 28600 6274 28656
rect 6330 28600 13542 28656
rect 13598 28600 13603 28656
rect 6269 28598 13603 28600
rect 6269 28595 6335 28598
rect 13537 28595 13603 28598
rect 16573 28658 16639 28661
rect 18270 28658 18276 28660
rect 16573 28656 18276 28658
rect 16573 28600 16578 28656
rect 16634 28600 18276 28656
rect 16573 28598 18276 28600
rect 16573 28595 16639 28598
rect 18270 28596 18276 28598
rect 18340 28596 18346 28660
rect 18462 28658 18522 28734
rect 22093 28792 27219 28794
rect 22093 28736 22098 28792
rect 22154 28736 27158 28792
rect 27214 28736 27219 28792
rect 22093 28734 27219 28736
rect 22093 28731 22159 28734
rect 27153 28731 27219 28734
rect 30281 28794 30347 28797
rect 30598 28794 30604 28796
rect 30281 28792 30604 28794
rect 30281 28736 30286 28792
rect 30342 28736 30604 28792
rect 30281 28734 30604 28736
rect 30281 28731 30347 28734
rect 30598 28732 30604 28734
rect 30668 28732 30674 28796
rect 30782 28732 30788 28796
rect 30852 28794 30858 28796
rect 32489 28794 32555 28797
rect 30852 28792 32555 28794
rect 30852 28736 32494 28792
rect 32550 28736 32555 28792
rect 30852 28734 32555 28736
rect 30852 28732 30858 28734
rect 32489 28731 32555 28734
rect 33317 28794 33383 28797
rect 34789 28794 34855 28797
rect 39200 28794 40000 28824
rect 33317 28792 34855 28794
rect 33317 28736 33322 28792
rect 33378 28736 34794 28792
rect 34850 28736 34855 28792
rect 33317 28734 34855 28736
rect 33317 28731 33383 28734
rect 34789 28731 34855 28734
rect 35436 28734 40000 28794
rect 30649 28658 30715 28661
rect 18462 28656 30715 28658
rect 18462 28600 30654 28656
rect 30710 28600 30715 28656
rect 18462 28598 30715 28600
rect 30649 28595 30715 28598
rect 31518 28596 31524 28660
rect 31588 28658 31594 28660
rect 31588 28598 34024 28658
rect 31588 28596 31594 28598
rect 11053 28522 11119 28525
rect 16113 28522 16179 28525
rect 11053 28520 16179 28522
rect 11053 28464 11058 28520
rect 11114 28464 16118 28520
rect 16174 28464 16179 28520
rect 11053 28462 16179 28464
rect 11053 28459 11119 28462
rect 16113 28459 16179 28462
rect 18270 28460 18276 28524
rect 18340 28522 18346 28524
rect 23841 28522 23907 28525
rect 18340 28520 23907 28522
rect 18340 28464 23846 28520
rect 23902 28464 23907 28520
rect 18340 28462 23907 28464
rect 18340 28460 18346 28462
rect 23841 28459 23907 28462
rect 24485 28522 24551 28525
rect 26049 28522 26115 28525
rect 24485 28520 26115 28522
rect 24485 28464 24490 28520
rect 24546 28464 26054 28520
rect 26110 28464 26115 28520
rect 24485 28462 26115 28464
rect 24485 28459 24551 28462
rect 26049 28459 26115 28462
rect 26233 28522 26299 28525
rect 33964 28522 34024 28598
rect 34094 28596 34100 28660
rect 34164 28658 34170 28660
rect 34881 28658 34947 28661
rect 34164 28656 34947 28658
rect 34164 28600 34886 28656
rect 34942 28600 34947 28656
rect 34164 28598 34947 28600
rect 34164 28596 34170 28598
rect 34881 28595 34947 28598
rect 35436 28522 35496 28734
rect 39200 28704 40000 28734
rect 35709 28660 35775 28661
rect 35709 28658 35756 28660
rect 35664 28656 35756 28658
rect 35664 28600 35714 28656
rect 35664 28598 35756 28600
rect 35709 28596 35756 28598
rect 35820 28596 35826 28660
rect 35709 28595 35775 28596
rect 26233 28520 33610 28522
rect 26233 28464 26238 28520
rect 26294 28464 33610 28520
rect 26233 28462 33610 28464
rect 33964 28462 35496 28522
rect 26233 28459 26299 28462
rect 11237 28386 11303 28389
rect 18781 28386 18847 28389
rect 11237 28384 18847 28386
rect 11237 28328 11242 28384
rect 11298 28328 18786 28384
rect 18842 28328 18847 28384
rect 11237 28326 18847 28328
rect 11237 28323 11303 28326
rect 18781 28323 18847 28326
rect 23238 28324 23244 28388
rect 23308 28386 23314 28388
rect 26182 28386 26188 28388
rect 23308 28326 26188 28386
rect 23308 28324 23314 28326
rect 26182 28324 26188 28326
rect 26252 28386 26258 28388
rect 27797 28386 27863 28389
rect 26252 28384 27863 28386
rect 26252 28328 27802 28384
rect 27858 28328 27863 28384
rect 26252 28326 27863 28328
rect 33550 28386 33610 28462
rect 34605 28386 34671 28389
rect 33550 28384 34671 28386
rect 33550 28328 34610 28384
rect 34666 28328 34671 28384
rect 33550 28326 34671 28328
rect 26252 28324 26258 28326
rect 27797 28323 27863 28326
rect 34605 28323 34671 28326
rect 35750 28324 35756 28388
rect 35820 28386 35826 28388
rect 35985 28386 36051 28389
rect 35820 28384 36051 28386
rect 35820 28328 35990 28384
rect 36046 28328 36051 28384
rect 35820 28326 36051 28328
rect 35820 28324 35826 28326
rect 35985 28323 36051 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 13670 28188 13676 28252
rect 13740 28250 13746 28252
rect 16757 28250 16823 28253
rect 13740 28248 16823 28250
rect 13740 28192 16762 28248
rect 16818 28192 16823 28248
rect 13740 28190 16823 28192
rect 13740 28188 13746 28190
rect 16757 28187 16823 28190
rect 20713 28250 20779 28253
rect 23749 28250 23815 28253
rect 20713 28248 23815 28250
rect 20713 28192 20718 28248
rect 20774 28192 23754 28248
rect 23810 28192 23815 28248
rect 20713 28190 23815 28192
rect 20713 28187 20779 28190
rect 23749 28187 23815 28190
rect 23933 28250 23999 28253
rect 26550 28250 26556 28252
rect 23933 28248 26556 28250
rect 23933 28192 23938 28248
rect 23994 28192 26556 28248
rect 23933 28190 26556 28192
rect 23933 28187 23999 28190
rect 26550 28188 26556 28190
rect 26620 28188 26626 28252
rect 34421 28250 34487 28253
rect 28950 28248 34487 28250
rect 28950 28192 34426 28248
rect 34482 28192 34487 28248
rect 28950 28190 34487 28192
rect 20437 28114 20503 28117
rect 14782 28112 20503 28114
rect 14782 28056 20442 28112
rect 20498 28056 20503 28112
rect 14782 28054 20503 28056
rect 1761 27978 1827 27981
rect 14782 27978 14842 28054
rect 20437 28051 20503 28054
rect 21449 28114 21515 28117
rect 27470 28114 27476 28116
rect 21449 28112 27476 28114
rect 21449 28056 21454 28112
rect 21510 28056 27476 28112
rect 21449 28054 27476 28056
rect 21449 28051 21515 28054
rect 27470 28052 27476 28054
rect 27540 28052 27546 28116
rect 28206 28052 28212 28116
rect 28276 28114 28282 28116
rect 28950 28114 29010 28190
rect 34421 28187 34487 28190
rect 34789 28250 34855 28253
rect 35934 28250 35940 28252
rect 34789 28248 35940 28250
rect 34789 28192 34794 28248
rect 34850 28192 35940 28248
rect 34789 28190 35940 28192
rect 34789 28187 34855 28190
rect 35934 28188 35940 28190
rect 36004 28188 36010 28252
rect 31661 28116 31727 28117
rect 31661 28114 31708 28116
rect 28276 28054 29010 28114
rect 31616 28112 31708 28114
rect 31616 28056 31666 28112
rect 31616 28054 31708 28056
rect 28276 28052 28282 28054
rect 31661 28052 31708 28054
rect 31772 28052 31778 28116
rect 33041 28114 33107 28117
rect 37457 28114 37523 28117
rect 33041 28112 37523 28114
rect 33041 28056 33046 28112
rect 33102 28056 37462 28112
rect 37518 28056 37523 28112
rect 33041 28054 37523 28056
rect 31661 28051 31727 28052
rect 33041 28051 33107 28054
rect 37457 28051 37523 28054
rect 21633 27978 21699 27981
rect 24485 27978 24551 27981
rect 1761 27976 14842 27978
rect 1761 27920 1766 27976
rect 1822 27920 14842 27976
rect 1761 27918 14842 27920
rect 14966 27976 24551 27978
rect 14966 27920 21638 27976
rect 21694 27920 24490 27976
rect 24546 27920 24551 27976
rect 14966 27918 24551 27920
rect 1761 27915 1827 27918
rect 6729 27842 6795 27845
rect 14966 27842 15026 27918
rect 21633 27915 21699 27918
rect 24485 27915 24551 27918
rect 24710 27916 24716 27980
rect 24780 27978 24786 27980
rect 24780 27918 29194 27978
rect 24780 27916 24786 27918
rect 6729 27840 15026 27842
rect 6729 27784 6734 27840
rect 6790 27784 15026 27840
rect 6729 27782 15026 27784
rect 15101 27844 15167 27845
rect 19425 27844 19491 27845
rect 15101 27840 15148 27844
rect 15212 27842 15218 27844
rect 19374 27842 19380 27844
rect 15101 27784 15106 27840
rect 6729 27779 6795 27782
rect 15101 27780 15148 27784
rect 15212 27782 15258 27842
rect 19334 27782 19380 27842
rect 19444 27840 19491 27844
rect 24025 27842 24091 27845
rect 19486 27784 19491 27840
rect 15212 27780 15218 27782
rect 19374 27780 19380 27782
rect 19444 27780 19491 27784
rect 15101 27779 15167 27780
rect 19425 27779 19491 27780
rect 22050 27840 24091 27842
rect 22050 27784 24030 27840
rect 24086 27784 24091 27840
rect 22050 27782 24091 27784
rect 29134 27842 29194 27918
rect 29678 27916 29684 27980
rect 29748 27978 29754 27980
rect 30005 27978 30071 27981
rect 30373 27980 30439 27981
rect 30373 27978 30420 27980
rect 29748 27976 30071 27978
rect 29748 27920 30010 27976
rect 30066 27920 30071 27976
rect 29748 27918 30071 27920
rect 30328 27976 30420 27978
rect 30328 27920 30378 27976
rect 30328 27918 30420 27920
rect 29748 27916 29754 27918
rect 30005 27915 30071 27918
rect 30373 27916 30420 27918
rect 30484 27916 30490 27980
rect 30833 27978 30899 27981
rect 34421 27980 34487 27981
rect 30966 27978 30972 27980
rect 30833 27976 30972 27978
rect 30833 27920 30838 27976
rect 30894 27920 30972 27976
rect 30833 27918 30972 27920
rect 30373 27915 30439 27916
rect 30833 27915 30899 27918
rect 30966 27916 30972 27918
rect 31036 27916 31042 27980
rect 34421 27978 34468 27980
rect 34376 27976 34468 27978
rect 34376 27920 34426 27976
rect 34376 27918 34468 27920
rect 34421 27916 34468 27918
rect 34532 27916 34538 27980
rect 34421 27915 34487 27916
rect 31661 27842 31727 27845
rect 29134 27840 31727 27842
rect 29134 27784 31666 27840
rect 31722 27784 31727 27840
rect 29134 27782 31727 27784
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 7649 27706 7715 27709
rect 22050 27706 22110 27782
rect 24025 27779 24091 27782
rect 31661 27779 31727 27782
rect 33910 27780 33916 27844
rect 33980 27842 33986 27844
rect 34278 27842 34284 27844
rect 33980 27782 34284 27842
rect 33980 27780 33986 27782
rect 34278 27780 34284 27782
rect 34348 27842 34354 27844
rect 34421 27842 34487 27845
rect 34348 27840 34487 27842
rect 34348 27784 34426 27840
rect 34482 27784 34487 27840
rect 34348 27782 34487 27784
rect 34348 27780 34354 27782
rect 34421 27779 34487 27782
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 7649 27704 22110 27706
rect 7649 27648 7654 27704
rect 7710 27648 22110 27704
rect 7649 27646 22110 27648
rect 22645 27708 22711 27709
rect 22645 27704 22692 27708
rect 22756 27706 22762 27708
rect 22921 27706 22987 27709
rect 26325 27706 26391 27709
rect 22645 27648 22650 27704
rect 7649 27643 7715 27646
rect 22645 27644 22692 27648
rect 22756 27646 22802 27706
rect 22921 27704 26391 27706
rect 22921 27648 22926 27704
rect 22982 27648 26330 27704
rect 26386 27648 26391 27704
rect 22921 27646 26391 27648
rect 22756 27644 22762 27646
rect 22645 27643 22711 27644
rect 22921 27643 22987 27646
rect 26325 27643 26391 27646
rect 26509 27706 26575 27709
rect 34605 27706 34671 27709
rect 26509 27704 34671 27706
rect 26509 27648 26514 27704
rect 26570 27648 34610 27704
rect 34666 27648 34671 27704
rect 26509 27646 34671 27648
rect 26509 27643 26575 27646
rect 34605 27643 34671 27646
rect 8753 27570 8819 27573
rect 17861 27572 17927 27573
rect 26049 27572 26115 27573
rect 13670 27570 13676 27572
rect 8753 27568 13676 27570
rect 8753 27512 8758 27568
rect 8814 27512 13676 27568
rect 8753 27510 13676 27512
rect 8753 27507 8819 27510
rect 13670 27508 13676 27510
rect 13740 27508 13746 27572
rect 17861 27568 17908 27572
rect 17972 27570 17978 27572
rect 23422 27570 23428 27572
rect 17861 27512 17866 27568
rect 17861 27508 17908 27512
rect 17972 27510 18018 27570
rect 18094 27510 23428 27570
rect 17972 27508 17978 27510
rect 17861 27507 17927 27508
rect 8661 27434 8727 27437
rect 15745 27434 15811 27437
rect 8661 27432 15811 27434
rect 8661 27376 8666 27432
rect 8722 27376 15750 27432
rect 15806 27376 15811 27432
rect 8661 27374 15811 27376
rect 8661 27371 8727 27374
rect 15745 27371 15811 27374
rect 17677 27434 17743 27437
rect 18094 27434 18154 27510
rect 23422 27508 23428 27510
rect 23492 27508 23498 27572
rect 25998 27508 26004 27572
rect 26068 27570 26115 27572
rect 27061 27572 27127 27573
rect 27521 27572 27587 27573
rect 27061 27570 27108 27572
rect 26068 27568 26160 27570
rect 26110 27512 26160 27568
rect 26068 27510 26160 27512
rect 27016 27568 27108 27570
rect 27016 27512 27066 27568
rect 27016 27510 27108 27512
rect 26068 27508 26115 27510
rect 26049 27507 26115 27508
rect 27061 27508 27108 27510
rect 27172 27508 27178 27572
rect 27470 27570 27476 27572
rect 27430 27510 27476 27570
rect 27540 27568 27587 27572
rect 27582 27512 27587 27568
rect 27470 27508 27476 27510
rect 27540 27508 27587 27512
rect 27061 27507 27127 27508
rect 27521 27507 27587 27508
rect 29637 27570 29703 27573
rect 29913 27570 29979 27573
rect 29637 27568 29979 27570
rect 29637 27512 29642 27568
rect 29698 27512 29918 27568
rect 29974 27512 29979 27568
rect 29637 27510 29979 27512
rect 29637 27507 29703 27510
rect 29913 27507 29979 27510
rect 30373 27570 30439 27573
rect 31334 27570 31340 27572
rect 30373 27568 31340 27570
rect 30373 27512 30378 27568
rect 30434 27512 31340 27568
rect 30373 27510 31340 27512
rect 30373 27507 30439 27510
rect 31334 27508 31340 27510
rect 31404 27570 31410 27572
rect 31569 27570 31635 27573
rect 31404 27568 31635 27570
rect 31404 27512 31574 27568
rect 31630 27512 31635 27568
rect 31404 27510 31635 27512
rect 31404 27508 31410 27510
rect 31569 27507 31635 27510
rect 32213 27570 32279 27573
rect 34094 27570 34100 27572
rect 32213 27568 34100 27570
rect 32213 27512 32218 27568
rect 32274 27512 34100 27568
rect 32213 27510 34100 27512
rect 32213 27507 32279 27510
rect 34094 27508 34100 27510
rect 34164 27508 34170 27572
rect 34278 27508 34284 27572
rect 34348 27570 34354 27572
rect 34513 27570 34579 27573
rect 34348 27568 34579 27570
rect 34348 27512 34518 27568
rect 34574 27512 34579 27568
rect 34348 27510 34579 27512
rect 34348 27508 34354 27510
rect 34513 27507 34579 27510
rect 35157 27570 35223 27573
rect 35433 27570 35499 27573
rect 35157 27568 35499 27570
rect 35157 27512 35162 27568
rect 35218 27512 35438 27568
rect 35494 27512 35499 27568
rect 35157 27510 35499 27512
rect 35157 27507 35223 27510
rect 35433 27507 35499 27510
rect 31518 27434 31524 27436
rect 17677 27432 18154 27434
rect 17677 27376 17682 27432
rect 17738 27376 18154 27432
rect 17677 27374 18154 27376
rect 18278 27374 31524 27434
rect 17677 27371 17743 27374
rect 6361 27298 6427 27301
rect 15837 27298 15903 27301
rect 6361 27296 15903 27298
rect 6361 27240 6366 27296
rect 6422 27240 15842 27296
rect 15898 27240 15903 27296
rect 6361 27238 15903 27240
rect 6361 27235 6427 27238
rect 15837 27235 15903 27238
rect 17350 27236 17356 27300
rect 17420 27298 17426 27300
rect 18278 27298 18338 27374
rect 31518 27372 31524 27374
rect 31588 27372 31594 27436
rect 31661 27434 31727 27437
rect 39200 27434 40000 27464
rect 31661 27432 40000 27434
rect 31661 27376 31666 27432
rect 31722 27376 40000 27432
rect 31661 27374 40000 27376
rect 31661 27371 31727 27374
rect 39200 27344 40000 27374
rect 17420 27238 18338 27298
rect 17420 27236 17426 27238
rect 20294 27236 20300 27300
rect 20364 27298 20370 27300
rect 23105 27298 23171 27301
rect 23606 27298 23612 27300
rect 20364 27238 22708 27298
rect 20364 27236 20370 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 11053 27162 11119 27165
rect 18270 27162 18276 27164
rect 11053 27160 18276 27162
rect 11053 27104 11058 27160
rect 11114 27104 18276 27160
rect 11053 27102 18276 27104
rect 11053 27099 11119 27102
rect 18270 27100 18276 27102
rect 18340 27100 18346 27164
rect 22648 27162 22708 27238
rect 23105 27296 23612 27298
rect 23105 27240 23110 27296
rect 23166 27240 23612 27296
rect 23105 27238 23612 27240
rect 23105 27235 23171 27238
rect 23606 27236 23612 27238
rect 23676 27236 23682 27300
rect 23841 27298 23907 27301
rect 27153 27298 27219 27301
rect 23841 27296 27219 27298
rect 23841 27240 23846 27296
rect 23902 27240 27158 27296
rect 27214 27240 27219 27296
rect 23841 27238 27219 27240
rect 23841 27235 23907 27238
rect 27153 27235 27219 27238
rect 27797 27298 27863 27301
rect 32213 27298 32279 27301
rect 27797 27296 32279 27298
rect 27797 27240 27802 27296
rect 27858 27240 32218 27296
rect 32274 27240 32279 27296
rect 27797 27238 32279 27240
rect 27797 27235 27863 27238
rect 32213 27235 32279 27238
rect 32397 27298 32463 27301
rect 34881 27298 34947 27301
rect 32397 27296 34947 27298
rect 32397 27240 32402 27296
rect 32458 27240 34886 27296
rect 34942 27240 34947 27296
rect 32397 27238 34947 27240
rect 32397 27235 32463 27238
rect 34881 27235 34947 27238
rect 24526 27162 24532 27164
rect 22648 27102 24532 27162
rect 24526 27100 24532 27102
rect 24596 27100 24602 27164
rect 25814 27100 25820 27164
rect 25884 27162 25890 27164
rect 30097 27162 30163 27165
rect 33501 27162 33567 27165
rect 36169 27162 36235 27165
rect 36353 27164 36419 27165
rect 25884 27160 30163 27162
rect 25884 27104 30102 27160
rect 30158 27104 30163 27160
rect 25884 27102 30163 27104
rect 25884 27100 25890 27102
rect 30097 27099 30163 27102
rect 30422 27160 36235 27162
rect 30422 27104 33506 27160
rect 33562 27104 36174 27160
rect 36230 27104 36235 27160
rect 30422 27102 36235 27104
rect 9857 27026 9923 27029
rect 11973 27026 12039 27029
rect 13445 27028 13511 27029
rect 13445 27026 13492 27028
rect 9857 27024 12039 27026
rect 9857 26968 9862 27024
rect 9918 26968 11978 27024
rect 12034 26968 12039 27024
rect 9857 26966 12039 26968
rect 13400 27024 13492 27026
rect 13400 26968 13450 27024
rect 13400 26966 13492 26968
rect 9857 26963 9923 26966
rect 11973 26963 12039 26966
rect 13445 26964 13492 26966
rect 13556 26964 13562 27028
rect 14549 27026 14615 27029
rect 15285 27026 15351 27029
rect 17401 27026 17467 27029
rect 14549 27024 17467 27026
rect 14549 26968 14554 27024
rect 14610 26968 15290 27024
rect 15346 26968 17406 27024
rect 17462 26968 17467 27024
rect 14549 26966 17467 26968
rect 13445 26963 13511 26964
rect 14549 26963 14615 26966
rect 15285 26963 15351 26966
rect 17401 26963 17467 26966
rect 17953 27026 18019 27029
rect 28993 27026 29059 27029
rect 17953 27024 29059 27026
rect 17953 26968 17958 27024
rect 18014 26968 28998 27024
rect 29054 26968 29059 27024
rect 17953 26966 29059 26968
rect 17953 26963 18019 26966
rect 28993 26963 29059 26966
rect 29269 27026 29335 27029
rect 29494 27026 29500 27028
rect 29269 27024 29500 27026
rect 29269 26968 29274 27024
rect 29330 26968 29500 27024
rect 29269 26966 29500 26968
rect 29269 26963 29335 26966
rect 29494 26964 29500 26966
rect 29564 26964 29570 27028
rect 29637 27026 29703 27029
rect 30422 27026 30482 27102
rect 33501 27099 33567 27102
rect 36169 27099 36235 27102
rect 36302 27100 36308 27164
rect 36372 27162 36419 27164
rect 36372 27160 36464 27162
rect 36414 27104 36464 27160
rect 36372 27102 36464 27104
rect 36372 27100 36419 27102
rect 36353 27099 36419 27100
rect 29637 27024 30482 27026
rect 29637 26968 29642 27024
rect 29698 26968 30482 27024
rect 29637 26966 30482 26968
rect 30557 27026 30623 27029
rect 31150 27026 31156 27028
rect 30557 27024 31156 27026
rect 30557 26968 30562 27024
rect 30618 26968 31156 27024
rect 30557 26966 31156 26968
rect 29637 26963 29703 26966
rect 30557 26963 30623 26966
rect 31150 26964 31156 26966
rect 31220 26964 31226 27028
rect 31753 27026 31819 27029
rect 32990 27026 32996 27028
rect 31753 27024 32996 27026
rect 31753 26968 31758 27024
rect 31814 26968 32996 27024
rect 31753 26966 32996 26968
rect 31753 26963 31819 26966
rect 32990 26964 32996 26966
rect 33060 26964 33066 27028
rect 34646 26964 34652 27028
rect 34716 27026 34722 27028
rect 34973 27026 35039 27029
rect 36629 27026 36695 27029
rect 34716 27024 35039 27026
rect 34716 26968 34978 27024
rect 35034 26968 35039 27024
rect 34716 26966 35039 26968
rect 34716 26964 34722 26966
rect 34973 26963 35039 26966
rect 35758 27024 36695 27026
rect 35758 26968 36634 27024
rect 36690 26968 36695 27024
rect 35758 26966 36695 26968
rect 13261 26890 13327 26893
rect 20662 26890 20668 26892
rect 13261 26888 20668 26890
rect 13261 26832 13266 26888
rect 13322 26832 20668 26888
rect 13261 26830 20668 26832
rect 13261 26827 13327 26830
rect 20662 26828 20668 26830
rect 20732 26828 20738 26892
rect 22921 26890 22987 26893
rect 32070 26890 32076 26892
rect 22921 26888 32076 26890
rect 22921 26832 22926 26888
rect 22982 26832 32076 26888
rect 22921 26830 32076 26832
rect 22921 26827 22987 26830
rect 32070 26828 32076 26830
rect 32140 26828 32146 26892
rect 34976 26890 35036 26963
rect 35758 26893 35818 26966
rect 36629 26963 36695 26966
rect 35709 26890 35818 26893
rect 34976 26888 35818 26890
rect 34976 26832 35714 26888
rect 35770 26832 35818 26888
rect 34976 26830 35818 26832
rect 35709 26827 35775 26830
rect 4889 26754 4955 26757
rect 18045 26756 18111 26757
rect 15326 26754 15332 26756
rect 4889 26752 15332 26754
rect 4889 26696 4894 26752
rect 4950 26696 15332 26752
rect 4889 26694 15332 26696
rect 4889 26691 4955 26694
rect 15326 26692 15332 26694
rect 15396 26692 15402 26756
rect 18045 26754 18092 26756
rect 18000 26752 18092 26754
rect 18000 26696 18050 26752
rect 18000 26694 18092 26696
rect 18045 26692 18092 26694
rect 18156 26692 18162 26756
rect 18781 26754 18847 26757
rect 24577 26754 24643 26757
rect 25221 26756 25287 26757
rect 25221 26754 25268 26756
rect 18781 26752 24643 26754
rect 18781 26696 18786 26752
rect 18842 26696 24582 26752
rect 24638 26696 24643 26752
rect 18781 26694 24643 26696
rect 25176 26752 25268 26754
rect 25176 26696 25226 26752
rect 25176 26694 25268 26696
rect 18045 26691 18111 26692
rect 18781 26691 18847 26694
rect 24577 26691 24643 26694
rect 25221 26692 25268 26694
rect 25332 26692 25338 26756
rect 29545 26754 29611 26757
rect 33041 26756 33107 26757
rect 32990 26754 32996 26756
rect 29545 26752 32996 26754
rect 33060 26752 33107 26756
rect 29545 26696 29550 26752
rect 29606 26696 32996 26752
rect 33102 26696 33107 26752
rect 29545 26694 32996 26696
rect 25221 26691 25287 26692
rect 29545 26691 29611 26694
rect 32990 26692 32996 26694
rect 33060 26692 33107 26696
rect 33041 26691 33107 26692
rect 35341 26754 35407 26757
rect 35341 26752 35450 26754
rect 35341 26696 35346 26752
rect 35402 26696 35450 26752
rect 35341 26691 35450 26696
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 8150 26556 8156 26620
rect 8220 26618 8226 26620
rect 26366 26618 26372 26620
rect 8220 26558 26372 26618
rect 8220 26556 8226 26558
rect 26366 26556 26372 26558
rect 26436 26556 26442 26620
rect 27654 26556 27660 26620
rect 27724 26618 27730 26620
rect 32397 26618 32463 26621
rect 34646 26618 34652 26620
rect 27724 26558 31770 26618
rect 27724 26556 27730 26558
rect 6310 26420 6316 26484
rect 6380 26482 6386 26484
rect 20846 26482 20852 26484
rect 6380 26422 20852 26482
rect 6380 26420 6386 26422
rect 20846 26420 20852 26422
rect 20916 26420 20922 26484
rect 21030 26420 21036 26484
rect 21100 26482 21106 26484
rect 24853 26482 24919 26485
rect 21100 26480 24919 26482
rect 21100 26424 24858 26480
rect 24914 26424 24919 26480
rect 21100 26422 24919 26424
rect 21100 26420 21106 26422
rect 24853 26419 24919 26422
rect 25129 26482 25195 26485
rect 28901 26482 28967 26485
rect 25129 26480 28967 26482
rect 25129 26424 25134 26480
rect 25190 26424 28906 26480
rect 28962 26424 28967 26480
rect 25129 26422 28967 26424
rect 25129 26419 25195 26422
rect 28901 26419 28967 26422
rect 30230 26420 30236 26484
rect 30300 26482 30306 26484
rect 30925 26482 30991 26485
rect 30300 26480 30991 26482
rect 30300 26424 30930 26480
rect 30986 26424 30991 26480
rect 30300 26422 30991 26424
rect 31710 26482 31770 26558
rect 32397 26616 34652 26618
rect 32397 26560 32402 26616
rect 32458 26560 34652 26616
rect 32397 26558 34652 26560
rect 32397 26555 32463 26558
rect 34646 26556 34652 26558
rect 34716 26556 34722 26620
rect 34881 26482 34947 26485
rect 31710 26480 34947 26482
rect 31710 26424 34886 26480
rect 34942 26424 34947 26480
rect 31710 26422 34947 26424
rect 30300 26420 30306 26422
rect 30925 26419 30991 26422
rect 34881 26419 34947 26422
rect 35157 26482 35223 26485
rect 35390 26482 35450 26691
rect 35157 26480 35450 26482
rect 35157 26424 35162 26480
rect 35218 26424 35450 26480
rect 35157 26422 35450 26424
rect 35157 26419 35223 26422
rect 16430 26284 16436 26348
rect 16500 26346 16506 26348
rect 17953 26346 18019 26349
rect 16500 26344 18019 26346
rect 16500 26288 17958 26344
rect 18014 26288 18019 26344
rect 16500 26286 18019 26288
rect 16500 26284 16506 26286
rect 17953 26283 18019 26286
rect 18597 26346 18663 26349
rect 20529 26346 20595 26349
rect 23289 26346 23355 26349
rect 18597 26344 20132 26346
rect 18597 26288 18602 26344
rect 18658 26288 20132 26344
rect 18597 26286 20132 26288
rect 18597 26283 18663 26286
rect 4981 26210 5047 26213
rect 18597 26210 18663 26213
rect 19006 26210 19012 26212
rect 4981 26208 17970 26210
rect 4981 26152 4986 26208
rect 5042 26152 17970 26208
rect 4981 26150 17970 26152
rect 4981 26147 5047 26150
rect 5441 26074 5507 26077
rect 13302 26074 13308 26076
rect 5441 26072 13308 26074
rect 5441 26016 5446 26072
rect 5502 26016 13308 26072
rect 5441 26014 13308 26016
rect 5441 26011 5507 26014
rect 13302 26012 13308 26014
rect 13372 26012 13378 26076
rect 17910 26074 17970 26150
rect 18597 26208 19012 26210
rect 18597 26152 18602 26208
rect 18658 26152 19012 26208
rect 18597 26150 19012 26152
rect 18597 26147 18663 26150
rect 19006 26148 19012 26150
rect 19076 26148 19082 26212
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 19057 26074 19123 26077
rect 17910 26072 19123 26074
rect 17910 26016 19062 26072
rect 19118 26016 19123 26072
rect 17910 26014 19123 26016
rect 20072 26074 20132 26286
rect 20529 26344 23355 26346
rect 20529 26288 20534 26344
rect 20590 26288 23294 26344
rect 23350 26288 23355 26344
rect 20529 26286 23355 26288
rect 20529 26283 20595 26286
rect 23289 26283 23355 26286
rect 23841 26346 23907 26349
rect 24158 26346 24164 26348
rect 23841 26344 24164 26346
rect 23841 26288 23846 26344
rect 23902 26288 24164 26344
rect 23841 26286 24164 26288
rect 23841 26283 23907 26286
rect 24158 26284 24164 26286
rect 24228 26284 24234 26348
rect 26141 26346 26207 26349
rect 29126 26346 29132 26348
rect 26141 26344 29132 26346
rect 26141 26288 26146 26344
rect 26202 26288 29132 26344
rect 26141 26286 29132 26288
rect 26141 26283 26207 26286
rect 29126 26284 29132 26286
rect 29196 26284 29202 26348
rect 29545 26346 29611 26349
rect 30281 26346 30347 26349
rect 29545 26344 30347 26346
rect 29545 26288 29550 26344
rect 29606 26288 30286 26344
rect 30342 26288 30347 26344
rect 29545 26286 30347 26288
rect 29545 26283 29611 26286
rect 30281 26283 30347 26286
rect 30598 26284 30604 26348
rect 30668 26346 30674 26348
rect 30925 26346 30991 26349
rect 30668 26344 30991 26346
rect 30668 26288 30930 26344
rect 30986 26288 30991 26344
rect 30668 26286 30991 26288
rect 30668 26284 30674 26286
rect 30925 26283 30991 26286
rect 31845 26348 31911 26349
rect 31845 26344 31892 26348
rect 31956 26346 31962 26348
rect 31845 26288 31850 26344
rect 31845 26284 31892 26288
rect 31956 26286 32002 26346
rect 31956 26284 31962 26286
rect 31845 26283 31911 26284
rect 20529 26212 20595 26213
rect 20478 26148 20484 26212
rect 20548 26210 20595 26212
rect 22461 26210 22527 26213
rect 24209 26210 24275 26213
rect 26785 26210 26851 26213
rect 20548 26208 20640 26210
rect 20590 26152 20640 26208
rect 20548 26150 20640 26152
rect 22461 26208 26851 26210
rect 22461 26152 22466 26208
rect 22522 26152 24214 26208
rect 24270 26152 26790 26208
rect 26846 26152 26851 26208
rect 22461 26150 26851 26152
rect 20548 26148 20595 26150
rect 20529 26147 20595 26148
rect 22461 26147 22527 26150
rect 24209 26147 24275 26150
rect 26785 26147 26851 26150
rect 27705 26210 27771 26213
rect 28758 26210 28764 26212
rect 27705 26208 28764 26210
rect 27705 26152 27710 26208
rect 27766 26152 28764 26208
rect 27705 26150 28764 26152
rect 27705 26147 27771 26150
rect 28758 26148 28764 26150
rect 28828 26148 28834 26212
rect 28993 26210 29059 26213
rect 32949 26210 33015 26213
rect 28993 26208 33015 26210
rect 28993 26152 28998 26208
rect 29054 26152 32954 26208
rect 33010 26152 33015 26208
rect 28993 26150 33015 26152
rect 28993 26147 29059 26150
rect 32949 26147 33015 26150
rect 20478 26074 20484 26076
rect 20072 26014 20484 26074
rect 19057 26011 19123 26014
rect 20478 26012 20484 26014
rect 20548 26012 20554 26076
rect 20989 26074 21055 26077
rect 30097 26074 30163 26077
rect 33225 26074 33291 26077
rect 20989 26072 29010 26074
rect 20989 26016 20994 26072
rect 21050 26016 29010 26072
rect 20989 26014 29010 26016
rect 20989 26011 21055 26014
rect 15142 25876 15148 25940
rect 15212 25938 15218 25940
rect 25589 25938 25655 25941
rect 26509 25938 26575 25941
rect 28809 25938 28875 25941
rect 15212 25878 24778 25938
rect 15212 25876 15218 25878
rect 12985 25802 13051 25805
rect 19425 25802 19491 25805
rect 12985 25800 19491 25802
rect 12985 25744 12990 25800
rect 13046 25744 19430 25800
rect 19486 25744 19491 25800
rect 12985 25742 19491 25744
rect 12985 25739 13051 25742
rect 19425 25739 19491 25742
rect 20161 25802 20227 25805
rect 24301 25802 24367 25805
rect 20161 25800 24367 25802
rect 20161 25744 20166 25800
rect 20222 25744 24306 25800
rect 24362 25744 24367 25800
rect 20161 25742 24367 25744
rect 24718 25802 24778 25878
rect 25589 25936 28875 25938
rect 25589 25880 25594 25936
rect 25650 25880 26514 25936
rect 26570 25880 28814 25936
rect 28870 25880 28875 25936
rect 25589 25878 28875 25880
rect 28950 25938 29010 26014
rect 30097 26072 33291 26074
rect 30097 26016 30102 26072
rect 30158 26016 33230 26072
rect 33286 26016 33291 26072
rect 30097 26014 33291 26016
rect 30097 26011 30163 26014
rect 33225 26011 33291 26014
rect 34278 26012 34284 26076
rect 34348 26074 34354 26076
rect 37365 26074 37431 26077
rect 34348 26072 37431 26074
rect 34348 26016 37370 26072
rect 37426 26016 37431 26072
rect 34348 26014 37431 26016
rect 34348 26012 34354 26014
rect 37365 26011 37431 26014
rect 38469 26074 38535 26077
rect 39200 26074 40000 26104
rect 38469 26072 40000 26074
rect 38469 26016 38474 26072
rect 38530 26016 40000 26072
rect 38469 26014 40000 26016
rect 38469 26011 38535 26014
rect 39200 25984 40000 26014
rect 30557 25938 30623 25941
rect 28950 25936 30623 25938
rect 28950 25880 30562 25936
rect 30618 25880 30623 25936
rect 28950 25878 30623 25880
rect 25589 25875 25655 25878
rect 26509 25875 26575 25878
rect 28809 25875 28875 25878
rect 30557 25875 30623 25878
rect 31201 25938 31267 25941
rect 31518 25938 31524 25940
rect 31201 25936 31524 25938
rect 31201 25880 31206 25936
rect 31262 25880 31524 25936
rect 31201 25878 31524 25880
rect 31201 25875 31267 25878
rect 31518 25876 31524 25878
rect 31588 25938 31594 25940
rect 34513 25938 34579 25941
rect 31588 25936 34579 25938
rect 31588 25880 34518 25936
rect 34574 25880 34579 25936
rect 31588 25878 34579 25880
rect 31588 25876 31594 25878
rect 34513 25875 34579 25878
rect 25957 25804 26023 25805
rect 25957 25802 26004 25804
rect 24718 25800 26004 25802
rect 24718 25744 25962 25800
rect 24718 25742 26004 25744
rect 20161 25739 20227 25742
rect 24301 25739 24367 25742
rect 25957 25740 26004 25742
rect 26068 25740 26074 25804
rect 26550 25740 26556 25804
rect 26620 25802 26626 25804
rect 29637 25802 29703 25805
rect 26620 25800 29703 25802
rect 26620 25744 29642 25800
rect 29698 25744 29703 25800
rect 26620 25742 29703 25744
rect 26620 25740 26626 25742
rect 25957 25739 26023 25740
rect 29637 25739 29703 25742
rect 30281 25802 30347 25805
rect 36077 25802 36143 25805
rect 30281 25800 36143 25802
rect 30281 25744 30286 25800
rect 30342 25744 36082 25800
rect 36138 25744 36143 25800
rect 30281 25742 36143 25744
rect 30281 25739 30347 25742
rect 36077 25739 36143 25742
rect 18413 25666 18479 25669
rect 23933 25666 23999 25669
rect 18413 25664 23999 25666
rect 18413 25608 18418 25664
rect 18474 25608 23938 25664
rect 23994 25608 23999 25664
rect 18413 25606 23999 25608
rect 18413 25603 18479 25606
rect 23933 25603 23999 25606
rect 24945 25666 25011 25669
rect 25957 25666 26023 25669
rect 24945 25664 26023 25666
rect 24945 25608 24950 25664
rect 25006 25608 25962 25664
rect 26018 25608 26023 25664
rect 24945 25606 26023 25608
rect 24945 25603 25011 25606
rect 25957 25603 26023 25606
rect 28533 25666 28599 25669
rect 28717 25666 28783 25669
rect 30189 25666 30255 25669
rect 28533 25664 30255 25666
rect 28533 25608 28538 25664
rect 28594 25608 28722 25664
rect 28778 25608 30194 25664
rect 30250 25608 30255 25664
rect 28533 25606 30255 25608
rect 28533 25603 28599 25606
rect 28717 25603 28783 25606
rect 30189 25603 30255 25606
rect 30925 25666 30991 25669
rect 31109 25666 31175 25669
rect 30925 25664 31175 25666
rect 30925 25608 30930 25664
rect 30986 25608 31114 25664
rect 31170 25608 31175 25664
rect 30925 25606 31175 25608
rect 30925 25603 30991 25606
rect 31109 25603 31175 25606
rect 31385 25666 31451 25669
rect 33777 25666 33843 25669
rect 31385 25664 33843 25666
rect 31385 25608 31390 25664
rect 31446 25608 33782 25664
rect 33838 25608 33843 25664
rect 31385 25606 33843 25608
rect 31385 25603 31451 25606
rect 33777 25603 33843 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 6126 25468 6132 25532
rect 6196 25530 6202 25532
rect 20621 25530 20687 25533
rect 6196 25528 20687 25530
rect 6196 25472 20626 25528
rect 20682 25472 20687 25528
rect 6196 25470 20687 25472
rect 6196 25468 6202 25470
rect 20621 25467 20687 25470
rect 22645 25530 22711 25533
rect 28206 25530 28212 25532
rect 22645 25528 28212 25530
rect 22645 25472 22650 25528
rect 22706 25472 28212 25528
rect 22645 25470 28212 25472
rect 22645 25467 22711 25470
rect 28206 25468 28212 25470
rect 28276 25468 28282 25532
rect 28349 25530 28415 25533
rect 28901 25530 28967 25533
rect 28349 25528 28967 25530
rect 28349 25472 28354 25528
rect 28410 25472 28906 25528
rect 28962 25472 28967 25528
rect 28349 25470 28967 25472
rect 28349 25467 28415 25470
rect 28901 25467 28967 25470
rect 29729 25530 29795 25533
rect 29862 25530 29868 25532
rect 29729 25528 29868 25530
rect 29729 25472 29734 25528
rect 29790 25472 29868 25528
rect 29729 25470 29868 25472
rect 29729 25467 29795 25470
rect 29862 25468 29868 25470
rect 29932 25468 29938 25532
rect 30005 25530 30071 25533
rect 31937 25530 32003 25533
rect 30005 25528 32003 25530
rect 30005 25472 30010 25528
rect 30066 25472 31942 25528
rect 31998 25472 32003 25528
rect 30005 25470 32003 25472
rect 30005 25467 30071 25470
rect 31937 25467 32003 25470
rect 4797 25394 4863 25397
rect 19425 25394 19491 25397
rect 20294 25394 20300 25396
rect 4797 25392 20300 25394
rect 4797 25336 4802 25392
rect 4858 25336 19430 25392
rect 19486 25336 20300 25392
rect 4797 25334 20300 25336
rect 4797 25331 4863 25334
rect 19425 25331 19491 25334
rect 20294 25332 20300 25334
rect 20364 25332 20370 25396
rect 20478 25332 20484 25396
rect 20548 25394 20554 25396
rect 26550 25394 26556 25396
rect 20548 25334 26556 25394
rect 20548 25332 20554 25334
rect 26550 25332 26556 25334
rect 26620 25332 26626 25396
rect 27521 25394 27587 25397
rect 33174 25394 33180 25396
rect 27521 25392 33180 25394
rect 27521 25336 27526 25392
rect 27582 25336 33180 25392
rect 27521 25334 33180 25336
rect 27521 25331 27587 25334
rect 33174 25332 33180 25334
rect 33244 25332 33250 25396
rect 33726 25332 33732 25396
rect 33796 25394 33802 25396
rect 35801 25394 35867 25397
rect 33796 25392 35867 25394
rect 33796 25336 35806 25392
rect 35862 25336 35867 25392
rect 33796 25334 35867 25336
rect 33796 25332 33802 25334
rect 35801 25331 35867 25334
rect 14457 25258 14523 25261
rect 22921 25258 22987 25261
rect 14457 25256 22987 25258
rect 14457 25200 14462 25256
rect 14518 25200 22926 25256
rect 22982 25200 22987 25256
rect 14457 25198 22987 25200
rect 14457 25195 14523 25198
rect 22921 25195 22987 25198
rect 25262 25196 25268 25260
rect 25332 25258 25338 25260
rect 25589 25258 25655 25261
rect 25332 25256 25655 25258
rect 25332 25200 25594 25256
rect 25650 25200 25655 25256
rect 25332 25198 25655 25200
rect 25332 25196 25338 25198
rect 25589 25195 25655 25198
rect 27613 25258 27679 25261
rect 30005 25258 30071 25261
rect 27613 25256 30071 25258
rect 27613 25200 27618 25256
rect 27674 25200 30010 25256
rect 30066 25200 30071 25256
rect 27613 25198 30071 25200
rect 27613 25195 27679 25198
rect 30005 25195 30071 25198
rect 30966 25196 30972 25260
rect 31036 25258 31042 25260
rect 35249 25258 35315 25261
rect 31036 25256 35315 25258
rect 31036 25200 35254 25256
rect 35310 25200 35315 25256
rect 31036 25198 35315 25200
rect 31036 25196 31042 25198
rect 35249 25195 35315 25198
rect 3785 25122 3851 25125
rect 18413 25122 18479 25125
rect 19425 25124 19491 25125
rect 19374 25122 19380 25124
rect 3785 25120 18479 25122
rect 3785 25064 3790 25120
rect 3846 25064 18418 25120
rect 18474 25064 18479 25120
rect 3785 25062 18479 25064
rect 19334 25062 19380 25122
rect 19444 25120 19491 25124
rect 19486 25064 19491 25120
rect 3785 25059 3851 25062
rect 18413 25059 18479 25062
rect 19374 25060 19380 25062
rect 19444 25060 19491 25064
rect 19425 25059 19491 25060
rect 19977 25122 20043 25125
rect 22461 25122 22527 25125
rect 19977 25120 22527 25122
rect 19977 25064 19982 25120
rect 20038 25064 22466 25120
rect 22522 25064 22527 25120
rect 19977 25062 22527 25064
rect 19977 25059 20043 25062
rect 22461 25059 22527 25062
rect 25405 25122 25471 25125
rect 32673 25122 32739 25125
rect 25405 25120 30988 25122
rect 25405 25064 25410 25120
rect 25466 25064 30988 25120
rect 25405 25062 30988 25064
rect 25405 25059 25471 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 15193 24986 15259 24989
rect 21725 24986 21791 24989
rect 22737 24986 22803 24989
rect 24853 24986 24919 24989
rect 15193 24984 16498 24986
rect 15193 24928 15198 24984
rect 15254 24928 16498 24984
rect 15193 24926 16498 24928
rect 15193 24923 15259 24926
rect 4061 24850 4127 24853
rect 16246 24850 16252 24852
rect 4061 24848 16252 24850
rect 4061 24792 4066 24848
rect 4122 24792 16252 24848
rect 4061 24790 16252 24792
rect 4061 24787 4127 24790
rect 16246 24788 16252 24790
rect 16316 24788 16322 24852
rect 16438 24850 16498 24926
rect 21725 24984 24919 24986
rect 21725 24928 21730 24984
rect 21786 24928 22742 24984
rect 22798 24928 24858 24984
rect 24914 24928 24919 24984
rect 21725 24926 24919 24928
rect 21725 24923 21791 24926
rect 22737 24923 22803 24926
rect 24853 24923 24919 24926
rect 25221 24986 25287 24989
rect 27889 24986 27955 24989
rect 25221 24984 27955 24986
rect 25221 24928 25226 24984
rect 25282 24928 27894 24984
rect 27950 24928 27955 24984
rect 25221 24926 27955 24928
rect 25221 24923 25287 24926
rect 27889 24923 27955 24926
rect 28625 24986 28691 24989
rect 28758 24986 28764 24988
rect 28625 24984 28764 24986
rect 28625 24928 28630 24984
rect 28686 24928 28764 24984
rect 28625 24926 28764 24928
rect 28625 24923 28691 24926
rect 28758 24924 28764 24926
rect 28828 24924 28834 24988
rect 29177 24986 29243 24989
rect 30465 24986 30531 24989
rect 29177 24984 30531 24986
rect 29177 24928 29182 24984
rect 29238 24928 30470 24984
rect 30526 24928 30531 24984
rect 29177 24926 30531 24928
rect 30928 24986 30988 25062
rect 31710 25120 32739 25122
rect 31710 25064 32678 25120
rect 32734 25064 32739 25120
rect 31710 25062 32739 25064
rect 31710 24986 31770 25062
rect 32673 25059 32739 25062
rect 33593 25122 33659 25125
rect 36077 25122 36143 25125
rect 33593 25120 36143 25122
rect 33593 25064 33598 25120
rect 33654 25064 36082 25120
rect 36138 25064 36143 25120
rect 33593 25062 36143 25064
rect 33593 25059 33659 25062
rect 36077 25059 36143 25062
rect 30928 24926 31770 24986
rect 32857 24986 32923 24989
rect 34053 24986 34119 24989
rect 32857 24984 34119 24986
rect 32857 24928 32862 24984
rect 32918 24928 34058 24984
rect 34114 24928 34119 24984
rect 32857 24926 34119 24928
rect 29177 24923 29243 24926
rect 30465 24923 30531 24926
rect 32857 24923 32923 24926
rect 34053 24923 34119 24926
rect 34881 24986 34947 24989
rect 35750 24986 35756 24988
rect 34881 24984 35756 24986
rect 34881 24928 34886 24984
rect 34942 24928 35756 24984
rect 34881 24926 35756 24928
rect 34881 24923 34947 24926
rect 35750 24924 35756 24926
rect 35820 24924 35826 24988
rect 23790 24850 23796 24852
rect 16438 24790 23796 24850
rect 23790 24788 23796 24790
rect 23860 24788 23866 24852
rect 23933 24850 23999 24853
rect 27797 24850 27863 24853
rect 23933 24848 27863 24850
rect 23933 24792 23938 24848
rect 23994 24792 27802 24848
rect 27858 24792 27863 24848
rect 23933 24790 27863 24792
rect 23933 24787 23999 24790
rect 27797 24787 27863 24790
rect 28625 24850 28691 24853
rect 28942 24850 28948 24852
rect 28625 24848 28948 24850
rect 28625 24792 28630 24848
rect 28686 24792 28948 24848
rect 28625 24790 28948 24792
rect 28625 24787 28691 24790
rect 28942 24788 28948 24790
rect 29012 24788 29018 24852
rect 29085 24850 29151 24853
rect 30782 24850 30788 24852
rect 29085 24848 30788 24850
rect 29085 24792 29090 24848
rect 29146 24792 30788 24848
rect 29085 24790 30788 24792
rect 29085 24787 29151 24790
rect 30782 24788 30788 24790
rect 30852 24788 30858 24852
rect 30925 24850 30991 24853
rect 32438 24850 32444 24852
rect 30925 24848 32444 24850
rect 30925 24792 30930 24848
rect 30986 24792 32444 24848
rect 30925 24790 32444 24792
rect 30925 24787 30991 24790
rect 32438 24788 32444 24790
rect 32508 24788 32514 24852
rect 32622 24788 32628 24852
rect 32692 24850 32698 24852
rect 35709 24850 35775 24853
rect 32692 24848 35775 24850
rect 32692 24792 35714 24848
rect 35770 24792 35775 24848
rect 32692 24790 35775 24792
rect 32692 24788 32698 24790
rect 35709 24787 35775 24790
rect 18045 24714 18111 24717
rect 20345 24714 20411 24717
rect 18045 24712 20411 24714
rect 18045 24656 18050 24712
rect 18106 24656 20350 24712
rect 20406 24656 20411 24712
rect 18045 24654 20411 24656
rect 18045 24651 18111 24654
rect 20345 24651 20411 24654
rect 20897 24714 20963 24717
rect 25497 24714 25563 24717
rect 20897 24712 25563 24714
rect 20897 24656 20902 24712
rect 20958 24656 25502 24712
rect 25558 24656 25563 24712
rect 20897 24654 25563 24656
rect 20897 24651 20963 24654
rect 25497 24651 25563 24654
rect 25957 24714 26023 24717
rect 26233 24714 26299 24717
rect 27981 24714 28047 24717
rect 35801 24714 35867 24717
rect 25957 24712 35867 24714
rect 25957 24656 25962 24712
rect 26018 24656 26238 24712
rect 26294 24656 27986 24712
rect 28042 24656 35806 24712
rect 35862 24656 35867 24712
rect 25957 24654 35867 24656
rect 25957 24651 26023 24654
rect 26233 24651 26299 24654
rect 27981 24651 28047 24654
rect 35801 24651 35867 24654
rect 38929 24714 38995 24717
rect 39200 24714 40000 24744
rect 38929 24712 40000 24714
rect 38929 24656 38934 24712
rect 38990 24656 40000 24712
rect 38929 24654 40000 24656
rect 38929 24651 38995 24654
rect 39200 24624 40000 24654
rect 5206 24516 5212 24580
rect 5276 24578 5282 24580
rect 20713 24578 20779 24581
rect 5276 24576 20779 24578
rect 5276 24520 20718 24576
rect 20774 24520 20779 24576
rect 5276 24518 20779 24520
rect 5276 24516 5282 24518
rect 20713 24515 20779 24518
rect 28073 24578 28139 24581
rect 30373 24578 30439 24581
rect 28073 24576 30439 24578
rect 28073 24520 28078 24576
rect 28134 24520 30378 24576
rect 30434 24520 30439 24576
rect 28073 24518 30439 24520
rect 28073 24515 28139 24518
rect 30373 24515 30439 24518
rect 30741 24578 30807 24581
rect 32949 24578 33015 24581
rect 30741 24576 33015 24578
rect 30741 24520 30746 24576
rect 30802 24520 32954 24576
rect 33010 24520 33015 24576
rect 30741 24518 33015 24520
rect 30741 24515 30807 24518
rect 32949 24515 33015 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 17769 24442 17835 24445
rect 31753 24442 31819 24445
rect 32397 24442 32463 24445
rect 33501 24444 33567 24445
rect 32806 24442 32812 24444
rect 17769 24440 32812 24442
rect 17769 24384 17774 24440
rect 17830 24384 31758 24440
rect 31814 24384 32402 24440
rect 32458 24384 32812 24440
rect 17769 24382 32812 24384
rect 17769 24379 17835 24382
rect 31753 24379 31819 24382
rect 32397 24379 32463 24382
rect 32806 24380 32812 24382
rect 32876 24380 32882 24444
rect 33501 24440 33548 24444
rect 33612 24442 33618 24444
rect 33501 24384 33506 24440
rect 33501 24380 33548 24384
rect 33612 24382 33658 24442
rect 33612 24380 33618 24382
rect 33501 24379 33567 24380
rect 19057 24306 19123 24309
rect 21725 24306 21791 24309
rect 19057 24304 21791 24306
rect 19057 24248 19062 24304
rect 19118 24248 21730 24304
rect 21786 24248 21791 24304
rect 19057 24246 21791 24248
rect 19057 24243 19123 24246
rect 21725 24243 21791 24246
rect 25037 24306 25103 24309
rect 27797 24306 27863 24309
rect 25037 24304 29010 24306
rect 25037 24248 25042 24304
rect 25098 24248 27802 24304
rect 27858 24248 29010 24304
rect 25037 24246 29010 24248
rect 25037 24243 25103 24246
rect 27797 24243 27863 24246
rect 19517 24170 19583 24173
rect 22185 24170 22251 24173
rect 19517 24168 22251 24170
rect 19517 24112 19522 24168
rect 19578 24112 22190 24168
rect 22246 24112 22251 24168
rect 19517 24110 22251 24112
rect 19517 24107 19583 24110
rect 22185 24107 22251 24110
rect 26141 24170 26207 24173
rect 27613 24170 27679 24173
rect 26141 24168 27679 24170
rect 26141 24112 26146 24168
rect 26202 24112 27618 24168
rect 27674 24112 27679 24168
rect 26141 24110 27679 24112
rect 28950 24170 29010 24246
rect 29126 24244 29132 24308
rect 29196 24306 29202 24308
rect 29453 24306 29519 24309
rect 29196 24304 29519 24306
rect 29196 24248 29458 24304
rect 29514 24248 29519 24304
rect 29196 24246 29519 24248
rect 29196 24244 29202 24246
rect 29453 24243 29519 24246
rect 31702 24244 31708 24308
rect 31772 24306 31778 24308
rect 39389 24306 39455 24309
rect 31772 24304 39455 24306
rect 31772 24248 39394 24304
rect 39450 24248 39455 24304
rect 31772 24246 39455 24248
rect 31772 24244 31778 24246
rect 39389 24243 39455 24246
rect 32857 24170 32923 24173
rect 28950 24168 32923 24170
rect 28950 24112 32862 24168
rect 32918 24112 32923 24168
rect 28950 24110 32923 24112
rect 26141 24107 26207 24110
rect 27613 24107 27679 24110
rect 32857 24107 32923 24110
rect 33593 24170 33659 24173
rect 34513 24170 34579 24173
rect 33593 24168 34579 24170
rect 33593 24112 33598 24168
rect 33654 24112 34518 24168
rect 34574 24112 34579 24168
rect 33593 24110 34579 24112
rect 33593 24107 33659 24110
rect 34513 24107 34579 24110
rect 26509 24034 26575 24037
rect 27429 24034 27495 24037
rect 26509 24032 27495 24034
rect 26509 23976 26514 24032
rect 26570 23976 27434 24032
rect 27490 23976 27495 24032
rect 26509 23974 27495 23976
rect 26509 23971 26575 23974
rect 27429 23971 27495 23974
rect 29085 24034 29151 24037
rect 29821 24034 29887 24037
rect 31753 24034 31819 24037
rect 29085 24032 31819 24034
rect 29085 23976 29090 24032
rect 29146 23976 29826 24032
rect 29882 23976 31758 24032
rect 31814 23976 31819 24032
rect 29085 23974 31819 23976
rect 29085 23971 29151 23974
rect 29821 23971 29887 23974
rect 31753 23971 31819 23974
rect 32857 24034 32923 24037
rect 32990 24034 32996 24036
rect 32857 24032 32996 24034
rect 32857 23976 32862 24032
rect 32918 23976 32996 24032
rect 32857 23974 32996 23976
rect 32857 23971 32923 23974
rect 32990 23972 32996 23974
rect 33060 23972 33066 24036
rect 33501 24034 33567 24037
rect 34053 24034 34119 24037
rect 35065 24034 35131 24037
rect 33501 24032 35131 24034
rect 33501 23976 33506 24032
rect 33562 23976 34058 24032
rect 34114 23976 35070 24032
rect 35126 23976 35131 24032
rect 33501 23974 35131 23976
rect 33501 23971 33567 23974
rect 34053 23971 34119 23974
rect 35065 23971 35131 23974
rect 35249 24034 35315 24037
rect 35750 24034 35756 24036
rect 35249 24032 35756 24034
rect 35249 23976 35254 24032
rect 35310 23976 35756 24032
rect 35249 23974 35756 23976
rect 35249 23971 35315 23974
rect 35750 23972 35756 23974
rect 35820 23972 35826 24036
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 28993 23898 29059 23901
rect 22050 23896 29059 23898
rect 22050 23840 28998 23896
rect 29054 23840 29059 23896
rect 22050 23838 29059 23840
rect 17677 23762 17743 23765
rect 22050 23762 22110 23838
rect 28993 23835 29059 23838
rect 29494 23836 29500 23900
rect 29564 23898 29570 23900
rect 30833 23898 30899 23901
rect 29564 23896 30899 23898
rect 29564 23840 30838 23896
rect 30894 23840 30899 23896
rect 29564 23838 30899 23840
rect 29564 23836 29570 23838
rect 30833 23835 30899 23838
rect 31937 23898 32003 23901
rect 36169 23898 36235 23901
rect 31937 23896 36235 23898
rect 31937 23840 31942 23896
rect 31998 23840 36174 23896
rect 36230 23840 36235 23896
rect 31937 23838 36235 23840
rect 31937 23835 32003 23838
rect 32492 23765 32552 23838
rect 36169 23835 36235 23838
rect 17677 23760 22110 23762
rect 17677 23704 17682 23760
rect 17738 23704 22110 23760
rect 17677 23702 22110 23704
rect 27153 23762 27219 23765
rect 29729 23762 29795 23765
rect 27153 23760 29795 23762
rect 27153 23704 27158 23760
rect 27214 23704 29734 23760
rect 29790 23704 29795 23760
rect 27153 23702 29795 23704
rect 17677 23699 17743 23702
rect 27153 23699 27219 23702
rect 29729 23699 29795 23702
rect 30741 23762 30807 23765
rect 30966 23762 30972 23764
rect 30741 23760 30972 23762
rect 30741 23704 30746 23760
rect 30802 23704 30972 23760
rect 30741 23702 30972 23704
rect 30741 23699 30807 23702
rect 30966 23700 30972 23702
rect 31036 23762 31042 23764
rect 31293 23762 31359 23765
rect 31036 23760 31359 23762
rect 31036 23704 31298 23760
rect 31354 23704 31359 23760
rect 31036 23702 31359 23704
rect 31036 23700 31042 23702
rect 31293 23699 31359 23702
rect 32489 23760 32555 23765
rect 32489 23704 32494 23760
rect 32550 23704 32555 23760
rect 32489 23699 32555 23704
rect 34646 23700 34652 23764
rect 34716 23762 34722 23764
rect 35433 23762 35499 23765
rect 34716 23760 35499 23762
rect 34716 23704 35438 23760
rect 35494 23704 35499 23760
rect 34716 23702 35499 23704
rect 34716 23700 34722 23702
rect 35433 23699 35499 23702
rect 18781 23626 18847 23629
rect 20713 23626 20779 23629
rect 18781 23624 20779 23626
rect 18781 23568 18786 23624
rect 18842 23568 20718 23624
rect 20774 23568 20779 23624
rect 18781 23566 20779 23568
rect 18781 23563 18847 23566
rect 20713 23563 20779 23566
rect 23197 23626 23263 23629
rect 27521 23626 27587 23629
rect 23197 23624 27587 23626
rect 23197 23568 23202 23624
rect 23258 23568 27526 23624
rect 27582 23568 27587 23624
rect 23197 23566 27587 23568
rect 23197 23563 23263 23566
rect 27521 23563 27587 23566
rect 29453 23626 29519 23629
rect 32857 23626 32923 23629
rect 37273 23626 37339 23629
rect 29453 23624 32923 23626
rect 29453 23568 29458 23624
rect 29514 23568 32862 23624
rect 32918 23568 32923 23624
rect 29453 23566 32923 23568
rect 29453 23563 29519 23566
rect 32857 23563 32923 23566
rect 33182 23624 37339 23626
rect 33182 23568 37278 23624
rect 37334 23568 37339 23624
rect 33182 23566 37339 23568
rect 17309 23490 17375 23493
rect 18965 23490 19031 23493
rect 17309 23488 19031 23490
rect 17309 23432 17314 23488
rect 17370 23432 18970 23488
rect 19026 23432 19031 23488
rect 17309 23430 19031 23432
rect 17309 23427 17375 23430
rect 18965 23427 19031 23430
rect 19241 23490 19307 23493
rect 24301 23490 24367 23493
rect 27654 23490 27660 23492
rect 19241 23488 24367 23490
rect 19241 23432 19246 23488
rect 19302 23432 24306 23488
rect 24362 23432 24367 23488
rect 19241 23430 24367 23432
rect 19241 23427 19307 23430
rect 24301 23427 24367 23430
rect 26926 23430 27660 23490
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 19149 23354 19215 23357
rect 20437 23354 20503 23357
rect 19149 23352 20503 23354
rect 19149 23296 19154 23352
rect 19210 23296 20442 23352
rect 20498 23296 20503 23352
rect 19149 23294 20503 23296
rect 19149 23291 19215 23294
rect 20437 23291 20503 23294
rect 20713 23354 20779 23357
rect 26926 23354 26986 23430
rect 27654 23428 27660 23430
rect 27724 23428 27730 23492
rect 28206 23428 28212 23492
rect 28276 23490 28282 23492
rect 28441 23490 28507 23493
rect 28276 23488 28507 23490
rect 28276 23432 28446 23488
rect 28502 23432 28507 23488
rect 28276 23430 28507 23432
rect 28276 23428 28282 23430
rect 28441 23427 28507 23430
rect 28574 23428 28580 23492
rect 28644 23490 28650 23492
rect 29085 23490 29151 23493
rect 28644 23488 29151 23490
rect 28644 23432 29090 23488
rect 29146 23432 29151 23488
rect 28644 23430 29151 23432
rect 28644 23428 28650 23430
rect 29085 23427 29151 23430
rect 31753 23490 31819 23493
rect 33182 23490 33242 23566
rect 37273 23563 37339 23566
rect 31753 23488 33242 23490
rect 31753 23432 31758 23488
rect 31814 23432 33242 23488
rect 31753 23430 33242 23432
rect 31753 23427 31819 23430
rect 33542 23428 33548 23492
rect 33612 23490 33618 23492
rect 34145 23490 34211 23493
rect 33612 23488 34211 23490
rect 33612 23432 34150 23488
rect 34206 23432 34211 23488
rect 33612 23430 34211 23432
rect 33612 23428 33618 23430
rect 34145 23427 34211 23430
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 20713 23352 26986 23354
rect 20713 23296 20718 23352
rect 20774 23296 26986 23352
rect 20713 23294 26986 23296
rect 28257 23354 28323 23357
rect 33685 23354 33751 23357
rect 28257 23352 33751 23354
rect 28257 23296 28262 23352
rect 28318 23296 33690 23352
rect 33746 23296 33751 23352
rect 28257 23294 33751 23296
rect 20713 23291 20779 23294
rect 28257 23291 28323 23294
rect 33685 23291 33751 23294
rect 38837 23354 38903 23357
rect 39200 23354 40000 23384
rect 38837 23352 40000 23354
rect 38837 23296 38842 23352
rect 38898 23296 40000 23352
rect 38837 23294 40000 23296
rect 38837 23291 38903 23294
rect 39200 23264 40000 23294
rect 7005 23218 7071 23221
rect 25405 23218 25471 23221
rect 7005 23216 25471 23218
rect 7005 23160 7010 23216
rect 7066 23160 25410 23216
rect 25466 23160 25471 23216
rect 7005 23158 25471 23160
rect 7005 23155 7071 23158
rect 25405 23155 25471 23158
rect 26182 23156 26188 23220
rect 26252 23218 26258 23220
rect 26785 23218 26851 23221
rect 26252 23216 26851 23218
rect 26252 23160 26790 23216
rect 26846 23160 26851 23216
rect 26252 23158 26851 23160
rect 26252 23156 26258 23158
rect 26785 23155 26851 23158
rect 27102 23156 27108 23220
rect 27172 23218 27178 23220
rect 29453 23218 29519 23221
rect 27172 23216 29519 23218
rect 27172 23160 29458 23216
rect 29514 23160 29519 23216
rect 27172 23158 29519 23160
rect 27172 23156 27178 23158
rect 29453 23155 29519 23158
rect 30005 23218 30071 23221
rect 30649 23218 30715 23221
rect 30005 23216 30715 23218
rect 30005 23160 30010 23216
rect 30066 23160 30654 23216
rect 30710 23160 30715 23216
rect 30005 23158 30715 23160
rect 30005 23155 30071 23158
rect 30649 23155 30715 23158
rect 31293 23218 31359 23221
rect 34646 23218 34652 23220
rect 31293 23216 34652 23218
rect 31293 23160 31298 23216
rect 31354 23160 34652 23216
rect 31293 23158 34652 23160
rect 31293 23155 31359 23158
rect 34646 23156 34652 23158
rect 34716 23156 34722 23220
rect 35934 23156 35940 23220
rect 36004 23218 36010 23220
rect 37457 23218 37523 23221
rect 36004 23216 37523 23218
rect 36004 23160 37462 23216
rect 37518 23160 37523 23216
rect 36004 23158 37523 23160
rect 36004 23156 36010 23158
rect 37457 23155 37523 23158
rect 10358 23020 10364 23084
rect 10428 23082 10434 23084
rect 22737 23082 22803 23085
rect 10428 23080 22803 23082
rect 10428 23024 22742 23080
rect 22798 23024 22803 23080
rect 10428 23022 22803 23024
rect 10428 23020 10434 23022
rect 22737 23019 22803 23022
rect 23657 23082 23723 23085
rect 24577 23082 24643 23085
rect 23657 23080 24643 23082
rect 23657 23024 23662 23080
rect 23718 23024 24582 23080
rect 24638 23024 24643 23080
rect 23657 23022 24643 23024
rect 23657 23019 23723 23022
rect 24577 23019 24643 23022
rect 30649 23082 30715 23085
rect 32489 23082 32555 23085
rect 30649 23080 32555 23082
rect 30649 23024 30654 23080
rect 30710 23024 32494 23080
rect 32550 23024 32555 23080
rect 30649 23022 32555 23024
rect 30649 23019 30715 23022
rect 32489 23019 32555 23022
rect 32857 23082 32923 23085
rect 33225 23082 33291 23085
rect 36997 23082 37063 23085
rect 32857 23080 37063 23082
rect 32857 23024 32862 23080
rect 32918 23024 33230 23080
rect 33286 23024 37002 23080
rect 37058 23024 37063 23080
rect 32857 23022 37063 23024
rect 32857 23019 32923 23022
rect 33225 23019 33291 23022
rect 36997 23019 37063 23022
rect 20253 22946 20319 22949
rect 22277 22946 22343 22949
rect 20253 22944 22343 22946
rect 20253 22888 20258 22944
rect 20314 22888 22282 22944
rect 22338 22888 22343 22944
rect 20253 22886 22343 22888
rect 20253 22883 20319 22886
rect 22277 22883 22343 22886
rect 22829 22946 22895 22949
rect 23422 22946 23428 22948
rect 22829 22944 23428 22946
rect 22829 22888 22834 22944
rect 22890 22888 23428 22944
rect 22829 22886 23428 22888
rect 22829 22883 22895 22886
rect 23422 22884 23428 22886
rect 23492 22884 23498 22948
rect 30281 22946 30347 22949
rect 32397 22946 32463 22949
rect 30281 22944 32463 22946
rect 30281 22888 30286 22944
rect 30342 22888 32402 22944
rect 32458 22888 32463 22944
rect 30281 22886 32463 22888
rect 30281 22883 30347 22886
rect 32397 22883 32463 22886
rect 33133 22946 33199 22949
rect 33358 22946 33364 22948
rect 33133 22944 33364 22946
rect 33133 22888 33138 22944
rect 33194 22888 33364 22944
rect 33133 22886 33364 22888
rect 33133 22883 33199 22886
rect 33358 22884 33364 22886
rect 33428 22884 33434 22948
rect 33777 22946 33843 22949
rect 34421 22946 34487 22949
rect 33777 22944 34487 22946
rect 33777 22888 33782 22944
rect 33838 22888 34426 22944
rect 34482 22888 34487 22944
rect 33777 22886 34487 22888
rect 33777 22883 33843 22886
rect 34421 22883 34487 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 27470 22748 27476 22812
rect 27540 22810 27546 22812
rect 28441 22810 28507 22813
rect 27540 22808 28507 22810
rect 27540 22752 28446 22808
rect 28502 22752 28507 22808
rect 27540 22750 28507 22752
rect 27540 22748 27546 22750
rect 28441 22747 28507 22750
rect 29729 22810 29795 22813
rect 36813 22810 36879 22813
rect 29729 22808 36879 22810
rect 29729 22752 29734 22808
rect 29790 22752 36818 22808
rect 36874 22752 36879 22808
rect 29729 22750 36879 22752
rect 29729 22747 29795 22750
rect 36813 22747 36879 22750
rect 3693 22674 3759 22677
rect 23197 22674 23263 22677
rect 3693 22672 23263 22674
rect 3693 22616 3698 22672
rect 3754 22616 23202 22672
rect 23258 22616 23263 22672
rect 3693 22614 23263 22616
rect 3693 22611 3759 22614
rect 23197 22611 23263 22614
rect 26366 22612 26372 22676
rect 26436 22674 26442 22676
rect 28993 22674 29059 22677
rect 26436 22672 29059 22674
rect 26436 22616 28998 22672
rect 29054 22616 29059 22672
rect 26436 22614 29059 22616
rect 26436 22612 26442 22614
rect 28993 22611 29059 22614
rect 30414 22612 30420 22676
rect 30484 22674 30490 22676
rect 30833 22674 30899 22677
rect 30484 22672 30899 22674
rect 30484 22616 30838 22672
rect 30894 22616 30899 22672
rect 30484 22614 30899 22616
rect 30484 22612 30490 22614
rect 30833 22611 30899 22614
rect 32489 22674 32555 22677
rect 33910 22674 33916 22676
rect 32489 22672 33916 22674
rect 32489 22616 32494 22672
rect 32550 22616 33916 22672
rect 32489 22614 33916 22616
rect 32489 22611 32555 22614
rect 33910 22612 33916 22614
rect 33980 22612 33986 22676
rect 35382 22674 35388 22676
rect 34102 22614 35388 22674
rect 18045 22538 18111 22541
rect 19793 22538 19859 22541
rect 18045 22536 19859 22538
rect 18045 22480 18050 22536
rect 18106 22480 19798 22536
rect 19854 22480 19859 22536
rect 18045 22478 19859 22480
rect 18045 22475 18111 22478
rect 19793 22475 19859 22478
rect 21950 22476 21956 22540
rect 22020 22538 22026 22540
rect 25221 22538 25287 22541
rect 25957 22538 26023 22541
rect 28993 22538 29059 22541
rect 22020 22536 29059 22538
rect 22020 22480 25226 22536
rect 25282 22480 25962 22536
rect 26018 22480 28998 22536
rect 29054 22480 29059 22536
rect 22020 22478 29059 22480
rect 22020 22476 22026 22478
rect 25221 22475 25287 22478
rect 25957 22475 26023 22478
rect 28993 22475 29059 22478
rect 29545 22538 29611 22541
rect 29862 22538 29868 22540
rect 29545 22536 29868 22538
rect 29545 22480 29550 22536
rect 29606 22480 29868 22536
rect 29545 22478 29868 22480
rect 29545 22475 29611 22478
rect 29862 22476 29868 22478
rect 29932 22476 29938 22540
rect 30189 22538 30255 22541
rect 32254 22538 32260 22540
rect 30189 22536 32260 22538
rect 30189 22480 30194 22536
rect 30250 22480 32260 22536
rect 30189 22478 32260 22480
rect 30189 22475 30255 22478
rect 32254 22476 32260 22478
rect 32324 22476 32330 22540
rect 32397 22538 32463 22541
rect 34102 22538 34162 22614
rect 35382 22612 35388 22614
rect 35452 22612 35458 22676
rect 34881 22538 34947 22541
rect 32397 22536 34162 22538
rect 32397 22480 32402 22536
rect 32458 22480 34162 22536
rect 32397 22478 34162 22480
rect 34516 22536 34947 22538
rect 34516 22480 34886 22536
rect 34942 22480 34947 22536
rect 34516 22478 34947 22480
rect 32397 22475 32463 22478
rect 34516 22405 34576 22478
rect 34881 22475 34947 22478
rect 20161 22402 20227 22405
rect 25681 22402 25747 22405
rect 33869 22404 33935 22405
rect 33869 22402 33916 22404
rect 20161 22400 25747 22402
rect 20161 22344 20166 22400
rect 20222 22344 25686 22400
rect 25742 22344 25747 22400
rect 20161 22342 25747 22344
rect 33824 22400 33916 22402
rect 33824 22344 33874 22400
rect 33824 22342 33916 22344
rect 20161 22339 20227 22342
rect 25681 22339 25747 22342
rect 33869 22340 33916 22342
rect 33980 22340 33986 22404
rect 34513 22400 34579 22405
rect 34513 22344 34518 22400
rect 34574 22344 34579 22400
rect 33869 22339 33935 22340
rect 34513 22339 34579 22344
rect 35341 22402 35407 22405
rect 35617 22402 35683 22405
rect 35341 22400 35683 22402
rect 35341 22344 35346 22400
rect 35402 22344 35622 22400
rect 35678 22344 35683 22400
rect 35341 22342 35683 22344
rect 35341 22339 35407 22342
rect 35617 22339 35683 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 9622 22204 9628 22268
rect 9692 22266 9698 22268
rect 34605 22266 34671 22269
rect 9692 22206 27860 22266
rect 9692 22204 9698 22206
rect 25814 22130 25820 22132
rect 23614 22070 25820 22130
rect 5073 21994 5139 21997
rect 19885 21994 19951 21997
rect 21950 21994 21956 21996
rect 5073 21992 6930 21994
rect 5073 21936 5078 21992
rect 5134 21936 6930 21992
rect 5073 21934 6930 21936
rect 5073 21931 5139 21934
rect 6870 21586 6930 21934
rect 19885 21992 21956 21994
rect 19885 21936 19890 21992
rect 19946 21936 21956 21992
rect 19885 21934 21956 21936
rect 19885 21931 19951 21934
rect 21950 21932 21956 21934
rect 22020 21932 22026 21996
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 20069 21722 20135 21725
rect 21633 21722 21699 21725
rect 20069 21720 21699 21722
rect 20069 21664 20074 21720
rect 20130 21664 21638 21720
rect 21694 21664 21699 21720
rect 20069 21662 21699 21664
rect 20069 21659 20135 21662
rect 21633 21659 21699 21662
rect 23614 21586 23674 22070
rect 25814 22068 25820 22070
rect 25884 22068 25890 22132
rect 27800 22130 27860 22206
rect 30054 22264 34671 22266
rect 30054 22208 34610 22264
rect 34666 22208 34671 22264
rect 30054 22206 34671 22208
rect 29545 22130 29611 22133
rect 29678 22130 29684 22132
rect 27800 22128 29684 22130
rect 27800 22072 29550 22128
rect 29606 22072 29684 22128
rect 27800 22070 29684 22072
rect 29545 22067 29611 22070
rect 29678 22068 29684 22070
rect 29748 22068 29754 22132
rect 24117 21994 24183 21997
rect 24342 21994 24348 21996
rect 24117 21992 24348 21994
rect 24117 21936 24122 21992
rect 24178 21936 24348 21992
rect 24117 21934 24348 21936
rect 24117 21931 24183 21934
rect 24342 21932 24348 21934
rect 24412 21932 24418 21996
rect 28993 21994 29059 21997
rect 30054 21994 30114 22206
rect 34605 22203 34671 22206
rect 30373 22130 30439 22133
rect 32070 22130 32076 22132
rect 30373 22128 32076 22130
rect 30373 22072 30378 22128
rect 30434 22072 32076 22128
rect 30373 22070 32076 22072
rect 30373 22067 30439 22070
rect 32070 22068 32076 22070
rect 32140 22068 32146 22132
rect 34462 22068 34468 22132
rect 34532 22130 34538 22132
rect 35433 22130 35499 22133
rect 34532 22128 35499 22130
rect 34532 22072 35438 22128
rect 35494 22072 35499 22128
rect 34532 22070 35499 22072
rect 34532 22068 34538 22070
rect 35433 22067 35499 22070
rect 28993 21992 30114 21994
rect 28993 21936 28998 21992
rect 29054 21936 30114 21992
rect 28993 21934 30114 21936
rect 30465 21994 30531 21997
rect 35065 21994 35131 21997
rect 35566 21994 35572 21996
rect 30465 21992 35572 21994
rect 30465 21936 30470 21992
rect 30526 21936 35070 21992
rect 35126 21936 35572 21992
rect 30465 21934 35572 21936
rect 28993 21931 29059 21934
rect 30465 21931 30531 21934
rect 35065 21931 35131 21934
rect 35566 21932 35572 21934
rect 35636 21932 35642 21996
rect 39021 21994 39087 21997
rect 39200 21994 40000 22024
rect 39021 21992 40000 21994
rect 39021 21936 39026 21992
rect 39082 21936 40000 21992
rect 39021 21934 40000 21936
rect 39021 21931 39087 21934
rect 39200 21904 40000 21934
rect 27286 21796 27292 21860
rect 27356 21858 27362 21860
rect 30097 21858 30163 21861
rect 27356 21856 30163 21858
rect 27356 21800 30102 21856
rect 30158 21800 30163 21856
rect 27356 21798 30163 21800
rect 27356 21796 27362 21798
rect 30097 21795 30163 21798
rect 30966 21796 30972 21860
rect 31036 21858 31042 21860
rect 31109 21858 31175 21861
rect 31036 21856 31175 21858
rect 31036 21800 31114 21856
rect 31170 21800 31175 21856
rect 31036 21798 31175 21800
rect 31036 21796 31042 21798
rect 31109 21795 31175 21798
rect 31518 21796 31524 21860
rect 31588 21858 31594 21860
rect 32305 21858 32371 21861
rect 31588 21856 32371 21858
rect 31588 21800 32310 21856
rect 32366 21800 32371 21856
rect 31588 21798 32371 21800
rect 31588 21796 31594 21798
rect 32305 21795 32371 21798
rect 25998 21660 26004 21724
rect 26068 21722 26074 21724
rect 34237 21722 34303 21725
rect 26068 21720 34303 21722
rect 26068 21664 34242 21720
rect 34298 21664 34303 21720
rect 26068 21662 34303 21664
rect 26068 21660 26074 21662
rect 34237 21659 34303 21662
rect 6870 21526 23674 21586
rect 24158 21524 24164 21588
rect 24228 21586 24234 21588
rect 28901 21586 28967 21589
rect 29310 21586 29316 21588
rect 24228 21584 29316 21586
rect 24228 21528 28906 21584
rect 28962 21528 29316 21584
rect 24228 21526 29316 21528
rect 24228 21524 24234 21526
rect 28901 21523 28967 21526
rect 29310 21524 29316 21526
rect 29380 21524 29386 21588
rect 30281 21586 30347 21589
rect 36629 21586 36695 21589
rect 37038 21586 37044 21588
rect 30281 21584 37044 21586
rect 30281 21528 30286 21584
rect 30342 21528 36634 21584
rect 36690 21528 37044 21584
rect 30281 21526 37044 21528
rect 30281 21523 30347 21526
rect 36629 21523 36695 21526
rect 37038 21524 37044 21526
rect 37108 21524 37114 21588
rect 19885 21450 19951 21453
rect 25037 21450 25103 21453
rect 19885 21448 25103 21450
rect 19885 21392 19890 21448
rect 19946 21392 25042 21448
rect 25098 21392 25103 21448
rect 19885 21390 25103 21392
rect 19885 21387 19951 21390
rect 25037 21387 25103 21390
rect 31201 21450 31267 21453
rect 39205 21450 39271 21453
rect 31201 21448 39271 21450
rect 31201 21392 31206 21448
rect 31262 21392 39210 21448
rect 39266 21392 39271 21448
rect 31201 21390 39271 21392
rect 31201 21387 31267 21390
rect 39205 21387 39271 21390
rect 22502 21252 22508 21316
rect 22572 21314 22578 21316
rect 24301 21314 24367 21317
rect 22572 21312 24367 21314
rect 22572 21256 24306 21312
rect 24362 21256 24367 21312
rect 22572 21254 24367 21256
rect 22572 21252 22578 21254
rect 24301 21251 24367 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 22461 21178 22527 21181
rect 24485 21178 24551 21181
rect 22461 21176 24551 21178
rect 22461 21120 22466 21176
rect 22522 21120 24490 21176
rect 24546 21120 24551 21176
rect 22461 21118 24551 21120
rect 22461 21115 22527 21118
rect 24485 21115 24551 21118
rect 27153 21178 27219 21181
rect 32213 21178 32279 21181
rect 33726 21178 33732 21180
rect 27153 21176 29010 21178
rect 27153 21120 27158 21176
rect 27214 21120 29010 21176
rect 27153 21118 29010 21120
rect 27153 21115 27219 21118
rect 18229 21042 18295 21045
rect 22829 21042 22895 21045
rect 18229 21040 22895 21042
rect 18229 20984 18234 21040
rect 18290 20984 22834 21040
rect 22890 20984 22895 21040
rect 18229 20982 22895 20984
rect 28950 21042 29010 21118
rect 32213 21176 33732 21178
rect 32213 21120 32218 21176
rect 32274 21120 33732 21176
rect 32213 21118 33732 21120
rect 32213 21115 32279 21118
rect 33726 21116 33732 21118
rect 33796 21116 33802 21180
rect 33777 21042 33843 21045
rect 28950 21040 33843 21042
rect 28950 20984 33782 21040
rect 33838 20984 33843 21040
rect 28950 20982 33843 20984
rect 18229 20979 18295 20982
rect 22829 20979 22895 20982
rect 33777 20979 33843 20982
rect 17125 20906 17191 20909
rect 26601 20906 26667 20909
rect 17125 20904 26667 20906
rect 17125 20848 17130 20904
rect 17186 20848 26606 20904
rect 26662 20848 26667 20904
rect 17125 20846 26667 20848
rect 17125 20843 17191 20846
rect 26601 20843 26667 20846
rect 28533 20906 28599 20909
rect 30046 20906 30052 20908
rect 28533 20904 30052 20906
rect 28533 20848 28538 20904
rect 28594 20848 30052 20904
rect 28533 20846 30052 20848
rect 28533 20843 28599 20846
rect 30046 20844 30052 20846
rect 30116 20906 30122 20908
rect 37641 20906 37707 20909
rect 30116 20904 37707 20906
rect 30116 20848 37646 20904
rect 37702 20848 37707 20904
rect 30116 20846 37707 20848
rect 30116 20844 30122 20846
rect 37641 20843 37707 20846
rect 32305 20770 32371 20773
rect 32949 20772 33015 20773
rect 32622 20770 32628 20772
rect 32305 20768 32628 20770
rect 32305 20712 32310 20768
rect 32366 20712 32628 20768
rect 32305 20710 32628 20712
rect 32305 20707 32371 20710
rect 32622 20708 32628 20710
rect 32692 20708 32698 20772
rect 32949 20768 32996 20772
rect 33060 20770 33066 20772
rect 33961 20770 34027 20773
rect 38285 20770 38351 20773
rect 32949 20712 32954 20768
rect 32949 20708 32996 20712
rect 33060 20710 33106 20770
rect 33961 20768 38351 20770
rect 33961 20712 33966 20768
rect 34022 20712 38290 20768
rect 38346 20712 38351 20768
rect 33961 20710 38351 20712
rect 33060 20708 33066 20710
rect 32949 20707 33015 20708
rect 33961 20707 34027 20710
rect 38285 20707 38351 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 12433 20634 12499 20637
rect 13997 20634 14063 20637
rect 12433 20632 14063 20634
rect 12433 20576 12438 20632
rect 12494 20576 14002 20632
rect 14058 20576 14063 20632
rect 12433 20574 14063 20576
rect 12433 20571 12499 20574
rect 13997 20571 14063 20574
rect 22645 20634 22711 20637
rect 23105 20634 23171 20637
rect 27337 20634 27403 20637
rect 22645 20632 27403 20634
rect 22645 20576 22650 20632
rect 22706 20576 23110 20632
rect 23166 20576 27342 20632
rect 27398 20576 27403 20632
rect 22645 20574 27403 20576
rect 22645 20571 22711 20574
rect 23105 20571 23171 20574
rect 27337 20571 27403 20574
rect 28349 20636 28415 20637
rect 28349 20632 28396 20636
rect 28460 20634 28466 20636
rect 28993 20634 29059 20637
rect 29729 20634 29795 20637
rect 28349 20576 28354 20632
rect 28349 20572 28396 20576
rect 28460 20574 28506 20634
rect 28993 20632 29795 20634
rect 28993 20576 28998 20632
rect 29054 20576 29734 20632
rect 29790 20576 29795 20632
rect 28993 20574 29795 20576
rect 28460 20572 28466 20574
rect 28349 20571 28415 20572
rect 28993 20571 29059 20574
rect 29729 20571 29795 20574
rect 33225 20634 33291 20637
rect 34237 20634 34303 20637
rect 33225 20632 34303 20634
rect 33225 20576 33230 20632
rect 33286 20576 34242 20632
rect 34298 20576 34303 20632
rect 33225 20574 34303 20576
rect 33225 20571 33291 20574
rect 34237 20571 34303 20574
rect 38929 20634 38995 20637
rect 39200 20634 40000 20664
rect 38929 20632 40000 20634
rect 38929 20576 38934 20632
rect 38990 20576 40000 20632
rect 38929 20574 40000 20576
rect 38929 20571 38995 20574
rect 39200 20544 40000 20574
rect 18045 20498 18111 20501
rect 22921 20498 22987 20501
rect 18045 20496 22987 20498
rect 18045 20440 18050 20496
rect 18106 20440 22926 20496
rect 22982 20440 22987 20496
rect 18045 20438 22987 20440
rect 18045 20435 18111 20438
rect 22921 20435 22987 20438
rect 24025 20498 24091 20501
rect 29545 20498 29611 20501
rect 24025 20496 29611 20498
rect 24025 20440 24030 20496
rect 24086 20440 29550 20496
rect 29606 20440 29611 20496
rect 24025 20438 29611 20440
rect 24025 20435 24091 20438
rect 29545 20435 29611 20438
rect 31845 20498 31911 20501
rect 32438 20498 32444 20500
rect 31845 20496 32444 20498
rect 31845 20440 31850 20496
rect 31906 20440 32444 20496
rect 31845 20438 32444 20440
rect 31845 20435 31911 20438
rect 32438 20436 32444 20438
rect 32508 20436 32514 20500
rect 32622 20436 32628 20500
rect 32692 20498 32698 20500
rect 32806 20498 32812 20500
rect 32692 20438 32812 20498
rect 32692 20436 32698 20438
rect 32806 20436 32812 20438
rect 32876 20498 32882 20500
rect 32949 20498 33015 20501
rect 32876 20496 33015 20498
rect 32876 20440 32954 20496
rect 33010 20440 33015 20496
rect 32876 20438 33015 20440
rect 32876 20436 32882 20438
rect 32949 20435 33015 20438
rect 34278 20436 34284 20500
rect 34348 20498 34354 20500
rect 34421 20498 34487 20501
rect 34348 20496 34487 20498
rect 34348 20440 34426 20496
rect 34482 20440 34487 20496
rect 34348 20438 34487 20440
rect 34348 20436 34354 20438
rect 34421 20435 34487 20438
rect 34973 20498 35039 20501
rect 38469 20498 38535 20501
rect 34973 20496 38535 20498
rect 34973 20440 34978 20496
rect 35034 20440 38474 20496
rect 38530 20440 38535 20496
rect 34973 20438 38535 20440
rect 34973 20435 35039 20438
rect 38469 20435 38535 20438
rect 18137 20362 18203 20365
rect 28349 20362 28415 20365
rect 18137 20360 28415 20362
rect 18137 20304 18142 20360
rect 18198 20304 28354 20360
rect 28410 20304 28415 20360
rect 18137 20302 28415 20304
rect 18137 20299 18203 20302
rect 28349 20299 28415 20302
rect 29177 20362 29243 20365
rect 32765 20362 32831 20365
rect 35985 20362 36051 20365
rect 29177 20360 32831 20362
rect 29177 20304 29182 20360
rect 29238 20304 32770 20360
rect 32826 20304 32831 20360
rect 29177 20302 32831 20304
rect 29177 20299 29243 20302
rect 32765 20299 32831 20302
rect 33964 20360 36051 20362
rect 33964 20304 35990 20360
rect 36046 20304 36051 20360
rect 33964 20302 36051 20304
rect 33964 20229 34024 20302
rect 35985 20299 36051 20302
rect 28758 20164 28764 20228
rect 28828 20226 28834 20228
rect 30373 20226 30439 20229
rect 28828 20224 30439 20226
rect 28828 20168 30378 20224
rect 30434 20168 30439 20224
rect 28828 20166 30439 20168
rect 28828 20164 28834 20166
rect 30373 20163 30439 20166
rect 30598 20164 30604 20228
rect 30668 20226 30674 20228
rect 33961 20226 34027 20229
rect 30668 20224 34027 20226
rect 30668 20168 33966 20224
rect 34022 20168 34027 20224
rect 30668 20166 34027 20168
rect 30668 20164 30674 20166
rect 33961 20163 34027 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 20069 20090 20135 20093
rect 25129 20090 25195 20093
rect 20069 20088 25195 20090
rect 20069 20032 20074 20088
rect 20130 20032 25134 20088
rect 25190 20032 25195 20088
rect 20069 20030 25195 20032
rect 20069 20027 20135 20030
rect 25129 20027 25195 20030
rect 26049 20090 26115 20093
rect 26550 20090 26556 20092
rect 26049 20088 26556 20090
rect 26049 20032 26054 20088
rect 26110 20032 26556 20088
rect 26049 20030 26556 20032
rect 26049 20027 26115 20030
rect 26550 20028 26556 20030
rect 26620 20090 26626 20092
rect 33593 20090 33659 20093
rect 34278 20090 34284 20092
rect 26620 20030 33288 20090
rect 26620 20028 26626 20030
rect 33228 19957 33288 20030
rect 33593 20088 34284 20090
rect 33593 20032 33598 20088
rect 33654 20032 34284 20088
rect 33593 20030 34284 20032
rect 33593 20027 33659 20030
rect 34278 20028 34284 20030
rect 34348 20028 34354 20092
rect 22185 19954 22251 19957
rect 23197 19954 23263 19957
rect 24025 19954 24091 19957
rect 22185 19952 24091 19954
rect 22185 19896 22190 19952
rect 22246 19896 23202 19952
rect 23258 19896 24030 19952
rect 24086 19896 24091 19952
rect 22185 19894 24091 19896
rect 22185 19891 22251 19894
rect 23197 19891 23263 19894
rect 24025 19891 24091 19894
rect 28993 19954 29059 19957
rect 32489 19954 32555 19957
rect 28993 19952 32555 19954
rect 28993 19896 28998 19952
rect 29054 19896 32494 19952
rect 32550 19896 32555 19952
rect 28993 19894 32555 19896
rect 28993 19891 29059 19894
rect 32489 19891 32555 19894
rect 33225 19952 33291 19957
rect 33225 19896 33230 19952
rect 33286 19896 33291 19952
rect 33225 19891 33291 19896
rect 22093 19818 22159 19821
rect 28257 19818 28323 19821
rect 22093 19816 28323 19818
rect 22093 19760 22098 19816
rect 22154 19760 28262 19816
rect 28318 19760 28323 19816
rect 22093 19758 28323 19760
rect 22093 19755 22159 19758
rect 28257 19755 28323 19758
rect 29453 19818 29519 19821
rect 30598 19818 30604 19820
rect 29453 19816 30604 19818
rect 29453 19760 29458 19816
rect 29514 19760 30604 19816
rect 29453 19758 30604 19760
rect 29453 19755 29519 19758
rect 30598 19756 30604 19758
rect 30668 19756 30674 19820
rect 35065 19818 35131 19821
rect 31756 19816 35131 19818
rect 31756 19760 35070 19816
rect 35126 19760 35131 19816
rect 31756 19758 35131 19760
rect 27429 19682 27495 19685
rect 30230 19682 30236 19684
rect 27429 19680 30236 19682
rect 27429 19624 27434 19680
rect 27490 19624 30236 19680
rect 27429 19622 30236 19624
rect 27429 19619 27495 19622
rect 30230 19620 30236 19622
rect 30300 19620 30306 19684
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 25957 19546 26023 19549
rect 28993 19546 29059 19549
rect 29126 19546 29132 19548
rect 25957 19544 29132 19546
rect 25957 19488 25962 19544
rect 26018 19488 28998 19544
rect 29054 19488 29132 19544
rect 25957 19486 29132 19488
rect 25957 19483 26023 19486
rect 28993 19483 29059 19486
rect 29126 19484 29132 19486
rect 29196 19546 29202 19548
rect 31756 19546 31816 19758
rect 35065 19755 35131 19758
rect 32213 19682 32279 19685
rect 32622 19682 32628 19684
rect 32213 19680 32628 19682
rect 32213 19624 32218 19680
rect 32274 19624 32628 19680
rect 32213 19622 32628 19624
rect 32213 19619 32279 19622
rect 32622 19620 32628 19622
rect 32692 19620 32698 19684
rect 32765 19682 32831 19685
rect 33910 19682 33916 19684
rect 32765 19680 33916 19682
rect 32765 19624 32770 19680
rect 32826 19624 33916 19680
rect 32765 19622 33916 19624
rect 32765 19619 32831 19622
rect 33910 19620 33916 19622
rect 33980 19682 33986 19684
rect 36721 19682 36787 19685
rect 33980 19680 36787 19682
rect 33980 19624 36726 19680
rect 36782 19624 36787 19680
rect 33980 19622 36787 19624
rect 33980 19620 33986 19622
rect 36721 19619 36787 19622
rect 29196 19486 31816 19546
rect 31937 19546 32003 19549
rect 32806 19546 32812 19548
rect 31937 19544 32812 19546
rect 31937 19488 31942 19544
rect 31998 19488 32812 19544
rect 31937 19486 32812 19488
rect 29196 19484 29202 19486
rect 31937 19483 32003 19486
rect 32806 19484 32812 19486
rect 32876 19484 32882 19548
rect 33225 19546 33291 19549
rect 33869 19546 33935 19549
rect 34605 19546 34671 19549
rect 33225 19544 33935 19546
rect 33225 19488 33230 19544
rect 33286 19488 33874 19544
rect 33930 19488 33935 19544
rect 33225 19486 33935 19488
rect 33225 19483 33291 19486
rect 33869 19483 33935 19486
rect 34286 19544 34671 19546
rect 34286 19488 34610 19544
rect 34666 19488 34671 19544
rect 34286 19486 34671 19488
rect 23749 19410 23815 19413
rect 24945 19410 25011 19413
rect 31753 19410 31819 19413
rect 23749 19408 25011 19410
rect 23749 19352 23754 19408
rect 23810 19352 24950 19408
rect 25006 19352 25011 19408
rect 23749 19350 25011 19352
rect 23749 19347 23815 19350
rect 24945 19347 25011 19350
rect 26190 19408 31819 19410
rect 26190 19352 31758 19408
rect 31814 19352 31819 19408
rect 26190 19350 31819 19352
rect 22461 19274 22527 19277
rect 22461 19272 23306 19274
rect 22461 19216 22466 19272
rect 22522 19216 23306 19272
rect 22461 19214 23306 19216
rect 22461 19211 22527 19214
rect 8385 19138 8451 19141
rect 22686 19138 22692 19140
rect 8385 19136 22692 19138
rect 8385 19080 8390 19136
rect 8446 19080 22692 19136
rect 8385 19078 22692 19080
rect 8385 19075 8451 19078
rect 22686 19076 22692 19078
rect 22756 19076 22762 19140
rect 23246 19138 23306 19214
rect 23422 19212 23428 19276
rect 23492 19274 23498 19276
rect 26190 19274 26250 19350
rect 31753 19347 31819 19350
rect 32489 19410 32555 19413
rect 34286 19410 34346 19486
rect 34605 19483 34671 19486
rect 32489 19408 34346 19410
rect 32489 19352 32494 19408
rect 32550 19352 34346 19408
rect 32489 19350 34346 19352
rect 34973 19410 35039 19413
rect 35249 19410 35315 19413
rect 35801 19412 35867 19413
rect 34973 19408 35315 19410
rect 34973 19352 34978 19408
rect 35034 19352 35254 19408
rect 35310 19352 35315 19408
rect 34973 19350 35315 19352
rect 32489 19347 32555 19350
rect 34973 19347 35039 19350
rect 35249 19347 35315 19350
rect 35750 19348 35756 19412
rect 35820 19410 35867 19412
rect 35820 19408 35912 19410
rect 35862 19352 35912 19408
rect 35820 19350 35912 19352
rect 35820 19348 35867 19350
rect 35801 19347 35867 19348
rect 23492 19214 26250 19274
rect 23492 19212 23498 19214
rect 26366 19212 26372 19276
rect 26436 19274 26442 19276
rect 26509 19274 26575 19277
rect 26436 19272 26575 19274
rect 26436 19216 26514 19272
rect 26570 19216 26575 19272
rect 26436 19214 26575 19216
rect 26436 19212 26442 19214
rect 26509 19211 26575 19214
rect 31201 19274 31267 19277
rect 38837 19274 38903 19277
rect 39200 19274 40000 19304
rect 31201 19272 35450 19274
rect 31201 19216 31206 19272
rect 31262 19216 35450 19272
rect 31201 19214 35450 19216
rect 31201 19211 31267 19214
rect 24025 19138 24091 19141
rect 23246 19136 24091 19138
rect 23246 19080 24030 19136
rect 24086 19080 24091 19136
rect 23246 19078 24091 19080
rect 24025 19075 24091 19078
rect 24577 19138 24643 19141
rect 25681 19138 25747 19141
rect 24577 19136 25747 19138
rect 24577 19080 24582 19136
rect 24638 19080 25686 19136
rect 25742 19080 25747 19136
rect 24577 19078 25747 19080
rect 24577 19075 24643 19078
rect 25681 19075 25747 19078
rect 25865 19138 25931 19141
rect 26877 19138 26943 19141
rect 25865 19136 26943 19138
rect 25865 19080 25870 19136
rect 25926 19080 26882 19136
rect 26938 19080 26943 19136
rect 25865 19078 26943 19080
rect 25865 19075 25931 19078
rect 26877 19075 26943 19078
rect 30281 19138 30347 19141
rect 33041 19138 33107 19141
rect 30281 19136 33107 19138
rect 30281 19080 30286 19136
rect 30342 19080 33046 19136
rect 33102 19080 33107 19136
rect 30281 19078 33107 19080
rect 35390 19138 35450 19214
rect 38837 19272 40000 19274
rect 38837 19216 38842 19272
rect 38898 19216 40000 19272
rect 38837 19214 40000 19216
rect 38837 19211 38903 19214
rect 39200 19184 40000 19214
rect 39021 19138 39087 19141
rect 35390 19136 39087 19138
rect 35390 19080 39026 19136
rect 39082 19080 39087 19136
rect 35390 19078 39087 19080
rect 30281 19075 30347 19078
rect 33041 19075 33107 19078
rect 39021 19075 39087 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 8886 18940 8892 19004
rect 8956 19002 8962 19004
rect 27429 19002 27495 19005
rect 8956 19000 27495 19002
rect 8956 18944 27434 19000
rect 27490 18944 27495 19000
rect 8956 18942 27495 18944
rect 8956 18940 8962 18942
rect 27429 18939 27495 18942
rect 29913 19002 29979 19005
rect 30465 19002 30531 19005
rect 29913 19000 30531 19002
rect 29913 18944 29918 19000
rect 29974 18944 30470 19000
rect 30526 18944 30531 19000
rect 29913 18942 30531 18944
rect 29913 18939 29979 18942
rect 30465 18939 30531 18942
rect 24117 18866 24183 18869
rect 28625 18866 28691 18869
rect 24117 18864 28691 18866
rect 24117 18808 24122 18864
rect 24178 18808 28630 18864
rect 28686 18808 28691 18864
rect 24117 18806 28691 18808
rect 24117 18803 24183 18806
rect 28625 18803 28691 18806
rect 29361 18866 29427 18869
rect 30925 18866 30991 18869
rect 31569 18866 31635 18869
rect 37365 18866 37431 18869
rect 29361 18864 31635 18866
rect 29361 18808 29366 18864
rect 29422 18808 30930 18864
rect 30986 18808 31574 18864
rect 31630 18808 31635 18864
rect 29361 18806 31635 18808
rect 29361 18803 29427 18806
rect 30925 18803 30991 18806
rect 31569 18803 31635 18806
rect 32446 18864 37431 18866
rect 32446 18808 37370 18864
rect 37426 18808 37431 18864
rect 32446 18806 37431 18808
rect 26233 18730 26299 18733
rect 27337 18730 27403 18733
rect 26233 18728 27403 18730
rect 26233 18672 26238 18728
rect 26294 18672 27342 18728
rect 27398 18672 27403 18728
rect 26233 18670 27403 18672
rect 26233 18667 26299 18670
rect 27337 18667 27403 18670
rect 28165 18730 28231 18733
rect 32446 18730 32506 18806
rect 37365 18803 37431 18806
rect 28165 18728 32506 18730
rect 28165 18672 28170 18728
rect 28226 18672 32506 18728
rect 28165 18670 32506 18672
rect 32581 18730 32647 18733
rect 35617 18730 35683 18733
rect 32581 18728 35683 18730
rect 32581 18672 32586 18728
rect 32642 18672 35622 18728
rect 35678 18672 35683 18728
rect 32581 18670 35683 18672
rect 28165 18667 28231 18670
rect 32581 18667 32647 18670
rect 35617 18667 35683 18670
rect 30005 18594 30071 18597
rect 30557 18594 30623 18597
rect 30005 18592 30623 18594
rect 30005 18536 30010 18592
rect 30066 18536 30562 18592
rect 30618 18536 30623 18592
rect 30005 18534 30623 18536
rect 30005 18531 30071 18534
rect 30557 18531 30623 18534
rect 32581 18594 32647 18597
rect 35801 18594 35867 18597
rect 32581 18592 35867 18594
rect 32581 18536 32586 18592
rect 32642 18536 35806 18592
rect 35862 18536 35867 18592
rect 32581 18534 35867 18536
rect 32581 18531 32647 18534
rect 35801 18531 35867 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 25681 18458 25747 18461
rect 26049 18458 26115 18461
rect 32673 18458 32739 18461
rect 25681 18456 32739 18458
rect 25681 18400 25686 18456
rect 25742 18400 26054 18456
rect 26110 18400 32678 18456
rect 32734 18400 32739 18456
rect 25681 18398 32739 18400
rect 25681 18395 25747 18398
rect 26049 18395 26115 18398
rect 32673 18395 32739 18398
rect 19793 18322 19859 18325
rect 24301 18322 24367 18325
rect 26417 18322 26483 18325
rect 19793 18320 26483 18322
rect 19793 18264 19798 18320
rect 19854 18264 24306 18320
rect 24362 18264 26422 18320
rect 26478 18264 26483 18320
rect 19793 18262 26483 18264
rect 19793 18259 19859 18262
rect 24301 18259 24367 18262
rect 26417 18259 26483 18262
rect 28349 18322 28415 18325
rect 32213 18322 32279 18325
rect 28349 18320 32279 18322
rect 28349 18264 28354 18320
rect 28410 18264 32218 18320
rect 32274 18264 32279 18320
rect 28349 18262 32279 18264
rect 28349 18259 28415 18262
rect 32213 18259 32279 18262
rect 20897 18186 20963 18189
rect 26233 18186 26299 18189
rect 20897 18184 26299 18186
rect 20897 18128 20902 18184
rect 20958 18128 26238 18184
rect 26294 18128 26299 18184
rect 20897 18126 26299 18128
rect 20897 18123 20963 18126
rect 26233 18123 26299 18126
rect 26509 18186 26575 18189
rect 28533 18186 28599 18189
rect 29085 18186 29151 18189
rect 26509 18184 29151 18186
rect 26509 18128 26514 18184
rect 26570 18128 28538 18184
rect 28594 18128 29090 18184
rect 29146 18128 29151 18184
rect 26509 18126 29151 18128
rect 26509 18123 26575 18126
rect 28533 18123 28599 18126
rect 29085 18123 29151 18126
rect 30966 18124 30972 18188
rect 31036 18186 31042 18188
rect 33133 18186 33199 18189
rect 31036 18184 33199 18186
rect 31036 18128 33138 18184
rect 33194 18128 33199 18184
rect 31036 18126 33199 18128
rect 31036 18124 31042 18126
rect 33133 18123 33199 18126
rect 34145 18186 34211 18189
rect 35249 18186 35315 18189
rect 34145 18184 35315 18186
rect 34145 18128 34150 18184
rect 34206 18128 35254 18184
rect 35310 18128 35315 18184
rect 34145 18126 35315 18128
rect 34145 18123 34211 18126
rect 35249 18123 35315 18126
rect 30005 18052 30071 18053
rect 30005 18048 30052 18052
rect 30116 18050 30122 18052
rect 33133 18050 33199 18053
rect 33317 18050 33383 18053
rect 30005 17992 30010 18048
rect 30005 17988 30052 17992
rect 30116 17990 30162 18050
rect 33133 18048 33383 18050
rect 33133 17992 33138 18048
rect 33194 17992 33322 18048
rect 33378 17992 33383 18048
rect 33133 17990 33383 17992
rect 30116 17988 30122 17990
rect 30005 17987 30071 17988
rect 33133 17987 33199 17990
rect 33317 17987 33383 17990
rect 33501 18050 33567 18053
rect 33869 18050 33935 18053
rect 33501 18048 33935 18050
rect 33501 17992 33506 18048
rect 33562 17992 33874 18048
rect 33930 17992 33935 18048
rect 33501 17990 33935 17992
rect 33501 17987 33567 17990
rect 33869 17987 33935 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 30649 17914 30715 17917
rect 31702 17914 31708 17916
rect 30649 17912 31708 17914
rect 30649 17856 30654 17912
rect 30710 17856 31708 17912
rect 30649 17854 31708 17856
rect 30649 17851 30715 17854
rect 31702 17852 31708 17854
rect 31772 17852 31778 17916
rect 39021 17914 39087 17917
rect 39200 17914 40000 17944
rect 39021 17912 40000 17914
rect 39021 17856 39026 17912
rect 39082 17856 40000 17912
rect 39021 17854 40000 17856
rect 39021 17851 39087 17854
rect 39200 17824 40000 17854
rect 27981 17778 28047 17781
rect 33409 17778 33475 17781
rect 27981 17776 33475 17778
rect 27981 17720 27986 17776
rect 28042 17720 33414 17776
rect 33470 17720 33475 17776
rect 27981 17718 33475 17720
rect 27981 17715 28047 17718
rect 33409 17715 33475 17718
rect 33685 17778 33751 17781
rect 37825 17778 37891 17781
rect 33685 17776 37891 17778
rect 33685 17720 33690 17776
rect 33746 17720 37830 17776
rect 37886 17720 37891 17776
rect 33685 17718 37891 17720
rect 33685 17715 33751 17718
rect 37825 17715 37891 17718
rect 23105 17642 23171 17645
rect 24761 17642 24827 17645
rect 23105 17640 24827 17642
rect 23105 17584 23110 17640
rect 23166 17584 24766 17640
rect 24822 17584 24827 17640
rect 23105 17582 24827 17584
rect 23105 17579 23171 17582
rect 24761 17579 24827 17582
rect 25773 17642 25839 17645
rect 30557 17642 30623 17645
rect 25773 17640 30623 17642
rect 25773 17584 25778 17640
rect 25834 17584 30562 17640
rect 30618 17584 30623 17640
rect 25773 17582 30623 17584
rect 25773 17579 25839 17582
rect 30557 17579 30623 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 23197 17370 23263 17373
rect 28349 17370 28415 17373
rect 23197 17368 28415 17370
rect 23197 17312 23202 17368
rect 23258 17312 28354 17368
rect 28410 17312 28415 17368
rect 23197 17310 28415 17312
rect 23197 17307 23263 17310
rect 28349 17307 28415 17310
rect 30741 17370 30807 17373
rect 33685 17370 33751 17373
rect 30741 17368 33751 17370
rect 30741 17312 30746 17368
rect 30802 17312 33690 17368
rect 33746 17312 33751 17368
rect 30741 17310 33751 17312
rect 30741 17307 30807 17310
rect 33685 17307 33751 17310
rect 22185 17234 22251 17237
rect 28257 17234 28323 17237
rect 22185 17232 28323 17234
rect 22185 17176 22190 17232
rect 22246 17176 28262 17232
rect 28318 17176 28323 17232
rect 22185 17174 28323 17176
rect 22185 17171 22251 17174
rect 28257 17171 28323 17174
rect 3877 17098 3943 17101
rect 39297 17098 39363 17101
rect 3877 17096 39363 17098
rect 3877 17040 3882 17096
rect 3938 17040 39302 17096
rect 39358 17040 39363 17096
rect 3877 17038 39363 17040
rect 3877 17035 3943 17038
rect 39297 17035 39363 17038
rect 28574 16900 28580 16964
rect 28644 16962 28650 16964
rect 34605 16962 34671 16965
rect 28644 16960 34671 16962
rect 28644 16904 34610 16960
rect 34666 16904 34671 16960
rect 28644 16902 34671 16904
rect 28644 16900 28650 16902
rect 34605 16899 34671 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 24853 16826 24919 16829
rect 35801 16826 35867 16829
rect 36302 16826 36308 16828
rect 24853 16824 29010 16826
rect 24853 16768 24858 16824
rect 24914 16768 29010 16824
rect 24853 16766 29010 16768
rect 24853 16763 24919 16766
rect 28950 16693 29010 16766
rect 35801 16824 36308 16826
rect 35801 16768 35806 16824
rect 35862 16768 36308 16824
rect 35801 16766 36308 16768
rect 35801 16763 35867 16766
rect 36302 16764 36308 16766
rect 36372 16764 36378 16828
rect 25773 16690 25839 16693
rect 26141 16690 26207 16693
rect 25773 16688 26207 16690
rect 25773 16632 25778 16688
rect 25834 16632 26146 16688
rect 26202 16632 26207 16688
rect 25773 16630 26207 16632
rect 28950 16688 29059 16693
rect 28950 16632 28998 16688
rect 29054 16632 29059 16688
rect 28950 16630 29059 16632
rect 25773 16627 25839 16630
rect 26141 16627 26207 16630
rect 28993 16627 29059 16630
rect 29177 16690 29243 16693
rect 30097 16690 30163 16693
rect 29177 16688 30163 16690
rect 29177 16632 29182 16688
rect 29238 16632 30102 16688
rect 30158 16632 30163 16688
rect 29177 16630 30163 16632
rect 29177 16627 29243 16630
rect 30097 16627 30163 16630
rect 36261 16690 36327 16693
rect 36486 16690 36492 16692
rect 36261 16688 36492 16690
rect 36261 16632 36266 16688
rect 36322 16632 36492 16688
rect 36261 16630 36492 16632
rect 36261 16627 36327 16630
rect 36486 16628 36492 16630
rect 36556 16628 36562 16692
rect 24342 16492 24348 16556
rect 24412 16554 24418 16556
rect 24577 16554 24643 16557
rect 24412 16552 24643 16554
rect 24412 16496 24582 16552
rect 24638 16496 24643 16552
rect 24412 16494 24643 16496
rect 24412 16492 24418 16494
rect 24577 16491 24643 16494
rect 30281 16554 30347 16557
rect 30966 16554 30972 16556
rect 30281 16552 30972 16554
rect 30281 16496 30286 16552
rect 30342 16496 30972 16552
rect 30281 16494 30972 16496
rect 30281 16491 30347 16494
rect 30966 16492 30972 16494
rect 31036 16492 31042 16556
rect 39021 16554 39087 16557
rect 39200 16554 40000 16584
rect 39021 16552 40000 16554
rect 39021 16496 39026 16552
rect 39082 16496 40000 16552
rect 39021 16494 40000 16496
rect 39021 16491 39087 16494
rect 39200 16464 40000 16494
rect 30189 16418 30255 16421
rect 37365 16418 37431 16421
rect 30189 16416 37431 16418
rect 30189 16360 30194 16416
rect 30250 16360 37370 16416
rect 37426 16360 37431 16416
rect 30189 16358 37431 16360
rect 30189 16355 30255 16358
rect 37365 16355 37431 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 28809 16282 28875 16285
rect 30097 16282 30163 16285
rect 30741 16282 30807 16285
rect 28809 16280 30807 16282
rect 28809 16224 28814 16280
rect 28870 16224 30102 16280
rect 30158 16224 30746 16280
rect 30802 16224 30807 16280
rect 28809 16222 30807 16224
rect 28809 16219 28875 16222
rect 30097 16219 30163 16222
rect 30741 16219 30807 16222
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 14733 15602 14799 15605
rect 38745 15602 38811 15605
rect 14733 15600 38811 15602
rect 14733 15544 14738 15600
rect 14794 15544 38750 15600
rect 38806 15544 38811 15600
rect 14733 15542 38811 15544
rect 14733 15539 14799 15542
rect 38745 15539 38811 15542
rect 35525 15468 35591 15469
rect 35525 15466 35572 15468
rect 35480 15464 35572 15466
rect 35480 15408 35530 15464
rect 35480 15406 35572 15408
rect 35525 15404 35572 15406
rect 35636 15404 35642 15468
rect 35525 15403 35591 15404
rect 30782 15268 30788 15332
rect 30852 15330 30858 15332
rect 36813 15330 36879 15333
rect 30852 15328 36879 15330
rect 30852 15272 36818 15328
rect 36874 15272 36879 15328
rect 30852 15270 36879 15272
rect 30852 15268 30858 15270
rect 36813 15267 36879 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 38101 15194 38167 15197
rect 39200 15194 40000 15224
rect 38101 15192 40000 15194
rect 38101 15136 38106 15192
rect 38162 15136 40000 15192
rect 38101 15134 40000 15136
rect 38101 15131 38167 15134
rect 39200 15104 40000 15134
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 25078 14316 25084 14380
rect 25148 14378 25154 14380
rect 37549 14378 37615 14381
rect 25148 14376 37615 14378
rect 25148 14320 37554 14376
rect 37610 14320 37615 14376
rect 25148 14318 37615 14320
rect 25148 14316 25154 14318
rect 37549 14315 37615 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 39021 13834 39087 13837
rect 39200 13834 40000 13864
rect 39021 13832 40000 13834
rect 39021 13776 39026 13832
rect 39082 13776 40000 13832
rect 39021 13774 40000 13776
rect 39021 13771 39087 13774
rect 39200 13744 40000 13774
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 34278 13364 34284 13428
rect 34348 13426 34354 13428
rect 36077 13426 36143 13429
rect 34348 13424 36143 13426
rect 34348 13368 36082 13424
rect 36138 13368 36143 13424
rect 34348 13366 36143 13368
rect 34348 13364 34354 13366
rect 36077 13363 36143 13366
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 38285 12474 38351 12477
rect 39200 12474 40000 12504
rect 38285 12472 40000 12474
rect 38285 12416 38290 12472
rect 38346 12416 40000 12472
rect 38285 12414 40000 12416
rect 38285 12411 38351 12414
rect 39200 12384 40000 12414
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 38101 11114 38167 11117
rect 39200 11114 40000 11144
rect 38101 11112 40000 11114
rect 38101 11056 38106 11112
rect 38162 11056 40000 11112
rect 38101 11054 40000 11056
rect 38101 11051 38167 11054
rect 39200 11024 40000 11054
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 38101 9754 38167 9757
rect 39200 9754 40000 9784
rect 38101 9752 40000 9754
rect 38101 9696 38106 9752
rect 38162 9696 40000 9752
rect 38101 9694 40000 9696
rect 38101 9691 38167 9694
rect 39200 9664 40000 9694
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 30046 8468 30052 8532
rect 30116 8530 30122 8532
rect 37825 8530 37891 8533
rect 30116 8528 37891 8530
rect 30116 8472 37830 8528
rect 37886 8472 37891 8528
rect 30116 8470 37891 8472
rect 30116 8468 30122 8470
rect 37825 8467 37891 8470
rect 38101 8394 38167 8397
rect 39200 8394 40000 8424
rect 38101 8392 40000 8394
rect 38101 8336 38106 8392
rect 38162 8336 40000 8392
rect 38101 8334 40000 8336
rect 38101 8331 38167 8334
rect 39200 8304 40000 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 38101 7034 38167 7037
rect 39200 7034 40000 7064
rect 38101 7032 40000 7034
rect 38101 6976 38106 7032
rect 38162 6976 40000 7032
rect 38101 6974 40000 6976
rect 38101 6971 38167 6974
rect 39200 6944 40000 6974
rect 32990 6836 32996 6900
rect 33060 6898 33066 6900
rect 37825 6898 37891 6901
rect 33060 6896 37891 6898
rect 33060 6840 37830 6896
rect 37886 6840 37891 6896
rect 33060 6838 37891 6840
rect 33060 6836 33066 6838
rect 37825 6835 37891 6838
rect 32438 6700 32444 6764
rect 32508 6762 32514 6764
rect 37365 6762 37431 6765
rect 32508 6760 37431 6762
rect 32508 6704 37370 6760
rect 37426 6704 37431 6760
rect 32508 6702 37431 6704
rect 32508 6700 32514 6702
rect 37365 6699 37431 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 38101 5674 38167 5677
rect 39200 5674 40000 5704
rect 38101 5672 40000 5674
rect 38101 5616 38106 5672
rect 38162 5616 40000 5672
rect 38101 5614 40000 5616
rect 38101 5611 38167 5614
rect 39200 5584 40000 5614
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 38101 4314 38167 4317
rect 39200 4314 40000 4344
rect 38101 4312 40000 4314
rect 38101 4256 38106 4312
rect 38162 4256 40000 4312
rect 38101 4254 40000 4256
rect 38101 4251 38167 4254
rect 39200 4224 40000 4254
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 38101 2954 38167 2957
rect 39200 2954 40000 2984
rect 38101 2952 40000 2954
rect 38101 2896 38106 2952
rect 38162 2896 40000 2952
rect 38101 2894 40000 2896
rect 38101 2891 38167 2894
rect 39200 2864 40000 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 32806 2484 32812 2548
rect 32876 2546 32882 2548
rect 37825 2546 37891 2549
rect 32876 2544 37891 2546
rect 32876 2488 37830 2544
rect 37886 2488 37891 2544
rect 32876 2486 37891 2488
rect 32876 2484 32882 2486
rect 37825 2483 37891 2486
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 38101 1594 38167 1597
rect 39200 1594 40000 1624
rect 38101 1592 40000 1594
rect 38101 1536 38106 1592
rect 38162 1536 40000 1592
rect 38101 1534 40000 1536
rect 38101 1531 38167 1534
rect 39200 1504 40000 1534
<< via3 >>
rect 22140 39340 22204 39404
rect 27476 39204 27540 39268
rect 27292 39068 27356 39132
rect 12572 38932 12636 38996
rect 27844 38252 27908 38316
rect 9628 37980 9692 38044
rect 16436 37768 16500 37772
rect 16436 37712 16486 37768
rect 16486 37712 16500 37768
rect 16436 37708 16500 37712
rect 29316 37708 29380 37772
rect 23428 37572 23492 37636
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4844 37300 4908 37364
rect 23612 37436 23676 37500
rect 26924 37300 26988 37364
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 15332 36892 15396 36956
rect 21956 36620 22020 36684
rect 7236 36484 7300 36548
rect 19380 36484 19444 36548
rect 24900 36484 24964 36548
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 18276 36348 18340 36412
rect 20116 36408 20180 36412
rect 20116 36352 20166 36408
rect 20166 36352 20180 36408
rect 20116 36348 20180 36352
rect 17724 36212 17788 36276
rect 25268 36212 25332 36276
rect 17356 36136 17420 36140
rect 17356 36080 17370 36136
rect 17370 36080 17420 36136
rect 17356 36076 17420 36080
rect 6132 36000 6196 36004
rect 6132 35944 6146 36000
rect 6146 35944 6196 36000
rect 6132 35940 6196 35944
rect 12756 35940 12820 36004
rect 26188 36076 26252 36140
rect 33180 35940 33244 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 10364 35804 10428 35868
rect 18092 35804 18156 35868
rect 21036 35804 21100 35868
rect 27476 35804 27540 35868
rect 23980 35668 24044 35732
rect 34100 35592 34164 35596
rect 34100 35536 34150 35592
rect 34150 35536 34164 35592
rect 34100 35532 34164 35536
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 18276 35260 18340 35324
rect 29500 35260 29564 35324
rect 30420 35124 30484 35188
rect 19196 34988 19260 35052
rect 4844 34776 4908 34780
rect 4844 34720 4858 34776
rect 4858 34720 4908 34776
rect 4844 34716 4908 34720
rect 5212 34716 5276 34780
rect 12204 34776 12268 34780
rect 12204 34720 12218 34776
rect 12218 34720 12268 34776
rect 12204 34716 12268 34720
rect 17908 34852 17972 34916
rect 24900 34988 24964 35052
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 8156 34640 8220 34644
rect 8156 34584 8206 34640
rect 8206 34584 8220 34640
rect 8156 34580 8220 34584
rect 11100 34580 11164 34644
rect 11284 34580 11348 34644
rect 27844 34776 27908 34780
rect 27844 34720 27894 34776
rect 27894 34720 27908 34776
rect 27844 34716 27908 34720
rect 36124 34852 36188 34916
rect 23244 34580 23308 34644
rect 29684 34580 29748 34644
rect 37044 34580 37108 34644
rect 23428 34308 23492 34372
rect 30788 34308 30852 34372
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 9628 34172 9692 34236
rect 26188 34232 26252 34236
rect 26188 34176 26238 34232
rect 26238 34176 26252 34232
rect 26188 34172 26252 34176
rect 33732 34172 33796 34236
rect 34284 34172 34348 34236
rect 35572 34172 35636 34236
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 31340 33628 31404 33692
rect 35940 33628 36004 33692
rect 23980 33356 24044 33420
rect 6316 33220 6380 33284
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 20852 33280 20916 33284
rect 20852 33224 20866 33280
rect 20866 33224 20916 33280
rect 20852 33220 20916 33224
rect 26372 33280 26436 33284
rect 27292 33552 27356 33556
rect 27292 33496 27342 33552
rect 27342 33496 27356 33552
rect 27292 33492 27356 33496
rect 33916 33492 33980 33556
rect 27476 33356 27540 33420
rect 26372 33224 26386 33280
rect 26386 33224 26436 33280
rect 26372 33220 26436 33224
rect 28212 33220 28276 33284
rect 28948 33220 29012 33284
rect 33180 33220 33244 33284
rect 33548 33220 33612 33284
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 25268 32948 25332 33012
rect 28580 33008 28644 33012
rect 28580 32952 28630 33008
rect 28630 32952 28644 33008
rect 28580 32948 28644 32952
rect 29132 32948 29196 33012
rect 28028 32676 28092 32740
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 11284 32540 11348 32604
rect 12388 32600 12452 32604
rect 12388 32544 12402 32600
rect 12402 32544 12452 32600
rect 12388 32540 12452 32544
rect 28396 32540 28460 32604
rect 31892 32404 31956 32468
rect 4844 32268 4908 32332
rect 13492 32132 13556 32196
rect 13676 32132 13740 32196
rect 20668 32132 20732 32196
rect 34652 32268 34716 32332
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 29684 32132 29748 32196
rect 33364 32132 33428 32196
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 24716 31996 24780 32060
rect 28212 31996 28276 32060
rect 29500 32056 29564 32060
rect 29500 32000 29514 32056
rect 29514 32000 29564 32056
rect 29500 31996 29564 32000
rect 13308 31860 13372 31924
rect 21036 31860 21100 31924
rect 23980 31860 24044 31924
rect 4844 31512 4908 31516
rect 4844 31456 4894 31512
rect 4894 31456 4908 31512
rect 4844 31452 4908 31456
rect 12572 31588 12636 31652
rect 13492 31588 13556 31652
rect 9444 31512 9508 31516
rect 9444 31456 9458 31512
rect 9458 31456 9508 31512
rect 9444 31452 9508 31456
rect 12204 31316 12268 31380
rect 15148 31044 15212 31108
rect 18276 31724 18340 31788
rect 25084 31724 25148 31788
rect 26556 31724 26620 31788
rect 28396 31724 28460 31788
rect 29316 31724 29380 31788
rect 20116 31588 20180 31652
rect 27292 31588 27356 31652
rect 35388 31996 35452 32060
rect 34468 31784 34532 31788
rect 34468 31728 34518 31784
rect 34518 31728 34532 31784
rect 34468 31724 34532 31728
rect 33548 31588 33612 31652
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 20484 31452 20548 31516
rect 25452 31316 25516 31380
rect 30052 31316 30116 31380
rect 34652 31316 34716 31380
rect 35388 31316 35452 31380
rect 16252 31180 16316 31244
rect 34468 31180 34532 31244
rect 32996 31044 33060 31108
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 28396 30908 28460 30972
rect 35756 31240 35820 31244
rect 35756 31184 35770 31240
rect 35770 31184 35820 31240
rect 35756 31180 35820 31184
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 9628 30636 9692 30700
rect 30420 30636 30484 30700
rect 30604 30636 30668 30700
rect 35388 30636 35452 30700
rect 37044 30636 37108 30700
rect 7236 30364 7300 30428
rect 8892 30364 8956 30428
rect 15332 30500 15396 30564
rect 23612 30500 23676 30564
rect 28948 30500 29012 30564
rect 34652 30500 34716 30564
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 26004 30424 26068 30428
rect 26004 30368 26054 30424
rect 26054 30368 26068 30424
rect 26004 30364 26068 30368
rect 24532 30228 24596 30292
rect 28580 30228 28644 30292
rect 25452 30092 25516 30156
rect 25636 30152 25700 30156
rect 33180 30228 33244 30292
rect 33916 30228 33980 30292
rect 35388 30364 35452 30428
rect 35940 30364 36004 30428
rect 25636 30096 25650 30152
rect 25650 30096 25700 30152
rect 25636 30092 25700 30096
rect 33364 30092 33428 30156
rect 33548 30092 33612 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 31156 29956 31220 30020
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 32444 29820 32508 29884
rect 19012 29684 19076 29748
rect 26924 29684 26988 29748
rect 28948 29684 29012 29748
rect 34468 29684 34532 29748
rect 12388 29608 12452 29612
rect 12388 29552 12438 29608
rect 12438 29552 12452 29608
rect 12388 29548 12452 29552
rect 13308 29548 13372 29612
rect 22140 29548 22204 29612
rect 9444 29472 9508 29476
rect 9444 29416 9458 29472
rect 9458 29416 9508 29472
rect 9444 29412 9508 29416
rect 12756 29412 12820 29476
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 11100 29276 11164 29340
rect 19380 29276 19444 29340
rect 17724 29140 17788 29204
rect 28764 29412 28828 29476
rect 34284 29412 34348 29476
rect 33364 29276 33428 29340
rect 36308 29276 36372 29340
rect 32076 29200 32140 29204
rect 32076 29144 32126 29200
rect 32126 29144 32140 29200
rect 32076 29140 32140 29144
rect 32260 29140 32324 29204
rect 33732 29140 33796 29204
rect 34468 29140 34532 29204
rect 22508 29004 22572 29068
rect 24900 29004 24964 29068
rect 25636 29004 25700 29068
rect 29316 29004 29380 29068
rect 33364 29004 33428 29068
rect 19196 28868 19260 28932
rect 23796 28868 23860 28932
rect 28028 28868 28092 28932
rect 30788 28868 30852 28932
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 18276 28596 18340 28660
rect 30604 28732 30668 28796
rect 30788 28732 30852 28796
rect 31524 28596 31588 28660
rect 18276 28460 18340 28524
rect 34100 28596 34164 28660
rect 35756 28656 35820 28660
rect 35756 28600 35770 28656
rect 35770 28600 35820 28656
rect 35756 28596 35820 28600
rect 23244 28324 23308 28388
rect 26188 28324 26252 28388
rect 35756 28324 35820 28388
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 13676 28188 13740 28252
rect 26556 28188 26620 28252
rect 27476 28052 27540 28116
rect 28212 28052 28276 28116
rect 35940 28188 36004 28252
rect 31708 28112 31772 28116
rect 31708 28056 31722 28112
rect 31722 28056 31772 28112
rect 31708 28052 31772 28056
rect 24716 27916 24780 27980
rect 15148 27840 15212 27844
rect 15148 27784 15162 27840
rect 15162 27784 15212 27840
rect 15148 27780 15212 27784
rect 19380 27840 19444 27844
rect 19380 27784 19430 27840
rect 19430 27784 19444 27840
rect 19380 27780 19444 27784
rect 29684 27916 29748 27980
rect 30420 27976 30484 27980
rect 30420 27920 30434 27976
rect 30434 27920 30484 27976
rect 30420 27916 30484 27920
rect 30972 27916 31036 27980
rect 34468 27976 34532 27980
rect 34468 27920 34482 27976
rect 34482 27920 34532 27976
rect 34468 27916 34532 27920
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 33916 27780 33980 27844
rect 34284 27780 34348 27844
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 22692 27704 22756 27708
rect 22692 27648 22706 27704
rect 22706 27648 22756 27704
rect 22692 27644 22756 27648
rect 13676 27508 13740 27572
rect 17908 27568 17972 27572
rect 17908 27512 17922 27568
rect 17922 27512 17972 27568
rect 17908 27508 17972 27512
rect 23428 27508 23492 27572
rect 26004 27568 26068 27572
rect 26004 27512 26054 27568
rect 26054 27512 26068 27568
rect 26004 27508 26068 27512
rect 27108 27568 27172 27572
rect 27108 27512 27122 27568
rect 27122 27512 27172 27568
rect 27108 27508 27172 27512
rect 27476 27568 27540 27572
rect 27476 27512 27526 27568
rect 27526 27512 27540 27568
rect 27476 27508 27540 27512
rect 31340 27508 31404 27572
rect 34100 27508 34164 27572
rect 34284 27508 34348 27572
rect 17356 27236 17420 27300
rect 31524 27372 31588 27436
rect 20300 27236 20364 27300
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 18276 27100 18340 27164
rect 23612 27236 23676 27300
rect 24532 27100 24596 27164
rect 25820 27100 25884 27164
rect 13492 27024 13556 27028
rect 13492 26968 13506 27024
rect 13506 26968 13556 27024
rect 13492 26964 13556 26968
rect 29500 26964 29564 27028
rect 36308 27160 36372 27164
rect 36308 27104 36358 27160
rect 36358 27104 36372 27160
rect 36308 27100 36372 27104
rect 31156 26964 31220 27028
rect 32996 26964 33060 27028
rect 34652 26964 34716 27028
rect 20668 26828 20732 26892
rect 32076 26828 32140 26892
rect 15332 26692 15396 26756
rect 18092 26752 18156 26756
rect 18092 26696 18106 26752
rect 18106 26696 18156 26752
rect 18092 26692 18156 26696
rect 25268 26752 25332 26756
rect 25268 26696 25282 26752
rect 25282 26696 25332 26752
rect 25268 26692 25332 26696
rect 32996 26752 33060 26756
rect 32996 26696 33046 26752
rect 33046 26696 33060 26752
rect 32996 26692 33060 26696
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 8156 26556 8220 26620
rect 26372 26556 26436 26620
rect 27660 26556 27724 26620
rect 6316 26420 6380 26484
rect 20852 26420 20916 26484
rect 21036 26420 21100 26484
rect 30236 26420 30300 26484
rect 34652 26556 34716 26620
rect 16436 26284 16500 26348
rect 13308 26012 13372 26076
rect 19012 26148 19076 26212
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 24164 26284 24228 26348
rect 29132 26284 29196 26348
rect 30604 26284 30668 26348
rect 31892 26344 31956 26348
rect 31892 26288 31906 26344
rect 31906 26288 31956 26344
rect 31892 26284 31956 26288
rect 20484 26208 20548 26212
rect 20484 26152 20534 26208
rect 20534 26152 20548 26208
rect 20484 26148 20548 26152
rect 28764 26148 28828 26212
rect 20484 26012 20548 26076
rect 15148 25876 15212 25940
rect 34284 26012 34348 26076
rect 31524 25876 31588 25940
rect 26004 25800 26068 25804
rect 26004 25744 26018 25800
rect 26018 25744 26068 25800
rect 26004 25740 26068 25744
rect 26556 25740 26620 25804
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 6132 25468 6196 25532
rect 28212 25468 28276 25532
rect 29868 25468 29932 25532
rect 20300 25332 20364 25396
rect 20484 25332 20548 25396
rect 26556 25332 26620 25396
rect 33180 25332 33244 25396
rect 33732 25332 33796 25396
rect 25268 25196 25332 25260
rect 30972 25196 31036 25260
rect 19380 25120 19444 25124
rect 19380 25064 19430 25120
rect 19430 25064 19444 25120
rect 19380 25060 19444 25064
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 16252 24788 16316 24852
rect 28764 24924 28828 24988
rect 35756 24924 35820 24988
rect 23796 24788 23860 24852
rect 28948 24788 29012 24852
rect 30788 24788 30852 24852
rect 32444 24788 32508 24852
rect 32628 24788 32692 24852
rect 5212 24516 5276 24580
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 32812 24380 32876 24444
rect 33548 24440 33612 24444
rect 33548 24384 33562 24440
rect 33562 24384 33612 24440
rect 33548 24380 33612 24384
rect 29132 24244 29196 24308
rect 31708 24244 31772 24308
rect 32996 23972 33060 24036
rect 35756 23972 35820 24036
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 29500 23836 29564 23900
rect 30972 23700 31036 23764
rect 34652 23700 34716 23764
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 27660 23428 27724 23492
rect 28212 23428 28276 23492
rect 28580 23428 28644 23492
rect 33548 23428 33612 23492
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 26188 23156 26252 23220
rect 27108 23156 27172 23220
rect 34652 23156 34716 23220
rect 35940 23156 36004 23220
rect 10364 23020 10428 23084
rect 23428 22884 23492 22948
rect 33364 22884 33428 22948
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 27476 22748 27540 22812
rect 26372 22612 26436 22676
rect 30420 22612 30484 22676
rect 33916 22612 33980 22676
rect 21956 22476 22020 22540
rect 29868 22476 29932 22540
rect 32260 22476 32324 22540
rect 35388 22612 35452 22676
rect 33916 22400 33980 22404
rect 33916 22344 33930 22400
rect 33930 22344 33980 22400
rect 33916 22340 33980 22344
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 9628 22204 9692 22268
rect 21956 21932 22020 21996
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 25820 22068 25884 22132
rect 29684 22068 29748 22132
rect 24348 21932 24412 21996
rect 32076 22068 32140 22132
rect 34468 22068 34532 22132
rect 35572 21932 35636 21996
rect 27292 21796 27356 21860
rect 30972 21796 31036 21860
rect 31524 21796 31588 21860
rect 26004 21660 26068 21724
rect 24164 21524 24228 21588
rect 29316 21524 29380 21588
rect 37044 21524 37108 21588
rect 22508 21252 22572 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 33732 21116 33796 21180
rect 30052 20844 30116 20908
rect 32628 20708 32692 20772
rect 32996 20768 33060 20772
rect 32996 20712 33010 20768
rect 33010 20712 33060 20768
rect 32996 20708 33060 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 28396 20632 28460 20636
rect 28396 20576 28410 20632
rect 28410 20576 28460 20632
rect 28396 20572 28460 20576
rect 32444 20436 32508 20500
rect 32628 20436 32692 20500
rect 32812 20436 32876 20500
rect 34284 20436 34348 20500
rect 28764 20164 28828 20228
rect 30604 20164 30668 20228
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 26556 20028 26620 20092
rect 34284 20028 34348 20092
rect 30604 19756 30668 19820
rect 30236 19620 30300 19684
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 29132 19484 29196 19548
rect 32628 19620 32692 19684
rect 33916 19620 33980 19684
rect 32812 19484 32876 19548
rect 22692 19076 22756 19140
rect 23428 19212 23492 19276
rect 35756 19408 35820 19412
rect 35756 19352 35806 19408
rect 35806 19352 35820 19408
rect 35756 19348 35820 19352
rect 26372 19212 26436 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 8892 18940 8956 19004
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 30972 18124 31036 18188
rect 30052 18048 30116 18052
rect 30052 17992 30066 18048
rect 30066 17992 30116 18048
rect 30052 17988 30116 17992
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 31708 17852 31772 17916
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 28580 16900 28644 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 36308 16764 36372 16828
rect 36492 16628 36556 16692
rect 24348 16492 24412 16556
rect 30972 16492 31036 16556
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 35572 15464 35636 15468
rect 35572 15408 35586 15464
rect 35586 15408 35636 15464
rect 35572 15404 35636 15408
rect 30788 15268 30852 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 25084 14316 25148 14380
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 34284 13364 34348 13428
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 30052 8468 30116 8532
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 32996 6836 33060 6900
rect 32444 6700 32508 6764
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 32812 2484 32876 2548
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 22139 39404 22205 39405
rect 22139 39340 22140 39404
rect 22204 39340 22205 39404
rect 22139 39339 22205 39340
rect 12571 38996 12637 38997
rect 12571 38932 12572 38996
rect 12636 38932 12637 38996
rect 12571 38931 12637 38932
rect 9627 38044 9693 38045
rect 9627 37980 9628 38044
rect 9692 37980 9693 38044
rect 9627 37979 9693 37980
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4843 37364 4909 37365
rect 4843 37300 4844 37364
rect 4908 37300 4909 37364
rect 4843 37299 4909 37300
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4846 34781 4906 37299
rect 7235 36548 7301 36549
rect 7235 36484 7236 36548
rect 7300 36484 7301 36548
rect 7235 36483 7301 36484
rect 6131 36004 6197 36005
rect 6131 35940 6132 36004
rect 6196 35940 6197 36004
rect 6131 35939 6197 35940
rect 4843 34780 4909 34781
rect 4843 34716 4844 34780
rect 4908 34716 4909 34780
rect 4843 34715 4909 34716
rect 5211 34780 5277 34781
rect 5211 34716 5212 34780
rect 5276 34716 5277 34780
rect 5211 34715 5277 34716
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4843 32332 4909 32333
rect 4843 32268 4844 32332
rect 4908 32268 4909 32332
rect 4843 32267 4909 32268
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4846 31517 4906 32267
rect 4843 31516 4909 31517
rect 4843 31452 4844 31516
rect 4908 31452 4909 31516
rect 4843 31451 4909 31452
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 5214 24581 5274 34715
rect 6134 25533 6194 35939
rect 6315 33284 6381 33285
rect 6315 33220 6316 33284
rect 6380 33220 6381 33284
rect 6315 33219 6381 33220
rect 6318 26485 6378 33219
rect 7238 30429 7298 36483
rect 8155 34644 8221 34645
rect 8155 34580 8156 34644
rect 8220 34580 8221 34644
rect 8155 34579 8221 34580
rect 7235 30428 7301 30429
rect 7235 30364 7236 30428
rect 7300 30364 7301 30428
rect 7235 30363 7301 30364
rect 8158 26621 8218 34579
rect 9630 34237 9690 37979
rect 10363 35868 10429 35869
rect 10363 35804 10364 35868
rect 10428 35804 10429 35868
rect 10363 35803 10429 35804
rect 9627 34236 9693 34237
rect 9627 34172 9628 34236
rect 9692 34172 9693 34236
rect 9627 34171 9693 34172
rect 9443 31516 9509 31517
rect 9443 31452 9444 31516
rect 9508 31452 9509 31516
rect 9443 31451 9509 31452
rect 8891 30428 8957 30429
rect 8891 30364 8892 30428
rect 8956 30364 8957 30428
rect 8891 30363 8957 30364
rect 8155 26620 8221 26621
rect 8155 26556 8156 26620
rect 8220 26556 8221 26620
rect 8155 26555 8221 26556
rect 6315 26484 6381 26485
rect 6315 26420 6316 26484
rect 6380 26420 6381 26484
rect 6315 26419 6381 26420
rect 6131 25532 6197 25533
rect 6131 25468 6132 25532
rect 6196 25468 6197 25532
rect 6131 25467 6197 25468
rect 5211 24580 5277 24581
rect 5211 24516 5212 24580
rect 5276 24516 5277 24580
rect 5211 24515 5277 24516
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 8894 19005 8954 30363
rect 9446 29477 9506 31451
rect 9627 30700 9693 30701
rect 9627 30636 9628 30700
rect 9692 30636 9693 30700
rect 9627 30635 9693 30636
rect 9443 29476 9509 29477
rect 9443 29412 9444 29476
rect 9508 29412 9509 29476
rect 9443 29411 9509 29412
rect 9630 22269 9690 30635
rect 10366 23085 10426 35803
rect 12203 34780 12269 34781
rect 12203 34716 12204 34780
rect 12268 34716 12269 34780
rect 12203 34715 12269 34716
rect 11099 34644 11165 34645
rect 11099 34580 11100 34644
rect 11164 34580 11165 34644
rect 11099 34579 11165 34580
rect 11283 34644 11349 34645
rect 11283 34580 11284 34644
rect 11348 34580 11349 34644
rect 11283 34579 11349 34580
rect 11102 29341 11162 34579
rect 11286 32605 11346 34579
rect 11283 32604 11349 32605
rect 11283 32540 11284 32604
rect 11348 32540 11349 32604
rect 11283 32539 11349 32540
rect 12206 31381 12266 34715
rect 12387 32604 12453 32605
rect 12387 32540 12388 32604
rect 12452 32540 12453 32604
rect 12387 32539 12453 32540
rect 12203 31380 12269 31381
rect 12203 31316 12204 31380
rect 12268 31316 12269 31380
rect 12203 31315 12269 31316
rect 12390 29613 12450 32539
rect 12574 31653 12634 38931
rect 16435 37772 16501 37773
rect 16435 37708 16436 37772
rect 16500 37708 16501 37772
rect 16435 37707 16501 37708
rect 15331 36956 15397 36957
rect 15331 36892 15332 36956
rect 15396 36892 15397 36956
rect 15331 36891 15397 36892
rect 12755 36004 12821 36005
rect 12755 35940 12756 36004
rect 12820 35940 12821 36004
rect 12755 35939 12821 35940
rect 12571 31652 12637 31653
rect 12571 31588 12572 31652
rect 12636 31588 12637 31652
rect 12571 31587 12637 31588
rect 12387 29612 12453 29613
rect 12387 29548 12388 29612
rect 12452 29548 12453 29612
rect 12387 29547 12453 29548
rect 12758 29477 12818 35939
rect 15334 33690 15394 36891
rect 15150 33630 15394 33690
rect 13310 32270 13738 32330
rect 13310 31925 13370 32270
rect 13678 32197 13738 32270
rect 13491 32196 13557 32197
rect 13491 32132 13492 32196
rect 13556 32132 13557 32196
rect 13491 32131 13557 32132
rect 13675 32196 13741 32197
rect 13675 32132 13676 32196
rect 13740 32132 13741 32196
rect 13675 32131 13741 32132
rect 13307 31924 13373 31925
rect 13307 31860 13308 31924
rect 13372 31860 13373 31924
rect 13307 31859 13373 31860
rect 13494 31653 13554 32131
rect 13491 31652 13557 31653
rect 13491 31588 13492 31652
rect 13556 31588 13557 31652
rect 13491 31587 13557 31588
rect 13307 29612 13373 29613
rect 13307 29548 13308 29612
rect 13372 29548 13373 29612
rect 13307 29547 13373 29548
rect 12755 29476 12821 29477
rect 12755 29412 12756 29476
rect 12820 29412 12821 29476
rect 12755 29411 12821 29412
rect 11099 29340 11165 29341
rect 11099 29276 11100 29340
rect 11164 29276 11165 29340
rect 11099 29275 11165 29276
rect 13310 26077 13370 29547
rect 13494 27029 13554 31587
rect 15150 31109 15210 33630
rect 16251 31244 16317 31245
rect 16251 31180 16252 31244
rect 16316 31180 16317 31244
rect 16251 31179 16317 31180
rect 15147 31108 15213 31109
rect 15147 31044 15148 31108
rect 15212 31044 15213 31108
rect 15147 31043 15213 31044
rect 15331 30564 15397 30565
rect 15331 30500 15332 30564
rect 15396 30500 15397 30564
rect 15331 30499 15397 30500
rect 13675 28252 13741 28253
rect 13675 28188 13676 28252
rect 13740 28188 13741 28252
rect 13675 28187 13741 28188
rect 13678 27573 13738 28187
rect 15147 27844 15213 27845
rect 15147 27780 15148 27844
rect 15212 27780 15213 27844
rect 15147 27779 15213 27780
rect 13675 27572 13741 27573
rect 13675 27508 13676 27572
rect 13740 27508 13741 27572
rect 13675 27507 13741 27508
rect 13491 27028 13557 27029
rect 13491 26964 13492 27028
rect 13556 26964 13557 27028
rect 13491 26963 13557 26964
rect 13307 26076 13373 26077
rect 13307 26012 13308 26076
rect 13372 26012 13373 26076
rect 13307 26011 13373 26012
rect 15150 25941 15210 27779
rect 15334 26757 15394 30499
rect 15331 26756 15397 26757
rect 15331 26692 15332 26756
rect 15396 26692 15397 26756
rect 15331 26691 15397 26692
rect 15147 25940 15213 25941
rect 15147 25876 15148 25940
rect 15212 25876 15213 25940
rect 15147 25875 15213 25876
rect 16254 24853 16314 31179
rect 16438 26349 16498 37707
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19379 36548 19445 36549
rect 19379 36484 19380 36548
rect 19444 36484 19445 36548
rect 19379 36483 19445 36484
rect 18275 36412 18341 36413
rect 18275 36348 18276 36412
rect 18340 36348 18341 36412
rect 18275 36347 18341 36348
rect 17723 36276 17789 36277
rect 17723 36212 17724 36276
rect 17788 36212 17789 36276
rect 17723 36211 17789 36212
rect 17355 36140 17421 36141
rect 17355 36076 17356 36140
rect 17420 36076 17421 36140
rect 17355 36075 17421 36076
rect 17358 27301 17418 36075
rect 17726 29205 17786 36211
rect 18091 35868 18157 35869
rect 18091 35804 18092 35868
rect 18156 35804 18157 35868
rect 18091 35803 18157 35804
rect 17907 34916 17973 34917
rect 17907 34852 17908 34916
rect 17972 34852 17973 34916
rect 17907 34851 17973 34852
rect 17723 29204 17789 29205
rect 17723 29140 17724 29204
rect 17788 29140 17789 29204
rect 17723 29139 17789 29140
rect 17910 27573 17970 34851
rect 17907 27572 17973 27573
rect 17907 27508 17908 27572
rect 17972 27508 17973 27572
rect 17907 27507 17973 27508
rect 17355 27300 17421 27301
rect 17355 27236 17356 27300
rect 17420 27236 17421 27300
rect 17355 27235 17421 27236
rect 18094 26757 18154 35803
rect 18278 35325 18338 36347
rect 18275 35324 18341 35325
rect 18275 35260 18276 35324
rect 18340 35260 18341 35324
rect 18275 35259 18341 35260
rect 19195 35052 19261 35053
rect 19195 34988 19196 35052
rect 19260 34988 19261 35052
rect 19195 34987 19261 34988
rect 18275 31788 18341 31789
rect 18275 31724 18276 31788
rect 18340 31724 18341 31788
rect 18275 31723 18341 31724
rect 18278 28661 18338 31723
rect 19011 29748 19077 29749
rect 19011 29684 19012 29748
rect 19076 29684 19077 29748
rect 19011 29683 19077 29684
rect 18275 28660 18341 28661
rect 18275 28596 18276 28660
rect 18340 28596 18341 28660
rect 18275 28595 18341 28596
rect 18275 28524 18341 28525
rect 18275 28460 18276 28524
rect 18340 28460 18341 28524
rect 18275 28459 18341 28460
rect 18278 27165 18338 28459
rect 18275 27164 18341 27165
rect 18275 27100 18276 27164
rect 18340 27100 18341 27164
rect 18275 27099 18341 27100
rect 18091 26756 18157 26757
rect 18091 26692 18092 26756
rect 18156 26692 18157 26756
rect 18091 26691 18157 26692
rect 16435 26348 16501 26349
rect 16435 26284 16436 26348
rect 16500 26284 16501 26348
rect 16435 26283 16501 26284
rect 19014 26213 19074 29683
rect 19198 28933 19258 34987
rect 19382 29341 19442 36483
rect 19568 35936 19888 36960
rect 21955 36684 22021 36685
rect 21955 36620 21956 36684
rect 22020 36620 22021 36684
rect 21955 36619 22021 36620
rect 20115 36412 20181 36413
rect 20115 36348 20116 36412
rect 20180 36348 20181 36412
rect 20115 36347 20181 36348
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 20118 31653 20178 36347
rect 21035 35868 21101 35869
rect 21035 35804 21036 35868
rect 21100 35804 21101 35868
rect 21035 35803 21101 35804
rect 20851 33284 20917 33285
rect 20851 33220 20852 33284
rect 20916 33220 20917 33284
rect 20851 33219 20917 33220
rect 20667 32196 20733 32197
rect 20667 32132 20668 32196
rect 20732 32132 20733 32196
rect 20667 32131 20733 32132
rect 20115 31652 20181 31653
rect 20115 31588 20116 31652
rect 20180 31588 20181 31652
rect 20115 31587 20181 31588
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 20483 31516 20549 31517
rect 20483 31452 20484 31516
rect 20548 31452 20549 31516
rect 20483 31451 20549 31452
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19379 29340 19445 29341
rect 19379 29276 19380 29340
rect 19444 29276 19445 29340
rect 19379 29275 19445 29276
rect 19195 28932 19261 28933
rect 19195 28868 19196 28932
rect 19260 28868 19261 28932
rect 19195 28867 19261 28868
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19379 27844 19445 27845
rect 19379 27780 19380 27844
rect 19444 27780 19445 27844
rect 19379 27779 19445 27780
rect 19011 26212 19077 26213
rect 19011 26148 19012 26212
rect 19076 26148 19077 26212
rect 19011 26147 19077 26148
rect 19382 25125 19442 27779
rect 19568 27232 19888 28256
rect 20299 27300 20365 27301
rect 20299 27236 20300 27300
rect 20364 27236 20365 27300
rect 20299 27235 20365 27236
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19379 25124 19445 25125
rect 19379 25060 19380 25124
rect 19444 25060 19445 25124
rect 19379 25059 19445 25060
rect 19568 25056 19888 26080
rect 20302 25397 20362 27235
rect 20486 26213 20546 31451
rect 20670 26893 20730 32131
rect 20667 26892 20733 26893
rect 20667 26828 20668 26892
rect 20732 26828 20733 26892
rect 20667 26827 20733 26828
rect 20854 26485 20914 33219
rect 21038 31925 21098 35803
rect 21035 31924 21101 31925
rect 21035 31860 21036 31924
rect 21100 31860 21101 31924
rect 21035 31859 21101 31860
rect 21038 26485 21098 31859
rect 20851 26484 20917 26485
rect 20851 26420 20852 26484
rect 20916 26420 20917 26484
rect 20851 26419 20917 26420
rect 21035 26484 21101 26485
rect 21035 26420 21036 26484
rect 21100 26420 21101 26484
rect 21035 26419 21101 26420
rect 20483 26212 20549 26213
rect 20483 26148 20484 26212
rect 20548 26148 20549 26212
rect 20483 26147 20549 26148
rect 20483 26076 20549 26077
rect 20483 26012 20484 26076
rect 20548 26012 20549 26076
rect 20483 26011 20549 26012
rect 20486 25397 20546 26011
rect 20299 25396 20365 25397
rect 20299 25332 20300 25396
rect 20364 25332 20365 25396
rect 20299 25331 20365 25332
rect 20483 25396 20549 25397
rect 20483 25332 20484 25396
rect 20548 25332 20549 25396
rect 20483 25331 20549 25332
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 16251 24852 16317 24853
rect 16251 24788 16252 24852
rect 16316 24788 16317 24852
rect 16251 24787 16317 24788
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 10363 23084 10429 23085
rect 10363 23020 10364 23084
rect 10428 23020 10429 23084
rect 10363 23019 10429 23020
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 9627 22268 9693 22269
rect 9627 22204 9628 22268
rect 9692 22204 9693 22268
rect 9627 22203 9693 22204
rect 19568 21792 19888 22816
rect 21958 22541 22018 36619
rect 22142 29613 22202 39339
rect 27475 39268 27541 39269
rect 27475 39204 27476 39268
rect 27540 39204 27541 39268
rect 27475 39203 27541 39204
rect 27291 39132 27357 39133
rect 27291 39068 27292 39132
rect 27356 39068 27357 39132
rect 27291 39067 27357 39068
rect 23427 37636 23493 37637
rect 23427 37572 23428 37636
rect 23492 37572 23493 37636
rect 23427 37571 23493 37572
rect 23243 34644 23309 34645
rect 23243 34580 23244 34644
rect 23308 34580 23309 34644
rect 23243 34579 23309 34580
rect 22139 29612 22205 29613
rect 22139 29548 22140 29612
rect 22204 29548 22205 29612
rect 22139 29547 22205 29548
rect 22507 29068 22573 29069
rect 22507 29004 22508 29068
rect 22572 29004 22573 29068
rect 22507 29003 22573 29004
rect 21955 22540 22021 22541
rect 21955 22476 21956 22540
rect 22020 22476 22021 22540
rect 21955 22475 22021 22476
rect 21958 21997 22018 22475
rect 21955 21996 22021 21997
rect 21955 21932 21956 21996
rect 22020 21932 22021 21996
rect 21955 21931 22021 21932
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 22510 21317 22570 29003
rect 23246 28389 23306 34579
rect 23430 34373 23490 37571
rect 23611 37500 23677 37501
rect 23611 37436 23612 37500
rect 23676 37436 23677 37500
rect 23611 37435 23677 37436
rect 23427 34372 23493 34373
rect 23427 34308 23428 34372
rect 23492 34308 23493 34372
rect 23427 34307 23493 34308
rect 23614 31770 23674 37435
rect 26923 37364 26989 37365
rect 26923 37300 26924 37364
rect 26988 37300 26989 37364
rect 26923 37299 26989 37300
rect 24899 36548 24965 36549
rect 24899 36484 24900 36548
rect 24964 36484 24965 36548
rect 24899 36483 24965 36484
rect 23979 35732 24045 35733
rect 23979 35668 23980 35732
rect 24044 35668 24045 35732
rect 23979 35667 24045 35668
rect 23982 33421 24042 35667
rect 24902 35053 24962 36483
rect 25267 36276 25333 36277
rect 25267 36212 25268 36276
rect 25332 36212 25333 36276
rect 25267 36211 25333 36212
rect 24899 35052 24965 35053
rect 24899 34988 24900 35052
rect 24964 34988 24965 35052
rect 24899 34987 24965 34988
rect 23979 33420 24045 33421
rect 23979 33356 23980 33420
rect 24044 33356 24045 33420
rect 23979 33355 24045 33356
rect 23982 31925 24042 33355
rect 24715 32060 24781 32061
rect 24715 31996 24716 32060
rect 24780 31996 24781 32060
rect 24715 31995 24781 31996
rect 23979 31924 24045 31925
rect 23979 31860 23980 31924
rect 24044 31860 24045 31924
rect 23979 31859 24045 31860
rect 23430 31710 23674 31770
rect 23243 28388 23309 28389
rect 23243 28324 23244 28388
rect 23308 28324 23309 28388
rect 23243 28323 23309 28324
rect 22691 27708 22757 27709
rect 22691 27644 22692 27708
rect 22756 27644 22757 27708
rect 22691 27643 22757 27644
rect 22507 21316 22573 21317
rect 22507 21252 22508 21316
rect 22572 21252 22573 21316
rect 22507 21251 22573 21252
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 8891 19004 8957 19005
rect 8891 18940 8892 19004
rect 8956 18940 8957 19004
rect 8891 18939 8957 18940
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 18528 19888 19552
rect 22694 19141 22754 27643
rect 23430 27573 23490 31710
rect 23611 30564 23677 30565
rect 23611 30500 23612 30564
rect 23676 30500 23677 30564
rect 23611 30499 23677 30500
rect 23427 27572 23493 27573
rect 23427 27508 23428 27572
rect 23492 27508 23493 27572
rect 23427 27507 23493 27508
rect 23614 27301 23674 30499
rect 24531 30292 24597 30293
rect 24531 30228 24532 30292
rect 24596 30228 24597 30292
rect 24531 30227 24597 30228
rect 23795 28932 23861 28933
rect 23795 28868 23796 28932
rect 23860 28868 23861 28932
rect 23795 28867 23861 28868
rect 23611 27300 23677 27301
rect 23611 27236 23612 27300
rect 23676 27236 23677 27300
rect 23611 27235 23677 27236
rect 23798 24853 23858 28867
rect 24534 27165 24594 30227
rect 24718 27981 24778 31995
rect 24902 29069 24962 34987
rect 25270 33013 25330 36211
rect 26187 36140 26253 36141
rect 26187 36076 26188 36140
rect 26252 36076 26253 36140
rect 26187 36075 26253 36076
rect 26190 34237 26250 36075
rect 26187 34236 26253 34237
rect 26187 34172 26188 34236
rect 26252 34172 26253 34236
rect 26187 34171 26253 34172
rect 26371 33284 26437 33285
rect 26371 33220 26372 33284
rect 26436 33220 26437 33284
rect 26371 33219 26437 33220
rect 25267 33012 25333 33013
rect 25267 32948 25268 33012
rect 25332 32948 25333 33012
rect 25267 32947 25333 32948
rect 25083 31788 25149 31789
rect 25083 31724 25084 31788
rect 25148 31724 25149 31788
rect 25083 31723 25149 31724
rect 24899 29068 24965 29069
rect 24899 29004 24900 29068
rect 24964 29004 24965 29068
rect 24899 29003 24965 29004
rect 24715 27980 24781 27981
rect 24715 27916 24716 27980
rect 24780 27916 24781 27980
rect 24715 27915 24781 27916
rect 24531 27164 24597 27165
rect 24531 27100 24532 27164
rect 24596 27100 24597 27164
rect 24531 27099 24597 27100
rect 24163 26348 24229 26349
rect 24163 26284 24164 26348
rect 24228 26284 24229 26348
rect 24163 26283 24229 26284
rect 23795 24852 23861 24853
rect 23795 24788 23796 24852
rect 23860 24788 23861 24852
rect 23795 24787 23861 24788
rect 23427 22948 23493 22949
rect 23427 22884 23428 22948
rect 23492 22884 23493 22948
rect 23427 22883 23493 22884
rect 23430 19277 23490 22883
rect 24166 21589 24226 26283
rect 24347 21996 24413 21997
rect 24347 21932 24348 21996
rect 24412 21932 24413 21996
rect 24347 21931 24413 21932
rect 24163 21588 24229 21589
rect 24163 21524 24164 21588
rect 24228 21524 24229 21588
rect 24163 21523 24229 21524
rect 23427 19276 23493 19277
rect 23427 19212 23428 19276
rect 23492 19212 23493 19276
rect 23427 19211 23493 19212
rect 22691 19140 22757 19141
rect 22691 19076 22692 19140
rect 22756 19076 22757 19140
rect 22691 19075 22757 19076
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 24350 16557 24410 21931
rect 24347 16556 24413 16557
rect 24347 16492 24348 16556
rect 24412 16492 24413 16556
rect 24347 16491 24413 16492
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 25086 14381 25146 31723
rect 25451 31380 25517 31381
rect 25451 31316 25452 31380
rect 25516 31316 25517 31380
rect 25451 31315 25517 31316
rect 25454 30157 25514 31315
rect 26003 30428 26069 30429
rect 26003 30364 26004 30428
rect 26068 30364 26069 30428
rect 26003 30363 26069 30364
rect 25451 30156 25517 30157
rect 25451 30092 25452 30156
rect 25516 30092 25517 30156
rect 25451 30091 25517 30092
rect 25635 30156 25701 30157
rect 25635 30092 25636 30156
rect 25700 30092 25701 30156
rect 25635 30091 25701 30092
rect 25638 29069 25698 30091
rect 25635 29068 25701 29069
rect 25635 29004 25636 29068
rect 25700 29004 25701 29068
rect 25635 29003 25701 29004
rect 26006 27573 26066 30363
rect 26187 28388 26253 28389
rect 26187 28324 26188 28388
rect 26252 28324 26253 28388
rect 26187 28323 26253 28324
rect 26003 27572 26069 27573
rect 26003 27508 26004 27572
rect 26068 27508 26069 27572
rect 26003 27507 26069 27508
rect 25819 27164 25885 27165
rect 25819 27100 25820 27164
rect 25884 27100 25885 27164
rect 25819 27099 25885 27100
rect 25267 26756 25333 26757
rect 25267 26692 25268 26756
rect 25332 26692 25333 26756
rect 25267 26691 25333 26692
rect 25270 25261 25330 26691
rect 25267 25260 25333 25261
rect 25267 25196 25268 25260
rect 25332 25196 25333 25260
rect 25267 25195 25333 25196
rect 25822 22133 25882 27099
rect 26003 25804 26069 25805
rect 26003 25740 26004 25804
rect 26068 25740 26069 25804
rect 26003 25739 26069 25740
rect 25819 22132 25885 22133
rect 25819 22068 25820 22132
rect 25884 22068 25885 22132
rect 25819 22067 25885 22068
rect 26006 21725 26066 25739
rect 26190 23221 26250 28323
rect 26374 26621 26434 33219
rect 26555 31788 26621 31789
rect 26555 31724 26556 31788
rect 26620 31724 26621 31788
rect 26555 31723 26621 31724
rect 26558 28253 26618 31723
rect 26926 29749 26986 37299
rect 27294 33557 27354 39067
rect 27478 35869 27538 39203
rect 27843 38316 27909 38317
rect 27843 38252 27844 38316
rect 27908 38252 27909 38316
rect 27843 38251 27909 38252
rect 27475 35868 27541 35869
rect 27475 35804 27476 35868
rect 27540 35804 27541 35868
rect 27475 35803 27541 35804
rect 27846 34781 27906 38251
rect 29315 37772 29381 37773
rect 29315 37708 29316 37772
rect 29380 37708 29381 37772
rect 29315 37707 29381 37708
rect 27843 34780 27909 34781
rect 27843 34716 27844 34780
rect 27908 34716 27909 34780
rect 27843 34715 27909 34716
rect 27291 33556 27357 33557
rect 27291 33492 27292 33556
rect 27356 33492 27357 33556
rect 27291 33491 27357 33492
rect 27475 33420 27541 33421
rect 27475 33356 27476 33420
rect 27540 33356 27541 33420
rect 27475 33355 27541 33356
rect 27291 31652 27357 31653
rect 27291 31588 27292 31652
rect 27356 31588 27357 31652
rect 27291 31587 27357 31588
rect 26923 29748 26989 29749
rect 26923 29684 26924 29748
rect 26988 29684 26989 29748
rect 26923 29683 26989 29684
rect 26555 28252 26621 28253
rect 26555 28188 26556 28252
rect 26620 28188 26621 28252
rect 26555 28187 26621 28188
rect 27107 27572 27173 27573
rect 27107 27508 27108 27572
rect 27172 27508 27173 27572
rect 27107 27507 27173 27508
rect 26371 26620 26437 26621
rect 26371 26556 26372 26620
rect 26436 26556 26437 26620
rect 26371 26555 26437 26556
rect 26555 25804 26621 25805
rect 26555 25740 26556 25804
rect 26620 25740 26621 25804
rect 26555 25739 26621 25740
rect 26558 25397 26618 25739
rect 26555 25396 26621 25397
rect 26555 25332 26556 25396
rect 26620 25332 26621 25396
rect 26555 25331 26621 25332
rect 26187 23220 26253 23221
rect 26187 23156 26188 23220
rect 26252 23156 26253 23220
rect 26187 23155 26253 23156
rect 26371 22676 26437 22677
rect 26371 22612 26372 22676
rect 26436 22612 26437 22676
rect 26371 22611 26437 22612
rect 26003 21724 26069 21725
rect 26003 21660 26004 21724
rect 26068 21660 26069 21724
rect 26003 21659 26069 21660
rect 26374 19277 26434 22611
rect 26558 20093 26618 25331
rect 27110 23221 27170 27507
rect 27107 23220 27173 23221
rect 27107 23156 27108 23220
rect 27172 23156 27173 23220
rect 27107 23155 27173 23156
rect 27294 21861 27354 31587
rect 27478 28117 27538 33355
rect 28211 33284 28277 33285
rect 28211 33220 28212 33284
rect 28276 33220 28277 33284
rect 28211 33219 28277 33220
rect 28947 33284 29013 33285
rect 28947 33220 28948 33284
rect 29012 33220 29013 33284
rect 28947 33219 29013 33220
rect 28027 32740 28093 32741
rect 28027 32676 28028 32740
rect 28092 32676 28093 32740
rect 28027 32675 28093 32676
rect 28030 28933 28090 32675
rect 28214 32061 28274 33219
rect 28579 33012 28645 33013
rect 28579 32948 28580 33012
rect 28644 32948 28645 33012
rect 28579 32947 28645 32948
rect 28395 32604 28461 32605
rect 28395 32540 28396 32604
rect 28460 32540 28461 32604
rect 28395 32539 28461 32540
rect 28211 32060 28277 32061
rect 28211 31996 28212 32060
rect 28276 31996 28277 32060
rect 28211 31995 28277 31996
rect 28398 31789 28458 32539
rect 28395 31788 28461 31789
rect 28395 31724 28396 31788
rect 28460 31724 28461 31788
rect 28395 31723 28461 31724
rect 28395 30972 28461 30973
rect 28395 30908 28396 30972
rect 28460 30908 28461 30972
rect 28395 30907 28461 30908
rect 28027 28932 28093 28933
rect 28027 28868 28028 28932
rect 28092 28868 28093 28932
rect 28027 28867 28093 28868
rect 27475 28116 27541 28117
rect 27475 28052 27476 28116
rect 27540 28052 27541 28116
rect 27475 28051 27541 28052
rect 28211 28116 28277 28117
rect 28211 28052 28212 28116
rect 28276 28052 28277 28116
rect 28211 28051 28277 28052
rect 27475 27572 27541 27573
rect 27475 27508 27476 27572
rect 27540 27508 27541 27572
rect 27475 27507 27541 27508
rect 27478 22813 27538 27507
rect 27659 26620 27725 26621
rect 27659 26556 27660 26620
rect 27724 26556 27725 26620
rect 27659 26555 27725 26556
rect 27662 23493 27722 26555
rect 28214 25533 28274 28051
rect 28211 25532 28277 25533
rect 28211 25468 28212 25532
rect 28276 25468 28277 25532
rect 28211 25467 28277 25468
rect 28214 23493 28274 25467
rect 27659 23492 27725 23493
rect 27659 23428 27660 23492
rect 27724 23428 27725 23492
rect 27659 23427 27725 23428
rect 28211 23492 28277 23493
rect 28211 23428 28212 23492
rect 28276 23428 28277 23492
rect 28211 23427 28277 23428
rect 27475 22812 27541 22813
rect 27475 22748 27476 22812
rect 27540 22748 27541 22812
rect 27475 22747 27541 22748
rect 27291 21860 27357 21861
rect 27291 21796 27292 21860
rect 27356 21796 27357 21860
rect 27291 21795 27357 21796
rect 28398 20637 28458 30907
rect 28582 30293 28642 32947
rect 28950 30565 29010 33219
rect 29131 33012 29197 33013
rect 29131 32948 29132 33012
rect 29196 32948 29197 33012
rect 29131 32947 29197 32948
rect 28947 30564 29013 30565
rect 28947 30500 28948 30564
rect 29012 30500 29013 30564
rect 28947 30499 29013 30500
rect 28579 30292 28645 30293
rect 28579 30228 28580 30292
rect 28644 30228 28645 30292
rect 28579 30227 28645 30228
rect 28947 29748 29013 29749
rect 28947 29684 28948 29748
rect 29012 29684 29013 29748
rect 28947 29683 29013 29684
rect 28763 29476 28829 29477
rect 28763 29412 28764 29476
rect 28828 29412 28829 29476
rect 28763 29411 28829 29412
rect 28766 26213 28826 29411
rect 28763 26212 28829 26213
rect 28763 26148 28764 26212
rect 28828 26148 28829 26212
rect 28763 26147 28829 26148
rect 28763 24988 28829 24989
rect 28763 24924 28764 24988
rect 28828 24924 28829 24988
rect 28763 24923 28829 24924
rect 28579 23492 28645 23493
rect 28579 23428 28580 23492
rect 28644 23428 28645 23492
rect 28579 23427 28645 23428
rect 28395 20636 28461 20637
rect 28395 20572 28396 20636
rect 28460 20572 28461 20636
rect 28395 20571 28461 20572
rect 26555 20092 26621 20093
rect 26555 20028 26556 20092
rect 26620 20028 26621 20092
rect 26555 20027 26621 20028
rect 26371 19276 26437 19277
rect 26371 19212 26372 19276
rect 26436 19212 26437 19276
rect 26371 19211 26437 19212
rect 28582 16965 28642 23427
rect 28766 20229 28826 24923
rect 28950 24853 29010 29683
rect 29134 26349 29194 32947
rect 29318 31789 29378 37707
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 33179 36004 33245 36005
rect 33179 35940 33180 36004
rect 33244 35940 33245 36004
rect 33179 35939 33245 35940
rect 29499 35324 29565 35325
rect 29499 35260 29500 35324
rect 29564 35260 29565 35324
rect 29499 35259 29565 35260
rect 29502 32061 29562 35259
rect 30419 35188 30485 35189
rect 30419 35124 30420 35188
rect 30484 35124 30485 35188
rect 30419 35123 30485 35124
rect 29683 34644 29749 34645
rect 29683 34580 29684 34644
rect 29748 34580 29749 34644
rect 29683 34579 29749 34580
rect 29686 32197 29746 34579
rect 29683 32196 29749 32197
rect 29683 32132 29684 32196
rect 29748 32132 29749 32196
rect 29683 32131 29749 32132
rect 29499 32060 29565 32061
rect 29499 31996 29500 32060
rect 29564 31996 29565 32060
rect 29499 31995 29565 31996
rect 29315 31788 29381 31789
rect 29315 31724 29316 31788
rect 29380 31724 29381 31788
rect 29315 31723 29381 31724
rect 30051 31380 30117 31381
rect 30051 31316 30052 31380
rect 30116 31316 30117 31380
rect 30051 31315 30117 31316
rect 29315 29068 29381 29069
rect 29315 29004 29316 29068
rect 29380 29004 29381 29068
rect 29315 29003 29381 29004
rect 29131 26348 29197 26349
rect 29131 26284 29132 26348
rect 29196 26284 29197 26348
rect 29131 26283 29197 26284
rect 28947 24852 29013 24853
rect 28947 24788 28948 24852
rect 29012 24788 29013 24852
rect 28947 24787 29013 24788
rect 29131 24308 29197 24309
rect 29131 24244 29132 24308
rect 29196 24244 29197 24308
rect 29131 24243 29197 24244
rect 28763 20228 28829 20229
rect 28763 20164 28764 20228
rect 28828 20164 28829 20228
rect 28763 20163 28829 20164
rect 29134 19549 29194 24243
rect 29318 21589 29378 29003
rect 29683 27980 29749 27981
rect 29683 27916 29684 27980
rect 29748 27916 29749 27980
rect 29683 27915 29749 27916
rect 29499 27028 29565 27029
rect 29499 26964 29500 27028
rect 29564 26964 29565 27028
rect 29499 26963 29565 26964
rect 29502 23901 29562 26963
rect 29499 23900 29565 23901
rect 29499 23836 29500 23900
rect 29564 23836 29565 23900
rect 29499 23835 29565 23836
rect 29686 22133 29746 27915
rect 29867 25532 29933 25533
rect 29867 25468 29868 25532
rect 29932 25468 29933 25532
rect 29867 25467 29933 25468
rect 29870 22541 29930 25467
rect 29867 22540 29933 22541
rect 29867 22476 29868 22540
rect 29932 22476 29933 22540
rect 29867 22475 29933 22476
rect 29683 22132 29749 22133
rect 29683 22068 29684 22132
rect 29748 22068 29749 22132
rect 29683 22067 29749 22068
rect 29315 21588 29381 21589
rect 29315 21524 29316 21588
rect 29380 21524 29381 21588
rect 29315 21523 29381 21524
rect 30054 20909 30114 31315
rect 30422 30701 30482 35123
rect 30787 34372 30853 34373
rect 30787 34308 30788 34372
rect 30852 34308 30853 34372
rect 30787 34307 30853 34308
rect 30419 30700 30485 30701
rect 30419 30636 30420 30700
rect 30484 30636 30485 30700
rect 30419 30635 30485 30636
rect 30603 30700 30669 30701
rect 30603 30636 30604 30700
rect 30668 30636 30669 30700
rect 30603 30635 30669 30636
rect 30606 28797 30666 30635
rect 30790 28933 30850 34307
rect 31339 33692 31405 33693
rect 31339 33628 31340 33692
rect 31404 33628 31405 33692
rect 31339 33627 31405 33628
rect 31155 30020 31221 30021
rect 31155 29956 31156 30020
rect 31220 29956 31221 30020
rect 31155 29955 31221 29956
rect 30787 28932 30853 28933
rect 30787 28868 30788 28932
rect 30852 28868 30853 28932
rect 30787 28867 30853 28868
rect 30603 28796 30669 28797
rect 30603 28732 30604 28796
rect 30668 28732 30669 28796
rect 30603 28731 30669 28732
rect 30787 28796 30853 28797
rect 30787 28732 30788 28796
rect 30852 28732 30853 28796
rect 30787 28731 30853 28732
rect 30419 27980 30485 27981
rect 30419 27916 30420 27980
rect 30484 27916 30485 27980
rect 30419 27915 30485 27916
rect 30235 26484 30301 26485
rect 30235 26420 30236 26484
rect 30300 26420 30301 26484
rect 30235 26419 30301 26420
rect 30051 20908 30117 20909
rect 30051 20844 30052 20908
rect 30116 20844 30117 20908
rect 30051 20843 30117 20844
rect 30238 19685 30298 26419
rect 30422 22677 30482 27915
rect 30603 26348 30669 26349
rect 30603 26284 30604 26348
rect 30668 26284 30669 26348
rect 30603 26283 30669 26284
rect 30419 22676 30485 22677
rect 30419 22612 30420 22676
rect 30484 22612 30485 22676
rect 30419 22611 30485 22612
rect 30606 20229 30666 26283
rect 30790 24853 30850 28731
rect 30971 27980 31037 27981
rect 30971 27916 30972 27980
rect 31036 27916 31037 27980
rect 30971 27915 31037 27916
rect 30974 25261 31034 27915
rect 31158 27029 31218 29955
rect 31342 27573 31402 33627
rect 33182 33285 33242 35939
rect 34099 35596 34165 35597
rect 34099 35532 34100 35596
rect 34164 35532 34165 35596
rect 34099 35531 34165 35532
rect 33731 34236 33797 34237
rect 33731 34172 33732 34236
rect 33796 34172 33797 34236
rect 33731 34171 33797 34172
rect 33179 33284 33245 33285
rect 33179 33220 33180 33284
rect 33244 33220 33245 33284
rect 33179 33219 33245 33220
rect 33547 33284 33613 33285
rect 33547 33220 33548 33284
rect 33612 33220 33613 33284
rect 33547 33219 33613 33220
rect 31891 32468 31957 32469
rect 31891 32404 31892 32468
rect 31956 32404 31957 32468
rect 31891 32403 31957 32404
rect 31523 28660 31589 28661
rect 31523 28596 31524 28660
rect 31588 28596 31589 28660
rect 31523 28595 31589 28596
rect 31339 27572 31405 27573
rect 31339 27508 31340 27572
rect 31404 27508 31405 27572
rect 31339 27507 31405 27508
rect 31526 27437 31586 28595
rect 31707 28116 31773 28117
rect 31707 28052 31708 28116
rect 31772 28052 31773 28116
rect 31707 28051 31773 28052
rect 31523 27436 31589 27437
rect 31523 27372 31524 27436
rect 31588 27372 31589 27436
rect 31523 27371 31589 27372
rect 31155 27028 31221 27029
rect 31155 26964 31156 27028
rect 31220 26964 31221 27028
rect 31155 26963 31221 26964
rect 30971 25260 31037 25261
rect 30971 25196 30972 25260
rect 31036 25196 31037 25260
rect 30971 25195 31037 25196
rect 30787 24852 30853 24853
rect 30787 24788 30788 24852
rect 30852 24788 30853 24852
rect 30787 24787 30853 24788
rect 30974 23765 31034 25195
rect 30971 23764 31037 23765
rect 30971 23700 30972 23764
rect 31036 23700 31037 23764
rect 30971 23699 31037 23700
rect 31158 22110 31218 26963
rect 31523 25940 31589 25941
rect 31523 25876 31524 25940
rect 31588 25876 31589 25940
rect 31523 25875 31589 25876
rect 30790 22050 31218 22110
rect 30603 20228 30669 20229
rect 30603 20164 30604 20228
rect 30668 20164 30669 20228
rect 30603 20163 30669 20164
rect 30606 19821 30666 20163
rect 30603 19820 30669 19821
rect 30603 19756 30604 19820
rect 30668 19756 30669 19820
rect 30603 19755 30669 19756
rect 30235 19684 30301 19685
rect 30235 19620 30236 19684
rect 30300 19620 30301 19684
rect 30235 19619 30301 19620
rect 29131 19548 29197 19549
rect 29131 19484 29132 19548
rect 29196 19484 29197 19548
rect 29131 19483 29197 19484
rect 30051 18052 30117 18053
rect 30051 17988 30052 18052
rect 30116 17988 30117 18052
rect 30051 17987 30117 17988
rect 28579 16964 28645 16965
rect 28579 16900 28580 16964
rect 28644 16900 28645 16964
rect 28579 16899 28645 16900
rect 25083 14380 25149 14381
rect 25083 14316 25084 14380
rect 25148 14316 25149 14380
rect 25083 14315 25149 14316
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 30054 8533 30114 17987
rect 30790 15333 30850 22050
rect 31526 21861 31586 25875
rect 31710 24309 31770 28051
rect 31894 26618 31954 32403
rect 33363 32196 33429 32197
rect 33363 32132 33364 32196
rect 33428 32132 33429 32196
rect 33363 32131 33429 32132
rect 32995 31108 33061 31109
rect 32995 31044 32996 31108
rect 33060 31044 33061 31108
rect 32995 31043 33061 31044
rect 32443 29884 32509 29885
rect 32443 29820 32444 29884
rect 32508 29820 32509 29884
rect 32443 29819 32509 29820
rect 32075 29204 32141 29205
rect 32075 29140 32076 29204
rect 32140 29140 32141 29204
rect 32075 29139 32141 29140
rect 32259 29204 32325 29205
rect 32259 29140 32260 29204
rect 32324 29140 32325 29204
rect 32259 29139 32325 29140
rect 32078 26893 32138 29139
rect 32075 26892 32141 26893
rect 32075 26828 32076 26892
rect 32140 26828 32141 26892
rect 32075 26827 32141 26828
rect 31894 26558 32138 26618
rect 31891 26348 31957 26349
rect 31891 26284 31892 26348
rect 31956 26284 31957 26348
rect 31891 26283 31957 26284
rect 31707 24308 31773 24309
rect 31707 24244 31708 24308
rect 31772 24244 31773 24308
rect 31707 24243 31773 24244
rect 31894 22110 31954 26283
rect 32078 22133 32138 26558
rect 32262 22541 32322 29139
rect 32446 24853 32506 29819
rect 32998 27029 33058 31043
rect 33179 30292 33245 30293
rect 33179 30228 33180 30292
rect 33244 30228 33245 30292
rect 33179 30227 33245 30228
rect 32995 27028 33061 27029
rect 32995 26964 32996 27028
rect 33060 26964 33061 27028
rect 32995 26963 33061 26964
rect 32995 26756 33061 26757
rect 32995 26692 32996 26756
rect 33060 26692 33061 26756
rect 32995 26691 33061 26692
rect 32443 24852 32509 24853
rect 32443 24788 32444 24852
rect 32508 24788 32509 24852
rect 32443 24787 32509 24788
rect 32627 24852 32693 24853
rect 32627 24788 32628 24852
rect 32692 24788 32693 24852
rect 32627 24787 32693 24788
rect 32259 22540 32325 22541
rect 32259 22476 32260 22540
rect 32324 22476 32325 22540
rect 32259 22475 32325 22476
rect 31710 22050 31954 22110
rect 32075 22132 32141 22133
rect 32075 22068 32076 22132
rect 32140 22068 32141 22132
rect 32075 22067 32141 22068
rect 30971 21860 31037 21861
rect 30971 21796 30972 21860
rect 31036 21796 31037 21860
rect 30971 21795 31037 21796
rect 31523 21860 31589 21861
rect 31523 21796 31524 21860
rect 31588 21796 31589 21860
rect 31523 21795 31589 21796
rect 30974 18189 31034 21795
rect 31710 21722 31770 22050
rect 31710 21662 31954 21722
rect 30971 18188 31037 18189
rect 30971 18124 30972 18188
rect 31036 18124 31037 18188
rect 30971 18123 31037 18124
rect 30974 16557 31034 18123
rect 31894 18050 31954 21662
rect 32630 20773 32690 24787
rect 32811 24444 32877 24445
rect 32811 24380 32812 24444
rect 32876 24380 32877 24444
rect 32811 24379 32877 24380
rect 32627 20772 32693 20773
rect 32627 20708 32628 20772
rect 32692 20708 32693 20772
rect 32627 20707 32693 20708
rect 32814 20501 32874 24379
rect 32998 24037 33058 26691
rect 33182 25397 33242 30227
rect 33366 30157 33426 32131
rect 33550 31653 33610 33219
rect 33547 31652 33613 31653
rect 33547 31588 33548 31652
rect 33612 31588 33613 31652
rect 33547 31587 33613 31588
rect 33363 30156 33429 30157
rect 33363 30092 33364 30156
rect 33428 30092 33429 30156
rect 33363 30091 33429 30092
rect 33547 30156 33613 30157
rect 33547 30092 33548 30156
rect 33612 30092 33613 30156
rect 33547 30091 33613 30092
rect 33363 29340 33429 29341
rect 33363 29276 33364 29340
rect 33428 29338 33429 29340
rect 33550 29338 33610 30091
rect 33428 29278 33610 29338
rect 33428 29276 33429 29278
rect 33363 29275 33429 29276
rect 33734 29205 33794 34171
rect 33915 33556 33981 33557
rect 33915 33492 33916 33556
rect 33980 33492 33981 33556
rect 33915 33491 33981 33492
rect 33918 30293 33978 33491
rect 33915 30292 33981 30293
rect 33915 30228 33916 30292
rect 33980 30228 33981 30292
rect 33915 30227 33981 30228
rect 33731 29204 33797 29205
rect 33731 29140 33732 29204
rect 33796 29140 33797 29204
rect 33731 29139 33797 29140
rect 33363 29068 33429 29069
rect 33363 29004 33364 29068
rect 33428 29004 33429 29068
rect 33363 29003 33429 29004
rect 33179 25396 33245 25397
rect 33179 25332 33180 25396
rect 33244 25332 33245 25396
rect 33179 25331 33245 25332
rect 32995 24036 33061 24037
rect 32995 23972 32996 24036
rect 33060 23972 33061 24036
rect 32995 23971 33061 23972
rect 33366 22949 33426 29003
rect 34102 28661 34162 35531
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 36123 34916 36189 34917
rect 36123 34852 36124 34916
rect 36188 34852 36189 34916
rect 36123 34851 36189 34852
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34283 34236 34349 34237
rect 34283 34172 34284 34236
rect 34348 34172 34349 34236
rect 34283 34171 34349 34172
rect 34286 29477 34346 34171
rect 34928 33216 35248 34240
rect 35571 34236 35637 34237
rect 35571 34172 35572 34236
rect 35636 34172 35637 34236
rect 35571 34171 35637 34172
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34651 32332 34717 32333
rect 34651 32268 34652 32332
rect 34716 32268 34717 32332
rect 34651 32267 34717 32268
rect 34467 31788 34533 31789
rect 34467 31724 34468 31788
rect 34532 31724 34533 31788
rect 34467 31723 34533 31724
rect 34470 31245 34530 31723
rect 34654 31381 34714 32267
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34651 31380 34717 31381
rect 34651 31316 34652 31380
rect 34716 31316 34717 31380
rect 34651 31315 34717 31316
rect 34467 31244 34533 31245
rect 34467 31180 34468 31244
rect 34532 31180 34533 31244
rect 34467 31179 34533 31180
rect 34928 31040 35248 32064
rect 35387 32060 35453 32061
rect 35387 31996 35388 32060
rect 35452 31996 35453 32060
rect 35387 31995 35453 31996
rect 35390 31381 35450 31995
rect 35387 31380 35453 31381
rect 35387 31316 35388 31380
rect 35452 31316 35453 31380
rect 35387 31315 35453 31316
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34651 30564 34717 30565
rect 34651 30500 34652 30564
rect 34716 30500 34717 30564
rect 34651 30499 34717 30500
rect 34467 29748 34533 29749
rect 34467 29684 34468 29748
rect 34532 29684 34533 29748
rect 34467 29683 34533 29684
rect 34283 29476 34349 29477
rect 34283 29412 34284 29476
rect 34348 29412 34349 29476
rect 34283 29411 34349 29412
rect 34099 28660 34165 28661
rect 34099 28596 34100 28660
rect 34164 28596 34165 28660
rect 34099 28595 34165 28596
rect 33915 27844 33981 27845
rect 33915 27780 33916 27844
rect 33980 27780 33981 27844
rect 33915 27779 33981 27780
rect 33731 25396 33797 25397
rect 33731 25332 33732 25396
rect 33796 25332 33797 25396
rect 33731 25331 33797 25332
rect 33547 24444 33613 24445
rect 33547 24380 33548 24444
rect 33612 24380 33613 24444
rect 33547 24379 33613 24380
rect 33550 23493 33610 24379
rect 33547 23492 33613 23493
rect 33547 23428 33548 23492
rect 33612 23428 33613 23492
rect 33547 23427 33613 23428
rect 33363 22948 33429 22949
rect 33363 22884 33364 22948
rect 33428 22884 33429 22948
rect 33363 22883 33429 22884
rect 33734 21181 33794 25331
rect 33918 22677 33978 27779
rect 34102 27573 34162 28595
rect 34286 27845 34346 29411
rect 34470 29205 34530 29683
rect 34467 29204 34533 29205
rect 34467 29140 34468 29204
rect 34532 29140 34533 29204
rect 34467 29139 34533 29140
rect 34467 27980 34533 27981
rect 34467 27916 34468 27980
rect 34532 27916 34533 27980
rect 34467 27915 34533 27916
rect 34283 27844 34349 27845
rect 34283 27780 34284 27844
rect 34348 27780 34349 27844
rect 34283 27779 34349 27780
rect 34099 27572 34165 27573
rect 34099 27508 34100 27572
rect 34164 27508 34165 27572
rect 34099 27507 34165 27508
rect 34283 27572 34349 27573
rect 34283 27508 34284 27572
rect 34348 27508 34349 27572
rect 34283 27507 34349 27508
rect 34286 26077 34346 27507
rect 34283 26076 34349 26077
rect 34283 26012 34284 26076
rect 34348 26012 34349 26076
rect 34283 26011 34349 26012
rect 33915 22676 33981 22677
rect 33915 22612 33916 22676
rect 33980 22612 33981 22676
rect 33915 22611 33981 22612
rect 33915 22404 33981 22405
rect 33915 22340 33916 22404
rect 33980 22340 33981 22404
rect 33915 22339 33981 22340
rect 33731 21180 33797 21181
rect 33731 21116 33732 21180
rect 33796 21116 33797 21180
rect 33731 21115 33797 21116
rect 32995 20772 33061 20773
rect 32995 20708 32996 20772
rect 33060 20708 33061 20772
rect 32995 20707 33061 20708
rect 32443 20500 32509 20501
rect 32443 20436 32444 20500
rect 32508 20436 32509 20500
rect 32443 20435 32509 20436
rect 32627 20500 32693 20501
rect 32627 20436 32628 20500
rect 32692 20436 32693 20500
rect 32627 20435 32693 20436
rect 32811 20500 32877 20501
rect 32811 20436 32812 20500
rect 32876 20436 32877 20500
rect 32811 20435 32877 20436
rect 31710 17990 31954 18050
rect 31710 17917 31770 17990
rect 31707 17916 31773 17917
rect 31707 17852 31708 17916
rect 31772 17852 31773 17916
rect 31707 17851 31773 17852
rect 30971 16556 31037 16557
rect 30971 16492 30972 16556
rect 31036 16492 31037 16556
rect 30971 16491 31037 16492
rect 30787 15332 30853 15333
rect 30787 15268 30788 15332
rect 30852 15268 30853 15332
rect 30787 15267 30853 15268
rect 30051 8532 30117 8533
rect 30051 8468 30052 8532
rect 30116 8468 30117 8532
rect 30051 8467 30117 8468
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 32446 6765 32506 20435
rect 32630 19685 32690 20435
rect 32627 19684 32693 19685
rect 32627 19620 32628 19684
rect 32692 19620 32693 19684
rect 32627 19619 32693 19620
rect 32811 19548 32877 19549
rect 32811 19484 32812 19548
rect 32876 19484 32877 19548
rect 32811 19483 32877 19484
rect 32443 6764 32509 6765
rect 32443 6700 32444 6764
rect 32508 6700 32509 6764
rect 32443 6699 32509 6700
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 32814 2549 32874 19483
rect 32998 6901 33058 20707
rect 33918 19685 33978 22339
rect 34286 20501 34346 26011
rect 34470 22133 34530 27915
rect 34654 27029 34714 30499
rect 34928 29952 35248 30976
rect 35390 30701 35450 31315
rect 35387 30700 35453 30701
rect 35387 30636 35388 30700
rect 35452 30636 35453 30700
rect 35387 30635 35453 30636
rect 35387 30428 35453 30429
rect 35387 30364 35388 30428
rect 35452 30364 35453 30428
rect 35387 30363 35453 30364
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34651 27028 34717 27029
rect 34651 26964 34652 27028
rect 34716 26964 34717 27028
rect 34651 26963 34717 26964
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34651 26620 34717 26621
rect 34651 26556 34652 26620
rect 34716 26556 34717 26620
rect 34651 26555 34717 26556
rect 34654 23765 34714 26555
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34651 23764 34717 23765
rect 34651 23700 34652 23764
rect 34716 23700 34717 23764
rect 34651 23699 34717 23700
rect 34654 23221 34714 23699
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34651 23220 34717 23221
rect 34651 23156 34652 23220
rect 34716 23156 34717 23220
rect 34651 23155 34717 23156
rect 34928 22336 35248 23360
rect 35390 22677 35450 30363
rect 35387 22676 35453 22677
rect 35387 22612 35388 22676
rect 35452 22612 35453 22676
rect 35387 22611 35453 22612
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34467 22132 34533 22133
rect 34467 22068 34468 22132
rect 34532 22068 34533 22132
rect 34467 22067 34533 22068
rect 34928 21248 35248 22272
rect 35574 21997 35634 34171
rect 35939 33692 36005 33693
rect 35939 33628 35940 33692
rect 36004 33628 36005 33692
rect 35939 33627 36005 33628
rect 35755 31244 35821 31245
rect 35755 31180 35756 31244
rect 35820 31180 35821 31244
rect 35755 31179 35821 31180
rect 35758 28661 35818 31179
rect 35942 30429 36002 33627
rect 35939 30428 36005 30429
rect 35939 30364 35940 30428
rect 36004 30364 36005 30428
rect 35939 30363 36005 30364
rect 35755 28660 35821 28661
rect 35755 28596 35756 28660
rect 35820 28596 35821 28660
rect 35755 28595 35821 28596
rect 35755 28388 35821 28389
rect 35755 28324 35756 28388
rect 35820 28324 35821 28388
rect 35755 28323 35821 28324
rect 35758 24989 35818 28323
rect 35939 28252 36005 28253
rect 35939 28188 35940 28252
rect 36004 28188 36005 28252
rect 35939 28187 36005 28188
rect 35755 24988 35821 24989
rect 35755 24924 35756 24988
rect 35820 24924 35821 24988
rect 35755 24923 35821 24924
rect 35755 24036 35821 24037
rect 35755 23972 35756 24036
rect 35820 23972 35821 24036
rect 35755 23971 35821 23972
rect 35571 21996 35637 21997
rect 35571 21932 35572 21996
rect 35636 21932 35637 21996
rect 35571 21931 35637 21932
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34283 20500 34349 20501
rect 34283 20436 34284 20500
rect 34348 20436 34349 20500
rect 34283 20435 34349 20436
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34283 20092 34349 20093
rect 34283 20028 34284 20092
rect 34348 20028 34349 20092
rect 34283 20027 34349 20028
rect 33915 19684 33981 19685
rect 33915 19620 33916 19684
rect 33980 19620 33981 19684
rect 33915 19619 33981 19620
rect 34286 13429 34346 20027
rect 34928 19072 35248 20096
rect 35758 19413 35818 23971
rect 35942 23221 36002 28187
rect 35939 23220 36005 23221
rect 35939 23156 35940 23220
rect 36004 23156 36005 23220
rect 35939 23155 36005 23156
rect 36126 22110 36186 34851
rect 37043 34644 37109 34645
rect 37043 34580 37044 34644
rect 37108 34580 37109 34644
rect 37043 34579 37109 34580
rect 37046 30701 37106 34579
rect 37043 30700 37109 30701
rect 37043 30636 37044 30700
rect 37108 30636 37109 30700
rect 37043 30635 37109 30636
rect 36307 29340 36373 29341
rect 36307 29276 36308 29340
rect 36372 29276 36373 29340
rect 36307 29275 36373 29276
rect 36310 27165 36370 29275
rect 36307 27164 36373 27165
rect 36307 27100 36308 27164
rect 36372 27100 36373 27164
rect 36307 27099 36373 27100
rect 36310 26210 36370 27099
rect 36310 26150 36554 26210
rect 36126 22050 36370 22110
rect 35755 19412 35821 19413
rect 35755 19350 35756 19412
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 35574 19348 35756 19350
rect 35820 19348 35821 19412
rect 35574 19347 35821 19348
rect 35574 19290 35818 19347
rect 35574 15469 35634 19290
rect 36310 16829 36370 22050
rect 36307 16828 36373 16829
rect 36307 16764 36308 16828
rect 36372 16764 36373 16828
rect 36307 16763 36373 16764
rect 36494 16693 36554 26150
rect 37046 21589 37106 30635
rect 37043 21588 37109 21589
rect 37043 21524 37044 21588
rect 37108 21524 37109 21588
rect 37043 21523 37109 21524
rect 36491 16692 36557 16693
rect 36491 16628 36492 16692
rect 36556 16628 36557 16692
rect 36491 16627 36557 16628
rect 35571 15468 35637 15469
rect 35571 15404 35572 15468
rect 35636 15404 35637 15468
rect 35571 15403 35637 15404
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34283 13428 34349 13429
rect 34283 13364 34284 13428
rect 34348 13364 34349 13428
rect 34283 13363 34349 13364
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 32995 6900 33061 6901
rect 32995 6836 32996 6900
rect 33060 6836 33061 6900
rect 32995 6835 33061 6836
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 32811 2548 32877 2549
rect 32811 2484 32812 2548
rect 32876 2484 32877 2548
rect 32811 2483 32877 2484
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36616 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 4784 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 4140 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 30544 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 4784 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 37536 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 25668 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 4692 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 32752 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 29716 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 28980 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 16928 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 33120 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 33948 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 21252 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 37536 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 3956 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 36800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 3128 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 10580 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 4784 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 5612 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 35512 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 22908 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 5336 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 30176 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1676037725
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_389 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_397
timestamp 1676037725
transform 1 0 37628 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1676037725
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_397
timestamp 1676037725
transform 1 0 37628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1676037725
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1676037725
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_292
timestamp 1676037725
transform 1 0 27968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_307
timestamp 1676037725
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_316
timestamp 1676037725
transform 1 0 30176 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_330
timestamp 1676037725
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1676037725
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1676037725
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_230
timestamp 1676037725
transform 1 0 22264 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_238
timestamp 1676037725
transform 1 0 23000 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_271
timestamp 1676037725
transform 1 0 26036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_288
timestamp 1676037725
transform 1 0 27600 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_315
timestamp 1676037725
transform 1 0 30084 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_325
timestamp 1676037725
transform 1 0 31004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_334
timestamp 1676037725
transform 1 0 31832 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_349
timestamp 1676037725
transform 1 0 33212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 1676037725
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_397
timestamp 1676037725
transform 1 0 37628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1676037725
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_201
timestamp 1676037725
transform 1 0 19596 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1676037725
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_231
timestamp 1676037725
transform 1 0 22356 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_251
timestamp 1676037725
transform 1 0 24196 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_259
timestamp 1676037725
transform 1 0 24932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1676037725
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_309
timestamp 1676037725
transform 1 0 29532 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_355
timestamp 1676037725
transform 1 0 33764 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_367
timestamp 1676037725
transform 1 0 34868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_379
timestamp 1676037725
transform 1 0 35972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1676037725
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1676037725
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_215
timestamp 1676037725
transform 1 0 20884 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_232
timestamp 1676037725
transform 1 0 22448 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_240
timestamp 1676037725
transform 1 0 23184 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_271
timestamp 1676037725
transform 1 0 26036 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_284
timestamp 1676037725
transform 1 0 27232 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1676037725
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_317
timestamp 1676037725
transform 1 0 30268 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_334
timestamp 1676037725
transform 1 0 31832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_354
timestamp 1676037725
transform 1 0 33672 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1676037725
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_376
timestamp 1676037725
transform 1 0 35696 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_388
timestamp 1676037725
transform 1 0 36800 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_396
timestamp 1676037725
transform 1 0 37536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1676037725
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_205
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_211
timestamp 1676037725
transform 1 0 20516 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1676037725
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_236
timestamp 1676037725
transform 1 0 22816 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_246
timestamp 1676037725
transform 1 0 23736 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_268
timestamp 1676037725
transform 1 0 25760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1676037725
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_292
timestamp 1676037725
transform 1 0 27968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_318
timestamp 1676037725
transform 1 0 30360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_331
timestamp 1676037725
transform 1 0 31556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_356
timestamp 1676037725
transform 1 0 33856 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_376
timestamp 1676037725
transform 1 0 35696 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_388
timestamp 1676037725
transform 1 0 36800 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1676037725
transform 1 0 20884 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_228
timestamp 1676037725
transform 1 0 22080 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1676037725
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_268
timestamp 1676037725
transform 1 0 25760 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_286
timestamp 1676037725
transform 1 0 27416 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_316
timestamp 1676037725
transform 1 0 30176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_328
timestamp 1676037725
transform 1 0 31280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_335
timestamp 1676037725
transform 1 0 31924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_339
timestamp 1676037725
transform 1 0 32292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_361
timestamp 1676037725
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_383
timestamp 1676037725
transform 1 0 36340 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_395
timestamp 1676037725
transform 1 0 37444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_212
timestamp 1676037725
transform 1 0 20608 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_240
timestamp 1676037725
transform 1 0 23184 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_253
timestamp 1676037725
transform 1 0 24380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_264
timestamp 1676037725
transform 1 0 25392 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_270
timestamp 1676037725
transform 1 0 25944 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1676037725
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1676037725
transform 1 0 28244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_308
timestamp 1676037725
transform 1 0 29440 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_316
timestamp 1676037725
transform 1 0 30176 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_326
timestamp 1676037725
transform 1 0 31096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_330
timestamp 1676037725
transform 1 0 31464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1676037725
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_360
timestamp 1676037725
transform 1 0 34224 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_373
timestamp 1676037725
transform 1 0 35420 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_380
timestamp 1676037725
transform 1 0 36064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1676037725
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_401
timestamp 1676037725
transform 1 0 37996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_202
timestamp 1676037725
transform 1 0 19688 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1676037725
transform 1 0 20424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1676037725
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_259
timestamp 1676037725
transform 1 0 24932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_272
timestamp 1676037725
transform 1 0 26128 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1676037725
transform 1 0 26496 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1676037725
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1676037725
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_328
timestamp 1676037725
transform 1 0 31280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_334
timestamp 1676037725
transform 1 0 31832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_344
timestamp 1676037725
transform 1 0 32752 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_352
timestamp 1676037725
transform 1 0 33488 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1676037725
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_376
timestamp 1676037725
transform 1 0 35696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_383
timestamp 1676037725
transform 1 0 36340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_390
timestamp 1676037725
transform 1 0 36984 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_397
timestamp 1676037725
transform 1 0 37628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_401
timestamp 1676037725
transform 1 0 37996 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1676037725
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_189
timestamp 1676037725
transform 1 0 18492 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_195
timestamp 1676037725
transform 1 0 19044 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_201
timestamp 1676037725
transform 1 0 19596 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1676037725
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_236
timestamp 1676037725
transform 1 0 22816 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_251
timestamp 1676037725
transform 1 0 24196 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1676037725
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1676037725
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_305
timestamp 1676037725
transform 1 0 29164 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_309
timestamp 1676037725
transform 1 0 29532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_315
timestamp 1676037725
transform 1 0 30084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_327
timestamp 1676037725
transform 1 0 31188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_361
timestamp 1676037725
transform 1 0 34316 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_381
timestamp 1676037725
transform 1 0 36156 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_386
timestamp 1676037725
transform 1 0 36616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1676037725
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_398
timestamp 1676037725
transform 1 0 37720 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1676037725
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_185
timestamp 1676037725
transform 1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_221
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_241
timestamp 1676037725
transform 1 0 23276 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_259
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_268
timestamp 1676037725
transform 1 0 25760 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_288
timestamp 1676037725
transform 1 0 27600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1676037725
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_331
timestamp 1676037725
transform 1 0 31556 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_351
timestamp 1676037725
transform 1 0 33396 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1676037725
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_383
timestamp 1676037725
transform 1 0 36340 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_392
timestamp 1676037725
transform 1 0 37168 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_398
timestamp 1676037725
transform 1 0 37720 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1676037725
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_177
timestamp 1676037725
transform 1 0 17388 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_186
timestamp 1676037725
transform 1 0 18216 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_207
timestamp 1676037725
transform 1 0 20148 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_247
timestamp 1676037725
transform 1 0 23828 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_255
timestamp 1676037725
transform 1 0 24564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1676037725
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1676037725
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_306
timestamp 1676037725
transform 1 0 29256 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_319
timestamp 1676037725
transform 1 0 30452 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1676037725
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_360
timestamp 1676037725
transform 1 0 34224 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_367
timestamp 1676037725
transform 1 0 34868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_376
timestamp 1676037725
transform 1 0 35696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1676037725
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_184
timestamp 1676037725
transform 1 0 18032 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_216
timestamp 1676037725
transform 1 0 20976 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_227
timestamp 1676037725
transform 1 0 21988 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_235
timestamp 1676037725
transform 1 0 22724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1676037725
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_275
timestamp 1676037725
transform 1 0 26404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_281
timestamp 1676037725
transform 1 0 26956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_298
timestamp 1676037725
transform 1 0 28520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_305
timestamp 1676037725
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_327
timestamp 1676037725
transform 1 0 31188 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_337
timestamp 1676037725
transform 1 0 32108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_369
timestamp 1676037725
transform 1 0 35052 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_375
timestamp 1676037725
transform 1 0 35604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_395
timestamp 1676037725
transform 1 0 37444 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1676037725
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp 1676037725
transform 1 0 15180 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_157
timestamp 1676037725
transform 1 0 15548 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_174
timestamp 1676037725
transform 1 0 17112 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_200
timestamp 1676037725
transform 1 0 19504 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1676037725
transform 1 0 20884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_246
timestamp 1676037725
transform 1 0 23736 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_256
timestamp 1676037725
transform 1 0 24656 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1676037725
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_297
timestamp 1676037725
transform 1 0 28428 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_314
timestamp 1676037725
transform 1 0 29992 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_327
timestamp 1676037725
transform 1 0 31188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_348
timestamp 1676037725
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_352
timestamp 1676037725
transform 1 0 33488 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_362
timestamp 1676037725
transform 1 0 34408 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1676037725
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_404
timestamp 1676037725
transform 1 0 38272 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1676037725
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_175
timestamp 1676037725
transform 1 0 17204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1676037725
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_217
timestamp 1676037725
transform 1 0 21068 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_223
timestamp 1676037725
transform 1 0 21620 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_243
timestamp 1676037725
transform 1 0 23460 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_260
timestamp 1676037725
transform 1 0 25024 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_272
timestamp 1676037725
transform 1 0 26128 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_287
timestamp 1676037725
transform 1 0 27508 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_298
timestamp 1676037725
transform 1 0 28520 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1676037725
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_318
timestamp 1676037725
transform 1 0 30360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_322
timestamp 1676037725
transform 1 0 30728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_340
timestamp 1676037725
transform 1 0 32384 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1676037725
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_372
timestamp 1676037725
transform 1 0 35328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_376
timestamp 1676037725
transform 1 0 35696 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_383
timestamp 1676037725
transform 1 0 36340 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_387
timestamp 1676037725
transform 1 0 36708 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_404
timestamp 1676037725
transform 1 0 38272 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_154
timestamp 1676037725
transform 1 0 15272 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1676037725
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1676037725
transform 1 0 17572 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_196
timestamp 1676037725
transform 1 0 19136 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_208
timestamp 1676037725
transform 1 0 20240 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1676037725
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1676037725
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_231
timestamp 1676037725
transform 1 0 22356 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_239
timestamp 1676037725
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_259
timestamp 1676037725
transform 1 0 24932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_272
timestamp 1676037725
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_290
timestamp 1676037725
transform 1 0 27784 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1676037725
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_316
timestamp 1676037725
transform 1 0 30176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_320
timestamp 1676037725
transform 1 0 30544 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1676037725
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1676037725
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_346
timestamp 1676037725
transform 1 0 32936 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_357
timestamp 1676037725
transform 1 0 33948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_368
timestamp 1676037725
transform 1 0 34960 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_380
timestamp 1676037725
transform 1 0 36064 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_390
timestamp 1676037725
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_404
timestamp 1676037725
transform 1 0 38272 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1676037725
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1676037725
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_176
timestamp 1676037725
transform 1 0 17296 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_187
timestamp 1676037725
transform 1 0 18308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_204
timestamp 1676037725
transform 1 0 19872 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_217
timestamp 1676037725
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_226
timestamp 1676037725
transform 1 0 21896 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_240
timestamp 1676037725
transform 1 0 23184 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_259
timestamp 1676037725
transform 1 0 24932 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_267
timestamp 1676037725
transform 1 0 25668 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_279
timestamp 1676037725
transform 1 0 26772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_291
timestamp 1676037725
transform 1 0 27876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1676037725
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_316
timestamp 1676037725
transform 1 0 30176 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_331
timestamp 1676037725
transform 1 0 31556 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_342
timestamp 1676037725
transform 1 0 32568 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1676037725
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_374
timestamp 1676037725
transform 1 0 35512 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_385
timestamp 1676037725
transform 1 0 36524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_405
timestamp 1676037725
transform 1 0 38364 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_145
timestamp 1676037725
transform 1 0 14444 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_158
timestamp 1676037725
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1676037725
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_192
timestamp 1676037725
transform 1 0 18768 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_205
timestamp 1676037725
transform 1 0 19964 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_218
timestamp 1676037725
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_235
timestamp 1676037725
transform 1 0 22724 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_246
timestamp 1676037725
transform 1 0 23736 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_257
timestamp 1676037725
transform 1 0 24748 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_271
timestamp 1676037725
transform 1 0 26036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_291
timestamp 1676037725
transform 1 0 27876 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_299
timestamp 1676037725
transform 1 0 28612 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_308
timestamp 1676037725
transform 1 0 29440 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_319
timestamp 1676037725
transform 1 0 30452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1676037725
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_347
timestamp 1676037725
transform 1 0 33028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_359
timestamp 1676037725
transform 1 0 34132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_365
timestamp 1676037725
transform 1 0 34684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_374
timestamp 1676037725
transform 1 0 35512 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1676037725
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_404
timestamp 1676037725
transform 1 0 38272 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_127
timestamp 1676037725
transform 1 0 12788 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_131
timestamp 1676037725
transform 1 0 13156 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1676037725
transform 1 0 14444 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1676037725
transform 1 0 15088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_160
timestamp 1676037725
transform 1 0 15824 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_206
timestamp 1676037725
transform 1 0 20056 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_210
timestamp 1676037725
transform 1 0 20424 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1676037725
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_227
timestamp 1676037725
transform 1 0 21988 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_241
timestamp 1676037725
transform 1 0 23276 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_268
timestamp 1676037725
transform 1 0 25760 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_274
timestamp 1676037725
transform 1 0 26312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_286
timestamp 1676037725
transform 1 0 27416 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_290
timestamp 1676037725
transform 1 0 27784 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_298
timestamp 1676037725
transform 1 0 28520 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_320
timestamp 1676037725
transform 1 0 30544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_334
timestamp 1676037725
transform 1 0 31832 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_350
timestamp 1676037725
transform 1 0 33304 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_354
timestamp 1676037725
transform 1 0 33672 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1676037725
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_375
timestamp 1676037725
transform 1 0 35604 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_383
timestamp 1676037725
transform 1 0 36340 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_402
timestamp 1676037725
transform 1 0 38088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1676037725
transform 1 0 38456 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_121
timestamp 1676037725
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_142
timestamp 1676037725
transform 1 0 14168 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_155
timestamp 1676037725
transform 1 0 15364 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_159
timestamp 1676037725
transform 1 0 15732 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_177
timestamp 1676037725
transform 1 0 17388 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_190
timestamp 1676037725
transform 1 0 18584 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_203
timestamp 1676037725
transform 1 0 19780 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_211
timestamp 1676037725
transform 1 0 20516 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_233
timestamp 1676037725
transform 1 0 22540 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_245
timestamp 1676037725
transform 1 0 23644 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_251
timestamp 1676037725
transform 1 0 24196 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_259
timestamp 1676037725
transform 1 0 24932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_266
timestamp 1676037725
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_291
timestamp 1676037725
transform 1 0 27876 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_306
timestamp 1676037725
transform 1 0 29256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_317
timestamp 1676037725
transform 1 0 30268 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_323
timestamp 1676037725
transform 1 0 30820 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_331
timestamp 1676037725
transform 1 0 31556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1676037725
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_353
timestamp 1676037725
transform 1 0 33580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_373
timestamp 1676037725
transform 1 0 35420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_383
timestamp 1676037725
transform 1 0 36340 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1676037725
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_126
timestamp 1676037725
transform 1 0 12696 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 1676037725
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_167
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_177
timestamp 1676037725
transform 1 0 17388 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1676037725
transform 1 0 20056 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_218
timestamp 1676037725
transform 1 0 21160 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_233
timestamp 1676037725
transform 1 0 22540 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_242
timestamp 1676037725
transform 1 0 23368 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_268
timestamp 1676037725
transform 1 0 25760 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_300
timestamp 1676037725
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_328
timestamp 1676037725
transform 1 0 31280 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_336
timestamp 1676037725
transform 1 0 32016 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_345
timestamp 1676037725
transform 1 0 32844 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_358
timestamp 1676037725
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_376
timestamp 1676037725
transform 1 0 35696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_385
timestamp 1676037725
transform 1 0 36524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1676037725
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1676037725
transform 1 0 12236 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_148
timestamp 1676037725
transform 1 0 14720 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_158
timestamp 1676037725
transform 1 0 15640 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_176
timestamp 1676037725
transform 1 0 17296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_184
timestamp 1676037725
transform 1 0 18032 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_202
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_215
timestamp 1676037725
transform 1 0 20884 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_244
timestamp 1676037725
transform 1 0 23552 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_248
timestamp 1676037725
transform 1 0 23920 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_257
timestamp 1676037725
transform 1 0 24748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1676037725
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1676037725
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1676037725
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_300
timestamp 1676037725
transform 1 0 28704 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_311
timestamp 1676037725
transform 1 0 29716 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_324
timestamp 1676037725
transform 1 0 30912 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1676037725
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_348
timestamp 1676037725
transform 1 0 33120 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_361
timestamp 1676037725
transform 1 0 34316 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_371
timestamp 1676037725
transform 1 0 35236 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_382
timestamp 1676037725
transform 1 0 36248 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1676037725
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_404
timestamp 1676037725
transform 1 0 38272 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_126
timestamp 1676037725
transform 1 0 12696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_137
timestamp 1676037725
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_152
timestamp 1676037725
transform 1 0 15088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_175
timestamp 1676037725
transform 1 0 17204 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_183
timestamp 1676037725
transform 1 0 17940 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_216
timestamp 1676037725
transform 1 0 20976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_224
timestamp 1676037725
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1676037725
transform 1 0 22632 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1676037725
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_264
timestamp 1676037725
transform 1 0 25392 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_273
timestamp 1676037725
transform 1 0 26220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_282
timestamp 1676037725
transform 1 0 27048 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_291
timestamp 1676037725
transform 1 0 27876 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_322
timestamp 1676037725
transform 1 0 30728 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_330
timestamp 1676037725
transform 1 0 31464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_342
timestamp 1676037725
transform 1 0 32568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_354
timestamp 1676037725
transform 1 0 33672 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1676037725
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_378
timestamp 1676037725
transform 1 0 35880 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_399
timestamp 1676037725
transform 1 0 37812 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_138
timestamp 1676037725
transform 1 0 13800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1676037725
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_177
timestamp 1676037725
transform 1 0 17388 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1676037725
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1676037725
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_214
timestamp 1676037725
transform 1 0 20792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_235
timestamp 1676037725
transform 1 0 22724 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_243
timestamp 1676037725
transform 1 0 23460 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_251
timestamp 1676037725
transform 1 0 24196 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_261
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_269
timestamp 1676037725
transform 1 0 25852 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_289
timestamp 1676037725
transform 1 0 27692 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_300
timestamp 1676037725
transform 1 0 28704 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_311
timestamp 1676037725
transform 1 0 29716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_319
timestamp 1676037725
transform 1 0 30452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_330
timestamp 1676037725
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_346
timestamp 1676037725
transform 1 0 32936 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_356
timestamp 1676037725
transform 1 0 33856 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_362
timestamp 1676037725
transform 1 0 34408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_371
timestamp 1676037725
transform 1 0 35236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_380
timestamp 1676037725
transform 1 0 36064 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1676037725
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_404
timestamp 1676037725
transform 1 0 38272 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_105
timestamp 1676037725
transform 1 0 10764 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_123
timestamp 1676037725
transform 1 0 12420 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_147
timestamp 1676037725
transform 1 0 14628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_155
timestamp 1676037725
transform 1 0 15364 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_178
timestamp 1676037725
transform 1 0 17480 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_186
timestamp 1676037725
transform 1 0 18216 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_205
timestamp 1676037725
transform 1 0 19964 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_212
timestamp 1676037725
transform 1 0 20608 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_216
timestamp 1676037725
transform 1 0 20976 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_230
timestamp 1676037725
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_243
timestamp 1676037725
transform 1 0 23460 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_261
timestamp 1676037725
transform 1 0 25116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_269
timestamp 1676037725
transform 1 0 25852 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_277
timestamp 1676037725
transform 1 0 26588 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_291
timestamp 1676037725
transform 1 0 27876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1676037725
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_316
timestamp 1676037725
transform 1 0 30176 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_324
timestamp 1676037725
transform 1 0 30912 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_333
timestamp 1676037725
transform 1 0 31740 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_345
timestamp 1676037725
transform 1 0 32844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1676037725
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1676037725
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_375
timestamp 1676037725
transform 1 0 35604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_385
timestamp 1676037725
transform 1 0 36524 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1676037725
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_144
timestamp 1676037725
transform 1 0 14352 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_159
timestamp 1676037725
transform 1 0 15732 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_173
timestamp 1676037725
transform 1 0 17020 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_182
timestamp 1676037725
transform 1 0 17848 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_214
timestamp 1676037725
transform 1 0 20792 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_218
timestamp 1676037725
transform 1 0 21160 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_240
timestamp 1676037725
transform 1 0 23184 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_250
timestamp 1676037725
transform 1 0 24104 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_258
timestamp 1676037725
transform 1 0 24840 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_266
timestamp 1676037725
transform 1 0 25576 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_291
timestamp 1676037725
transform 1 0 27876 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_300
timestamp 1676037725
transform 1 0 28704 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_309
timestamp 1676037725
transform 1 0 29532 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1676037725
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_350
timestamp 1676037725
transform 1 0 33304 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_362
timestamp 1676037725
transform 1 0 34408 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_377
timestamp 1676037725
transform 1 0 35788 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1676037725
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_401
timestamp 1676037725
transform 1 0 37996 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_128
timestamp 1676037725
transform 1 0 12880 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_174
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_205
timestamp 1676037725
transform 1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_229
timestamp 1676037725
transform 1 0 22172 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_239
timestamp 1676037725
transform 1 0 23092 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_268
timestamp 1676037725
transform 1 0 25760 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_279
timestamp 1676037725
transform 1 0 26772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_289
timestamp 1676037725
transform 1 0 27692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_298
timestamp 1676037725
transform 1 0 28520 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1676037725
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_319
timestamp 1676037725
transform 1 0 30452 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_327
timestamp 1676037725
transform 1 0 31188 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_340
timestamp 1676037725
transform 1 0 32384 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_352
timestamp 1676037725
transform 1 0 33488 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1676037725
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_375
timestamp 1676037725
transform 1 0 35604 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_398
timestamp 1676037725
transform 1 0 37720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_405
timestamp 1676037725
transform 1 0 38364 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_89
timestamp 1676037725
transform 1 0 9292 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_107
timestamp 1676037725
transform 1 0 10948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_117
timestamp 1676037725
transform 1 0 11868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_127
timestamp 1676037725
transform 1 0 12788 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_133
timestamp 1676037725
transform 1 0 13340 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_151
timestamp 1676037725
transform 1 0 14996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_162
timestamp 1676037725
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_173
timestamp 1676037725
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_177
timestamp 1676037725
transform 1 0 17388 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_190
timestamp 1676037725
transform 1 0 18584 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_198
timestamp 1676037725
transform 1 0 19320 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_216
timestamp 1676037725
transform 1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_232
timestamp 1676037725
transform 1 0 22448 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_256
timestamp 1676037725
transform 1 0 24656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1676037725
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_289
timestamp 1676037725
transform 1 0 27692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_297
timestamp 1676037725
transform 1 0 28428 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_307
timestamp 1676037725
transform 1 0 29348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_319
timestamp 1676037725
transform 1 0 30452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_330
timestamp 1676037725
transform 1 0 31464 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_352
timestamp 1676037725
transform 1 0 33488 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_364
timestamp 1676037725
transform 1 0 34592 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_376
timestamp 1676037725
transform 1 0 35696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_387
timestamp 1676037725
transform 1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1676037725
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_404
timestamp 1676037725
transform 1 0 38272 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_121
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_129
timestamp 1676037725
transform 1 0 12972 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_147
timestamp 1676037725
transform 1 0 14628 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_167
timestamp 1676037725
transform 1 0 16468 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_180
timestamp 1676037725
transform 1 0 17664 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_184
timestamp 1676037725
transform 1 0 18032 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_217
timestamp 1676037725
transform 1 0 21068 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_235
timestamp 1676037725
transform 1 0 22724 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1676037725
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_263
timestamp 1676037725
transform 1 0 25300 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_280
timestamp 1676037725
transform 1 0 26864 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_298
timestamp 1676037725
transform 1 0 28520 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1676037725
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_318
timestamp 1676037725
transform 1 0 30360 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_326
timestamp 1676037725
transform 1 0 31096 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_337
timestamp 1676037725
transform 1 0 32108 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_346
timestamp 1676037725
transform 1 0 32936 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1676037725
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_371
timestamp 1676037725
transform 1 0 35236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_382
timestamp 1676037725
transform 1 0 36248 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_388
timestamp 1676037725
transform 1 0 36800 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1676037725
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1676037725
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1676037725
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_122
timestamp 1676037725
transform 1 0 12328 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_144
timestamp 1676037725
transform 1 0 14352 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_157
timestamp 1676037725
transform 1 0 15548 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1676037725
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_174
timestamp 1676037725
transform 1 0 17112 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_185
timestamp 1676037725
transform 1 0 18124 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_207
timestamp 1676037725
transform 1 0 20148 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1676037725
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_243
timestamp 1676037725
transform 1 0 23460 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_247
timestamp 1676037725
transform 1 0 23828 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_264
timestamp 1676037725
transform 1 0 25392 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1676037725
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_285
timestamp 1676037725
transform 1 0 27324 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_301
timestamp 1676037725
transform 1 0 28796 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_305
timestamp 1676037725
transform 1 0 29164 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_314
timestamp 1676037725
transform 1 0 29992 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_322
timestamp 1676037725
transform 1 0 30728 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 1676037725
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_347
timestamp 1676037725
transform 1 0 33028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_359
timestamp 1676037725
transform 1 0 34132 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_363
timestamp 1676037725
transform 1 0 34500 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_372
timestamp 1676037725
transform 1 0 35328 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_384
timestamp 1676037725
transform 1 0 36432 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_404
timestamp 1676037725
transform 1 0 38272 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_96
timestamp 1676037725
transform 1 0 9936 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_100
timestamp 1676037725
transform 1 0 10304 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_104
timestamp 1676037725
transform 1 0 10672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_112
timestamp 1676037725
transform 1 0 11408 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_116
timestamp 1676037725
transform 1 0 11776 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_128
timestamp 1676037725
transform 1 0 12880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 1676037725
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_147
timestamp 1676037725
transform 1 0 14628 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_158
timestamp 1676037725
transform 1 0 15640 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_166
timestamp 1676037725
transform 1 0 16376 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_174
timestamp 1676037725
transform 1 0 17112 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_187
timestamp 1676037725
transform 1 0 18308 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_206
timestamp 1676037725
transform 1 0 20056 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_214
timestamp 1676037725
transform 1 0 20792 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_225
timestamp 1676037725
transform 1 0 21804 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_236
timestamp 1676037725
transform 1 0 22816 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_242
timestamp 1676037725
transform 1 0 23368 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1676037725
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_262
timestamp 1676037725
transform 1 0 25208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_271
timestamp 1676037725
transform 1 0 26036 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_280
timestamp 1676037725
transform 1 0 26864 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_290
timestamp 1676037725
transform 1 0 27784 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1676037725
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1676037725
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_318
timestamp 1676037725
transform 1 0 30360 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_329
timestamp 1676037725
transform 1 0 31372 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_348
timestamp 1676037725
transform 1 0 33120 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1676037725
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_374
timestamp 1676037725
transform 1 0 35512 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_385
timestamp 1676037725
transform 1 0 36524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1676037725
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_77
timestamp 1676037725
transform 1 0 8188 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_95
timestamp 1676037725
transform 1 0 9844 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1676037725
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_131
timestamp 1676037725
transform 1 0 13156 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_138
timestamp 1676037725
transform 1 0 13800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_145
timestamp 1676037725
transform 1 0 14444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1676037725
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_183
timestamp 1676037725
transform 1 0 17940 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_187
timestamp 1676037725
transform 1 0 18308 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_202
timestamp 1676037725
transform 1 0 19688 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_211
timestamp 1676037725
transform 1 0 20516 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1676037725
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_231
timestamp 1676037725
transform 1 0 22356 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_242
timestamp 1676037725
transform 1 0 23368 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_252
timestamp 1676037725
transform 1 0 24288 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_269
timestamp 1676037725
transform 1 0 25852 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1676037725
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_297
timestamp 1676037725
transform 1 0 28428 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_308
timestamp 1676037725
transform 1 0 29440 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1676037725
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1676037725
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_351
timestamp 1676037725
transform 1 0 33396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_364
timestamp 1676037725
transform 1 0 34592 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_372
timestamp 1676037725
transform 1 0 35328 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1676037725
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_404
timestamp 1676037725
transform 1 0 38272 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_93
timestamp 1676037725
transform 1 0 9660 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_112
timestamp 1676037725
transform 1 0 11408 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_132
timestamp 1676037725
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_147
timestamp 1676037725
transform 1 0 14628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_155
timestamp 1676037725
transform 1 0 15364 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_175
timestamp 1676037725
transform 1 0 17204 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_179
timestamp 1676037725
transform 1 0 17572 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_185
timestamp 1676037725
transform 1 0 18124 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1676037725
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_213
timestamp 1676037725
transform 1 0 20700 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_228
timestamp 1676037725
transform 1 0 22080 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1676037725
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_263
timestamp 1676037725
transform 1 0 25300 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_271
timestamp 1676037725
transform 1 0 26036 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_281
timestamp 1676037725
transform 1 0 26956 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_289
timestamp 1676037725
transform 1 0 27692 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_299
timestamp 1676037725
transform 1 0 28612 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1676037725
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_316
timestamp 1676037725
transform 1 0 30176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_328
timestamp 1676037725
transform 1 0 31280 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_337
timestamp 1676037725
transform 1 0 32108 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_352
timestamp 1676037725
transform 1 0 33488 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1676037725
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_374
timestamp 1676037725
transform 1 0 35512 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_385
timestamp 1676037725
transform 1 0 36524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1676037725
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_84
timestamp 1676037725
transform 1 0 8832 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_99
timestamp 1676037725
transform 1 0 10212 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1676037725
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_127
timestamp 1676037725
transform 1 0 12788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_131
timestamp 1676037725
transform 1 0 13156 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_135
timestamp 1676037725
transform 1 0 13524 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_155
timestamp 1676037725
transform 1 0 15364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1676037725
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_189
timestamp 1676037725
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_200
timestamp 1676037725
transform 1 0 19504 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_216
timestamp 1676037725
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_238
timestamp 1676037725
transform 1 0 23000 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_247
timestamp 1676037725
transform 1 0 23828 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_258
timestamp 1676037725
transform 1 0 24840 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_264
timestamp 1676037725
transform 1 0 25392 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1676037725
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_291
timestamp 1676037725
transform 1 0 27876 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_313
timestamp 1676037725
transform 1 0 29900 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_321
timestamp 1676037725
transform 1 0 30636 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_330
timestamp 1676037725
transform 1 0 31464 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_341
timestamp 1676037725
transform 1 0 32476 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_351
timestamp 1676037725
transform 1 0 33396 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_364
timestamp 1676037725
transform 1 0 34592 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_375
timestamp 1676037725
transform 1 0 35604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_386
timestamp 1676037725
transform 1 0 36616 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_404
timestamp 1676037725
transform 1 0 38272 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1676037725
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_90
timestamp 1676037725
transform 1 0 9384 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_99
timestamp 1676037725
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_122
timestamp 1676037725
transform 1 0 12328 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_150
timestamp 1676037725
transform 1 0 14904 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_174
timestamp 1676037725
transform 1 0 17112 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_191
timestamp 1676037725
transform 1 0 18676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_218
timestamp 1676037725
transform 1 0 21160 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_224
timestamp 1676037725
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_234
timestamp 1676037725
transform 1 0 22632 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_243
timestamp 1676037725
transform 1 0 23460 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_263
timestamp 1676037725
transform 1 0 25300 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_277
timestamp 1676037725
transform 1 0 26588 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_285
timestamp 1676037725
transform 1 0 27324 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_294
timestamp 1676037725
transform 1 0 28152 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1676037725
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_324
timestamp 1676037725
transform 1 0 30912 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_328
timestamp 1676037725
transform 1 0 31280 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_340
timestamp 1676037725
transform 1 0 32384 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_355
timestamp 1676037725
transform 1 0 33764 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1676037725
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_375
timestamp 1676037725
transform 1 0 35604 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_383
timestamp 1676037725
transform 1 0 36340 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_404
timestamp 1676037725
transform 1 0 38272 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_84
timestamp 1676037725
transform 1 0 8832 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_98
timestamp 1676037725
transform 1 0 10120 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1676037725
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_124
timestamp 1676037725
transform 1 0 12512 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_144
timestamp 1676037725
transform 1 0 14352 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_151
timestamp 1676037725
transform 1 0 14996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_162
timestamp 1676037725
transform 1 0 16008 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_174
timestamp 1676037725
transform 1 0 17112 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_187
timestamp 1676037725
transform 1 0 18308 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_200
timestamp 1676037725
transform 1 0 19504 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1676037725
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1676037725
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1676037725
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_247
timestamp 1676037725
transform 1 0 23828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_253
timestamp 1676037725
transform 1 0 24380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_260
timestamp 1676037725
transform 1 0 25024 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1676037725
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1676037725
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_299
timestamp 1676037725
transform 1 0 28612 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_312
timestamp 1676037725
transform 1 0 29808 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1676037725
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_350
timestamp 1676037725
transform 1 0 33304 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_363
timestamp 1676037725
transform 1 0 34500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_370
timestamp 1676037725
transform 1 0 35144 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_390
timestamp 1676037725
transform 1 0 36984 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_404
timestamp 1676037725
transform 1 0 38272 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1676037725
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_94
timestamp 1676037725
transform 1 0 9752 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_100
timestamp 1676037725
transform 1 0 10304 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_108
timestamp 1676037725
transform 1 0 11040 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_119
timestamp 1676037725
transform 1 0 12052 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_130
timestamp 1676037725
transform 1 0 13064 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1676037725
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_154
timestamp 1676037725
transform 1 0 15272 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_174
timestamp 1676037725
transform 1 0 17112 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_187
timestamp 1676037725
transform 1 0 18308 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1676037725
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1676037725
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_219
timestamp 1676037725
transform 1 0 21252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_225
timestamp 1676037725
transform 1 0 21804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_243
timestamp 1676037725
transform 1 0 23460 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1676037725
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_264
timestamp 1676037725
transform 1 0 25392 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_268
timestamp 1676037725
transform 1 0 25760 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_275
timestamp 1676037725
transform 1 0 26404 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_284
timestamp 1676037725
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_294
timestamp 1676037725
transform 1 0 28152 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_298
timestamp 1676037725
transform 1 0 28520 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1676037725
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_327
timestamp 1676037725
transform 1 0 31188 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_347
timestamp 1676037725
transform 1 0 33028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1676037725
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_383
timestamp 1676037725
transform 1 0 36340 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_387
timestamp 1676037725
transform 1 0 36708 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_405
timestamp 1676037725
transform 1 0 38364 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_65
timestamp 1676037725
transform 1 0 7084 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_70
timestamp 1676037725
transform 1 0 7544 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_77
timestamp 1676037725
transform 1 0 8188 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_84
timestamp 1676037725
transform 1 0 8832 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_95
timestamp 1676037725
transform 1 0 9844 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1676037725
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_117
timestamp 1676037725
transform 1 0 11868 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_124
timestamp 1676037725
transform 1 0 12512 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_132
timestamp 1676037725
transform 1 0 13248 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_152
timestamp 1676037725
transform 1 0 15088 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_163
timestamp 1676037725
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_177
timestamp 1676037725
transform 1 0 17388 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_191
timestamp 1676037725
transform 1 0 18676 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_195
timestamp 1676037725
transform 1 0 19044 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_212
timestamp 1676037725
transform 1 0 20608 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1676037725
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_236
timestamp 1676037725
transform 1 0 22816 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_244
timestamp 1676037725
transform 1 0 23552 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_252
timestamp 1676037725
transform 1 0 24288 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_264
timestamp 1676037725
transform 1 0 25392 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_269
timestamp 1676037725
transform 1 0 25852 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1676037725
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_288
timestamp 1676037725
transform 1 0 27600 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_299
timestamp 1676037725
transform 1 0 28612 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_303
timestamp 1676037725
transform 1 0 28980 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_312
timestamp 1676037725
transform 1 0 29808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_324
timestamp 1676037725
transform 1 0 30912 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1676037725
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_350
timestamp 1676037725
transform 1 0 33304 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_362
timestamp 1676037725
transform 1 0 34408 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_373
timestamp 1676037725
transform 1 0 35420 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1676037725
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_404
timestamp 1676037725
transform 1 0 38272 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_61
timestamp 1676037725
transform 1 0 6716 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_72
timestamp 1676037725
transform 1 0 7728 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1676037725
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_95
timestamp 1676037725
transform 1 0 9844 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_107
timestamp 1676037725
transform 1 0 10948 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_111
timestamp 1676037725
transform 1 0 11316 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_119
timestamp 1676037725
transform 1 0 12052 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_128
timestamp 1676037725
transform 1 0 12880 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_132
timestamp 1676037725
transform 1 0 13248 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1676037725
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_154
timestamp 1676037725
transform 1 0 15272 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_173
timestamp 1676037725
transform 1 0 17020 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_191
timestamp 1676037725
transform 1 0 18676 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_210
timestamp 1676037725
transform 1 0 20424 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_237
timestamp 1676037725
transform 1 0 22908 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1676037725
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_264
timestamp 1676037725
transform 1 0 25392 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_270
timestamp 1676037725
transform 1 0 25944 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_281
timestamp 1676037725
transform 1 0 26956 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_291
timestamp 1676037725
transform 1 0 27876 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1676037725
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_313
timestamp 1676037725
transform 1 0 29900 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_323
timestamp 1676037725
transform 1 0 30820 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_343
timestamp 1676037725
transform 1 0 32660 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_355
timestamp 1676037725
transform 1 0 33764 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1676037725
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_372
timestamp 1676037725
transform 1 0 35328 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_384
timestamp 1676037725
transform 1 0 36432 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1676037725
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_64
timestamp 1676037725
transform 1 0 6992 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_84
timestamp 1676037725
transform 1 0 8832 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_99
timestamp 1676037725
transform 1 0 10212 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1676037725
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_118
timestamp 1676037725
transform 1 0 11960 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_129
timestamp 1676037725
transform 1 0 12972 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_139
timestamp 1676037725
transform 1 0 13892 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_146
timestamp 1676037725
transform 1 0 14536 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1676037725
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_178
timestamp 1676037725
transform 1 0 17480 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_184
timestamp 1676037725
transform 1 0 18032 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_204
timestamp 1676037725
transform 1 0 19872 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_244
timestamp 1676037725
transform 1 0 23552 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_251
timestamp 1676037725
transform 1 0 24196 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_262
timestamp 1676037725
transform 1 0 25208 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_272
timestamp 1676037725
transform 1 0 26128 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_290
timestamp 1676037725
transform 1 0 27784 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_305
timestamp 1676037725
transform 1 0 29164 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_321
timestamp 1676037725
transform 1 0 30636 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1676037725
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_348
timestamp 1676037725
transform 1 0 33120 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_361
timestamp 1676037725
transform 1 0 34316 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1676037725
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_404
timestamp 1676037725
transform 1 0 38272 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_37
timestamp 1676037725
transform 1 0 4508 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_42
timestamp 1676037725
transform 1 0 4968 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_47
timestamp 1676037725
transform 1 0 5428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_54
timestamp 1676037725
transform 1 0 6072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_62
timestamp 1676037725
transform 1 0 6808 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1676037725
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_93
timestamp 1676037725
transform 1 0 9660 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_106
timestamp 1676037725
transform 1 0 10856 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_110
timestamp 1676037725
transform 1 0 11224 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_116
timestamp 1676037725
transform 1 0 11776 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_125
timestamp 1676037725
transform 1 0 12604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_137
timestamp 1676037725
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_150
timestamp 1676037725
transform 1 0 14904 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_159
timestamp 1676037725
transform 1 0 15732 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_179
timestamp 1676037725
transform 1 0 17572 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1676037725
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_203
timestamp 1676037725
transform 1 0 19780 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_216
timestamp 1676037725
transform 1 0 20976 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_222
timestamp 1676037725
transform 1 0 21528 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_230
timestamp 1676037725
transform 1 0 22264 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1676037725
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_264
timestamp 1676037725
transform 1 0 25392 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_275
timestamp 1676037725
transform 1 0 26404 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_289
timestamp 1676037725
transform 1 0 27692 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1676037725
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_320
timestamp 1676037725
transform 1 0 30544 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_340
timestamp 1676037725
transform 1 0 32384 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_352
timestamp 1676037725
transform 1 0 33488 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1676037725
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_374
timestamp 1676037725
transform 1 0 35512 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_386
timestamp 1676037725
transform 1 0 36616 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_397
timestamp 1676037725
transform 1 0 37628 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1676037725
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_43
timestamp 1676037725
transform 1 0 5060 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_47
timestamp 1676037725
transform 1 0 5428 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1676037725
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_63
timestamp 1676037725
transform 1 0 6900 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_78
timestamp 1676037725
transform 1 0 8280 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_87
timestamp 1676037725
transform 1 0 9108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_99
timestamp 1676037725
transform 1 0 10212 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1676037725
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_119
timestamp 1676037725
transform 1 0 12052 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_129
timestamp 1676037725
transform 1 0 12972 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_143
timestamp 1676037725
transform 1 0 14260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_158
timestamp 1676037725
transform 1 0 15640 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1676037725
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_177
timestamp 1676037725
transform 1 0 17388 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_201
timestamp 1676037725
transform 1 0 19596 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 1676037725
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_231
timestamp 1676037725
transform 1 0 22356 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_237
timestamp 1676037725
transform 1 0 22908 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_257
timestamp 1676037725
transform 1 0 24748 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_263
timestamp 1676037725
transform 1 0 25300 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1676037725
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1676037725
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_289
timestamp 1676037725
transform 1 0 27692 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_313
timestamp 1676037725
transform 1 0 29900 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_321
timestamp 1676037725
transform 1 0 30636 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1676037725
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_353
timestamp 1676037725
transform 1 0 33580 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_365
timestamp 1676037725
transform 1 0 34684 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_376
timestamp 1676037725
transform 1 0 35696 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_380
timestamp 1676037725
transform 1 0 36064 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1676037725
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_404
timestamp 1676037725
transform 1 0 38272 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_38
timestamp 1676037725
transform 1 0 4600 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_42
timestamp 1676037725
transform 1 0 4968 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_47
timestamp 1676037725
transform 1 0 5428 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_54
timestamp 1676037725
transform 1 0 6072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_63
timestamp 1676037725
transform 1 0 6900 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_72
timestamp 1676037725
transform 1 0 7728 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1676037725
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_95
timestamp 1676037725
transform 1 0 9844 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_108
timestamp 1676037725
transform 1 0 11040 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_112
timestamp 1676037725
transform 1 0 11408 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_118
timestamp 1676037725
transform 1 0 11960 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1676037725
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_146
timestamp 1676037725
transform 1 0 14536 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_156
timestamp 1676037725
transform 1 0 15456 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_162
timestamp 1676037725
transform 1 0 16008 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_168
timestamp 1676037725
transform 1 0 16560 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1676037725
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_210
timestamp 1676037725
transform 1 0 20424 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_225
timestamp 1676037725
transform 1 0 21804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_231
timestamp 1676037725
transform 1 0 22356 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_242
timestamp 1676037725
transform 1 0 23368 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1676037725
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_264
timestamp 1676037725
transform 1 0 25392 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_279
timestamp 1676037725
transform 1 0 26772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_285
timestamp 1676037725
transform 1 0 27324 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_292
timestamp 1676037725
transform 1 0 27968 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1676037725
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_320
timestamp 1676037725
transform 1 0 30544 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_342
timestamp 1676037725
transform 1 0 32568 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_354
timestamp 1676037725
transform 1 0 33672 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 1676037725
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_384
timestamp 1676037725
transform 1 0 36432 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1676037725
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_31
timestamp 1676037725
transform 1 0 3956 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_35
timestamp 1676037725
transform 1 0 4324 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_42
timestamp 1676037725
transform 1 0 4968 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_50
timestamp 1676037725
transform 1 0 5704 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1676037725
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_66
timestamp 1676037725
transform 1 0 7176 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_87
timestamp 1676037725
transform 1 0 9108 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_101
timestamp 1676037725
transform 1 0 10396 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1676037725
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_122
timestamp 1676037725
transform 1 0 12328 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_134
timestamp 1676037725
transform 1 0 13432 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_147
timestamp 1676037725
transform 1 0 14628 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_160
timestamp 1676037725
transform 1 0 15824 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_177
timestamp 1676037725
transform 1 0 17388 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_188
timestamp 1676037725
transform 1 0 18400 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_196
timestamp 1676037725
transform 1 0 19136 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_203
timestamp 1676037725
transform 1 0 19780 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_210
timestamp 1676037725
transform 1 0 20424 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1676037725
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_229
timestamp 1676037725
transform 1 0 22172 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_238
timestamp 1676037725
transform 1 0 23000 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_246
timestamp 1676037725
transform 1 0 23736 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_253
timestamp 1676037725
transform 1 0 24380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_267
timestamp 1676037725
transform 1 0 25668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_271
timestamp 1676037725
transform 1 0 26036 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1676037725
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_287
timestamp 1676037725
transform 1 0 27508 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_294
timestamp 1676037725
transform 1 0 28152 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_307
timestamp 1676037725
transform 1 0 29348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_317
timestamp 1676037725
transform 1 0 30268 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1676037725
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_342
timestamp 1676037725
transform 1 0 32568 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_352
timestamp 1676037725
transform 1 0 33488 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_363
timestamp 1676037725
transform 1 0 34500 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_374
timestamp 1676037725
transform 1 0 35512 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1676037725
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1676037725
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_404
timestamp 1676037725
transform 1 0 38272 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_40
timestamp 1676037725
transform 1 0 4784 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_47
timestamp 1676037725
transform 1 0 5428 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_54
timestamp 1676037725
transform 1 0 6072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_58
timestamp 1676037725
transform 1 0 6440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_63
timestamp 1676037725
transform 1 0 6900 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_72
timestamp 1676037725
transform 1 0 7728 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1676037725
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_94
timestamp 1676037725
transform 1 0 9752 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_100
timestamp 1676037725
transform 1 0 10304 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_107
timestamp 1676037725
transform 1 0 10948 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_118
timestamp 1676037725
transform 1 0 11960 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_128
timestamp 1676037725
transform 1 0 12880 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1676037725
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_148
timestamp 1676037725
transform 1 0 14720 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_158
timestamp 1676037725
transform 1 0 15640 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_168
timestamp 1676037725
transform 1 0 16560 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_172
timestamp 1676037725
transform 1 0 16928 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_180
timestamp 1676037725
transform 1 0 17664 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_190
timestamp 1676037725
transform 1 0 18584 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_210
timestamp 1676037725
transform 1 0 20424 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_217
timestamp 1676037725
transform 1 0 21068 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_227
timestamp 1676037725
transform 1 0 21988 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_237
timestamp 1676037725
transform 1 0 22908 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_243
timestamp 1676037725
transform 1 0 23460 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1676037725
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_263
timestamp 1676037725
transform 1 0 25300 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_269
timestamp 1676037725
transform 1 0 25852 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_277
timestamp 1676037725
transform 1 0 26588 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_285
timestamp 1676037725
transform 1 0 27324 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_292
timestamp 1676037725
transform 1 0 27968 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1676037725
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_322
timestamp 1676037725
transform 1 0 30728 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_342
timestamp 1676037725
transform 1 0 32568 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_354
timestamp 1676037725
transform 1 0 33672 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1676037725
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_370
timestamp 1676037725
transform 1 0 35144 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_382
timestamp 1676037725
transform 1 0 36248 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1676037725
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_33
timestamp 1676037725
transform 1 0 4140 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_38
timestamp 1676037725
transform 1 0 4600 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_42
timestamp 1676037725
transform 1 0 4968 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_47
timestamp 1676037725
transform 1 0 5428 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1676037725
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_61
timestamp 1676037725
transform 1 0 6716 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_67
timestamp 1676037725
transform 1 0 7268 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_88
timestamp 1676037725
transform 1 0 9200 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_101
timestamp 1676037725
transform 1 0 10396 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1676037725
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_119
timestamp 1676037725
transform 1 0 12052 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_130
timestamp 1676037725
transform 1 0 13064 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_134
timestamp 1676037725
transform 1 0 13432 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_142
timestamp 1676037725
transform 1 0 14168 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_150
timestamp 1676037725
transform 1 0 14904 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_194
timestamp 1676037725
transform 1 0 18952 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_202
timestamp 1676037725
transform 1 0 19688 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_209
timestamp 1676037725
transform 1 0 20332 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_215
timestamp 1676037725
transform 1 0 20884 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1676037725
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_236
timestamp 1676037725
transform 1 0 22816 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_244
timestamp 1676037725
transform 1 0 23552 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_251
timestamp 1676037725
transform 1 0 24196 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_263
timestamp 1676037725
transform 1 0 25300 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 1676037725
transform 1 0 26404 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1676037725
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_289
timestamp 1676037725
transform 1 0 27692 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_300
timestamp 1676037725
transform 1 0 28704 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_306
timestamp 1676037725
transform 1 0 29256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_314
timestamp 1676037725
transform 1 0 29992 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_318
timestamp 1676037725
transform 1 0 30360 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_328
timestamp 1676037725
transform 1 0 31280 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_353
timestamp 1676037725
transform 1 0 33580 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_365
timestamp 1676037725
transform 1 0 34684 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_376
timestamp 1676037725
transform 1 0 35696 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_388
timestamp 1676037725
transform 1 0 36800 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_402
timestamp 1676037725
transform 1 0 38088 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_406
timestamp 1676037725
transform 1 0 38456 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_33
timestamp 1676037725
transform 1 0 4140 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_38
timestamp 1676037725
transform 1 0 4600 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_46
timestamp 1676037725
transform 1 0 5336 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_55
timestamp 1676037725
transform 1 0 6164 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_64
timestamp 1676037725
transform 1 0 6992 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_73
timestamp 1676037725
transform 1 0 7820 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1676037725
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_96
timestamp 1676037725
transform 1 0 9936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_117
timestamp 1676037725
transform 1 0 11868 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_127
timestamp 1676037725
transform 1 0 12788 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1676037725
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_150
timestamp 1676037725
transform 1 0 14904 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_173
timestamp 1676037725
transform 1 0 17020 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_184
timestamp 1676037725
transform 1 0 18032 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_188
timestamp 1676037725
transform 1 0 18400 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1676037725
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_206
timestamp 1676037725
transform 1 0 20056 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_214
timestamp 1676037725
transform 1 0 20792 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_222
timestamp 1676037725
transform 1 0 21528 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_232
timestamp 1676037725
transform 1 0 22448 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_240
timestamp 1676037725
transform 1 0 23184 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1676037725
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_263
timestamp 1676037725
transform 1 0 25300 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_276
timestamp 1676037725
transform 1 0 26496 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_286
timestamp 1676037725
transform 1 0 27416 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_290
timestamp 1676037725
transform 1 0 27784 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_299
timestamp 1676037725
transform 1 0 28612 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1676037725
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_318
timestamp 1676037725
transform 1 0 30360 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_322
timestamp 1676037725
transform 1 0 30728 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_337
timestamp 1676037725
transform 1 0 32108 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_345
timestamp 1676037725
transform 1 0 32844 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_355
timestamp 1676037725
transform 1 0 33764 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1676037725
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_375
timestamp 1676037725
transform 1 0 35604 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_384
timestamp 1676037725
transform 1 0 36432 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_405
timestamp 1676037725
transform 1 0 38364 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_21
timestamp 1676037725
transform 1 0 3036 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_24
timestamp 1676037725
transform 1 0 3312 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_29
timestamp 1676037725
transform 1 0 3772 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_36
timestamp 1676037725
transform 1 0 4416 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_45
timestamp 1676037725
transform 1 0 5244 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1676037725
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_64
timestamp 1676037725
transform 1 0 6992 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_73
timestamp 1676037725
transform 1 0 7820 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_82
timestamp 1676037725
transform 1 0 8648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_86
timestamp 1676037725
transform 1 0 9016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_104
timestamp 1676037725
transform 1 0 10672 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_122
timestamp 1676037725
transform 1 0 12328 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_130
timestamp 1676037725
transform 1 0 13064 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_138
timestamp 1676037725
transform 1 0 13800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_160
timestamp 1676037725
transform 1 0 15824 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_180
timestamp 1676037725
transform 1 0 17664 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_184
timestamp 1676037725
transform 1 0 18032 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_191
timestamp 1676037725
transform 1 0 18676 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_199
timestamp 1676037725
transform 1 0 19412 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_206
timestamp 1676037725
transform 1 0 20056 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_218
timestamp 1676037725
transform 1 0 21160 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_235
timestamp 1676037725
transform 1 0 22724 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_242
timestamp 1676037725
transform 1 0 23368 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_255
timestamp 1676037725
transform 1 0 24564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_263
timestamp 1676037725
transform 1 0 25300 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_272
timestamp 1676037725
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_292
timestamp 1676037725
transform 1 0 27968 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_312
timestamp 1676037725
transform 1 0 29808 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_320
timestamp 1676037725
transform 1 0 30544 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_328
timestamp 1676037725
transform 1 0 31280 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_345
timestamp 1676037725
transform 1 0 32844 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_351
timestamp 1676037725
transform 1 0 33396 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_361
timestamp 1676037725
transform 1 0 34316 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_373
timestamp 1676037725
transform 1 0 35420 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_381
timestamp 1676037725
transform 1 0 36156 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1676037725
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_404
timestamp 1676037725
transform 1 0 38272 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_33
timestamp 1676037725
transform 1 0 4140 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_37
timestamp 1676037725
transform 1 0 4508 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_46
timestamp 1676037725
transform 1 0 5336 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_55
timestamp 1676037725
transform 1 0 6164 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_64
timestamp 1676037725
transform 1 0 6992 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_73
timestamp 1676037725
transform 1 0 7820 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1676037725
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_96
timestamp 1676037725
transform 1 0 9936 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_107
timestamp 1676037725
transform 1 0 10948 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_111
timestamp 1676037725
transform 1 0 11316 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_128
timestamp 1676037725
transform 1 0 12880 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1676037725
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_149
timestamp 1676037725
transform 1 0 14812 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_160
timestamp 1676037725
transform 1 0 15824 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_185
timestamp 1676037725
transform 1 0 18124 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1676037725
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_206
timestamp 1676037725
transform 1 0 20056 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_216
timestamp 1676037725
transform 1 0 20976 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_229
timestamp 1676037725
transform 1 0 22172 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_239
timestamp 1676037725
transform 1 0 23092 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_249
timestamp 1676037725
transform 1 0 24012 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_267
timestamp 1676037725
transform 1 0 25668 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_275
timestamp 1676037725
transform 1 0 26404 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_288
timestamp 1676037725
transform 1 0 27600 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_292
timestamp 1676037725
transform 1 0 27968 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1676037725
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_324
timestamp 1676037725
transform 1 0 30912 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_335
timestamp 1676037725
transform 1 0 31924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_343
timestamp 1676037725
transform 1 0 32660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_351
timestamp 1676037725
transform 1 0 33396 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1676037725
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_370
timestamp 1676037725
transform 1 0 35144 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_391
timestamp 1676037725
transform 1 0 37076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_402
timestamp 1676037725
transform 1 0 38088 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1676037725
transform 1 0 38456 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_31
timestamp 1676037725
transform 1 0 3956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_38
timestamp 1676037725
transform 1 0 4600 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_44
timestamp 1676037725
transform 1 0 5152 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_48
timestamp 1676037725
transform 1 0 5520 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1676037725
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_62
timestamp 1676037725
transform 1 0 6808 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_71
timestamp 1676037725
transform 1 0 7636 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_91
timestamp 1676037725
transform 1 0 9476 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_104
timestamp 1676037725
transform 1 0 10672 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_127
timestamp 1676037725
transform 1 0 12788 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_131
timestamp 1676037725
transform 1 0 13156 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_150
timestamp 1676037725
transform 1 0 14904 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1676037725
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_180
timestamp 1676037725
transform 1 0 17664 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_188
timestamp 1676037725
transform 1 0 18400 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_208
timestamp 1676037725
transform 1 0 20240 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1676037725
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_233
timestamp 1676037725
transform 1 0 22540 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_243
timestamp 1676037725
transform 1 0 23460 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_266
timestamp 1676037725
transform 1 0 25576 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1676037725
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_301
timestamp 1676037725
transform 1 0 28796 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_309
timestamp 1676037725
transform 1 0 29532 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_323
timestamp 1676037725
transform 1 0 30820 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp 1676037725
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_346
timestamp 1676037725
transform 1 0 32936 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_355
timestamp 1676037725
transform 1 0 33764 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_376
timestamp 1676037725
transform 1 0 35696 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1676037725
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1676037725
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_19
timestamp 1676037725
transform 1 0 2852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1676037725
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_38
timestamp 1676037725
transform 1 0 4600 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_47
timestamp 1676037725
transform 1 0 5428 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_55
timestamp 1676037725
transform 1 0 6164 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_64
timestamp 1676037725
transform 1 0 6992 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_73
timestamp 1676037725
transform 1 0 7820 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1676037725
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_98
timestamp 1676037725
transform 1 0 10120 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_111
timestamp 1676037725
transform 1 0 11316 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_131
timestamp 1676037725
transform 1 0 13156 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1676037725
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_147
timestamp 1676037725
transform 1 0 14628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_157
timestamp 1676037725
transform 1 0 15548 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_181
timestamp 1676037725
transform 1 0 17756 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1676037725
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_208
timestamp 1676037725
transform 1 0 20240 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_218
timestamp 1676037725
transform 1 0 21160 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_243
timestamp 1676037725
transform 1 0 23460 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1676037725
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_260
timestamp 1676037725
transform 1 0 25024 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_272
timestamp 1676037725
transform 1 0 26128 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_278
timestamp 1676037725
transform 1 0 26680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_292
timestamp 1676037725
transform 1 0 27968 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1676037725
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_317
timestamp 1676037725
transform 1 0 30268 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_327
timestamp 1676037725
transform 1 0 31188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_333
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_351
timestamp 1676037725
transform 1 0 33396 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_361
timestamp 1676037725
transform 1 0 34316 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_373
timestamp 1676037725
transform 1 0 35420 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_379
timestamp 1676037725
transform 1 0 35972 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1676037725
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1676037725
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1676037725
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_16
timestamp 1676037725
transform 1 0 2576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_23
timestamp 1676037725
transform 1 0 3220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_30
timestamp 1676037725
transform 1 0 3864 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_37
timestamp 1676037725
transform 1 0 4508 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_45
timestamp 1676037725
transform 1 0 5244 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1676037725
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_70
timestamp 1676037725
transform 1 0 7544 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_90
timestamp 1676037725
transform 1 0 9384 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1676037725
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_145
timestamp 1676037725
transform 1 0 14444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_165
timestamp 1676037725
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_173
timestamp 1676037725
transform 1 0 17020 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_190
timestamp 1676037725
transform 1 0 18584 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_198
timestamp 1676037725
transform 1 0 19320 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1676037725
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_229
timestamp 1676037725
transform 1 0 22172 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_253
timestamp 1676037725
transform 1 0 24380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_277
timestamp 1676037725
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_293
timestamp 1676037725
transform 1 0 28060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_318
timestamp 1676037725
transform 1 0 30360 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_324
timestamp 1676037725
transform 1 0 30912 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1676037725
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_355
timestamp 1676037725
transform 1 0 33764 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_359
timestamp 1676037725
transform 1 0 34132 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_368
timestamp 1676037725
transform 1 0 34960 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_372
timestamp 1676037725
transform 1 0 35328 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1676037725
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_401
timestamp 1676037725
transform 1 0 37996 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1676037725
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_17
timestamp 1676037725
transform 1 0 2668 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1676037725
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_35
timestamp 1676037725
transform 1 0 4324 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_40
timestamp 1676037725
transform 1 0 4784 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_57
timestamp 1676037725
transform 1 0 6348 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_63
timestamp 1676037725
transform 1 0 6900 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_69
timestamp 1676037725
transform 1 0 7452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1676037725
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_96
timestamp 1676037725
transform 1 0 9936 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_100
timestamp 1676037725
transform 1 0 10304 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1676037725
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_113
timestamp 1676037725
transform 1 0 11500 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_125
timestamp 1676037725
transform 1 0 12604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1676037725
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_148
timestamp 1676037725
transform 1 0 14720 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_163
timestamp 1676037725
transform 1 0 16100 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1676037725
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_169
timestamp 1676037725
transform 1 0 16652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_179
timestamp 1676037725
transform 1 0 17572 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1676037725
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_219
timestamp 1676037725
transform 1 0 21252 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1676037725
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1676037725
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_236
timestamp 1676037725
transform 1 0 22816 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1676037725
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_259
timestamp 1676037725
transform 1 0 24932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_269
timestamp 1676037725
transform 1 0 25852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1676037725
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1676037725
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_289
timestamp 1676037725
transform 1 0 27692 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_299
timestamp 1676037725
transform 1 0 28612 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1676037725
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1676037725
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_345
timestamp 1676037725
transform 1 0 32844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_355
timestamp 1676037725
transform 1 0 33764 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1676037725
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1676037725
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_393
timestamp 1676037725
transform 1 0 37260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1676037725
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0828_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4324 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1676037725
transform 1 0 34132 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23736 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1676037725
transform 1 0 14352 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1676037725
transform 1 0 23920 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1676037725
transform 1 0 23828 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1676037725
transform 1 0 18676 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1676037725
transform 1 0 5152 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1676037725
transform 1 0 14260 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0838_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28612 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _0839_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17848 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _0840_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11960 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1676037725
transform 1 0 5796 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0843_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1676037725
transform 1 0 13524 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _0845_
timestamp 1676037725
transform 1 0 15272 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_8  _0846_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12328 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1676037725
transform 1 0 9936 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0848_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0849_
timestamp 1676037725
transform 1 0 7360 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0850_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25392 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28428 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0853_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31280 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0855_
timestamp 1676037725
transform 1 0 29716 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11500 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27968 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _0859_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35972 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31648 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1676037725
transform 1 0 23092 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _0862_
timestamp 1676037725
transform 1 0 30636 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28152 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_8  _0864_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28428 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _0865_
timestamp 1676037725
transform 1 0 27508 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0866_
timestamp 1676037725
transform 1 0 14260 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _0867_
timestamp 1676037725
transform 1 0 28060 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__or3b_4  _0868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0869_
timestamp 1676037725
transform 1 0 29072 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0870_
timestamp 1676037725
transform 1 0 29716 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0871_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28520 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0872_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7360 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0873_
timestamp 1676037725
transform 1 0 6532 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0874_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7360 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_4  _0875_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23828 0 -1 35904
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_1  _0876_
timestamp 1676037725
transform 1 0 14720 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0877_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31556 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0878_
timestamp 1676037725
transform 1 0 31464 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _0879_
timestamp 1676037725
transform 1 0 25760 0 1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _0880_
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0881_
timestamp 1676037725
transform 1 0 29900 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0882_
timestamp 1676037725
transform 1 0 21620 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0883_
timestamp 1676037725
transform 1 0 6992 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0884_
timestamp 1676037725
transform 1 0 20056 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0885_
timestamp 1676037725
transform 1 0 5152 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0887_
timestamp 1676037725
transform 1 0 28520 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1676037725
transform 1 0 34132 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0889_
timestamp 1676037725
transform 1 0 6808 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0890_
timestamp 1676037725
transform 1 0 3864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0891_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0892_
timestamp 1676037725
transform 1 0 17664 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1676037725
transform 1 0 1656 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0894_
timestamp 1676037725
transform 1 0 29348 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0895_
timestamp 1676037725
transform 1 0 21068 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0896_
timestamp 1676037725
transform 1 0 20240 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_4  _0897_
timestamp 1676037725
transform 1 0 24564 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _0898_
timestamp 1676037725
transform 1 0 24564 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0899_
timestamp 1676037725
transform 1 0 27140 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0900_
timestamp 1676037725
transform 1 0 25576 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0901_
timestamp 1676037725
transform 1 0 22356 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0902_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0903_
timestamp 1676037725
transform 1 0 15364 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0904_
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_4  _0905_
timestamp 1676037725
transform 1 0 29532 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0906_
timestamp 1676037725
transform 1 0 20792 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _0907_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _0908_
timestamp 1676037725
transform 1 0 26404 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0909_
timestamp 1676037725
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_2  _0910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25944 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _0911_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1676037725
transform 1 0 21896 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25760 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 1676037725
transform 1 0 28980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0915_
timestamp 1676037725
transform 1 0 4324 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_4  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22632 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_4  _0917_
timestamp 1676037725
transform 1 0 30084 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1676037725
transform 1 0 3496 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0919_
timestamp 1676037725
transform 1 0 28336 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0920_
timestamp 1676037725
transform 1 0 22448 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25392 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0922_
timestamp 1676037725
transform 1 0 34868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0923_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26128 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1676037725
transform 1 0 31556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0925_
timestamp 1676037725
transform 1 0 24564 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _0926_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26772 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_4  _0928_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__o22ai_1  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26772 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0930_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28152 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0931_
timestamp 1676037725
transform 1 0 28428 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _0932_
timestamp 1676037725
transform 1 0 29716 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0933_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26772 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_1  _0934_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25944 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _0935_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26036 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__nand4b_4  _0936_
timestamp 1676037725
transform 1 0 21160 0 1 29376
box -38 -48 1786 592
use sky130_fd_sc_hd__o31a_1  _0937_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21620 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0938_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20240 0 -1 30464
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _0939_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24748 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0940_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0941_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20608 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_4  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21896 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1676037725
transform 1 0 29716 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0944_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30544 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _0945_
timestamp 1676037725
transform 1 0 27692 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  _0946_
timestamp 1676037725
transform 1 0 30084 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__a221oi_4  _0947_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _0948_
timestamp 1676037725
transform 1 0 36708 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_8  _0949_
timestamp 1676037725
transform 1 0 27140 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _0950_
timestamp 1676037725
transform 1 0 24656 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _0951_
timestamp 1676037725
transform 1 0 27692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0953_
timestamp 1676037725
transform 1 0 27416 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _0954_
timestamp 1676037725
transform 1 0 29716 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0956_
timestamp 1676037725
transform 1 0 18400 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _0957_
timestamp 1676037725
transform 1 0 27784 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0958_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _0959_
timestamp 1676037725
transform 1 0 24932 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1676037725
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0961_
timestamp 1676037725
transform 1 0 29624 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0962_
timestamp 1676037725
transform 1 0 30452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _0963_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _0964_
timestamp 1676037725
transform 1 0 34592 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0965_
timestamp 1676037725
transform 1 0 29716 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _0966_
timestamp 1676037725
transform 1 0 26128 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0967_
timestamp 1676037725
transform 1 0 24564 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0968_
timestamp 1676037725
transform 1 0 24564 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0969_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34040 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0970_
timestamp 1676037725
transform 1 0 4324 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0971_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26864 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _0972_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0973_
timestamp 1676037725
transform 1 0 25852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_4  _0974_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0976_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25116 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _0977_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _0978_
timestamp 1676037725
transform 1 0 21068 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _0979_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24012 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _0980_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0981_
timestamp 1676037725
transform 1 0 19504 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0982_
timestamp 1676037725
transform 1 0 23644 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1676037725
transform 1 0 25300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0985_
timestamp 1676037725
transform 1 0 21252 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_2  _0987_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23552 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0988_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1676037725
transform 1 0 13524 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0990_
timestamp 1676037725
transform 1 0 14720 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0992_
timestamp 1676037725
transform 1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0993_
timestamp 1676037725
transform 1 0 18952 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0994_
timestamp 1676037725
transform 1 0 12880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0995_
timestamp 1676037725
transform 1 0 17296 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _0996_
timestamp 1676037725
transform 1 0 17664 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0997_
timestamp 1676037725
transform 1 0 29716 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0998_
timestamp 1676037725
transform 1 0 28520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _0999_
timestamp 1676037725
transform 1 0 32292 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1000_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1001_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28888 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1002_
timestamp 1676037725
transform 1 0 29624 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1003_
timestamp 1676037725
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1004_
timestamp 1676037725
transform 1 0 31556 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1005_
timestamp 1676037725
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24104 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1007_
timestamp 1676037725
transform 1 0 24288 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1008_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1009_
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1011_
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1012_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1013_
timestamp 1676037725
transform 1 0 17020 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1014_
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1015_
timestamp 1676037725
transform 1 0 31372 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1016_
timestamp 1676037725
transform 1 0 30728 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1017_
timestamp 1676037725
transform 1 0 32384 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1018_
timestamp 1676037725
transform 1 0 29348 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1019_
timestamp 1676037725
transform 1 0 30728 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1020_
timestamp 1676037725
transform 1 0 28796 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1021_
timestamp 1676037725
transform 1 0 26680 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1022_
timestamp 1676037725
transform 1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1023_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1024_
timestamp 1676037725
transform 1 0 26404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1025_
timestamp 1676037725
transform 1 0 23552 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1026_
timestamp 1676037725
transform 1 0 22724 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1027_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23092 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1028_
timestamp 1676037725
transform 1 0 20240 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1676037725
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1676037725
transform 1 0 21436 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _1031_
timestamp 1676037725
transform 1 0 19964 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_1  _1032_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23644 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1033_
timestamp 1676037725
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1034_
timestamp 1676037725
transform 1 0 23092 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1035_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1036_
timestamp 1676037725
transform 1 0 22448 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1037_
timestamp 1676037725
transform 1 0 29716 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1038_
timestamp 1676037725
transform 1 0 35972 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1039_
timestamp 1676037725
transform 1 0 27876 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1040_
timestamp 1676037725
transform 1 0 27140 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1041_
timestamp 1676037725
transform 1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1042_
timestamp 1676037725
transform 1 0 23092 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1043_
timestamp 1676037725
transform 1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1044_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1045_
timestamp 1676037725
transform 1 0 22632 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1046_
timestamp 1676037725
transform 1 0 22080 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1047_
timestamp 1676037725
transform 1 0 20332 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1048_
timestamp 1676037725
transform 1 0 20608 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1049_
timestamp 1676037725
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1051_
timestamp 1676037725
transform 1 0 28336 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1052_
timestamp 1676037725
transform 1 0 26312 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1053_
timestamp 1676037725
transform 1 0 28152 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1054_
timestamp 1676037725
transform 1 0 27232 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1055_
timestamp 1676037725
transform 1 0 28060 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1056_
timestamp 1676037725
transform 1 0 27140 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1057_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1058_
timestamp 1676037725
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1059_
timestamp 1676037725
transform 1 0 20516 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1060_
timestamp 1676037725
transform 1 0 20424 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1061_
timestamp 1676037725
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1062_
timestamp 1676037725
transform 1 0 17112 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1063_
timestamp 1676037725
transform 1 0 19596 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _1064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26128 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1066_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1067_
timestamp 1676037725
transform 1 0 24104 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1068_
timestamp 1676037725
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1069_
timestamp 1676037725
transform 1 0 23368 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1070_
timestamp 1676037725
transform 1 0 28796 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1071_
timestamp 1676037725
transform 1 0 30360 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1072_
timestamp 1676037725
transform 1 0 27324 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1073_
timestamp 1676037725
transform 1 0 21620 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21896 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _1075_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_2  _1076_
timestamp 1676037725
transform 1 0 20056 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _1077_
timestamp 1676037725
transform 1 0 18308 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__and2b_1  _1079_
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1080_
timestamp 1676037725
transform 1 0 19964 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1081_
timestamp 1676037725
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1082_
timestamp 1676037725
transform 1 0 20240 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1083_
timestamp 1676037725
transform 1 0 23828 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1084_
timestamp 1676037725
transform 1 0 20148 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1085_
timestamp 1676037725
transform 1 0 22724 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1086_
timestamp 1676037725
transform 1 0 24472 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1087_
timestamp 1676037725
transform 1 0 24196 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1089_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1090_
timestamp 1676037725
transform 1 0 20700 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1091_
timestamp 1676037725
transform 1 0 17112 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1092_
timestamp 1676037725
transform 1 0 17112 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_4  _1093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18400 0 -1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_2  _1094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _1095_
timestamp 1676037725
transform 1 0 17572 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _1096_
timestamp 1676037725
transform 1 0 17940 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_2  _1097_
timestamp 1676037725
transform 1 0 21344 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1098_
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1099_
timestamp 1676037725
transform 1 0 18400 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1100_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19504 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _1102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _1103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__o211ai_4  _1104_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _1105_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1106_
timestamp 1676037725
transform 1 0 18584 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1107_
timestamp 1676037725
transform 1 0 18768 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1108_
timestamp 1676037725
transform 1 0 17572 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_4  _1109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15916 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__o211ai_4  _1110_
timestamp 1676037725
transform 1 0 15640 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_1  _1111_
timestamp 1676037725
transform 1 0 26128 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1112_
timestamp 1676037725
transform 1 0 25024 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1113_
timestamp 1676037725
transform 1 0 27324 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _1114_
timestamp 1676037725
transform 1 0 38088 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1115_
timestamp 1676037725
transform 1 0 27416 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _1116_
timestamp 1676037725
transform 1 0 27232 0 1 23936
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _1117_
timestamp 1676037725
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1118_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1119_
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1120_
timestamp 1676037725
transform 1 0 21896 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1121_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1122_
timestamp 1676037725
transform 1 0 17572 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1123_
timestamp 1676037725
transform 1 0 16560 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1124_
timestamp 1676037725
transform 1 0 15824 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1126_
timestamp 1676037725
transform 1 0 16192 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1127_
timestamp 1676037725
transform 1 0 14996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1129_
timestamp 1676037725
transform 1 0 15180 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _1130_
timestamp 1676037725
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1131_
timestamp 1676037725
transform 1 0 21160 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1132_
timestamp 1676037725
transform 1 0 23736 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1133_
timestamp 1676037725
transform 1 0 23000 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1135_
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1136_
timestamp 1676037725
transform 1 0 16008 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp 1676037725
transform 1 0 14628 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1138_
timestamp 1676037725
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1139_
timestamp 1676037725
transform 1 0 12328 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1140_
timestamp 1676037725
transform 1 0 14536 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1141_
timestamp 1676037725
transform 1 0 15456 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1142_
timestamp 1676037725
transform 1 0 13984 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1143_
timestamp 1676037725
transform 1 0 15640 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1144_
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1145_
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15088 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1148_
timestamp 1676037725
transform 1 0 13248 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1149_
timestamp 1676037725
transform 1 0 18216 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18308 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1151_
timestamp 1676037725
transform 1 0 4692 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1676037725
transform 1 0 19228 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1153_
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1154_
timestamp 1676037725
transform 1 0 31004 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1155_
timestamp 1676037725
transform 1 0 31096 0 1 30464
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_2  _1156_
timestamp 1676037725
transform 1 0 35604 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_8  _1157_
timestamp 1676037725
transform 1 0 29716 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__o31ai_4  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_8  _1159_
timestamp 1676037725
transform 1 0 30360 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _1160_
timestamp 1676037725
transform 1 0 30912 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1161_
timestamp 1676037725
transform 1 0 31096 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1162_
timestamp 1676037725
transform 1 0 5704 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1163_
timestamp 1676037725
transform 1 0 5152 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1164_
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1165_
timestamp 1676037725
transform 1 0 34868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1166_
timestamp 1676037725
transform 1 0 37904 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1167_
timestamp 1676037725
transform 1 0 29072 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1168_
timestamp 1676037725
transform 1 0 30176 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1169_
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29072 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30728 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _1172_
timestamp 1676037725
transform 1 0 31188 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_2  _1173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31188 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1174_
timestamp 1676037725
transform 1 0 30636 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1175_
timestamp 1676037725
transform 1 0 31280 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1176_
timestamp 1676037725
transform 1 0 31556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1177_
timestamp 1676037725
transform 1 0 33580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1178_
timestamp 1676037725
transform 1 0 33212 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1179_
timestamp 1676037725
transform 1 0 29900 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _1180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30912 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_2  _1181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31924 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1182_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _1184_
timestamp 1676037725
transform 1 0 34868 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1185_
timestamp 1676037725
transform 1 0 33764 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1186_
timestamp 1676037725
transform 1 0 33948 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1187_
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1188_
timestamp 1676037725
transform 1 0 34684 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1189_
timestamp 1676037725
transform 1 0 33948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1190_
timestamp 1676037725
transform 1 0 36708 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1191_
timestamp 1676037725
transform 1 0 35880 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1192_
timestamp 1676037725
transform 1 0 34500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1193_
timestamp 1676037725
transform 1 0 34040 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1194_
timestamp 1676037725
transform 1 0 35144 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1195_
timestamp 1676037725
transform 1 0 35236 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1196_
timestamp 1676037725
transform 1 0 34960 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1197_
timestamp 1676037725
transform 1 0 34868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 1676037725
transform 1 0 36064 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1199_
timestamp 1676037725
transform 1 0 36156 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1200_
timestamp 1676037725
transform 1 0 34592 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1201_
timestamp 1676037725
transform 1 0 36616 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1202_
timestamp 1676037725
transform 1 0 36064 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1203_
timestamp 1676037725
transform 1 0 35236 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1204_
timestamp 1676037725
transform 1 0 36432 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1205_
timestamp 1676037725
transform 1 0 33396 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1206_
timestamp 1676037725
transform 1 0 35788 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1207_
timestamp 1676037725
transform 1 0 34868 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33672 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1209_
timestamp 1676037725
transform 1 0 36984 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1210_
timestamp 1676037725
transform 1 0 33028 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1211_
timestamp 1676037725
transform 1 0 33672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32844 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1213_
timestamp 1676037725
transform 1 0 30084 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1214_
timestamp 1676037725
transform 1 0 37352 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1215_
timestamp 1676037725
transform 1 0 32752 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1216_
timestamp 1676037725
transform 1 0 33488 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1217_
timestamp 1676037725
transform 1 0 34868 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1218_
timestamp 1676037725
transform 1 0 32844 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1219_
timestamp 1676037725
transform 1 0 33948 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1220_
timestamp 1676037725
transform 1 0 30084 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1221_
timestamp 1676037725
transform 1 0 28336 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1222_
timestamp 1676037725
transform 1 0 5152 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1223_
timestamp 1676037725
transform 1 0 32936 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1224_
timestamp 1676037725
transform 1 0 33488 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1225_
timestamp 1676037725
transform 1 0 33764 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1226_
timestamp 1676037725
transform 1 0 32936 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1227_
timestamp 1676037725
transform 1 0 34868 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1228_
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1229_
timestamp 1676037725
transform 1 0 4784 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1230_
timestamp 1676037725
transform 1 0 3680 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1231_
timestamp 1676037725
transform 1 0 32844 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1232_
timestamp 1676037725
transform 1 0 33948 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1233_
timestamp 1676037725
transform 1 0 3220 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 1676037725
transform 1 0 7084 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1235_
timestamp 1676037725
transform 1 0 5612 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1236_
timestamp 1676037725
transform 1 0 33028 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1237_
timestamp 1676037725
transform 1 0 34684 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1238_
timestamp 1676037725
transform 1 0 34316 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1239_
timestamp 1676037725
transform 1 0 14812 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1240_
timestamp 1676037725
transform 1 0 15272 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1241_
timestamp 1676037725
transform 1 0 18400 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1242_
timestamp 1676037725
transform 1 0 14076 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1243_
timestamp 1676037725
transform 1 0 9108 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1244_
timestamp 1676037725
transform 1 0 4140 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1245_
timestamp 1676037725
transform 1 0 11776 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _1246_
timestamp 1676037725
transform 1 0 6532 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _1247_
timestamp 1676037725
transform 1 0 11684 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1248_
timestamp 1676037725
transform 1 0 9844 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1249_
timestamp 1676037725
transform 1 0 9292 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1250_
timestamp 1676037725
transform 1 0 10304 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1251_
timestamp 1676037725
transform 1 0 5704 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1252_
timestamp 1676037725
transform 1 0 4784 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2_4  _1253_
timestamp 1676037725
transform 1 0 10028 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1254_
timestamp 1676037725
transform 1 0 10304 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1676037725
transform 1 0 7176 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_8  _1256_
timestamp 1676037725
transform 1 0 11408 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _1257_
timestamp 1676037725
transform 1 0 12420 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1258_
timestamp 1676037725
transform 1 0 7360 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1259_
timestamp 1676037725
transform 1 0 12328 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1260_
timestamp 1676037725
transform 1 0 11684 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1261_
timestamp 1676037725
transform 1 0 18492 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22264 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1263_
timestamp 1676037725
transform 1 0 30544 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1264_
timestamp 1676037725
transform 1 0 21988 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_1  _1265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21436 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1266_
timestamp 1676037725
transform 1 0 22356 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1267_
timestamp 1676037725
transform 1 0 6532 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1268_
timestamp 1676037725
transform 1 0 15180 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1269_
timestamp 1676037725
transform 1 0 9200 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1270_
timestamp 1676037725
transform 1 0 15272 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1271_
timestamp 1676037725
transform 1 0 14260 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1272_
timestamp 1676037725
transform 1 0 14260 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1273_
timestamp 1676037725
transform 1 0 20976 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1274_
timestamp 1676037725
transform 1 0 7268 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1275_
timestamp 1676037725
transform 1 0 5796 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1276_
timestamp 1676037725
transform 1 0 5152 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1277_
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1278_
timestamp 1676037725
transform 1 0 10396 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1279_
timestamp 1676037725
transform 1 0 16928 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1280_
timestamp 1676037725
transform 1 0 14168 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1281_
timestamp 1676037725
transform 1 0 22816 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1282_
timestamp 1676037725
transform 1 0 5796 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1283_
timestamp 1676037725
transform 1 0 25576 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1284_
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1285_
timestamp 1676037725
transform 1 0 33304 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1286_
timestamp 1676037725
transform 1 0 23644 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1287_
timestamp 1676037725
transform 1 0 26220 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1288_
timestamp 1676037725
transform 1 0 16928 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1289_
timestamp 1676037725
transform 1 0 27232 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1290_
timestamp 1676037725
transform 1 0 24564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1291_
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1292_
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1293_
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1294_
timestamp 1676037725
transform 1 0 15088 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1295_
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1296_
timestamp 1676037725
transform 1 0 14904 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1297_
timestamp 1676037725
transform 1 0 19780 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1298_
timestamp 1676037725
transform 1 0 34132 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1676037725
transform 1 0 6716 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1676037725
transform 1 0 4048 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1301_
timestamp 1676037725
transform 1 0 8188 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1302_
timestamp 1676037725
transform 1 0 16008 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1303_
timestamp 1676037725
transform 1 0 13248 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1304_
timestamp 1676037725
transform 1 0 20792 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1305_
timestamp 1676037725
transform 1 0 14168 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1306_
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1307_
timestamp 1676037725
transform 1 0 12144 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1308_
timestamp 1676037725
transform 1 0 13248 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1309_
timestamp 1676037725
transform 1 0 17020 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1310_
timestamp 1676037725
transform 1 0 13248 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18492 0 -1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__xnor2_1  _1312_
timestamp 1676037725
transform 1 0 19596 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1313_
timestamp 1676037725
transform 1 0 23736 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1314_
timestamp 1676037725
transform 1 0 15180 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1315_
timestamp 1676037725
transform 1 0 24564 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20424 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1317_
timestamp 1676037725
transform 1 0 19412 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19504 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1319_
timestamp 1676037725
transform 1 0 4968 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1320_
timestamp 1676037725
transform 1 0 9476 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1321_
timestamp 1676037725
transform 1 0 13248 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1322_
timestamp 1676037725
transform 1 0 5612 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1323_
timestamp 1676037725
transform 1 0 7268 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1324_
timestamp 1676037725
transform 1 0 13156 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1325_
timestamp 1676037725
transform 1 0 13524 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1326_
timestamp 1676037725
transform 1 0 7268 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1327_
timestamp 1676037725
transform 1 0 11316 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17020 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1329_
timestamp 1676037725
transform 1 0 16928 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1330_
timestamp 1676037725
transform 1 0 15272 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1331_
timestamp 1676037725
transform 1 0 15088 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1332_
timestamp 1676037725
transform 1 0 15456 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1333_
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1334_
timestamp 1676037725
transform 1 0 24748 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _1336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24748 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _1337_
timestamp 1676037725
transform 1 0 25484 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1338_
timestamp 1676037725
transform 1 0 19780 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1339_
timestamp 1676037725
transform 1 0 24564 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1340_
timestamp 1676037725
transform 1 0 20976 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1341_
timestamp 1676037725
transform 1 0 16100 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1342_
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1343_
timestamp 1676037725
transform 1 0 17756 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1344_
timestamp 1676037725
transform 1 0 14260 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1345_
timestamp 1676037725
transform 1 0 4508 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1346_
timestamp 1676037725
transform 1 0 10948 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1347_
timestamp 1676037725
transform 1 0 21896 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1348_
timestamp 1676037725
transform 1 0 20424 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1349_
timestamp 1676037725
transform 1 0 13524 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1350_
timestamp 1676037725
transform 1 0 37996 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1351_
timestamp 1676037725
transform 1 0 27140 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1352_
timestamp 1676037725
transform 1 0 20976 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1353_
timestamp 1676037725
transform 1 0 21988 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 1676037725
transform 1 0 28336 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1355_
timestamp 1676037725
transform 1 0 27876 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _1356_
timestamp 1676037725
transform 1 0 25484 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1357_
timestamp 1676037725
transform 1 0 28980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1358_
timestamp 1676037725
transform 1 0 23552 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1359_
timestamp 1676037725
transform 1 0 4232 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1360_
timestamp 1676037725
transform 1 0 23552 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1361_
timestamp 1676037725
transform 1 0 18952 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_2  _1362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26772 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1363_
timestamp 1676037725
transform 1 0 34868 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1364_
timestamp 1676037725
transform 1 0 32292 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1365_
timestamp 1676037725
transform 1 0 25852 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1366_
timestamp 1676037725
transform 1 0 25668 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1367_
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _1368_
timestamp 1676037725
transform 1 0 31924 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_4  _1369_
timestamp 1676037725
transform 1 0 33764 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _1370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31096 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__o21ai_4  _1371_
timestamp 1676037725
transform 1 0 30636 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _1372_
timestamp 1676037725
transform 1 0 35880 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1373_
timestamp 1676037725
transform 1 0 14352 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1374_
timestamp 1676037725
transform 1 0 28336 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1375_
timestamp 1676037725
transform 1 0 32292 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1376_
timestamp 1676037725
transform 1 0 31280 0 1 32640
box -38 -48 1326 592
use sky130_fd_sc_hd__or3_4  _1377_
timestamp 1676037725
transform 1 0 32568 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_2  _1378_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28980 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1379_
timestamp 1676037725
transform 1 0 33396 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _1380_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33304 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _1381_
timestamp 1676037725
transform 1 0 33488 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1382_
timestamp 1676037725
transform 1 0 32108 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1383_
timestamp 1676037725
transform 1 0 33672 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1384_
timestamp 1676037725
transform 1 0 33304 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1385_
timestamp 1676037725
transform 1 0 33304 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1386_
timestamp 1676037725
transform 1 0 34868 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1387_
timestamp 1676037725
transform 1 0 33396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1388_
timestamp 1676037725
transform 1 0 32292 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1389_
timestamp 1676037725
transform 1 0 34316 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1390_
timestamp 1676037725
transform 1 0 34776 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1391_
timestamp 1676037725
transform 1 0 32568 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1392_
timestamp 1676037725
transform 1 0 35880 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1393_
timestamp 1676037725
transform 1 0 34960 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1394_
timestamp 1676037725
transform 1 0 32844 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1395_
timestamp 1676037725
transform 1 0 35604 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1396_
timestamp 1676037725
transform 1 0 34868 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1397_
timestamp 1676037725
transform 1 0 33212 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1398_
timestamp 1676037725
transform 1 0 35144 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1399_
timestamp 1676037725
transform 1 0 34868 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1400_
timestamp 1676037725
transform 1 0 33672 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1401_
timestamp 1676037725
transform 1 0 36064 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1402_
timestamp 1676037725
transform 1 0 35696 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1403_
timestamp 1676037725
transform 1 0 33396 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1404_
timestamp 1676037725
transform 1 0 35604 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1405_
timestamp 1676037725
transform 1 0 35972 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _1406_
timestamp 1676037725
transform 1 0 33764 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1407_
timestamp 1676037725
transform 1 0 35880 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1408_
timestamp 1676037725
transform 1 0 34776 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1409_
timestamp 1676037725
transform 1 0 34868 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1410_
timestamp 1676037725
transform 1 0 35880 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1411_
timestamp 1676037725
transform 1 0 36432 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1412_
timestamp 1676037725
transform 1 0 35052 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1413_
timestamp 1676037725
transform 1 0 35696 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1414_
timestamp 1676037725
transform 1 0 35880 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1415_
timestamp 1676037725
transform 1 0 35880 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1416_
timestamp 1676037725
transform 1 0 33856 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1417_
timestamp 1676037725
transform 1 0 36156 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1418_
timestamp 1676037725
transform 1 0 37444 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1419_
timestamp 1676037725
transform 1 0 35512 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1420_
timestamp 1676037725
transform 1 0 37444 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1421_
timestamp 1676037725
transform 1 0 36064 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1422_
timestamp 1676037725
transform 1 0 35052 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1423_
timestamp 1676037725
transform 1 0 36248 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _1424_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30728 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_4  _1425_
timestamp 1676037725
transform 1 0 29992 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _1426_
timestamp 1676037725
transform 1 0 34868 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1427_
timestamp 1676037725
transform 1 0 32292 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1428_
timestamp 1676037725
transform 1 0 35788 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1429_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31832 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1430_
timestamp 1676037725
transform 1 0 30084 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1431_
timestamp 1676037725
transform 1 0 32752 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _1432_
timestamp 1676037725
transform 1 0 32384 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1433_
timestamp 1676037725
transform 1 0 30268 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 1676037725
transform 1 0 34960 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1435_
timestamp 1676037725
transform 1 0 36708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1436_
timestamp 1676037725
transform 1 0 32936 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1437_
timestamp 1676037725
transform 1 0 30820 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1438_
timestamp 1676037725
transform 1 0 31004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_2  _1439_
timestamp 1676037725
transform 1 0 32292 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1440_
timestamp 1676037725
transform 1 0 33856 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1441_
timestamp 1676037725
transform 1 0 30544 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1442_
timestamp 1676037725
transform 1 0 30820 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_2  _1443_
timestamp 1676037725
transform 1 0 28520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _1444_
timestamp 1676037725
transform 1 0 29808 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1445_
timestamp 1676037725
transform 1 0 36064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1446_
timestamp 1676037725
transform 1 0 33856 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1447_
timestamp 1676037725
transform 1 0 32108 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1448_
timestamp 1676037725
transform 1 0 33304 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1449_
timestamp 1676037725
transform 1 0 30820 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1450_
timestamp 1676037725
transform 1 0 33856 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _1451_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32476 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1452_
timestamp 1676037725
transform 1 0 34868 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1453_
timestamp 1676037725
transform 1 0 32292 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _1454_
timestamp 1676037725
transform 1 0 31096 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _1455_
timestamp 1676037725
transform 1 0 22724 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_4  _1456_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 26112
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_4  _1457_
timestamp 1676037725
transform 1 0 26588 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1458_
timestamp 1676037725
transform 1 0 24932 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1459_
timestamp 1676037725
transform 1 0 23552 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1460_
timestamp 1676037725
transform 1 0 26588 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1461_
timestamp 1676037725
transform 1 0 26036 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1462_
timestamp 1676037725
transform 1 0 27416 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1463_
timestamp 1676037725
transform 1 0 25852 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1464_
timestamp 1676037725
transform 1 0 25484 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1465_
timestamp 1676037725
transform 1 0 31556 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1466_
timestamp 1676037725
transform 1 0 27140 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 1676037725
transform 1 0 27140 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1468_
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1469_
timestamp 1676037725
transform 1 0 31648 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1470_
timestamp 1676037725
transform 1 0 28888 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1471_
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_2  _1472_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25300 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1473_
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1474_
timestamp 1676037725
transform 1 0 25392 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1475_
timestamp 1676037725
transform 1 0 27876 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1476_
timestamp 1676037725
transform 1 0 29716 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1477_
timestamp 1676037725
transform 1 0 28244 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1478_
timestamp 1676037725
transform 1 0 29532 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1479_
timestamp 1676037725
transform 1 0 28428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1480_
timestamp 1676037725
transform 1 0 28520 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1481_
timestamp 1676037725
transform 1 0 25760 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1482_
timestamp 1676037725
transform 1 0 21252 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1483_
timestamp 1676037725
transform 1 0 27324 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1484_
timestamp 1676037725
transform 1 0 27232 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1485_
timestamp 1676037725
transform 1 0 29072 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1487_
timestamp 1676037725
transform 1 0 29624 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1488_
timestamp 1676037725
transform 1 0 28244 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1489_
timestamp 1676037725
transform 1 0 34132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1490_
timestamp 1676037725
transform 1 0 28888 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1491_
timestamp 1676037725
transform 1 0 28060 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_2  _1492_
timestamp 1676037725
transform 1 0 28244 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1493_
timestamp 1676037725
transform 1 0 28612 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1494_
timestamp 1676037725
transform 1 0 27140 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1495_
timestamp 1676037725
transform 1 0 25944 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1496_
timestamp 1676037725
transform 1 0 28980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1497_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_2  _1498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26036 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1499_
timestamp 1676037725
transform 1 0 25300 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1500_
timestamp 1676037725
transform 1 0 22540 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1501_
timestamp 1676037725
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1502_
timestamp 1676037725
transform 1 0 24932 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1503_
timestamp 1676037725
transform 1 0 21252 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1504_
timestamp 1676037725
transform 1 0 34592 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1505_
timestamp 1676037725
transform 1 0 32384 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1506_
timestamp 1676037725
transform 1 0 31924 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1507_
timestamp 1676037725
transform 1 0 33580 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1508_
timestamp 1676037725
transform 1 0 27968 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1509_
timestamp 1676037725
transform 1 0 34040 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1510_
timestamp 1676037725
transform 1 0 28060 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1511_
timestamp 1676037725
transform 1 0 5152 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1512_
timestamp 1676037725
transform 1 0 26036 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1513_
timestamp 1676037725
transform 1 0 27324 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1514_
timestamp 1676037725
transform 1 0 34868 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1515_
timestamp 1676037725
transform 1 0 23000 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1516_
timestamp 1676037725
transform 1 0 25852 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1517_
timestamp 1676037725
transform 1 0 30084 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1518_
timestamp 1676037725
transform 1 0 32476 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1519_
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1520_
timestamp 1676037725
transform 1 0 33580 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1522_
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1523_
timestamp 1676037725
transform 1 0 37444 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1524_
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1525_
timestamp 1676037725
transform 1 0 37444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1526_
timestamp 1676037725
transform 1 0 37444 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1527_
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1528_
timestamp 1676037725
transform 1 0 18124 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1529_
timestamp 1676037725
transform 1 0 19596 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1530_
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1531_
timestamp 1676037725
transform 1 0 18676 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1532_
timestamp 1676037725
transform 1 0 17480 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1533_
timestamp 1676037725
transform 1 0 17848 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1534_
timestamp 1676037725
transform 1 0 17480 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1535_
timestamp 1676037725
transform 1 0 23736 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1536_
timestamp 1676037725
transform 1 0 20884 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1537_
timestamp 1676037725
transform 1 0 22172 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1539_
timestamp 1676037725
transform 1 0 23460 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1540_
timestamp 1676037725
transform 1 0 24564 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1541_
timestamp 1676037725
transform 1 0 23828 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1542_
timestamp 1676037725
transform 1 0 23276 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1543_
timestamp 1676037725
transform 1 0 23092 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1544_
timestamp 1676037725
transform 1 0 21896 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1545_
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1546_
timestamp 1676037725
transform 1 0 20424 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1547_
timestamp 1676037725
transform 1 0 20976 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1548_
timestamp 1676037725
transform 1 0 20516 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1549_
timestamp 1676037725
transform 1 0 16560 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1550_
timestamp 1676037725
transform 1 0 17388 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1551_
timestamp 1676037725
transform 1 0 17480 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1552_
timestamp 1676037725
transform 1 0 17296 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1553_
timestamp 1676037725
transform 1 0 16836 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1554_
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _1555_
timestamp 1676037725
transform 1 0 23276 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1556_
timestamp 1676037725
transform 1 0 23184 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1557_
timestamp 1676037725
transform 1 0 21988 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1558_
timestamp 1676037725
transform 1 0 21804 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1559_
timestamp 1676037725
transform 1 0 23368 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1560_
timestamp 1676037725
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1562_
timestamp 1676037725
transform 1 0 13064 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1563_
timestamp 1676037725
transform 1 0 13156 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1564_
timestamp 1676037725
transform 1 0 14168 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1565_
timestamp 1676037725
transform 1 0 17112 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1566_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1567_
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1568_
timestamp 1676037725
transform 1 0 19412 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1569_
timestamp 1676037725
transform 1 0 9108 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1570_
timestamp 1676037725
transform 1 0 9108 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1571_
timestamp 1676037725
transform 1 0 10488 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1572_
timestamp 1676037725
transform 1 0 11776 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1573_
timestamp 1676037725
transform 1 0 12972 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1574_
timestamp 1676037725
transform 1 0 16560 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1575_
timestamp 1676037725
transform 1 0 14720 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1576_
timestamp 1676037725
transform 1 0 19412 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1577_
timestamp 1676037725
transform 1 0 4232 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1578_
timestamp 1676037725
transform 1 0 26036 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _1579_
timestamp 1676037725
transform 1 0 11776 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1580_
timestamp 1676037725
transform 1 0 4324 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1581_
timestamp 1676037725
transform 1 0 12144 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1582_
timestamp 1676037725
transform 1 0 7452 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1583_
timestamp 1676037725
transform 1 0 6992 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1584_
timestamp 1676037725
transform 1 0 10396 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1585_
timestamp 1676037725
transform 1 0 9108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1586_
timestamp 1676037725
transform 1 0 8096 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1587_
timestamp 1676037725
transform 1 0 11316 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1588_
timestamp 1676037725
transform 1 0 7912 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1589_
timestamp 1676037725
transform 1 0 6808 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1590_
timestamp 1676037725
transform 1 0 6440 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1591_
timestamp 1676037725
transform 1 0 8648 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1592_
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1593_
timestamp 1676037725
transform 1 0 10212 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1594_
timestamp 1676037725
transform 1 0 9108 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1595_
timestamp 1676037725
transform 1 0 37444 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1596_
timestamp 1676037725
transform 1 0 4508 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9384 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1598_
timestamp 1676037725
transform 1 0 9108 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1599_
timestamp 1676037725
transform 1 0 9200 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1600_
timestamp 1676037725
transform 1 0 20976 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1601_
timestamp 1676037725
transform 1 0 19228 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1602_
timestamp 1676037725
transform 1 0 10580 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1603_
timestamp 1676037725
transform 1 0 10212 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1604_
timestamp 1676037725
transform 1 0 9108 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1605_
timestamp 1676037725
transform 1 0 8004 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1606_
timestamp 1676037725
transform 1 0 12420 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1607_
timestamp 1676037725
transform 1 0 12880 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1608_
timestamp 1676037725
transform 1 0 11408 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1609_
timestamp 1676037725
transform 1 0 9200 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1610_
timestamp 1676037725
transform 1 0 8096 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1611_
timestamp 1676037725
transform 1 0 9752 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1612_
timestamp 1676037725
transform 1 0 9476 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1613_
timestamp 1676037725
transform 1 0 7820 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1614_
timestamp 1676037725
transform 1 0 4324 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1615_
timestamp 1676037725
transform 1 0 12972 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1616_
timestamp 1676037725
transform 1 0 20148 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1617_
timestamp 1676037725
transform 1 0 8096 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1618_
timestamp 1676037725
transform 1 0 9568 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1619_
timestamp 1676037725
transform 1 0 6440 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1620_
timestamp 1676037725
transform 1 0 9108 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1621_
timestamp 1676037725
transform 1 0 8004 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1622_
timestamp 1676037725
transform 1 0 9568 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1623_
timestamp 1676037725
transform 1 0 9568 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1624_
timestamp 1676037725
transform 1 0 13432 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1676037725
transform 1 0 14260 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1626_
timestamp 1676037725
transform 1 0 11408 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1627_
timestamp 1676037725
transform 1 0 12236 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1628_
timestamp 1676037725
transform 1 0 15732 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1629_
timestamp 1676037725
transform 1 0 15364 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1630_
timestamp 1676037725
transform 1 0 10580 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1631_
timestamp 1676037725
transform 1 0 10580 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1632_
timestamp 1676037725
transform 1 0 10396 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1633_
timestamp 1676037725
transform 1 0 6716 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1634_
timestamp 1676037725
transform 1 0 11776 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1635_
timestamp 1676037725
transform 1 0 12696 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1636_
timestamp 1676037725
transform 1 0 13340 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1637_
timestamp 1676037725
transform 1 0 11776 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1638_
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1639_
timestamp 1676037725
transform 1 0 10672 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1640_
timestamp 1676037725
transform 1 0 10396 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _1641_
timestamp 1676037725
transform 1 0 13340 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1642_
timestamp 1676037725
transform 1 0 12328 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1643_
timestamp 1676037725
transform 1 0 12420 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1644_
timestamp 1676037725
transform 1 0 11684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1645_
timestamp 1676037725
transform 1 0 11684 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1646_
timestamp 1676037725
transform 1 0 13064 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1647_
timestamp 1676037725
transform 1 0 11960 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1648_
timestamp 1676037725
transform 1 0 11500 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1676037725
transform 1 0 11684 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1650_
timestamp 1676037725
transform 1 0 14720 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1651_
timestamp 1676037725
transform 1 0 10028 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1652_
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1653_
timestamp 1676037725
transform 1 0 13248 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1654_
timestamp 1676037725
transform 1 0 16836 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1655_
timestamp 1676037725
transform 1 0 14444 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1656_
timestamp 1676037725
transform 1 0 15640 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1657_
timestamp 1676037725
transform 1 0 14996 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1658_
timestamp 1676037725
transform 1 0 14720 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1659_
timestamp 1676037725
transform 1 0 15364 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1660_
timestamp 1676037725
transform 1 0 15456 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1676037725
transform 1 0 17940 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1662_
timestamp 1676037725
transform 1 0 17756 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1663_
timestamp 1676037725
transform 1 0 32292 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1664_
timestamp 1676037725
transform 1 0 5704 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 1676037725
transform 1 0 37444 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1666_
timestamp 1676037725
transform 1 0 37444 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1667_
timestamp 1676037725
transform 1 0 37444 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1668_
timestamp 1676037725
transform 1 0 37444 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1669_
timestamp 1676037725
transform 1 0 37444 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1670_
timestamp 1676037725
transform 1 0 37444 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1671_
timestamp 1676037725
transform 1 0 37444 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1672_
timestamp 1676037725
transform 1 0 37536 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1673_
timestamp 1676037725
transform 1 0 27416 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1674_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1675_
timestamp 1676037725
transform 1 0 27968 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1676_
timestamp 1676037725
transform 1 0 21988 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1677_
timestamp 1676037725
transform 1 0 30728 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1678_
timestamp 1676037725
transform 1 0 30176 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1679_
timestamp 1676037725
transform 1 0 30360 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1680_
timestamp 1676037725
transform 1 0 30268 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1681_
timestamp 1676037725
transform 1 0 25392 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1682_
timestamp 1676037725
transform 1 0 26036 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1683_
timestamp 1676037725
transform 1 0 22908 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1684_
timestamp 1676037725
transform 1 0 26404 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1685_
timestamp 1676037725
transform 1 0 20608 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1686_
timestamp 1676037725
transform 1 0 34868 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1687_
timestamp 1676037725
transform 1 0 32384 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1688_
timestamp 1676037725
transform 1 0 31004 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 1676037725
transform 1 0 34868 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1690_
timestamp 1676037725
transform 1 0 27232 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1691_
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1676037725
transform 1 0 2944 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1676037725
transform 1 0 6532 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1694_
timestamp 1676037725
transform 1 0 3220 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1695_
timestamp 1676037725
transform 1 0 2300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19688 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1697_
timestamp 1676037725
transform 1 0 19412 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1698_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22264 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _1699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21528 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1700_
timestamp 1676037725
transform 1 0 24748 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1701_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28428 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1702_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1676037725
transform 1 0 26128 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1676037725
transform 1 0 22724 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1676037725
transform 1 0 27784 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1676037725
transform 1 0 28520 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1676037725
transform 1 0 27784 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1676037725
transform 1 0 24748 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1676037725
transform 1 0 21804 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1676037725
transform 1 0 24288 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1676037725
transform 1 0 34868 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1676037725
transform 1 0 32200 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1676037725
transform 1 0 31924 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1676037725
transform 1 0 34684 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1676037725
transform 1 0 26128 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12972 0 -1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1719_
timestamp 1676037725
transform 1 0 12420 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1676037725
transform 1 0 23460 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1721_
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1722_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1723_
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1724_
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1725_
timestamp 1676037725
transform 1 0 21712 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1726_
timestamp 1676037725
transform 1 0 15456 0 1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1727_
timestamp 1676037725
transform 1 0 15732 0 1 21760
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1676037725
transform 1 0 11224 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1731_
timestamp 1676037725
transform 1 0 28612 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1732_
timestamp 1676037725
transform 1 0 30820 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1733_
timestamp 1676037725
transform 1 0 34960 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1734_
timestamp 1676037725
transform 1 0 36524 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1735_
timestamp 1676037725
transform 1 0 36248 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1736_
timestamp 1676037725
transform 1 0 36156 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1737_
timestamp 1676037725
transform 1 0 35420 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1676037725
transform 1 0 35512 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1676037725
transform 1 0 34868 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1676037725
transform 1 0 35052 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1741_
timestamp 1676037725
transform 1 0 34868 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1742_
timestamp 1676037725
transform 1 0 35512 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1743_
timestamp 1676037725
transform 1 0 34132 0 -1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1744_
timestamp 1676037725
transform 1 0 35420 0 -1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1745_
timestamp 1676037725
transform 1 0 36064 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1676037725
transform 1 0 35972 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1676037725
transform 1 0 32936 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1676037725
transform 1 0 36800 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1676037725
transform 1 0 36892 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1676037725
transform 1 0 36892 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1754_
timestamp 1676037725
transform 1 0 16928 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1676037725
transform 1 0 20700 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1676037725
transform 1 0 23920 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1676037725
transform 1 0 21988 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1676037725
transform 1 0 19596 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1759_
timestamp 1676037725
transform 1 0 15548 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1760_
timestamp 1676037725
transform 1 0 22448 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1676037725
transform 1 0 17480 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1676037725
transform 1 0 7912 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1676037725
transform 1 0 8004 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1676037725
transform 1 0 9752 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1676037725
transform 1 0 11684 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1676037725
transform 1 0 12972 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1676037725
transform 1 0 15916 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1676037725
transform 1 0 17112 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1770_
timestamp 1676037725
transform 1 0 18492 0 -1 35904
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1676037725
transform 1 0 8188 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1676037725
transform 1 0 30268 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1676037725
transform 1 0 19136 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1676037725
transform 1 0 7176 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1676037725
transform 1 0 7360 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1676037725
transform 1 0 7176 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1676037725
transform 1 0 19964 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1778_
timestamp 1676037725
transform 1 0 7636 0 -1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1779_
timestamp 1676037725
transform 1 0 7544 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1780_
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1676037725
transform 1 0 8372 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1676037725
transform 1 0 13892 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1676037725
transform 1 0 11776 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1676037725
transform 1 0 14996 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1676037725
transform 1 0 9936 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1676037725
transform 1 0 10948 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1676037725
transform 1 0 12880 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1788_
timestamp 1676037725
transform 1 0 12788 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1789_
timestamp 1676037725
transform 1 0 13432 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1676037725
transform 1 0 11408 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1791_
timestamp 1676037725
transform 1 0 10764 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1676037725
transform 1 0 12880 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1676037725
transform 1 0 9476 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1676037725
transform 1 0 16100 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1676037725
transform 1 0 14904 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1676037725
transform 1 0 15732 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1676037725
transform 1 0 15640 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1676037725
transform 1 0 15640 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1800_
timestamp 1676037725
transform 1 0 18124 0 -1 30464
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1676037725
transform 1 0 18124 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1676037725
transform 1 0 13616 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1676037725
transform 1 0 11684 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1676037725
transform 1 0 17204 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1676037725
transform 1 0 32292 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1806_
timestamp 1676037725
transform 1 0 31832 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1807_
timestamp 1676037725
transform 1 0 36892 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1808_
timestamp 1676037725
transform 1 0 36708 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1809_
timestamp 1676037725
transform 1 0 36800 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1810_
timestamp 1676037725
transform 1 0 36800 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1811_
timestamp 1676037725
transform 1 0 36800 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1812_
timestamp 1676037725
transform 1 0 36800 0 1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1813_
timestamp 1676037725
transform 1 0 36800 0 1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1814_
timestamp 1676037725
transform 1 0 35420 0 1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1676037725
transform 1 0 20792 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1676037725
transform 1 0 25208 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1676037725
transform 1 0 20976 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1676037725
transform 1 0 30360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1676037725
transform 1 0 29900 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1676037725
transform 1 0 29716 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1676037725
transform 1 0 29808 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1676037725
transform 1 0 24748 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1676037725
transform 1 0 22356 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1676037725
transform 1 0 34224 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1676037725
transform 1 0 32292 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1676037725
transform 1 0 32476 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1676037725
transform 1 0 27048 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22816 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1676037725
transform 1 0 12788 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1676037725
transform 1 0 17940 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1676037725
transform 1 0 18676 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1676037725
transform 1 0 14260 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1676037725
transform 1 0 14260 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1676037725
transform 1 0 19412 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1676037725
transform 1 0 17940 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1676037725
transform 1 0 26496 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1676037725
transform 1 0 25760 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1676037725
transform 1 0 30544 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1676037725
transform 1 0 30820 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1676037725
transform 1 0 32476 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1676037725
transform 1 0 32384 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1676037725
transform 1 0 31372 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1676037725
transform 1 0 32752 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37444 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35788 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36248 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1676037725
transform 1 0 23552 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout43
timestamp 1676037725
transform 1 0 32292 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_16  fanout44
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout45
timestamp 1676037725
transform 1 0 23184 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout46
timestamp 1676037725
transform 1 0 20976 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout47
timestamp 1676037725
transform 1 0 15548 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout48
timestamp 1676037725
transform 1 0 10396 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout49
timestamp 1676037725
transform 1 0 31280 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout50
timestamp 1676037725
transform 1 0 37444 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout51
timestamp 1676037725
transform 1 0 13248 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout52
timestamp 1676037725
transform 1 0 28244 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout53
timestamp 1676037725
transform 1 0 12880 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout54
timestamp 1676037725
transform 1 0 33856 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp 1676037725
transform 1 0 16652 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout56
timestamp 1676037725
transform 1 0 16836 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout57
timestamp 1676037725
transform 1 0 16836 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout58
timestamp 1676037725
transform 1 0 18124 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16008 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout60
timestamp 1676037725
transform 1 0 19412 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout61
timestamp 1676037725
transform 1 0 31004 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout62
timestamp 1676037725
transform 1 0 11960 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout63
timestamp 1676037725
transform 1 0 6532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout64
timestamp 1676037725
transform 1 0 19780 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  fanout65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23276 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  fanout66
timestamp 1676037725
transform 1 0 26036 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout67
timestamp 1676037725
transform 1 0 27140 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout68
timestamp 1676037725
transform 1 0 27600 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout69
timestamp 1676037725
transform 1 0 32936 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout70
timestamp 1676037725
transform 1 0 32476 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout71
timestamp 1676037725
transform 1 0 13800 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  fanout72
timestamp 1676037725
transform 1 0 31556 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  fanout73
timestamp 1676037725
transform 1 0 14260 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout74 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout75
timestamp 1676037725
transform 1 0 33764 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  fanout76
timestamp 1676037725
transform 1 0 28336 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout77
timestamp 1676037725
transform 1 0 23736 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout78
timestamp 1676037725
transform 1 0 31188 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout79
timestamp 1676037725
transform 1 0 31280 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout80
timestamp 1676037725
transform 1 0 18032 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout81
timestamp 1676037725
transform 1 0 27232 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout82
timestamp 1676037725
transform 1 0 28060 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 1676037725
transform 1 0 30636 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout84
timestamp 1676037725
transform 1 0 23552 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout85
timestamp 1676037725
transform 1 0 34868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout86
timestamp 1676037725
transform 1 0 22540 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout87
timestamp 1676037725
transform 1 0 27140 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout88
timestamp 1676037725
transform 1 0 23460 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout89
timestamp 1676037725
transform 1 0 29716 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout90
timestamp 1676037725
transform 1 0 22908 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1676037725
transform 1 0 1840 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input2
timestamp 1676037725
transform 1 0 5152 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input3
timestamp 1676037725
transform 1 0 7820 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input4
timestamp 1676037725
transform 1 0 10396 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  input5
timestamp 1676037725
transform 1 0 15088 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input6
timestamp 1676037725
transform 1 0 17940 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  input7
timestamp 1676037725
transform 1 0 21988 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input8
timestamp 1676037725
transform 1 0 25024 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1676037725
transform 1 0 5796 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform 1 0 4876 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input11
timestamp 1676037725
transform 1 0 37536 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform 1 0 20976 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1676037725
transform 1 0 37812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1676037725
transform 1 0 37812 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1676037725
transform 1 0 37812 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output16
timestamp 1676037725
transform 1 0 35512 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output17
timestamp 1676037725
transform 1 0 36432 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output18
timestamp 1676037725
transform 1 0 37812 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output19
timestamp 1676037725
transform 1 0 37812 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output20
timestamp 1676037725
transform 1 0 35972 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output21
timestamp 1676037725
transform 1 0 36432 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output22
timestamp 1676037725
transform 1 0 34684 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output23
timestamp 1676037725
transform 1 0 23828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output24
timestamp 1676037725
transform 1 0 37812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output25
timestamp 1676037725
transform 1 0 17020 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output26
timestamp 1676037725
transform 1 0 21620 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output27
timestamp 1676037725
transform 1 0 26128 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output28
timestamp 1676037725
transform 1 0 27600 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output29
timestamp 1676037725
transform 1 0 27416 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output30
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output31
timestamp 1676037725
transform 1 0 20608 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output32
timestamp 1676037725
transform 1 0 37812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output33
timestamp 1676037725
transform 1 0 37812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output34
timestamp 1676037725
transform 1 0 37812 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output35
timestamp 1676037725
transform 1 0 37812 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output36
timestamp 1676037725
transform 1 0 37812 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output37
timestamp 1676037725
transform 1 0 37812 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_91 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_92
timestamp 1676037725
transform 1 0 38088 0 1 13056
box -38 -48 314 592
<< labels >>
flabel metal2 s 34886 39200 34942 40000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 1766 39200 1822 40000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 5078 39200 5134 40000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 8390 39200 8446 40000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 11702 39200 11758 40000 0 FreeSans 224 90 0 0 io_in[3]
port 4 nsew signal input
flabel metal2 s 15014 39200 15070 40000 0 FreeSans 224 90 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 18326 39200 18382 40000 0 FreeSans 224 90 0 0 io_in[5]
port 6 nsew signal input
flabel metal2 s 21638 39200 21694 40000 0 FreeSans 224 90 0 0 io_in[6]
port 7 nsew signal input
flabel metal2 s 24950 39200 25006 40000 0 FreeSans 224 90 0 0 io_in[7]
port 8 nsew signal input
flabel metal2 s 28262 39200 28318 40000 0 FreeSans 224 90 0 0 io_in[8]
port 9 nsew signal input
flabel metal2 s 31574 39200 31630 40000 0 FreeSans 224 90 0 0 io_in[9]
port 10 nsew signal input
flabel metal3 s 39200 38224 40000 38344 0 FreeSans 480 0 0 0 io_oeb
port 11 nsew signal tristate
flabel metal3 s 39200 1504 40000 1624 0 FreeSans 480 0 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal3 s 39200 15104 40000 15224 0 FreeSans 480 0 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal3 s 39200 16464 40000 16584 0 FreeSans 480 0 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal3 s 39200 17824 40000 17944 0 FreeSans 480 0 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal3 s 39200 19184 40000 19304 0 FreeSans 480 0 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal3 s 39200 20544 40000 20664 0 FreeSans 480 0 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal3 s 39200 21904 40000 22024 0 FreeSans 480 0 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal3 s 39200 23264 40000 23384 0 FreeSans 480 0 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal3 s 39200 24624 40000 24744 0 FreeSans 480 0 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal3 s 39200 25984 40000 26104 0 FreeSans 480 0 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal3 s 39200 27344 40000 27464 0 FreeSans 480 0 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal3 s 39200 2864 40000 2984 0 FreeSans 480 0 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal3 s 39200 28704 40000 28824 0 FreeSans 480 0 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal3 s 39200 30064 40000 30184 0 FreeSans 480 0 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal3 s 39200 31424 40000 31544 0 FreeSans 480 0 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal3 s 39200 32784 40000 32904 0 FreeSans 480 0 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal3 s 39200 34144 40000 34264 0 FreeSans 480 0 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal3 s 39200 35504 40000 35624 0 FreeSans 480 0 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal3 s 39200 36864 40000 36984 0 FreeSans 480 0 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal3 s 39200 4224 40000 4344 0 FreeSans 480 0 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal3 s 39200 5584 40000 5704 0 FreeSans 480 0 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal3 s 39200 6944 40000 7064 0 FreeSans 480 0 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal3 s 39200 8304 40000 8424 0 FreeSans 480 0 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal3 s 39200 9664 40000 9784 0 FreeSans 480 0 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal3 s 39200 11024 40000 11144 0 FreeSans 480 0 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal3 s 39200 12384 40000 12504 0 FreeSans 480 0 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal3 s 39200 13744 40000 13864 0 FreeSans 480 0 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal2 s 38198 39200 38254 40000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
