// This is the unpowered netlist.
module tt2_tholin_diceroll (clk,
    io_in,
    rst,
    io_out);
 input clk;
 input io_in;
 input rst;
 output [7:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire \dice.bcd[0] ;
 wire \dice.bcd[1] ;
 wire \dice.bcd[2] ;
 wire \dice.clkdiv[0] ;
 wire \dice.clkdiv[1] ;
 wire \dice.clkdiv[2] ;
 wire \dice.clkdiv[3] ;
 wire \dice.clkdiv[4] ;
 wire \dice.clkdiv[5] ;
 wire \dice.clkdiv[6] ;
 wire \dice.clkdiv[7] ;
 wire \dice.counter[0] ;
 wire \dice.counter[10] ;
 wire \dice.counter[11] ;
 wire \dice.counter[12] ;
 wire \dice.counter[13] ;
 wire \dice.counter[14] ;
 wire \dice.counter[15] ;
 wire \dice.counter[1] ;
 wire \dice.counter[2] ;
 wire \dice.counter[3] ;
 wire \dice.counter[4] ;
 wire \dice.counter[5] ;
 wire \dice.counter[6] ;
 wire \dice.counter[7] ;
 wire \dice.counter[8] ;
 wire \dice.counter[9] ;
 wire \dice.lfsr[0] ;
 wire \dice.lfsr[10] ;
 wire \dice.lfsr[11] ;
 wire \dice.lfsr[12] ;
 wire \dice.lfsr[13] ;
 wire \dice.lfsr[14] ;
 wire \dice.lfsr[15] ;
 wire \dice.lfsr[1] ;
 wire \dice.lfsr[2] ;
 wire \dice.lfsr[3] ;
 wire \dice.lfsr[4] ;
 wire \dice.lfsr[5] ;
 wire \dice.lfsr[6] ;
 wire \dice.lfsr[7] ;
 wire \dice.lfsr[8] ;
 wire \dice.lfsr[9] ;
 wire \dice.r_counter[0] ;
 wire \dice.r_counter[1] ;
 wire \dice.r_counter[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__nand2_1 _252_ (.A(\dice.r_counter[0] ),
    .B(\dice.lfsr[0] ),
    .Y(_054_));
 sky130_fd_sc_hd__xor2_1 _253_ (.A(\dice.lfsr[1] ),
    .B(\dice.r_counter[1] ),
    .X(_055_));
 sky130_fd_sc_hd__xnor2_1 _254_ (.A(_054_),
    .B(_055_),
    .Y(_056_));
 sky130_fd_sc_hd__and2_1 _255_ (.A(\dice.lfsr[1] ),
    .B(\dice.r_counter[1] ),
    .X(_057_));
 sky130_fd_sc_hd__a31o_1 _256_ (.A1(\dice.r_counter[0] ),
    .A2(\dice.lfsr[0] ),
    .A3(_055_),
    .B1(_057_),
    .X(_058_));
 sky130_fd_sc_hd__xor2_1 _257_ (.A(\dice.r_counter[2] ),
    .B(\dice.lfsr[2] ),
    .X(_059_));
 sky130_fd_sc_hd__xnor2_1 _258_ (.A(_058_),
    .B(_059_),
    .Y(_060_));
 sky130_fd_sc_hd__or2_1 _259_ (.A(_056_),
    .B(_060_),
    .X(_061_));
 sky130_fd_sc_hd__inv_2 _260_ (.A(net1),
    .Y(_062_));
 sky130_fd_sc_hd__and2_1 _261_ (.A(_062_),
    .B(\dice.clkdiv[3] ),
    .X(_063_));
 sky130_fd_sc_hd__and4b_1 _262_ (.A_N(net1),
    .B(\dice.counter[0] ),
    .C(\dice.counter[1] ),
    .D(\dice.counter[2] ),
    .X(_064_));
 sky130_fd_sc_hd__buf_2 _263_ (.A(net1),
    .X(_065_));
 sky130_fd_sc_hd__nor2b_1 _264_ (.A(_065_),
    .B_N(\dice.counter[3] ),
    .Y(_066_));
 sky130_fd_sc_hd__xnor2_1 _265_ (.A(_064_),
    .B(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__xnor2_1 _266_ (.A(_063_),
    .B(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__or2b_1 _267_ (.A(net1),
    .B_N(\dice.counter[2] ),
    .X(_069_));
 sky130_fd_sc_hd__and3b_1 _268_ (.A_N(net1),
    .B(\dice.counter[0] ),
    .C(\dice.counter[1] ),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _269_ (.A0(_069_),
    .A1(\dice.counter[2] ),
    .S(_070_),
    .X(_071_));
 sky130_fd_sc_hd__and2_1 _270_ (.A(_062_),
    .B(\dice.clkdiv[2] ),
    .X(_072_));
 sky130_fd_sc_hd__clkbuf_2 _271_ (.A(_072_),
    .X(_073_));
 sky130_fd_sc_hd__xnor2_1 _272_ (.A(_071_),
    .B(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__or2b_1 _273_ (.A(_065_),
    .B_N(\dice.counter[0] ),
    .X(_075_));
 sky130_fd_sc_hd__nor2b_2 _274_ (.A(_065_),
    .B_N(\dice.clkdiv[0] ),
    .Y(_076_));
 sky130_fd_sc_hd__mux2_1 _275_ (.A0(_075_),
    .A1(\dice.counter[0] ),
    .S(_076_),
    .X(_077_));
 sky130_fd_sc_hd__buf_2 _276_ (.A(_065_),
    .X(_078_));
 sky130_fd_sc_hd__or2_1 _277_ (.A(_078_),
    .B(\dice.clkdiv[1] ),
    .X(_079_));
 sky130_fd_sc_hd__nor2_1 _278_ (.A(\dice.counter[0] ),
    .B(\dice.counter[1] ),
    .Y(_080_));
 sky130_fd_sc_hd__or3_1 _279_ (.A(_078_),
    .B(_070_),
    .C(_080_),
    .X(_081_));
 sky130_fd_sc_hd__xnor2_1 _280_ (.A(_079_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__or4_1 _281_ (.A(_068_),
    .B(_074_),
    .C(_077_),
    .D(_082_),
    .X(_083_));
 sky130_fd_sc_hd__inv_2 _282_ (.A(\dice.counter[4] ),
    .Y(_084_));
 sky130_fd_sc_hd__clkinv_2 _283_ (.A(\dice.counter[5] ),
    .Y(_085_));
 sky130_fd_sc_hd__nand4b_1 _284_ (.A_N(net1),
    .B(\dice.counter[0] ),
    .C(\dice.counter[1] ),
    .D(\dice.counter[2] ),
    .Y(_086_));
 sky130_fd_sc_hd__or2b_1 _285_ (.A(_065_),
    .B_N(\dice.counter[3] ),
    .X(_087_));
 sky130_fd_sc_hd__or4_2 _286_ (.A(_084_),
    .B(_085_),
    .C(_086_),
    .D(_087_),
    .X(_088_));
 sky130_fd_sc_hd__buf_2 _287_ (.A(_062_),
    .X(_089_));
 sky130_fd_sc_hd__a32o_1 _288_ (.A1(\dice.counter[4] ),
    .A2(_064_),
    .A3(_066_),
    .B1(\dice.counter[5] ),
    .B2(_089_),
    .X(_090_));
 sky130_fd_sc_hd__nand2_1 _289_ (.A(_062_),
    .B(\dice.clkdiv[5] ),
    .Y(_091_));
 sky130_fd_sc_hd__a21oi_1 _290_ (.A1(_088_),
    .A2(_090_),
    .B1(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__and3_1 _291_ (.A(_088_),
    .B(_090_),
    .C(_091_),
    .X(_093_));
 sky130_fd_sc_hd__nor2_1 _292_ (.A(_092_),
    .B(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__or3_1 _293_ (.A(_084_),
    .B(_086_),
    .C(_087_),
    .X(_095_));
 sky130_fd_sc_hd__a22o_1 _294_ (.A1(_089_),
    .A2(\dice.counter[4] ),
    .B1(_064_),
    .B2(_066_),
    .X(_096_));
 sky130_fd_sc_hd__and2_1 _295_ (.A(_089_),
    .B(\dice.clkdiv[4] ),
    .X(_097_));
 sky130_fd_sc_hd__a21o_1 _296_ (.A1(_095_),
    .A2(_096_),
    .B1(_097_),
    .X(_098_));
 sky130_fd_sc_hd__nand3_1 _297_ (.A(\dice.clkdiv[4] ),
    .B(_095_),
    .C(_096_),
    .Y(_099_));
 sky130_fd_sc_hd__nand2_1 _298_ (.A(_098_),
    .B(_099_),
    .Y(_100_));
 sky130_fd_sc_hd__and2_1 _299_ (.A(_062_),
    .B(\dice.counter[12] ),
    .X(_101_));
 sky130_fd_sc_hd__nor2b_1 _300_ (.A(_078_),
    .B_N(\dice.counter[14] ),
    .Y(_102_));
 sky130_fd_sc_hd__and2b_1 _301_ (.A_N(_065_),
    .B(\dice.counter[13] ),
    .X(_103_));
 sky130_fd_sc_hd__and2b_1 _302_ (.A_N(_065_),
    .B(\dice.counter[8] ),
    .X(_104_));
 sky130_fd_sc_hd__o21ba_1 _303_ (.A1(\dice.counter[10] ),
    .A2(\dice.counter[15] ),
    .B1_N(_065_),
    .X(_105_));
 sky130_fd_sc_hd__o21ba_1 _304_ (.A1(\dice.counter[9] ),
    .A2(\dice.counter[11] ),
    .B1_N(_065_),
    .X(_106_));
 sky130_fd_sc_hd__or4_1 _305_ (.A(_103_),
    .B(_104_),
    .C(_105_),
    .D(_106_),
    .X(_107_));
 sky130_fd_sc_hd__nor3_1 _306_ (.A(_101_),
    .B(_102_),
    .C(_107_),
    .Y(_108_));
 sky130_fd_sc_hd__and4b_1 _307_ (.A_N(_078_),
    .B(\dice.counter[9] ),
    .C(\dice.counter[10] ),
    .D(\dice.counter[11] ),
    .X(_109_));
 sky130_fd_sc_hd__and3_1 _308_ (.A(\dice.counter[8] ),
    .B(\dice.counter[15] ),
    .C(_103_),
    .X(_110_));
 sky130_fd_sc_hd__and4_1 _309_ (.A(\dice.counter[12] ),
    .B(_102_),
    .C(_109_),
    .D(_110_),
    .X(_111_));
 sky130_fd_sc_hd__inv_2 _310_ (.A(\dice.counter[7] ),
    .Y(_112_));
 sky130_fd_sc_hd__and2b_1 _311_ (.A_N(_078_),
    .B(\dice.counter[6] ),
    .X(_113_));
 sky130_fd_sc_hd__nor3b_1 _312_ (.A(_112_),
    .B(_088_),
    .C_N(_113_),
    .Y(_114_));
 sky130_fd_sc_hd__mux2_1 _313_ (.A0(_108_),
    .A1(_111_),
    .S(_114_),
    .X(_115_));
 sky130_fd_sc_hd__and4b_1 _314_ (.A_N(_083_),
    .B(_094_),
    .C(_100_),
    .D(_115_),
    .X(_116_));
 sky130_fd_sc_hd__nand3b_1 _315_ (.A_N(_065_),
    .B(\dice.counter[5] ),
    .C(\dice.counter[6] ),
    .Y(_117_));
 sky130_fd_sc_hd__or4_2 _316_ (.A(_084_),
    .B(_086_),
    .C(_087_),
    .D(_117_),
    .X(_118_));
 sky130_fd_sc_hd__a41o_1 _317_ (.A1(\dice.counter[4] ),
    .A2(\dice.counter[5] ),
    .A3(_064_),
    .A4(_066_),
    .B1(_113_),
    .X(_119_));
 sky130_fd_sc_hd__nand3_1 _318_ (.A(\dice.clkdiv[6] ),
    .B(_118_),
    .C(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__and2_1 _319_ (.A(_089_),
    .B(\dice.clkdiv[6] ),
    .X(_121_));
 sky130_fd_sc_hd__a21o_1 _320_ (.A1(_118_),
    .A2(_119_),
    .B1(_121_),
    .X(_122_));
 sky130_fd_sc_hd__inv_2 _321_ (.A(\dice.clkdiv[7] ),
    .Y(_123_));
 sky130_fd_sc_hd__nor2_1 _322_ (.A(_078_),
    .B(_123_),
    .Y(_124_));
 sky130_fd_sc_hd__nand2_1 _323_ (.A(_089_),
    .B(\dice.counter[7] ),
    .Y(_125_));
 sky130_fd_sc_hd__mux2_1 _324_ (.A0(\dice.counter[7] ),
    .A1(_125_),
    .S(_118_),
    .X(_126_));
 sky130_fd_sc_hd__xnor2_1 _325_ (.A(_124_),
    .B(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__a21oi_2 _326_ (.A1(_120_),
    .A2(_122_),
    .B1(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__or3_1 _327_ (.A(\dice.clkdiv[1] ),
    .B(\dice.clkdiv[3] ),
    .C(_076_),
    .X(_129_));
 sky130_fd_sc_hd__or3_1 _328_ (.A(_091_),
    .B(_073_),
    .C(_129_),
    .X(_130_));
 sky130_fd_sc_hd__or4_1 _329_ (.A(\dice.clkdiv[4] ),
    .B(\dice.clkdiv[6] ),
    .C(_123_),
    .D(_130_),
    .X(_131_));
 sky130_fd_sc_hd__buf_2 _330_ (.A(_131_),
    .X(_132_));
 sky130_fd_sc_hd__or2_1 _331_ (.A(\dice.r_counter[0] ),
    .B(\dice.lfsr[0] ),
    .X(_133_));
 sky130_fd_sc_hd__and3_1 _332_ (.A(_054_),
    .B(_055_),
    .C(_133_),
    .X(_134_));
 sky130_fd_sc_hd__nand2_1 _333_ (.A(_060_),
    .B(_134_),
    .Y(_135_));
 sky130_fd_sc_hd__and4_1 _334_ (.A(_116_),
    .B(_128_),
    .C(_132_),
    .D(_135_),
    .X(_136_));
 sky130_fd_sc_hd__a31oi_2 _335_ (.A1(_116_),
    .A2(_128_),
    .A3(_132_),
    .B1(\dice.bcd[2] ),
    .Y(_137_));
 sky130_fd_sc_hd__clkbuf_4 _336_ (.A(net2),
    .X(_138_));
 sky130_fd_sc_hd__a211oi_4 _337_ (.A1(_061_),
    .A2(_136_),
    .B1(_137_),
    .C1(_138_),
    .Y(_052_));
 sky130_fd_sc_hd__and2_1 _338_ (.A(_054_),
    .B(_133_),
    .X(_139_));
 sky130_fd_sc_hd__nor2_1 _339_ (.A(_056_),
    .B(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__clkinv_2 _340_ (.A(_139_),
    .Y(_141_));
 sky130_fd_sc_hd__mux2_1 _341_ (.A0(_134_),
    .A1(_141_),
    .S(_060_),
    .X(_142_));
 sky130_fd_sc_hd__or2_1 _342_ (.A(_140_),
    .B(_142_),
    .X(_143_));
 sky130_fd_sc_hd__and3_1 _343_ (.A(_116_),
    .B(_128_),
    .C(_132_),
    .X(_144_));
 sky130_fd_sc_hd__mux2_1 _344_ (.A0(\dice.bcd[0] ),
    .A1(_143_),
    .S(_144_),
    .X(_145_));
 sky130_fd_sc_hd__inv_2 _345_ (.A(\dice.bcd[1] ),
    .Y(_146_));
 sky130_fd_sc_hd__a31o_1 _346_ (.A1(_116_),
    .A2(_128_),
    .A3(_132_),
    .B1(_146_),
    .X(_147_));
 sky130_fd_sc_hd__clkinv_2 _347_ (.A(_135_),
    .Y(_148_));
 sky130_fd_sc_hd__or3b_1 _348_ (.A(_097_),
    .B(_073_),
    .C_N(_124_),
    .X(_149_));
 sky130_fd_sc_hd__nor2_1 _349_ (.A(_091_),
    .B(_121_),
    .Y(_150_));
 sky130_fd_sc_hd__nor2_1 _350_ (.A(_063_),
    .B(_076_),
    .Y(_151_));
 sky130_fd_sc_hd__and4bb_2 _351_ (.A_N(_079_),
    .B_N(_149_),
    .C(_150_),
    .D(_151_),
    .X(_152_));
 sky130_fd_sc_hd__or3_1 _352_ (.A(_101_),
    .B(_102_),
    .C(_107_),
    .X(_153_));
 sky130_fd_sc_hd__nor4_1 _353_ (.A(_084_),
    .B(_086_),
    .C(_087_),
    .D(_117_),
    .Y(_154_));
 sky130_fd_sc_hd__nand2_1 _354_ (.A(\dice.counter[7] ),
    .B(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__nand2_1 _355_ (.A(\dice.counter[12] ),
    .B(_102_),
    .Y(_156_));
 sky130_fd_sc_hd__or2b_1 _356_ (.A(_078_),
    .B_N(\dice.counter[15] ),
    .X(_157_));
 sky130_fd_sc_hd__and3b_1 _357_ (.A_N(_078_),
    .B(\dice.counter[8] ),
    .C(\dice.counter[13] ),
    .X(_158_));
 sky130_fd_sc_hd__nand3b_1 _358_ (.A_N(_157_),
    .B(_109_),
    .C(_158_),
    .Y(_159_));
 sky130_fd_sc_hd__o211a_1 _359_ (.A1(_156_),
    .A2(_159_),
    .B1(\dice.counter[7] ),
    .C1(_154_),
    .X(_160_));
 sky130_fd_sc_hd__nor2_1 _360_ (.A(_071_),
    .B(_073_),
    .Y(_161_));
 sky130_fd_sc_hd__a2111o_1 _361_ (.A1(_153_),
    .A2(_155_),
    .B1(_160_),
    .C1(_161_),
    .D1(_082_),
    .X(_162_));
 sky130_fd_sc_hd__a31o_1 _362_ (.A1(_089_),
    .A2(\dice.clkdiv[2] ),
    .A3(_071_),
    .B1(_077_),
    .X(_163_));
 sky130_fd_sc_hd__a211o_1 _363_ (.A1(_098_),
    .A2(_099_),
    .B1(_068_),
    .C1(_163_),
    .X(_164_));
 sky130_fd_sc_hd__a211o_1 _364_ (.A1(_120_),
    .A2(_122_),
    .B1(_092_),
    .C1(_093_),
    .X(_165_));
 sky130_fd_sc_hd__nor4_2 _365_ (.A(_127_),
    .B(_162_),
    .C(_164_),
    .D(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__or4b_1 _366_ (.A(_148_),
    .B(_152_),
    .C(_140_),
    .D_N(_166_),
    .X(_167_));
 sky130_fd_sc_hd__a21oi_1 _367_ (.A1(_147_),
    .A2(_167_),
    .B1(_138_),
    .Y(_051_));
 sky130_fd_sc_hd__and2b_1 _368_ (.A_N(_052_),
    .B(_051_),
    .X(_168_));
 sky130_fd_sc_hd__clkbuf_4 _369_ (.A(_138_),
    .X(_169_));
 sky130_fd_sc_hd__nor3_1 _370_ (.A(_169_),
    .B(_052_),
    .C(_145_),
    .Y(_170_));
 sky130_fd_sc_hd__a211o_1 _371_ (.A1(_052_),
    .A2(_145_),
    .B1(_168_),
    .C1(_170_),
    .X(_000_));
 sky130_fd_sc_hd__a21boi_1 _372_ (.A1(_145_),
    .A2(_051_),
    .B1_N(_052_),
    .Y(_171_));
 sky130_fd_sc_hd__nand2_1 _373_ (.A(_147_),
    .B(_167_),
    .Y(_172_));
 sky130_fd_sc_hd__or3_1 _374_ (.A(_138_),
    .B(_145_),
    .C(_172_),
    .X(_173_));
 sky130_fd_sc_hd__a211o_1 _375_ (.A1(_171_),
    .A2(_173_),
    .B1(_168_),
    .C1(_170_),
    .X(_001_));
 sky130_fd_sc_hd__or2_1 _376_ (.A(_138_),
    .B(_145_),
    .X(_174_));
 sky130_fd_sc_hd__clkbuf_1 _377_ (.A(_174_),
    .X(_050_));
 sky130_fd_sc_hd__a31oi_1 _378_ (.A1(_052_),
    .A2(_147_),
    .A3(_167_),
    .B1(_050_),
    .Y(_002_));
 sky130_fd_sc_hd__a21bo_1 _379_ (.A1(_145_),
    .A2(_051_),
    .B1_N(_052_),
    .X(_175_));
 sky130_fd_sc_hd__nand2_1 _380_ (.A(_175_),
    .B(_173_),
    .Y(_003_));
 sky130_fd_sc_hd__or2b_1 _381_ (.A(_052_),
    .B_N(_051_),
    .X(_176_));
 sky130_fd_sc_hd__nand2_1 _382_ (.A(_176_),
    .B(_175_),
    .Y(_004_));
 sky130_fd_sc_hd__nand2_1 _383_ (.A(_171_),
    .B(_173_),
    .Y(_005_));
 sky130_fd_sc_hd__clkbuf_4 _384_ (.A(_169_),
    .X(_177_));
 sky130_fd_sc_hd__nor2_1 _385_ (.A(\dice.r_counter[0] ),
    .B(_177_),
    .Y(_006_));
 sky130_fd_sc_hd__clkbuf_4 _386_ (.A(_138_),
    .X(_178_));
 sky130_fd_sc_hd__a21oi_1 _387_ (.A1(\dice.r_counter[0] ),
    .A2(\dice.r_counter[1] ),
    .B1(_178_),
    .Y(_179_));
 sky130_fd_sc_hd__o21a_1 _388_ (.A1(\dice.r_counter[0] ),
    .A2(\dice.r_counter[1] ),
    .B1(_179_),
    .X(_007_));
 sky130_fd_sc_hd__a21oi_1 _389_ (.A1(\dice.r_counter[0] ),
    .A2(\dice.r_counter[1] ),
    .B1(\dice.r_counter[2] ),
    .Y(_180_));
 sky130_fd_sc_hd__a31o_1 _390_ (.A1(\dice.r_counter[0] ),
    .A2(\dice.r_counter[2] ),
    .A3(\dice.r_counter[1] ),
    .B1(_169_),
    .X(_181_));
 sky130_fd_sc_hd__nor2_1 _391_ (.A(_180_),
    .B(_181_),
    .Y(_008_));
 sky130_fd_sc_hd__a211o_1 _392_ (.A1(net10),
    .A2(_089_),
    .B1(_177_),
    .C1(_152_),
    .X(_009_));
 sky130_fd_sc_hd__and2_1 _393_ (.A(_116_),
    .B(_128_),
    .X(_182_));
 sky130_fd_sc_hd__a21oi_1 _394_ (.A1(_076_),
    .A2(_182_),
    .B1(_178_),
    .Y(_183_));
 sky130_fd_sc_hd__o21a_1 _395_ (.A1(_076_),
    .A2(_144_),
    .B1(_183_),
    .X(_010_));
 sky130_fd_sc_hd__a21oi_1 _396_ (.A1(_076_),
    .A2(_166_),
    .B1(_079_),
    .Y(_184_));
 sky130_fd_sc_hd__and3_1 _397_ (.A(_079_),
    .B(_076_),
    .C(_166_),
    .X(_185_));
 sky130_fd_sc_hd__nor3_1 _398_ (.A(_177_),
    .B(_184_),
    .C(_185_),
    .Y(_011_));
 sky130_fd_sc_hd__and4_1 _399_ (.A(\dice.clkdiv[1] ),
    .B(_073_),
    .C(_076_),
    .D(_182_),
    .X(_186_));
 sky130_fd_sc_hd__clkbuf_2 _400_ (.A(_186_),
    .X(_187_));
 sky130_fd_sc_hd__nor2_1 _401_ (.A(_178_),
    .B(_187_),
    .Y(_188_));
 sky130_fd_sc_hd__o21a_1 _402_ (.A1(_073_),
    .A2(_185_),
    .B1(_188_),
    .X(_012_));
 sky130_fd_sc_hd__nand2_1 _403_ (.A(\dice.clkdiv[3] ),
    .B(_187_),
    .Y(_189_));
 sky130_fd_sc_hd__inv_2 _404_ (.A(_138_),
    .Y(_190_));
 sky130_fd_sc_hd__buf_2 _405_ (.A(_190_),
    .X(_191_));
 sky130_fd_sc_hd__o211a_1 _406_ (.A1(_063_),
    .A2(_187_),
    .B1(_189_),
    .C1(_191_),
    .X(_013_));
 sky130_fd_sc_hd__a31o_1 _407_ (.A1(\dice.clkdiv[3] ),
    .A2(_073_),
    .A3(_185_),
    .B1(_097_),
    .X(_192_));
 sky130_fd_sc_hd__and2_1 _408_ (.A(\dice.clkdiv[4] ),
    .B(_063_),
    .X(_193_));
 sky130_fd_sc_hd__a21oi_1 _409_ (.A1(_187_),
    .A2(_193_),
    .B1(_138_),
    .Y(_194_));
 sky130_fd_sc_hd__and2_1 _410_ (.A(_192_),
    .B(_194_),
    .X(_195_));
 sky130_fd_sc_hd__clkbuf_1 _411_ (.A(_195_),
    .X(_014_));
 sky130_fd_sc_hd__and4_1 _412_ (.A(\dice.clkdiv[5] ),
    .B(_190_),
    .C(_187_),
    .D(_193_),
    .X(_196_));
 sky130_fd_sc_hd__a21oi_1 _413_ (.A1(_091_),
    .A2(_194_),
    .B1(_196_),
    .Y(_015_));
 sky130_fd_sc_hd__and4_1 _414_ (.A(\dice.clkdiv[5] ),
    .B(_073_),
    .C(_185_),
    .D(_193_),
    .X(_197_));
 sky130_fd_sc_hd__a41o_1 _415_ (.A1(\dice.clkdiv[5] ),
    .A2(_121_),
    .A3(_187_),
    .A4(_193_),
    .B1(_169_),
    .X(_198_));
 sky130_fd_sc_hd__o21ba_1 _416_ (.A1(_121_),
    .A2(_197_),
    .B1_N(_198_),
    .X(_016_));
 sky130_fd_sc_hd__a211oi_1 _417_ (.A1(\dice.clkdiv[6] ),
    .A2(_197_),
    .B1(_123_),
    .C1(_078_),
    .Y(_199_));
 sky130_fd_sc_hd__a31o_1 _418_ (.A1(_123_),
    .A2(_121_),
    .A3(_197_),
    .B1(_138_),
    .X(_200_));
 sky130_fd_sc_hd__or2_1 _419_ (.A(_199_),
    .B(_200_),
    .X(_201_));
 sky130_fd_sc_hd__clkbuf_1 _420_ (.A(_201_),
    .X(_017_));
 sky130_fd_sc_hd__nand2b_2 _421_ (.A_N(_182_),
    .B(_132_),
    .Y(_202_));
 sky130_fd_sc_hd__nand2_1 _422_ (.A(_075_),
    .B(_202_),
    .Y(_203_));
 sky130_fd_sc_hd__o211a_1 _423_ (.A1(_075_),
    .A2(_152_),
    .B1(_203_),
    .C1(_191_),
    .X(_018_));
 sky130_fd_sc_hd__nor2_1 _424_ (.A(_081_),
    .B(_166_),
    .Y(_204_));
 sky130_fd_sc_hd__inv_2 _425_ (.A(\dice.counter[0] ),
    .Y(_205_));
 sky130_fd_sc_hd__nor2_1 _426_ (.A(_205_),
    .B(_132_),
    .Y(_206_));
 sky130_fd_sc_hd__nand2_1 _427_ (.A(_204_),
    .B(_206_),
    .Y(_207_));
 sky130_fd_sc_hd__o211a_1 _428_ (.A1(_204_),
    .A2(_206_),
    .B1(_207_),
    .C1(_191_),
    .X(_019_));
 sky130_fd_sc_hd__or2_1 _429_ (.A(_069_),
    .B(_132_),
    .X(_208_));
 sky130_fd_sc_hd__o21a_1 _430_ (.A1(_071_),
    .A2(_202_),
    .B1(_208_),
    .X(_209_));
 sky130_fd_sc_hd__nor2_1 _431_ (.A(_177_),
    .B(_209_),
    .Y(_020_));
 sky130_fd_sc_hd__o2bb2a_1 _432_ (.A1_N(\dice.counter[3] ),
    .A2_N(_152_),
    .B1(_202_),
    .B2(_067_),
    .X(_210_));
 sky130_fd_sc_hd__nor2_1 _433_ (.A(_177_),
    .B(_210_),
    .Y(_021_));
 sky130_fd_sc_hd__nand2_1 _434_ (.A(_095_),
    .B(_096_),
    .Y(_211_));
 sky130_fd_sc_hd__o2bb2a_1 _435_ (.A1_N(\dice.counter[4] ),
    .A2_N(_152_),
    .B1(_202_),
    .B2(_211_),
    .X(_212_));
 sky130_fd_sc_hd__nor2_1 _436_ (.A(_177_),
    .B(_212_),
    .Y(_022_));
 sky130_fd_sc_hd__nand2_1 _437_ (.A(_088_),
    .B(_090_),
    .Y(_213_));
 sky130_fd_sc_hd__o2bb2a_1 _438_ (.A1_N(\dice.counter[5] ),
    .A2_N(_152_),
    .B1(_202_),
    .B2(_213_),
    .X(_214_));
 sky130_fd_sc_hd__nor2_1 _439_ (.A(_177_),
    .B(_214_),
    .Y(_023_));
 sky130_fd_sc_hd__nand2_1 _440_ (.A(_118_),
    .B(_119_),
    .Y(_215_));
 sky130_fd_sc_hd__o2bb2a_1 _441_ (.A1_N(\dice.counter[6] ),
    .A2_N(_152_),
    .B1(_202_),
    .B2(_215_),
    .X(_216_));
 sky130_fd_sc_hd__nor2_1 _442_ (.A(_177_),
    .B(_216_),
    .Y(_024_));
 sky130_fd_sc_hd__o2bb2a_1 _443_ (.A1_N(\dice.counter[7] ),
    .A2_N(_152_),
    .B1(_202_),
    .B2(_126_),
    .X(_217_));
 sky130_fd_sc_hd__nor2_1 _444_ (.A(_177_),
    .B(_217_),
    .Y(_025_));
 sky130_fd_sc_hd__a21oi_1 _445_ (.A1(_114_),
    .A2(_132_),
    .B1(_104_),
    .Y(_218_));
 sky130_fd_sc_hd__and4b_1 _446_ (.A_N(_152_),
    .B(_154_),
    .C(_104_),
    .D(\dice.counter[7] ),
    .X(_219_));
 sky130_fd_sc_hd__clkbuf_2 _447_ (.A(_219_),
    .X(_220_));
 sky130_fd_sc_hd__nor3_1 _448_ (.A(_178_),
    .B(_218_),
    .C(_220_),
    .Y(_026_));
 sky130_fd_sc_hd__a21o_1 _449_ (.A1(_089_),
    .A2(\dice.counter[9] ),
    .B1(_220_),
    .X(_221_));
 sky130_fd_sc_hd__nand2_1 _450_ (.A(\dice.counter[9] ),
    .B(_220_),
    .Y(_222_));
 sky130_fd_sc_hd__and3_1 _451_ (.A(_190_),
    .B(_221_),
    .C(_222_),
    .X(_223_));
 sky130_fd_sc_hd__clkbuf_1 _452_ (.A(_223_),
    .X(_027_));
 sky130_fd_sc_hd__a22o_1 _453_ (.A1(_089_),
    .A2(\dice.counter[10] ),
    .B1(_220_),
    .B2(\dice.counter[9] ),
    .X(_224_));
 sky130_fd_sc_hd__or3b_1 _454_ (.A(_222_),
    .B(_078_),
    .C_N(\dice.counter[10] ),
    .X(_225_));
 sky130_fd_sc_hd__and3_1 _455_ (.A(_190_),
    .B(_224_),
    .C(_225_),
    .X(_226_));
 sky130_fd_sc_hd__clkbuf_1 _456_ (.A(_226_),
    .X(_028_));
 sky130_fd_sc_hd__nand2_1 _457_ (.A(_089_),
    .B(\dice.counter[11] ),
    .Y(_227_));
 sky130_fd_sc_hd__a21o_1 _458_ (.A1(_109_),
    .A2(_220_),
    .B1(_169_),
    .X(_228_));
 sky130_fd_sc_hd__a21oi_1 _459_ (.A1(_227_),
    .A2(_225_),
    .B1(_228_),
    .Y(_029_));
 sky130_fd_sc_hd__a21oi_1 _460_ (.A1(_109_),
    .A2(_220_),
    .B1(_101_),
    .Y(_229_));
 sky130_fd_sc_hd__and3_1 _461_ (.A(_101_),
    .B(_109_),
    .C(_220_),
    .X(_230_));
 sky130_fd_sc_hd__nor3_1 _462_ (.A(_178_),
    .B(_229_),
    .C(_230_),
    .Y(_030_));
 sky130_fd_sc_hd__nor2_1 _463_ (.A(_103_),
    .B(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__a211oi_1 _464_ (.A1(\dice.counter[13] ),
    .A2(_230_),
    .B1(_231_),
    .C1(_178_),
    .Y(_031_));
 sky130_fd_sc_hd__a21oi_1 _465_ (.A1(\dice.counter[13] ),
    .A2(_230_),
    .B1(_102_),
    .Y(_232_));
 sky130_fd_sc_hd__and3_1 _466_ (.A(\dice.counter[13] ),
    .B(_102_),
    .C(_230_),
    .X(_233_));
 sky130_fd_sc_hd__nor3_1 _467_ (.A(_178_),
    .B(_232_),
    .C(_233_),
    .Y(_032_));
 sky130_fd_sc_hd__mux2_1 _468_ (.A0(_157_),
    .A1(\dice.counter[15] ),
    .S(_233_),
    .X(_234_));
 sky130_fd_sc_hd__nor2_1 _469_ (.A(_177_),
    .B(_234_),
    .Y(_033_));
 sky130_fd_sc_hd__and2_1 _470_ (.A(\dice.lfsr[1] ),
    .B(_191_),
    .X(_235_));
 sky130_fd_sc_hd__clkbuf_1 _471_ (.A(_235_),
    .X(_034_));
 sky130_fd_sc_hd__or2_1 _472_ (.A(\dice.lfsr[2] ),
    .B(_169_),
    .X(_236_));
 sky130_fd_sc_hd__clkbuf_1 _473_ (.A(_236_),
    .X(_035_));
 sky130_fd_sc_hd__and2_1 _474_ (.A(_191_),
    .B(\dice.lfsr[3] ),
    .X(_237_));
 sky130_fd_sc_hd__clkbuf_1 _475_ (.A(_237_),
    .X(_036_));
 sky130_fd_sc_hd__or2_1 _476_ (.A(_169_),
    .B(\dice.lfsr[4] ),
    .X(_238_));
 sky130_fd_sc_hd__clkbuf_1 _477_ (.A(_238_),
    .X(_037_));
 sky130_fd_sc_hd__or2_1 _478_ (.A(_169_),
    .B(\dice.lfsr[5] ),
    .X(_239_));
 sky130_fd_sc_hd__clkbuf_1 _479_ (.A(_239_),
    .X(_038_));
 sky130_fd_sc_hd__and2_1 _480_ (.A(_191_),
    .B(\dice.lfsr[6] ),
    .X(_240_));
 sky130_fd_sc_hd__clkbuf_1 _481_ (.A(_240_),
    .X(_039_));
 sky130_fd_sc_hd__or2_1 _482_ (.A(_169_),
    .B(\dice.lfsr[7] ),
    .X(_241_));
 sky130_fd_sc_hd__clkbuf_1 _483_ (.A(_241_),
    .X(_040_));
 sky130_fd_sc_hd__or2_1 _484_ (.A(_169_),
    .B(\dice.lfsr[8] ),
    .X(_242_));
 sky130_fd_sc_hd__clkbuf_1 _485_ (.A(_242_),
    .X(_041_));
 sky130_fd_sc_hd__and2_1 _486_ (.A(_191_),
    .B(\dice.lfsr[9] ),
    .X(_243_));
 sky130_fd_sc_hd__clkbuf_1 _487_ (.A(_243_),
    .X(_042_));
 sky130_fd_sc_hd__and2_1 _488_ (.A(_191_),
    .B(\dice.lfsr[10] ),
    .X(_244_));
 sky130_fd_sc_hd__clkbuf_1 _489_ (.A(_244_),
    .X(_043_));
 sky130_fd_sc_hd__a21oi_1 _490_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[11] ),
    .B1(_178_),
    .Y(_245_));
 sky130_fd_sc_hd__o21a_1 _491_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[11] ),
    .B1(_245_),
    .X(_044_));
 sky130_fd_sc_hd__and2_1 _492_ (.A(_191_),
    .B(\dice.lfsr[12] ),
    .X(_246_));
 sky130_fd_sc_hd__clkbuf_1 _493_ (.A(_246_),
    .X(_045_));
 sky130_fd_sc_hd__a21oi_1 _494_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[13] ),
    .B1(_178_),
    .Y(_247_));
 sky130_fd_sc_hd__o21a_1 _495_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[13] ),
    .B1(_247_),
    .X(_046_));
 sky130_fd_sc_hd__a21oi_1 _496_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[14] ),
    .B1(_178_),
    .Y(_248_));
 sky130_fd_sc_hd__o21a_1 _497_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[14] ),
    .B1(_248_),
    .X(_047_));
 sky130_fd_sc_hd__and2_1 _498_ (.A(_191_),
    .B(\dice.lfsr[15] ),
    .X(_249_));
 sky130_fd_sc_hd__clkbuf_1 _499_ (.A(_249_),
    .X(_048_));
 sky130_fd_sc_hd__and2_1 _500_ (.A(\dice.lfsr[0] ),
    .B(_190_),
    .X(_250_));
 sky130_fd_sc_hd__clkbuf_1 _501_ (.A(_250_),
    .X(_049_));
 sky130_fd_sc_hd__or2_1 _502_ (.A(_050_),
    .B(_176_),
    .X(_251_));
 sky130_fd_sc_hd__clkbuf_1 _503_ (.A(_251_),
    .X(_053_));
 sky130_fd_sc_hd__dfxtp_1 _504_ (.CLK(clknet_2_0__leaf_clk),
    .D(_005_),
    .Q(net4));
 sky130_fd_sc_hd__dfxtp_1 _505_ (.CLK(clknet_2_0__leaf_clk),
    .D(_000_),
    .Q(net3));
 sky130_fd_sc_hd__dfxtp_1 _506_ (.CLK(clknet_2_0__leaf_clk),
    .D(_001_),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_1 _507_ (.CLK(clknet_2_1__leaf_clk),
    .D(_002_),
    .Q(net7));
 sky130_fd_sc_hd__dfxtp_1 _508_ (.CLK(clknet_2_1__leaf_clk),
    .D(_003_),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_1 _509_ (.CLK(clknet_2_1__leaf_clk),
    .D(_004_),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_1 _510_ (.CLK(clknet_2_0__leaf_clk),
    .D(_006_),
    .Q(\dice.r_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _511_ (.CLK(clknet_2_0__leaf_clk),
    .D(_007_),
    .Q(\dice.r_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _512_ (.CLK(clknet_2_0__leaf_clk),
    .D(_008_),
    .Q(\dice.r_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _513_ (.CLK(clknet_2_1__leaf_clk),
    .D(_009_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _514_ (.CLK(clknet_2_1__leaf_clk),
    .D(_010_),
    .Q(\dice.clkdiv[0] ));
 sky130_fd_sc_hd__dfxtp_1 _515_ (.CLK(clknet_2_2__leaf_clk),
    .D(_011_),
    .Q(\dice.clkdiv[1] ));
 sky130_fd_sc_hd__dfxtp_1 _516_ (.CLK(clknet_2_2__leaf_clk),
    .D(_012_),
    .Q(\dice.clkdiv[2] ));
 sky130_fd_sc_hd__dfxtp_1 _517_ (.CLK(clknet_2_3__leaf_clk),
    .D(_013_),
    .Q(\dice.clkdiv[3] ));
 sky130_fd_sc_hd__dfxtp_1 _518_ (.CLK(clknet_2_2__leaf_clk),
    .D(_014_),
    .Q(\dice.clkdiv[4] ));
 sky130_fd_sc_hd__dfxtp_1 _519_ (.CLK(clknet_2_2__leaf_clk),
    .D(_015_),
    .Q(\dice.clkdiv[5] ));
 sky130_fd_sc_hd__dfxtp_1 _520_ (.CLK(clknet_2_3__leaf_clk),
    .D(_016_),
    .Q(\dice.clkdiv[6] ));
 sky130_fd_sc_hd__dfxtp_1 _521_ (.CLK(clknet_2_3__leaf_clk),
    .D(_017_),
    .Q(\dice.clkdiv[7] ));
 sky130_fd_sc_hd__dfxtp_1 _522_ (.CLK(clknet_2_3__leaf_clk),
    .D(_018_),
    .Q(\dice.counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _523_ (.CLK(clknet_2_3__leaf_clk),
    .D(_019_),
    .Q(\dice.counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _524_ (.CLK(clknet_2_3__leaf_clk),
    .D(_020_),
    .Q(\dice.counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _525_ (.CLK(clknet_2_3__leaf_clk),
    .D(_021_),
    .Q(\dice.counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _526_ (.CLK(clknet_2_3__leaf_clk),
    .D(_022_),
    .Q(\dice.counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _527_ (.CLK(clknet_2_3__leaf_clk),
    .D(_023_),
    .Q(\dice.counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _528_ (.CLK(clknet_2_1__leaf_clk),
    .D(_024_),
    .Q(\dice.counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _529_ (.CLK(clknet_2_1__leaf_clk),
    .D(_025_),
    .Q(\dice.counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _530_ (.CLK(clknet_2_1__leaf_clk),
    .D(_026_),
    .Q(\dice.counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _531_ (.CLK(clknet_2_1__leaf_clk),
    .D(_027_),
    .Q(\dice.counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _532_ (.CLK(clknet_2_1__leaf_clk),
    .D(_028_),
    .Q(\dice.counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _533_ (.CLK(clknet_2_1__leaf_clk),
    .D(_029_),
    .Q(\dice.counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _534_ (.CLK(clknet_2_1__leaf_clk),
    .D(_030_),
    .Q(\dice.counter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _535_ (.CLK(clknet_2_1__leaf_clk),
    .D(_031_),
    .Q(\dice.counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _536_ (.CLK(clknet_2_1__leaf_clk),
    .D(_032_),
    .Q(\dice.counter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _537_ (.CLK(clknet_2_1__leaf_clk),
    .D(_033_),
    .Q(\dice.counter[15] ));
 sky130_fd_sc_hd__dfxtp_2 _538_ (.CLK(clknet_2_2__leaf_clk),
    .D(_034_),
    .Q(\dice.lfsr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _539_ (.CLK(clknet_2_0__leaf_clk),
    .D(_035_),
    .Q(\dice.lfsr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _540_ (.CLK(clknet_2_2__leaf_clk),
    .D(_036_),
    .Q(\dice.lfsr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _541_ (.CLK(clknet_2_2__leaf_clk),
    .D(_037_),
    .Q(\dice.lfsr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _542_ (.CLK(clknet_2_2__leaf_clk),
    .D(_038_),
    .Q(\dice.lfsr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _543_ (.CLK(clknet_2_2__leaf_clk),
    .D(_039_),
    .Q(\dice.lfsr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _544_ (.CLK(clknet_2_3__leaf_clk),
    .D(_040_),
    .Q(\dice.lfsr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _545_ (.CLK(clknet_2_3__leaf_clk),
    .D(_041_),
    .Q(\dice.lfsr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _546_ (.CLK(clknet_2_3__leaf_clk),
    .D(_042_),
    .Q(\dice.lfsr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _547_ (.CLK(clknet_2_2__leaf_clk),
    .D(_043_),
    .Q(\dice.lfsr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _548_ (.CLK(clknet_2_2__leaf_clk),
    .D(_044_),
    .Q(\dice.lfsr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _549_ (.CLK(clknet_2_2__leaf_clk),
    .D(_045_),
    .Q(\dice.lfsr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _550_ (.CLK(clknet_2_2__leaf_clk),
    .D(_046_),
    .Q(\dice.lfsr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _551_ (.CLK(clknet_2_2__leaf_clk),
    .D(_047_),
    .Q(\dice.lfsr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _552_ (.CLK(clknet_2_2__leaf_clk),
    .D(_048_),
    .Q(\dice.lfsr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _553_ (.CLK(clknet_2_2__leaf_clk),
    .D(_049_),
    .Q(\dice.lfsr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _554_ (.CLK(clknet_2_0__leaf_clk),
    .D(_050_),
    .Q(\dice.bcd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _555_ (.CLK(clknet_2_0__leaf_clk),
    .D(_051_),
    .Q(\dice.bcd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _556_ (.CLK(clknet_2_0__leaf_clk),
    .D(_052_),
    .Q(\dice.bcd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _557_ (.CLK(clknet_2_0__leaf_clk),
    .D(_053_),
    .Q(net5));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(io_in),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(rst),
    .X(net2));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(io_out[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__454__B (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__417__C1 (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__357__A_N (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__356__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__322__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__311__A_N (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__307__A_N (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__300__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__279__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__277__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__484__A (.DIODE(_169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__482__A (.DIODE(_169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__478__A (.DIODE(_169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__476__A (.DIODE(_169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__472__B (.DIODE(_169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__458__B1 (.DIODE(_169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__415__B1 (.DIODE(_169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__390__B1 (.DIODE(_169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__384__A (.DIODE(_169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__370__A (.DIODE(_169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__469__A (.DIODE(_177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__444__A (.DIODE(_177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__442__A (.DIODE(_177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__439__A (.DIODE(_177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__436__A (.DIODE(_177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__433__A (.DIODE(_177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__431__A (.DIODE(_177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__398__A (.DIODE(_177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__392__B1 (.DIODE(_177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__385__B (.DIODE(_177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__496__B1 (.DIODE(_178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__494__B1 (.DIODE(_178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__490__B1 (.DIODE(_178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__467__A (.DIODE(_178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__464__C1 (.DIODE(_178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__462__A (.DIODE(_178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__448__A (.DIODE(_178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__401__A (.DIODE(_178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__394__B1 (.DIODE(_178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__387__B1 (.DIODE(_178_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(rst));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_189 ();
endmodule

