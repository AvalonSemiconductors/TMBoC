magic
tech sky130B
magscale 1 2
timestamp 1675277843
<< obsli1 >>
rect 1104 2159 83812 77809
<< obsm1 >>
rect 14 1640 84258 79280
<< metal2 >>
rect 4314 79200 4426 80000
rect 12778 79200 12890 80000
rect 21242 79200 21354 80000
rect 29706 79200 29818 80000
rect 38170 79200 38282 80000
rect 46634 79200 46746 80000
rect 55098 79200 55210 80000
rect 63562 79200 63674 80000
rect 72026 79200 72138 80000
rect 80490 79200 80602 80000
<< obsm2 >>
rect 18 79144 4258 79286
rect 4482 79144 12722 79286
rect 12946 79144 21186 79286
rect 21410 79144 29650 79286
rect 29874 79144 38114 79286
rect 38338 79144 46578 79286
rect 46802 79144 55042 79286
rect 55266 79144 63506 79286
rect 63730 79144 71970 79286
rect 72194 79144 80434 79286
rect 80658 79144 84252 79286
rect 18 1391 84252 79144
<< metal3 >>
rect 0 78420 800 78660
rect 0 75564 800 75804
rect 0 72708 800 72948
rect 0 69852 800 70092
rect 0 66996 800 67236
rect 0 64140 800 64380
rect 0 61284 800 61524
rect 0 58428 800 58668
rect 0 55572 800 55812
rect 0 52716 800 52956
rect 0 49860 800 50100
rect 0 47004 800 47244
rect 0 44148 800 44388
rect 0 41292 800 41532
rect 0 38436 800 38676
rect 0 35580 800 35820
rect 0 32724 800 32964
rect 0 29868 800 30108
rect 0 27012 800 27252
rect 0 24156 800 24396
rect 0 21300 800 21540
rect 0 18444 800 18684
rect 0 15588 800 15828
rect 0 12732 800 12972
rect 0 9876 800 10116
rect 0 7020 800 7260
rect 0 4164 800 4404
rect 0 1308 800 1548
<< obsm3 >>
rect 13 78740 83799 78981
rect 880 78340 83799 78740
rect 13 75884 83799 78340
rect 880 75484 83799 75884
rect 13 73028 83799 75484
rect 880 72628 83799 73028
rect 13 70172 83799 72628
rect 880 69772 83799 70172
rect 13 67316 83799 69772
rect 880 66916 83799 67316
rect 13 64460 83799 66916
rect 880 64060 83799 64460
rect 13 61604 83799 64060
rect 880 61204 83799 61604
rect 13 58748 83799 61204
rect 880 58348 83799 58748
rect 13 55892 83799 58348
rect 880 55492 83799 55892
rect 13 53036 83799 55492
rect 880 52636 83799 53036
rect 13 50180 83799 52636
rect 880 49780 83799 50180
rect 13 47324 83799 49780
rect 880 46924 83799 47324
rect 13 44468 83799 46924
rect 880 44068 83799 44468
rect 13 41612 83799 44068
rect 880 41212 83799 41612
rect 13 38756 83799 41212
rect 880 38356 83799 38756
rect 13 35900 83799 38356
rect 880 35500 83799 35900
rect 13 33044 83799 35500
rect 880 32644 83799 33044
rect 13 30188 83799 32644
rect 880 29788 83799 30188
rect 13 27332 83799 29788
rect 880 26932 83799 27332
rect 13 24476 83799 26932
rect 880 24076 83799 24476
rect 13 21620 83799 24076
rect 880 21220 83799 21620
rect 13 18764 83799 21220
rect 880 18364 83799 18764
rect 13 15908 83799 18364
rect 880 15508 83799 15908
rect 13 13052 83799 15508
rect 880 12652 83799 13052
rect 13 10196 83799 12652
rect 880 9796 83799 10196
rect 13 7340 83799 9796
rect 880 6940 83799 7340
rect 13 4484 83799 6940
rect 880 4084 83799 4484
rect 13 1628 83799 4084
rect 880 1395 83799 1628
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
rect 81008 2128 81328 77840
<< obsm4 >>
rect 59 77920 82741 78981
rect 59 30091 4128 77920
rect 4608 30091 19488 77920
rect 19968 30091 34848 77920
rect 35328 30091 50208 77920
rect 50688 30091 65568 77920
rect 66048 30091 80928 77920
rect 81408 30091 82741 77920
<< labels >>
rlabel metal2 s 72026 79200 72138 80000 6 clk
port 1 nsew signal input
rlabel metal2 s 4314 79200 4426 80000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 12778 79200 12890 80000 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 21242 79200 21354 80000 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 29706 79200 29818 80000 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 38170 79200 38282 80000 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 46634 79200 46746 80000 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 55098 79200 55210 80000 6 io_in[6]
port 8 nsew signal input
rlabel metal2 s 63562 79200 63674 80000 6 io_in[7]
port 9 nsew signal input
rlabel metal3 s 0 78420 800 78660 6 io_oeb
port 10 nsew signal output
rlabel metal3 s 0 1308 800 1548 6 io_out[0]
port 11 nsew signal output
rlabel metal3 s 0 29868 800 30108 6 io_out[10]
port 12 nsew signal output
rlabel metal3 s 0 32724 800 32964 6 io_out[11]
port 13 nsew signal output
rlabel metal3 s 0 35580 800 35820 6 io_out[12]
port 14 nsew signal output
rlabel metal3 s 0 38436 800 38676 6 io_out[13]
port 15 nsew signal output
rlabel metal3 s 0 41292 800 41532 6 io_out[14]
port 16 nsew signal output
rlabel metal3 s 0 44148 800 44388 6 io_out[15]
port 17 nsew signal output
rlabel metal3 s 0 47004 800 47244 6 io_out[16]
port 18 nsew signal output
rlabel metal3 s 0 49860 800 50100 6 io_out[17]
port 19 nsew signal output
rlabel metal3 s 0 52716 800 52956 6 io_out[18]
port 20 nsew signal output
rlabel metal3 s 0 55572 800 55812 6 io_out[19]
port 21 nsew signal output
rlabel metal3 s 0 4164 800 4404 6 io_out[1]
port 22 nsew signal output
rlabel metal3 s 0 58428 800 58668 6 io_out[20]
port 23 nsew signal output
rlabel metal3 s 0 61284 800 61524 6 io_out[21]
port 24 nsew signal output
rlabel metal3 s 0 64140 800 64380 6 io_out[22]
port 25 nsew signal output
rlabel metal3 s 0 66996 800 67236 6 io_out[23]
port 26 nsew signal output
rlabel metal3 s 0 69852 800 70092 6 io_out[24]
port 27 nsew signal output
rlabel metal3 s 0 72708 800 72948 6 io_out[25]
port 28 nsew signal output
rlabel metal3 s 0 75564 800 75804 6 io_out[26]
port 29 nsew signal output
rlabel metal3 s 0 7020 800 7260 6 io_out[2]
port 30 nsew signal output
rlabel metal3 s 0 9876 800 10116 6 io_out[3]
port 31 nsew signal output
rlabel metal3 s 0 12732 800 12972 6 io_out[4]
port 32 nsew signal output
rlabel metal3 s 0 15588 800 15828 6 io_out[5]
port 33 nsew signal output
rlabel metal3 s 0 18444 800 18684 6 io_out[6]
port 34 nsew signal output
rlabel metal3 s 0 21300 800 21540 6 io_out[7]
port 35 nsew signal output
rlabel metal3 s 0 24156 800 24396 6 io_out[8]
port 36 nsew signal output
rlabel metal3 s 0 27012 800 27252 6 io_out[9]
port 37 nsew signal output
rlabel metal2 s 80490 79200 80602 80000 6 rst
port 38 nsew signal input
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 77840 6 vssd1
port 40 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 85000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 18631904
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS2650/runs/23_02_01_19_43/results/signoff/wrapped_as2650.magic.gds
string GDS_START 1060172
<< end >>

