magic
tech sky130B
magscale 1 2
timestamp 1676307437
<< viali >>
rect 8585 53193 8619 53227
rect 9321 53193 9355 53227
rect 21097 53193 21131 53227
rect 26617 53193 26651 53227
rect 29193 53193 29227 53227
rect 31769 53193 31803 53227
rect 47133 53193 47167 53227
rect 49709 53193 49743 53227
rect 3157 53125 3191 53159
rect 4905 53125 4939 53159
rect 5457 53125 5491 53159
rect 6653 53125 6687 53159
rect 51825 53125 51859 53159
rect 2329 53057 2363 53091
rect 4169 53057 4203 53091
rect 7757 53057 7791 53091
rect 9137 53057 9171 53091
rect 10149 53057 10183 53091
rect 12081 53057 12115 53091
rect 12541 53057 12575 53091
rect 14841 53057 14875 53091
rect 16313 53057 16347 53091
rect 16865 53057 16899 53091
rect 18889 53057 18923 53091
rect 19717 53057 19751 53091
rect 20453 53057 20487 53091
rect 20913 53057 20947 53091
rect 22109 53057 22143 53091
rect 22845 53057 22879 53091
rect 23305 53057 23339 53091
rect 24041 53057 24075 53091
rect 24593 53057 24627 53091
rect 25697 53057 25731 53091
rect 27169 53057 27203 53091
rect 28273 53057 28307 53091
rect 29929 53057 29963 53091
rect 30665 53057 30699 53091
rect 31125 53057 31159 53091
rect 32505 53057 32539 53091
rect 33149 53057 33183 53091
rect 34253 53057 34287 53091
rect 35449 53057 35483 53091
rect 35909 53057 35943 53091
rect 36645 53057 36679 53091
rect 37841 53057 37875 53091
rect 38301 53057 38335 53091
rect 39037 53057 39071 53091
rect 40233 53057 40267 53091
rect 40693 53057 40727 53091
rect 41429 53057 41463 53091
rect 41889 53057 41923 53091
rect 42809 53057 42843 53091
rect 43637 53057 43671 53091
rect 45201 53057 45235 53091
rect 47777 53057 47811 53091
rect 50353 53057 50387 53091
rect 53205 53057 53239 53091
rect 2605 52989 2639 53023
rect 10425 52989 10459 53023
rect 12817 52989 12851 53023
rect 16037 52989 16071 53023
rect 18613 52989 18647 53023
rect 43913 52989 43947 53023
rect 45477 52989 45511 53023
rect 48053 52989 48087 53023
rect 50629 52989 50663 53023
rect 53481 52989 53515 53023
rect 4353 52921 4387 52955
rect 19901 52921 19935 52955
rect 24777 52921 24811 52955
rect 32965 52921 32999 52955
rect 37657 52921 37691 52955
rect 51641 52921 51675 52955
rect 3249 52853 3283 52887
rect 5549 52853 5583 52887
rect 6745 52853 6779 52887
rect 7941 52853 7975 52887
rect 15025 52853 15059 52887
rect 22293 52853 22327 52887
rect 23489 52853 23523 52887
rect 25881 52853 25915 52887
rect 27353 52853 27387 52887
rect 28089 52853 28123 52887
rect 29745 52853 29779 52887
rect 30481 52853 30515 52887
rect 32321 52853 32355 52887
rect 34069 52853 34103 52887
rect 35265 52853 35299 52887
rect 36461 52853 36495 52887
rect 38853 52853 38887 52887
rect 40049 52853 40083 52887
rect 41245 52853 41279 52887
rect 42625 52853 42659 52887
rect 3157 52649 3191 52683
rect 4077 52649 4111 52683
rect 6469 52649 6503 52683
rect 7665 52649 7699 52683
rect 10057 52649 10091 52683
rect 13645 52649 13679 52683
rect 15117 52649 15151 52683
rect 18797 52649 18831 52683
rect 19533 52649 19567 52683
rect 22017 52649 22051 52683
rect 26341 52649 26375 52683
rect 27997 52649 28031 52683
rect 32781 52649 32815 52683
rect 33977 52649 34011 52683
rect 36369 52649 36403 52683
rect 38761 52649 38795 52683
rect 42441 52649 42475 52683
rect 43545 52649 43579 52683
rect 45201 52649 45235 52683
rect 51549 52649 51583 52683
rect 53113 52649 53147 52683
rect 10885 52513 10919 52547
rect 11345 52513 11379 52547
rect 16865 52513 16899 52547
rect 17325 52513 17359 52547
rect 46029 52513 46063 52547
rect 47961 52513 47995 52547
rect 48421 52513 48455 52547
rect 48697 52513 48731 52547
rect 52009 52513 52043 52547
rect 1869 52445 1903 52479
rect 2605 52445 2639 52479
rect 11621 52445 11655 52479
rect 14473 52445 14507 52479
rect 17601 52445 17635 52479
rect 27169 52445 27203 52479
rect 46305 52445 46339 52479
rect 52193 52445 52227 52479
rect 54033 52445 54067 52479
rect 1685 52377 1719 52411
rect 2421 52377 2455 52411
rect 54217 52377 54251 52411
rect 14289 52309 14323 52343
rect 25789 52309 25823 52343
rect 2421 52105 2455 52139
rect 24593 52105 24627 52139
rect 45937 52105 45971 52139
rect 51457 52105 51491 52139
rect 54309 52105 54343 52139
rect 3433 52037 3467 52071
rect 25421 52037 25455 52071
rect 27721 52037 27755 52071
rect 27813 52037 27847 52071
rect 1685 51969 1719 52003
rect 2881 51969 2915 52003
rect 25145 51969 25179 52003
rect 25329 51969 25363 52003
rect 25513 51969 25547 52003
rect 26617 51969 26651 52003
rect 27537 51969 27571 52003
rect 27905 51969 27939 52003
rect 1869 51833 1903 51867
rect 25697 51765 25731 51799
rect 28089 51765 28123 51799
rect 2881 51561 2915 51595
rect 27353 51561 27387 51595
rect 1685 51289 1719 51323
rect 2329 51289 2363 51323
rect 53757 51289 53791 51323
rect 1777 51221 1811 51255
rect 26065 51221 26099 51255
rect 54309 51221 54343 51255
rect 54309 50881 54343 50915
rect 2145 50813 2179 50847
rect 2421 50813 2455 50847
rect 2881 50813 2915 50847
rect 53573 50677 53607 50711
rect 54125 50677 54159 50711
rect 54125 50405 54159 50439
rect 2145 50269 2179 50303
rect 2421 50269 2455 50303
rect 2881 50269 2915 50303
rect 54309 50269 54343 50303
rect 52653 50201 52687 50235
rect 53113 50133 53147 50167
rect 54125 49929 54159 49963
rect 1685 49793 1719 49827
rect 2329 49793 2363 49827
rect 52377 49793 52411 49827
rect 53665 49793 53699 49827
rect 54309 49793 54343 49827
rect 1869 49725 1903 49759
rect 53481 49657 53515 49691
rect 52929 49589 52963 49623
rect 53757 49249 53791 49283
rect 2145 49181 2179 49215
rect 2421 49181 2455 49215
rect 2881 49181 2915 49215
rect 52285 49181 52319 49215
rect 53021 49181 53055 49215
rect 53481 49181 53515 49215
rect 51825 49113 51859 49147
rect 32781 49045 32815 49079
rect 33333 49045 33367 49079
rect 52837 49045 52871 49079
rect 52929 48841 52963 48875
rect 51181 48773 51215 48807
rect 52377 48705 52411 48739
rect 53757 48705 53791 48739
rect 2145 48637 2179 48671
rect 2421 48637 2455 48671
rect 2881 48637 2915 48671
rect 53481 48637 53515 48671
rect 52193 48569 52227 48603
rect 32781 48501 32815 48535
rect 33241 48501 33275 48535
rect 33885 48501 33919 48535
rect 34437 48501 34471 48535
rect 51641 48501 51675 48535
rect 32321 48229 32355 48263
rect 34161 48161 34195 48195
rect 2145 48093 2179 48127
rect 2421 48093 2455 48127
rect 2881 48093 2915 48127
rect 33057 48093 33091 48127
rect 33150 48093 33184 48127
rect 33425 48093 33459 48127
rect 33563 48093 33597 48127
rect 35541 48093 35575 48127
rect 52193 48093 52227 48127
rect 52653 48093 52687 48127
rect 53297 48093 53331 48127
rect 53481 48093 53515 48127
rect 53665 48093 53699 48127
rect 33333 48025 33367 48059
rect 53573 48025 53607 48059
rect 31861 47957 31895 47991
rect 33701 47957 33735 47991
rect 34897 47957 34931 47991
rect 50997 47957 51031 47991
rect 51549 47957 51583 47991
rect 52009 47957 52043 47991
rect 52837 47957 52871 47991
rect 53849 47957 53883 47991
rect 29653 47753 29687 47787
rect 33425 47685 33459 47719
rect 34437 47685 34471 47719
rect 50169 47685 50203 47719
rect 52193 47685 52227 47719
rect 52929 47685 52963 47719
rect 2145 47617 2179 47651
rect 33057 47617 33091 47651
rect 33150 47617 33184 47651
rect 33333 47617 33367 47651
rect 33563 47617 33597 47651
rect 34345 47617 34379 47651
rect 34529 47617 34563 47651
rect 34713 47617 34747 47651
rect 50721 47617 50755 47651
rect 51181 47617 51215 47651
rect 51985 47617 52019 47651
rect 52109 47617 52143 47651
rect 52377 47617 52411 47651
rect 2421 47549 2455 47583
rect 2881 47549 2915 47583
rect 53481 47549 53515 47583
rect 53757 47549 53791 47583
rect 32321 47481 32355 47515
rect 34161 47481 34195 47515
rect 36369 47481 36403 47515
rect 51365 47481 51399 47515
rect 51825 47481 51859 47515
rect 30665 47413 30699 47447
rect 31677 47413 31711 47447
rect 33701 47413 33735 47447
rect 35173 47413 35207 47447
rect 35817 47413 35851 47447
rect 29101 47209 29135 47243
rect 52469 47209 52503 47243
rect 31493 47141 31527 47175
rect 33793 47141 33827 47175
rect 51457 47141 51491 47175
rect 2145 47073 2179 47107
rect 34989 47073 35023 47107
rect 2421 47005 2455 47039
rect 2881 47005 2915 47039
rect 29837 47005 29871 47039
rect 30113 47005 30147 47039
rect 30205 47005 30239 47039
rect 30849 47005 30883 47039
rect 30942 47005 30976 47039
rect 31217 47005 31251 47039
rect 31355 47005 31389 47039
rect 31953 47005 31987 47039
rect 32046 47005 32080 47039
rect 32321 47005 32355 47039
rect 32459 47005 32493 47039
rect 33149 47005 33183 47039
rect 33297 47005 33331 47039
rect 33655 47005 33689 47039
rect 34345 47005 34379 47039
rect 50905 47005 50939 47039
rect 51617 47005 51651 47039
rect 52009 47005 52043 47039
rect 52653 47005 52687 47039
rect 52837 47005 52871 47039
rect 53021 47005 53055 47039
rect 53481 47005 53515 47039
rect 53757 47005 53791 47039
rect 30021 46937 30055 46971
rect 31125 46937 31159 46971
rect 32229 46937 32263 46971
rect 33425 46937 33459 46971
rect 33517 46937 33551 46971
rect 49801 46937 49835 46971
rect 51733 46937 51767 46971
rect 51825 46937 51859 46971
rect 52745 46937 52779 46971
rect 30389 46869 30423 46903
rect 32597 46869 32631 46903
rect 35449 46869 35483 46903
rect 50445 46869 50479 46903
rect 30481 46665 30515 46699
rect 29469 46597 29503 46631
rect 34069 46597 34103 46631
rect 2145 46529 2179 46563
rect 32505 46529 32539 46563
rect 32597 46529 32631 46563
rect 32689 46529 32723 46563
rect 32873 46529 32907 46563
rect 33977 46529 34011 46563
rect 34161 46529 34195 46563
rect 34345 46529 34379 46563
rect 50537 46529 50571 46563
rect 53757 46529 53791 46563
rect 2421 46461 2455 46495
rect 2881 46461 2915 46495
rect 52101 46461 52135 46495
rect 52377 46461 52411 46495
rect 53481 46461 53515 46495
rect 31677 46393 31711 46427
rect 34805 46393 34839 46427
rect 31217 46325 31251 46359
rect 32321 46325 32355 46359
rect 33793 46325 33827 46359
rect 35449 46325 35483 46359
rect 51089 46325 51123 46359
rect 53021 46325 53055 46359
rect 32965 46121 32999 46155
rect 34989 46121 35023 46155
rect 31401 46053 31435 46087
rect 34069 46053 34103 46087
rect 31861 45985 31895 46019
rect 53757 45985 53791 46019
rect 2145 45917 2179 45951
rect 2421 45917 2455 45951
rect 2881 45917 2915 45951
rect 32413 45917 32447 45951
rect 32597 45917 32631 45951
rect 32781 45917 32815 45951
rect 51733 45917 51767 45951
rect 52193 45917 52227 45951
rect 52469 45917 52503 45951
rect 53481 45917 53515 45951
rect 32689 45849 32723 45883
rect 51181 45849 51215 45883
rect 33517 45781 33551 45815
rect 33425 45509 33459 45543
rect 51089 45441 51123 45475
rect 53757 45441 53791 45475
rect 2145 45373 2179 45407
rect 2421 45373 2455 45407
rect 2881 45373 2915 45407
rect 52101 45373 52135 45407
rect 52377 45373 52411 45407
rect 53481 45373 53515 45407
rect 32321 45237 32355 45271
rect 32873 45237 32907 45271
rect 53021 45237 53055 45271
rect 27445 45033 27479 45067
rect 28089 45033 28123 45067
rect 52469 44897 52503 44931
rect 2145 44829 2179 44863
rect 2421 44829 2455 44863
rect 2881 44829 2915 44863
rect 51733 44829 51767 44863
rect 52193 44829 52227 44863
rect 53481 44829 53515 44863
rect 53757 44829 53791 44863
rect 51181 44761 51215 44795
rect 26893 44693 26927 44727
rect 28641 44489 28675 44523
rect 51089 44489 51123 44523
rect 26249 44421 26283 44455
rect 26341 44421 26375 44455
rect 25513 44353 25547 44387
rect 26157 44353 26191 44387
rect 26525 44353 26559 44387
rect 53757 44353 53791 44387
rect 2145 44285 2179 44319
rect 2421 44285 2455 44319
rect 2881 44285 2915 44319
rect 27169 44285 27203 44319
rect 52101 44285 52135 44319
rect 52377 44285 52411 44319
rect 53481 44285 53515 44319
rect 25973 44217 26007 44251
rect 32321 44217 32355 44251
rect 27997 44149 28031 44183
rect 30481 44149 30515 44183
rect 31033 44149 31067 44183
rect 32873 44149 32907 44183
rect 53021 44149 53055 44183
rect 34161 43945 34195 43979
rect 29745 43877 29779 43911
rect 25973 43809 26007 43843
rect 2145 43741 2179 43775
rect 2421 43741 2455 43775
rect 2881 43741 2915 43775
rect 27215 43741 27249 43775
rect 27353 43741 27387 43775
rect 27445 43741 27479 43775
rect 27628 43741 27662 43775
rect 27721 43741 27755 43775
rect 28549 43741 28583 43775
rect 51733 43741 51767 43775
rect 53481 43741 53515 43775
rect 53757 43741 53791 43775
rect 31493 43673 31527 43707
rect 52285 43673 52319 43707
rect 52929 43673 52963 43707
rect 26525 43605 26559 43639
rect 27077 43605 27111 43639
rect 29009 43605 29043 43639
rect 30389 43605 30423 43639
rect 30849 43605 30883 43639
rect 31953 43605 31987 43639
rect 32597 43605 32631 43639
rect 33149 43605 33183 43639
rect 33701 43605 33735 43639
rect 52837 43605 52871 43639
rect 34621 43401 34655 43435
rect 25421 43333 25455 43367
rect 26065 43333 26099 43367
rect 26617 43333 26651 43367
rect 28273 43333 28307 43367
rect 2145 43265 2179 43299
rect 32873 43265 32907 43299
rect 2421 43197 2455 43231
rect 2881 43197 2915 43231
rect 29653 43197 29687 43231
rect 32413 43197 32447 43231
rect 52377 43197 52411 43231
rect 53481 43197 53515 43231
rect 53757 43197 53791 43231
rect 33517 43129 33551 43163
rect 27629 43061 27663 43095
rect 29101 43061 29135 43095
rect 30205 43061 30239 43095
rect 30757 43061 30791 43095
rect 31401 43061 31435 43095
rect 34069 43061 34103 43095
rect 35173 43061 35207 43095
rect 53021 43061 53055 43095
rect 25605 42857 25639 42891
rect 27169 42789 27203 42823
rect 27813 42789 27847 42823
rect 26157 42721 26191 42755
rect 28365 42721 28399 42755
rect 53757 42721 53791 42755
rect 2145 42653 2179 42687
rect 2421 42653 2455 42687
rect 2881 42653 2915 42687
rect 29193 42653 29227 42687
rect 29929 42653 29963 42687
rect 30021 42653 30055 42687
rect 30297 42653 30331 42687
rect 32505 42653 32539 42687
rect 32598 42653 32632 42687
rect 32873 42653 32907 42687
rect 32970 42653 33004 42687
rect 33977 42653 34011 42687
rect 53021 42653 53055 42687
rect 53481 42653 53515 42687
rect 25053 42585 25087 42619
rect 26709 42585 26743 42619
rect 30113 42585 30147 42619
rect 31309 42585 31343 42619
rect 31861 42585 31895 42619
rect 32781 42585 32815 42619
rect 33609 42585 33643 42619
rect 33793 42585 33827 42619
rect 51825 42585 51859 42619
rect 29745 42517 29779 42551
rect 30849 42517 30883 42551
rect 33149 42517 33183 42551
rect 34897 42517 34931 42551
rect 35541 42517 35575 42551
rect 52377 42517 52411 42551
rect 52837 42517 52871 42551
rect 29377 42313 29411 42347
rect 33149 42313 33183 42347
rect 35725 42313 35759 42347
rect 36369 42313 36403 42347
rect 26157 42245 26191 42279
rect 26249 42245 26283 42279
rect 30389 42245 30423 42279
rect 30481 42245 30515 42279
rect 32873 42245 32907 42279
rect 33885 42245 33919 42279
rect 24869 42177 24903 42211
rect 24961 42177 24995 42211
rect 25145 42177 25179 42211
rect 25237 42177 25271 42211
rect 25421 42177 25455 42211
rect 25881 42177 25915 42211
rect 25974 42177 26008 42211
rect 26387 42177 26421 42211
rect 28457 42177 28491 42211
rect 28549 42177 28583 42211
rect 28733 42177 28767 42211
rect 28825 42177 28859 42211
rect 30292 42177 30326 42211
rect 30664 42177 30698 42211
rect 30757 42177 30791 42211
rect 32505 42177 32539 42211
rect 32598 42177 32632 42211
rect 32781 42177 32815 42211
rect 32970 42177 33004 42211
rect 33793 42177 33827 42211
rect 33977 42177 34011 42211
rect 34161 42177 34195 42211
rect 53757 42177 53791 42211
rect 2145 42109 2179 42143
rect 2421 42109 2455 42143
rect 2881 42109 2915 42143
rect 31309 42109 31343 42143
rect 53481 42109 53515 42143
rect 33609 42041 33643 42075
rect 34713 42041 34747 42075
rect 51825 42041 51859 42075
rect 23857 41973 23891 42007
rect 24409 41973 24443 42007
rect 26525 41973 26559 42007
rect 27629 41973 27663 42007
rect 28273 41973 28307 42007
rect 30113 41973 30147 42007
rect 35265 41973 35299 42007
rect 52285 41973 52319 42007
rect 53021 41973 53055 42007
rect 28365 41769 28399 41803
rect 28825 41769 28859 41803
rect 30849 41769 30883 41803
rect 33517 41769 33551 41803
rect 54125 41769 54159 41803
rect 25973 41701 26007 41735
rect 52837 41701 52871 41735
rect 53481 41701 53515 41735
rect 2145 41633 2179 41667
rect 26433 41633 26467 41667
rect 2421 41565 2455 41599
rect 2881 41565 2915 41599
rect 27261 41565 27295 41599
rect 27721 41565 27755 41599
rect 27814 41565 27848 41599
rect 28089 41565 28123 41599
rect 28227 41565 28261 41599
rect 29885 41565 29919 41599
rect 30021 41565 30055 41599
rect 30296 41565 30330 41599
rect 30382 41565 30416 41599
rect 30987 41565 31021 41599
rect 31125 41565 31159 41599
rect 31400 41565 31434 41599
rect 31493 41565 31527 41599
rect 32592 41565 32626 41599
rect 32689 41565 32723 41599
rect 32964 41565 32998 41599
rect 33057 41565 33091 41599
rect 33701 41565 33735 41599
rect 33793 41565 33827 41599
rect 34069 41565 34103 41599
rect 34897 41565 34931 41599
rect 36369 41565 36403 41599
rect 51733 41565 51767 41599
rect 52377 41565 52411 41599
rect 53021 41565 53055 41599
rect 53665 41565 53699 41599
rect 54309 41565 54343 41599
rect 23489 41497 23523 41531
rect 24685 41497 24719 41531
rect 27997 41497 28031 41531
rect 30113 41497 30147 41531
rect 31217 41497 31251 41531
rect 32781 41497 32815 41531
rect 33885 41497 33919 41531
rect 35081 41497 35115 41531
rect 24041 41429 24075 41463
rect 24961 41429 24995 41463
rect 27077 41429 27111 41463
rect 29745 41429 29779 41463
rect 32413 41429 32447 41463
rect 35265 41429 35299 41463
rect 35725 41429 35759 41463
rect 36829 41429 36863 41463
rect 52193 41429 52227 41463
rect 24501 41225 24535 41259
rect 26341 41225 26375 41259
rect 28273 41225 28307 41259
rect 30941 41225 30975 41259
rect 31585 41225 31619 41259
rect 26249 41157 26283 41191
rect 27445 41157 27479 41191
rect 27537 41157 27571 41191
rect 28549 41157 28583 41191
rect 29653 41157 29687 41191
rect 33057 41157 33091 41191
rect 33149 41157 33183 41191
rect 33885 41157 33919 41191
rect 2145 41089 2179 41123
rect 24041 41089 24075 41123
rect 27353 41089 27387 41123
rect 27721 41089 27755 41123
rect 28457 41089 28491 41123
rect 28641 41089 28675 41123
rect 28825 41089 28859 41123
rect 29285 41089 29319 41123
rect 29433 41089 29467 41123
rect 29561 41089 29595 41123
rect 29791 41089 29825 41123
rect 32960 41089 32994 41123
rect 33332 41089 33366 41123
rect 33425 41089 33459 41123
rect 34069 41089 34103 41123
rect 35265 41089 35299 41123
rect 53757 41089 53791 41123
rect 2421 41021 2455 41055
rect 2881 41021 2915 41055
rect 25145 41021 25179 41055
rect 34713 41021 34747 41055
rect 35817 41021 35851 41055
rect 51825 41021 51859 41055
rect 53481 41021 53515 41055
rect 52377 40953 52411 40987
rect 25697 40885 25731 40919
rect 27169 40885 27203 40919
rect 29929 40885 29963 40919
rect 30389 40885 30423 40919
rect 32781 40885 32815 40919
rect 34253 40885 34287 40919
rect 52929 40885 52963 40919
rect 23397 40681 23431 40715
rect 24961 40681 24995 40715
rect 52193 40681 52227 40715
rect 53021 40681 53055 40715
rect 54125 40681 54159 40715
rect 27905 40613 27939 40647
rect 29009 40613 29043 40647
rect 30389 40613 30423 40647
rect 30849 40545 30883 40579
rect 2145 40477 2179 40511
rect 2421 40477 2455 40511
rect 2881 40477 2915 40511
rect 26157 40477 26191 40511
rect 26281 40477 26315 40511
rect 26433 40477 26467 40511
rect 26525 40477 26559 40511
rect 27261 40477 27295 40511
rect 27354 40477 27388 40511
rect 27629 40477 27663 40511
rect 27767 40477 27801 40511
rect 28365 40477 28399 40511
rect 28513 40477 28547 40511
rect 28641 40477 28675 40511
rect 28871 40477 28905 40511
rect 31769 40477 31803 40511
rect 32592 40477 32626 40511
rect 32781 40477 32815 40511
rect 32964 40477 32998 40511
rect 33057 40477 33091 40511
rect 33517 40477 33551 40511
rect 35081 40477 35115 40511
rect 51733 40477 51767 40511
rect 52377 40477 52411 40511
rect 52837 40477 52871 40511
rect 53665 40477 53699 40511
rect 54309 40477 54343 40511
rect 27537 40409 27571 40443
rect 28733 40409 28767 40443
rect 32689 40409 32723 40443
rect 33701 40409 33735 40443
rect 34897 40409 34931 40443
rect 36277 40409 36311 40443
rect 23949 40341 23983 40375
rect 25513 40341 25547 40375
rect 25973 40341 26007 40375
rect 29745 40341 29779 40375
rect 31861 40341 31895 40375
rect 32413 40341 32447 40375
rect 33885 40341 33919 40375
rect 35633 40341 35667 40375
rect 53481 40341 53515 40375
rect 24409 40137 24443 40171
rect 25053 40137 25087 40171
rect 35817 40137 35851 40171
rect 27537 40069 27571 40103
rect 30205 40069 30239 40103
rect 31309 40069 31343 40103
rect 32597 40069 32631 40103
rect 33425 40069 33459 40103
rect 33609 40069 33643 40103
rect 34253 40069 34287 40103
rect 2145 40001 2179 40035
rect 23857 40001 23891 40035
rect 25605 40001 25639 40035
rect 26433 40001 26467 40035
rect 26617 40001 26651 40035
rect 27169 40001 27203 40035
rect 27317 40001 27351 40035
rect 27445 40001 27479 40035
rect 27675 40001 27709 40035
rect 28733 40001 28767 40035
rect 28825 40001 28859 40035
rect 29009 40001 29043 40035
rect 29101 40001 29135 40035
rect 29837 40001 29871 40035
rect 29985 40001 30019 40035
rect 30113 40001 30147 40035
rect 30343 40001 30377 40035
rect 31493 40001 31527 40035
rect 32500 40001 32534 40035
rect 32689 40001 32723 40035
rect 32827 40001 32861 40035
rect 32976 40001 33010 40035
rect 34437 40001 34471 40035
rect 34621 40001 34655 40035
rect 35173 40001 35207 40035
rect 53757 40001 53791 40035
rect 2421 39933 2455 39967
rect 2881 39933 2915 39967
rect 51825 39933 51859 39967
rect 53481 39933 53515 39967
rect 23305 39865 23339 39899
rect 35357 39865 35391 39899
rect 52377 39865 52411 39899
rect 22845 39797 22879 39831
rect 25697 39797 25731 39831
rect 26249 39797 26283 39831
rect 27813 39797 27847 39831
rect 28549 39797 28583 39831
rect 30481 39797 30515 39831
rect 31677 39797 31711 39831
rect 32321 39797 32355 39831
rect 33793 39797 33827 39831
rect 53021 39797 53055 39831
rect 22293 39593 22327 39627
rect 25697 39593 25731 39627
rect 52837 39593 52871 39627
rect 2145 39457 2179 39491
rect 22937 39457 22971 39491
rect 34161 39457 34195 39491
rect 2421 39389 2455 39423
rect 2881 39389 2915 39423
rect 25053 39389 25087 39423
rect 25146 39389 25180 39423
rect 25421 39389 25455 39423
rect 25518 39389 25552 39423
rect 26157 39389 26191 39423
rect 26250 39389 26284 39423
rect 26525 39389 26559 39423
rect 26622 39389 26656 39423
rect 27537 39389 27571 39423
rect 27721 39389 27755 39423
rect 27905 39389 27939 39423
rect 28365 39389 28399 39423
rect 28549 39389 28583 39423
rect 30665 39389 30699 39423
rect 31585 39389 31619 39423
rect 32505 39389 32539 39423
rect 33701 39389 33735 39423
rect 34989 39389 35023 39423
rect 52377 39389 52411 39423
rect 53021 39389 53055 39423
rect 53481 39389 53515 39423
rect 53757 39389 53791 39423
rect 25329 39321 25363 39355
rect 26433 39321 26467 39355
rect 27629 39321 27663 39355
rect 31401 39321 31435 39355
rect 32689 39321 32723 39355
rect 33517 39321 33551 39355
rect 35173 39321 35207 39355
rect 51825 39321 51859 39355
rect 23489 39253 23523 39287
rect 23949 39253 23983 39287
rect 26801 39253 26835 39287
rect 27353 39253 27387 39287
rect 28733 39253 28767 39287
rect 29745 39253 29779 39287
rect 30573 39253 30607 39287
rect 31217 39253 31251 39287
rect 32873 39253 32907 39287
rect 33333 39253 33367 39287
rect 35633 39253 35667 39287
rect 16221 39049 16255 39083
rect 17417 39049 17451 39083
rect 22937 39049 22971 39083
rect 23581 39049 23615 39083
rect 25145 39049 25179 39083
rect 27169 39049 27203 39083
rect 27813 39049 27847 39083
rect 30481 39049 30515 39083
rect 17141 38981 17175 39015
rect 24593 38981 24627 39015
rect 29101 38981 29135 39015
rect 29193 38981 29227 39015
rect 31677 38981 31711 39015
rect 32873 38981 32907 39015
rect 33057 38981 33091 39015
rect 33885 38981 33919 39015
rect 2145 38913 2179 38947
rect 16865 38913 16899 38947
rect 17049 38913 17083 38947
rect 17233 38913 17267 38947
rect 26433 38913 26467 38947
rect 26617 38913 26651 38947
rect 27537 38913 27571 38947
rect 27905 38913 27939 38947
rect 28825 38913 28859 38947
rect 28918 38913 28952 38947
rect 29290 38913 29324 38947
rect 33241 38913 33275 38947
rect 34529 38913 34563 38947
rect 52101 38913 52135 38947
rect 53757 38913 53791 38947
rect 2421 38845 2455 38879
rect 2881 38845 2915 38879
rect 17969 38845 18003 38879
rect 52377 38845 52411 38879
rect 53481 38845 53515 38879
rect 34713 38777 34747 38811
rect 24133 38709 24167 38743
rect 25789 38709 25823 38743
rect 26249 38709 26283 38743
rect 26617 38709 26651 38743
rect 27445 38709 27479 38743
rect 27629 38709 27663 38743
rect 29469 38709 29503 38743
rect 29929 38709 29963 38743
rect 31585 38709 31619 38743
rect 32321 38709 32355 38743
rect 33793 38709 33827 38743
rect 53021 38709 53055 38743
rect 24869 38505 24903 38539
rect 26985 38505 27019 38539
rect 27537 38505 27571 38539
rect 31585 38505 31619 38539
rect 29193 38437 29227 38471
rect 25881 38369 25915 38403
rect 27629 38369 27663 38403
rect 52469 38369 52503 38403
rect 53757 38369 53791 38403
rect 23489 38301 23523 38335
rect 26433 38301 26467 38335
rect 26617 38301 26651 38335
rect 26801 38301 26835 38335
rect 27721 38301 27755 38335
rect 28457 38301 28491 38335
rect 28641 38301 28675 38335
rect 29837 38301 29871 38335
rect 30849 38301 30883 38335
rect 31407 38301 31441 38335
rect 32781 38301 32815 38335
rect 33517 38301 33551 38335
rect 51733 38301 51767 38335
rect 52193 38301 52227 38335
rect 53481 38301 53515 38335
rect 1685 38233 1719 38267
rect 2329 38233 2363 38267
rect 22845 38233 22879 38267
rect 26709 38233 26743 38267
rect 27445 38233 27479 38267
rect 30021 38233 30055 38267
rect 34069 38233 34103 38267
rect 51181 38233 51215 38267
rect 1777 38165 1811 38199
rect 17509 38165 17543 38199
rect 24041 38165 24075 38199
rect 25421 38165 25455 38199
rect 27905 38165 27939 38199
rect 30205 38165 30239 38199
rect 30757 38165 30791 38199
rect 32689 38165 32723 38199
rect 33425 38165 33459 38199
rect 24133 37961 24167 37995
rect 26617 37961 26651 37995
rect 27905 37961 27939 37995
rect 29009 37961 29043 37995
rect 30113 37961 30147 37995
rect 32689 37961 32723 37995
rect 34345 37961 34379 37995
rect 27537 37893 27571 37927
rect 29285 37893 29319 37927
rect 29377 37893 29411 37927
rect 30389 37893 30423 37927
rect 30481 37893 30515 37927
rect 33793 37893 33827 37927
rect 51089 37893 51123 37927
rect 1593 37825 1627 37859
rect 2789 37825 2823 37859
rect 24777 37825 24811 37859
rect 25421 37825 25455 37859
rect 25605 37825 25639 37859
rect 26065 37825 26099 37859
rect 26249 37825 26283 37859
rect 26341 37825 26375 37859
rect 26433 37825 26467 37859
rect 27353 37825 27387 37859
rect 27629 37825 27663 37859
rect 27767 37825 27801 37859
rect 29147 37825 29181 37859
rect 29560 37825 29594 37859
rect 29653 37825 29687 37859
rect 30251 37825 30285 37859
rect 30609 37825 30643 37859
rect 30757 37825 30791 37859
rect 31217 37825 31251 37859
rect 32413 37825 32447 37859
rect 33241 37825 33275 37859
rect 53757 37825 53791 37859
rect 52101 37757 52135 37791
rect 52377 37757 52411 37791
rect 53481 37757 53515 37791
rect 1777 37689 1811 37723
rect 23121 37689 23155 37723
rect 23673 37689 23707 37723
rect 2329 37621 2363 37655
rect 22569 37621 22603 37655
rect 25237 37621 25271 37655
rect 25605 37621 25639 37655
rect 28365 37621 28399 37655
rect 34897 37621 34931 37655
rect 53021 37621 53055 37655
rect 24041 37417 24075 37451
rect 24685 37417 24719 37451
rect 27629 37417 27663 37451
rect 28733 37417 28767 37451
rect 31585 37417 31619 37451
rect 32137 37417 32171 37451
rect 25237 37349 25271 37383
rect 2421 37281 2455 37315
rect 22385 37281 22419 37315
rect 28825 37281 28859 37315
rect 31125 37281 31159 37315
rect 33793 37281 33827 37315
rect 51733 37281 51767 37315
rect 53481 37281 53515 37315
rect 2145 37213 2179 37247
rect 25881 37213 25915 37247
rect 26663 37213 26697 37247
rect 26893 37213 26927 37247
rect 27076 37213 27110 37247
rect 27169 37213 27203 37247
rect 27767 37213 27801 37247
rect 27997 37213 28031 37247
rect 28180 37213 28214 37247
rect 28273 37213 28307 37247
rect 28733 37213 28767 37247
rect 29924 37213 29958 37247
rect 30296 37213 30330 37247
rect 30389 37213 30423 37247
rect 30941 37213 30975 37247
rect 52745 37213 52779 37247
rect 53021 37213 53055 37247
rect 53757 37213 53791 37247
rect 26065 37145 26099 37179
rect 26801 37145 26835 37179
rect 27908 37145 27942 37179
rect 30021 37145 30055 37179
rect 30113 37145 30147 37179
rect 32965 37145 32999 37179
rect 22937 37077 22971 37111
rect 23489 37077 23523 37111
rect 26525 37077 26559 37111
rect 29101 37077 29135 37111
rect 29745 37077 29779 37111
rect 33057 37077 33091 37111
rect 26433 36873 26467 36907
rect 27721 36873 27755 36907
rect 28733 36873 28767 36907
rect 32321 36873 32355 36907
rect 32965 36873 32999 36907
rect 53021 36873 53055 36907
rect 22109 36805 22143 36839
rect 26157 36805 26191 36839
rect 27445 36805 27479 36839
rect 29377 36805 29411 36839
rect 2145 36737 2179 36771
rect 25421 36737 25455 36771
rect 25881 36737 25915 36771
rect 26065 36737 26099 36771
rect 26249 36737 26283 36771
rect 27169 36737 27203 36771
rect 27353 36737 27387 36771
rect 27537 36737 27571 36771
rect 28171 36759 28205 36793
rect 28273 36737 28307 36771
rect 28457 36737 28491 36771
rect 28549 36737 28583 36771
rect 30297 36737 30331 36771
rect 31769 36737 31803 36771
rect 2421 36669 2455 36703
rect 2881 36669 2915 36703
rect 24317 36669 24351 36703
rect 52377 36669 52411 36703
rect 53481 36669 53515 36703
rect 53757 36669 53791 36703
rect 22569 36601 22603 36635
rect 24869 36601 24903 36635
rect 30481 36601 30515 36635
rect 31217 36601 31251 36635
rect 23121 36533 23155 36567
rect 23765 36533 23799 36567
rect 29285 36533 29319 36567
rect 33425 36533 33459 36567
rect 23489 36329 23523 36363
rect 26341 36329 26375 36363
rect 31953 36329 31987 36363
rect 22293 36261 22327 36295
rect 24777 36261 24811 36295
rect 29745 36261 29779 36295
rect 31493 36261 31527 36295
rect 51825 36261 51859 36295
rect 2145 36193 2179 36227
rect 21833 36193 21867 36227
rect 26709 36193 26743 36227
rect 53757 36193 53791 36227
rect 2421 36125 2455 36159
rect 2881 36125 2915 36159
rect 25237 36125 25271 36159
rect 25330 36125 25364 36159
rect 25605 36125 25639 36159
rect 25743 36125 25777 36159
rect 26525 36125 26559 36159
rect 27169 36125 27203 36159
rect 27353 36125 27387 36159
rect 27537 36125 27571 36159
rect 28365 36125 28399 36159
rect 28457 36125 28491 36159
rect 28549 36125 28583 36159
rect 28733 36125 28767 36159
rect 52377 36125 52411 36159
rect 53021 36125 53055 36159
rect 53481 36125 53515 36159
rect 21281 36057 21315 36091
rect 25513 36057 25547 36091
rect 27445 36057 27479 36091
rect 22937 35989 22971 36023
rect 24041 35989 24075 36023
rect 25881 35989 25915 36023
rect 27721 35989 27755 36023
rect 28181 35989 28215 36023
rect 30297 35989 30331 36023
rect 30941 35989 30975 36023
rect 32597 35989 32631 36023
rect 52837 35989 52871 36023
rect 23029 35785 23063 35819
rect 24225 35785 24259 35819
rect 26617 35785 26651 35819
rect 23857 35717 23891 35751
rect 23949 35717 23983 35751
rect 25053 35717 25087 35751
rect 26341 35717 26375 35751
rect 27537 35717 27571 35751
rect 28733 35717 28767 35751
rect 29377 35717 29411 35751
rect 2145 35649 2179 35683
rect 23581 35649 23615 35683
rect 23674 35649 23708 35683
rect 24046 35649 24080 35683
rect 24685 35649 24719 35683
rect 24778 35649 24812 35683
rect 24961 35649 24995 35683
rect 25150 35649 25184 35683
rect 26065 35649 26099 35683
rect 26249 35649 26283 35683
rect 26433 35649 26467 35683
rect 27307 35649 27341 35683
rect 27445 35649 27479 35683
rect 27720 35649 27754 35683
rect 27813 35649 27847 35683
rect 28365 35649 28399 35683
rect 29929 35649 29963 35683
rect 30021 35649 30055 35683
rect 30205 35649 30239 35683
rect 30297 35649 30331 35683
rect 32413 35649 32447 35683
rect 2421 35581 2455 35615
rect 2881 35581 2915 35615
rect 30481 35581 30515 35615
rect 52377 35581 52411 35615
rect 53481 35581 53515 35615
rect 53757 35581 53791 35615
rect 22569 35513 22603 35547
rect 32965 35513 32999 35547
rect 20269 35445 20303 35479
rect 20821 35445 20855 35479
rect 21465 35445 21499 35479
rect 25329 35445 25363 35479
rect 27169 35445 27203 35479
rect 29285 35445 29319 35479
rect 31033 35445 31067 35479
rect 31585 35445 31619 35479
rect 53021 35445 53055 35479
rect 16589 35241 16623 35275
rect 27997 35241 28031 35275
rect 29193 35241 29227 35275
rect 15485 35173 15519 35207
rect 27077 35173 27111 35207
rect 32229 35173 32263 35207
rect 32873 35173 32907 35207
rect 15945 35105 15979 35139
rect 21189 35105 21223 35139
rect 22293 35105 22327 35139
rect 53757 35105 53791 35139
rect 1593 35037 1627 35071
rect 2789 35037 2823 35071
rect 14841 35037 14875 35071
rect 14934 35037 14968 35071
rect 15209 35037 15243 35071
rect 15347 35037 15381 35071
rect 21741 35037 21775 35071
rect 22845 35037 22879 35071
rect 23465 35037 23499 35071
rect 23857 35037 23891 35071
rect 25145 35037 25179 35071
rect 25697 35037 25731 35071
rect 25881 35037 25915 35071
rect 26065 35037 26099 35071
rect 26525 35037 26559 35071
rect 26709 35037 26743 35071
rect 26801 35037 26835 35071
rect 26945 35037 26979 35071
rect 28641 35037 28675 35071
rect 29055 35037 29089 35071
rect 30113 35037 30147 35071
rect 30261 35037 30295 35071
rect 30619 35037 30653 35071
rect 31493 35037 31527 35071
rect 53021 35037 53055 35071
rect 53481 35037 53515 35071
rect 15117 34969 15151 35003
rect 23581 34969 23615 35003
rect 23673 34969 23707 35003
rect 28089 34969 28123 35003
rect 28825 34969 28859 35003
rect 28917 34969 28951 35003
rect 30389 34969 30423 35003
rect 30481 34969 30515 35003
rect 1777 34901 1811 34935
rect 2329 34901 2363 34935
rect 14381 34901 14415 34935
rect 23305 34901 23339 34935
rect 25053 34901 25087 34935
rect 30757 34901 30791 34935
rect 31677 34901 31711 34935
rect 33425 34901 33459 34935
rect 24593 34697 24627 34731
rect 25605 34697 25639 34731
rect 27353 34697 27387 34731
rect 32413 34697 32447 34731
rect 24225 34629 24259 34663
rect 25329 34629 25363 34663
rect 26249 34629 26283 34663
rect 51733 34629 51767 34663
rect 2145 34561 2179 34595
rect 14013 34561 14047 34595
rect 14197 34561 14231 34595
rect 14289 34561 14323 34595
rect 14427 34561 14461 34595
rect 15669 34561 15703 34595
rect 24041 34561 24075 34595
rect 24317 34561 24351 34595
rect 24455 34561 24489 34595
rect 27261 34561 27295 34595
rect 28273 34561 28307 34595
rect 28365 34561 28399 34595
rect 28549 34561 28583 34595
rect 28641 34561 28675 34595
rect 29285 34561 29319 34595
rect 29378 34561 29412 34595
rect 29561 34561 29595 34595
rect 29653 34561 29687 34595
rect 29791 34561 29825 34595
rect 30389 34561 30423 34595
rect 30481 34561 30515 34595
rect 30665 34561 30699 34595
rect 30757 34561 30791 34595
rect 52193 34561 52227 34595
rect 53481 34561 53515 34595
rect 53757 34561 53791 34595
rect 2421 34493 2455 34527
rect 13461 34493 13495 34527
rect 15025 34493 15059 34527
rect 21373 34493 21407 34527
rect 23581 34493 23615 34527
rect 31585 34493 31619 34527
rect 53021 34493 53055 34527
rect 14565 34425 14599 34459
rect 23029 34425 23063 34459
rect 29929 34425 29963 34459
rect 32873 34425 32907 34459
rect 52377 34425 52411 34459
rect 22477 34357 22511 34391
rect 26341 34357 26375 34391
rect 28825 34357 28859 34391
rect 30941 34357 30975 34391
rect 14749 34153 14783 34187
rect 22293 34153 22327 34187
rect 22845 34153 22879 34187
rect 23489 34153 23523 34187
rect 24041 34153 24075 34187
rect 24777 34153 24811 34187
rect 25789 34153 25823 34187
rect 31401 34153 31435 34187
rect 32045 34153 32079 34187
rect 26249 34085 26283 34119
rect 30849 34085 30883 34119
rect 53389 34085 53423 34119
rect 2145 34017 2179 34051
rect 26617 34017 26651 34051
rect 28181 34017 28215 34051
rect 28917 34017 28951 34051
rect 2421 33949 2455 33983
rect 2881 33949 2915 33983
rect 25329 33949 25363 33983
rect 25605 33949 25639 33983
rect 26893 33949 26927 33983
rect 27353 33949 27387 33983
rect 27537 33949 27571 33983
rect 27997 33949 28031 33983
rect 30021 33949 30055 33983
rect 30113 33949 30147 33983
rect 30297 33949 30331 33983
rect 30389 33949 30423 33983
rect 53521 33949 53555 33983
rect 53665 33949 53699 33983
rect 53941 33949 53975 33983
rect 26408 33881 26442 33915
rect 52745 33881 52779 33915
rect 53757 33881 53791 33915
rect 25421 33813 25455 33847
rect 26525 33813 26559 33847
rect 27445 33813 27479 33847
rect 29837 33813 29871 33847
rect 24225 33609 24259 33643
rect 27445 33609 27479 33643
rect 27813 33609 27847 33643
rect 53113 33609 53147 33643
rect 23857 33541 23891 33575
rect 27353 33541 27387 33575
rect 23673 33473 23707 33507
rect 23949 33473 23983 33507
rect 24041 33473 24075 33507
rect 24685 33473 24719 33507
rect 24961 33473 24995 33507
rect 25605 33473 25639 33507
rect 25789 33473 25823 33507
rect 26341 33473 26375 33507
rect 27261 33473 27295 33507
rect 29101 33473 29135 33507
rect 29745 33473 29779 33507
rect 2145 33405 2179 33439
rect 2421 33405 2455 33439
rect 2881 33405 2915 33439
rect 25513 33405 25547 33439
rect 27997 33405 28031 33439
rect 29377 33405 29411 33439
rect 29653 33405 29687 33439
rect 30573 33405 30607 33439
rect 24685 33337 24719 33371
rect 24777 33337 24811 33371
rect 30113 33337 30147 33371
rect 23121 33269 23155 33303
rect 31217 33269 31251 33303
rect 54309 33269 54343 33303
rect 23397 33065 23431 33099
rect 25605 33065 25639 33099
rect 26065 33065 26099 33099
rect 27905 33065 27939 33099
rect 29009 33065 29043 33099
rect 26801 32997 26835 33031
rect 25329 32929 25363 32963
rect 27445 32929 27479 32963
rect 1593 32861 1627 32895
rect 2789 32861 2823 32895
rect 25237 32861 25271 32895
rect 25421 32861 25455 32895
rect 28089 32861 28123 32895
rect 28181 32861 28215 32895
rect 28365 32861 28399 32895
rect 28457 32861 28491 32895
rect 54309 32861 54343 32895
rect 26801 32793 26835 32827
rect 1777 32725 1811 32759
rect 2329 32725 2363 32759
rect 24593 32725 24627 32759
rect 26249 32725 26283 32759
rect 26341 32725 26375 32759
rect 29837 32725 29871 32759
rect 25605 32521 25639 32555
rect 27261 32521 27295 32555
rect 24593 32453 24627 32487
rect 28365 32453 28399 32487
rect 25789 32385 25823 32419
rect 26341 32385 26375 32419
rect 27169 32385 27203 32419
rect 27353 32385 27387 32419
rect 2145 32317 2179 32351
rect 2421 32317 2455 32351
rect 26433 32317 26467 32351
rect 27813 32249 27847 32283
rect 24869 32181 24903 32215
rect 24961 31977 24995 32011
rect 26065 31977 26099 32011
rect 27261 31909 27295 31943
rect 2145 31773 2179 31807
rect 2421 31773 2455 31807
rect 2881 31773 2915 31807
rect 26617 31773 26651 31807
rect 26710 31773 26744 31807
rect 26985 31773 27019 31807
rect 27082 31773 27116 31807
rect 27905 31773 27939 31807
rect 54309 31773 54343 31807
rect 26893 31705 26927 31739
rect 27721 31705 27755 31739
rect 25605 31637 25639 31671
rect 28089 31637 28123 31671
rect 26433 31433 26467 31467
rect 26341 31365 26375 31399
rect 26525 31365 26559 31399
rect 2145 31297 2179 31331
rect 28365 31297 28399 31331
rect 2421 31229 2455 31263
rect 2881 31229 2915 31263
rect 25789 31229 25823 31263
rect 25973 31229 26007 31263
rect 28089 31229 28123 31263
rect 54309 31093 54343 31127
rect 27261 30889 27295 30923
rect 2145 30753 2179 30787
rect 2421 30685 2455 30719
rect 2881 30685 2915 30719
rect 26709 30685 26743 30719
rect 26893 30685 26927 30719
rect 27077 30685 27111 30719
rect 26985 30617 27019 30651
rect 26157 30549 26191 30583
rect 27813 30549 27847 30583
rect 26341 30345 26375 30379
rect 2145 30209 2179 30243
rect 54033 30209 54067 30243
rect 2421 30141 2455 30175
rect 53481 30005 53515 30039
rect 54217 30005 54251 30039
rect 2237 29801 2271 29835
rect 26893 29801 26927 29835
rect 1593 29597 1627 29631
rect 2789 29597 2823 29631
rect 53573 29597 53607 29631
rect 54217 29597 54251 29631
rect 27905 29529 27939 29563
rect 1777 29461 1811 29495
rect 54125 29461 54159 29495
rect 25973 29257 26007 29291
rect 28273 29257 28307 29291
rect 54217 29257 54251 29291
rect 14105 29189 14139 29223
rect 27445 29189 27479 29223
rect 2145 29121 2179 29155
rect 13829 29121 13863 29155
rect 14013 29121 14047 29155
rect 14197 29121 14231 29155
rect 26525 29121 26559 29155
rect 27169 29121 27203 29155
rect 27353 29121 27387 29155
rect 27537 29121 27571 29155
rect 54033 29121 54067 29155
rect 2421 29053 2455 29087
rect 2881 29053 2915 29087
rect 14841 29053 14875 29087
rect 14381 28985 14415 29019
rect 53481 28985 53515 29019
rect 27721 28917 27755 28951
rect 53021 28917 53055 28951
rect 27077 28713 27111 28747
rect 28917 28713 28951 28747
rect 28365 28645 28399 28679
rect 2145 28509 2179 28543
rect 2421 28509 2455 28543
rect 2881 28509 2915 28543
rect 25605 28509 25639 28543
rect 27077 28509 27111 28543
rect 28181 28509 28215 28543
rect 28365 28509 28399 28543
rect 29745 28509 29779 28543
rect 54217 28509 54251 28543
rect 26525 28441 26559 28475
rect 29929 28441 29963 28475
rect 52837 28441 52871 28475
rect 53481 28441 53515 28475
rect 14565 28373 14599 28407
rect 25145 28373 25179 28407
rect 26433 28373 26467 28407
rect 30113 28373 30147 28407
rect 53389 28373 53423 28407
rect 54125 28373 54159 28407
rect 24685 28169 24719 28203
rect 26617 28169 26651 28203
rect 27813 28169 27847 28203
rect 54217 28169 54251 28203
rect 25237 28101 25271 28135
rect 25881 28101 25915 28135
rect 27537 28101 27571 28135
rect 2145 28033 2179 28067
rect 26433 28033 26467 28067
rect 27169 28033 27203 28067
rect 27262 28033 27296 28067
rect 27445 28033 27479 28067
rect 27634 28033 27668 28067
rect 28273 28033 28307 28067
rect 53297 28033 53331 28067
rect 54033 28033 54067 28067
rect 2421 27965 2455 27999
rect 26341 27965 26375 27999
rect 28365 27965 28399 27999
rect 25881 27897 25915 27931
rect 29101 27897 29135 27931
rect 28273 27829 28307 27863
rect 28641 27829 28675 27863
rect 52285 27829 52319 27863
rect 53481 27829 53515 27863
rect 2237 27625 2271 27659
rect 25053 27625 25087 27659
rect 26433 27557 26467 27591
rect 27169 27557 27203 27591
rect 24041 27489 24075 27523
rect 28273 27489 28307 27523
rect 1593 27421 1627 27455
rect 2789 27421 2823 27455
rect 25053 27421 25087 27455
rect 25237 27421 25271 27455
rect 25881 27421 25915 27455
rect 26249 27421 26283 27455
rect 27307 27421 27341 27455
rect 27445 27421 27479 27455
rect 27720 27421 27754 27455
rect 27813 27421 27847 27455
rect 28549 27421 28583 27455
rect 29929 27421 29963 27455
rect 52469 27421 52503 27455
rect 53481 27421 53515 27455
rect 53757 27421 53791 27455
rect 26065 27353 26099 27387
rect 26157 27353 26191 27387
rect 27537 27353 27571 27387
rect 1777 27285 1811 27319
rect 25421 27285 25455 27319
rect 29837 27285 29871 27319
rect 52929 27285 52963 27319
rect 24409 27081 24443 27115
rect 25513 27081 25547 27115
rect 28825 27081 28859 27115
rect 34529 27081 34563 27115
rect 35909 27081 35943 27115
rect 51825 27013 51859 27047
rect 54217 27013 54251 27047
rect 26065 26945 26099 26979
rect 27537 26945 27571 26979
rect 28089 26945 28123 26979
rect 52377 26945 52411 26979
rect 53481 26945 53515 26979
rect 2145 26877 2179 26911
rect 2421 26877 2455 26911
rect 2881 26877 2915 26911
rect 25053 26877 25087 26911
rect 26525 26877 26559 26911
rect 27261 26809 27295 26843
rect 54033 26809 54067 26843
rect 26341 26741 26375 26775
rect 28273 26741 28307 26775
rect 35081 26741 35115 26775
rect 53389 26741 53423 26775
rect 26065 26537 26099 26571
rect 34345 26537 34379 26571
rect 36001 26537 36035 26571
rect 36553 26537 36587 26571
rect 37197 26537 37231 26571
rect 54217 26537 54251 26571
rect 26801 26469 26835 26503
rect 35541 26469 35575 26503
rect 53389 26469 53423 26503
rect 2145 26401 2179 26435
rect 25513 26401 25547 26435
rect 26249 26401 26283 26435
rect 2421 26333 2455 26367
rect 26341 26333 26375 26367
rect 28181 26333 28215 26367
rect 52837 26333 52871 26367
rect 53573 26333 53607 26367
rect 54033 26333 54067 26367
rect 26801 26265 26835 26299
rect 27353 26265 27387 26299
rect 27537 26265 27571 26299
rect 33333 26197 33367 26231
rect 34897 26197 34931 26231
rect 2237 25993 2271 26027
rect 26433 25993 26467 26027
rect 27261 25993 27295 26027
rect 32597 25993 32631 26027
rect 33609 25993 33643 26027
rect 35817 25993 35851 26027
rect 37473 25993 37507 26027
rect 38209 25993 38243 26027
rect 1593 25857 1627 25891
rect 25421 25857 25455 25891
rect 26249 25857 26283 25891
rect 27537 25857 27571 25891
rect 34529 25857 34563 25891
rect 35357 25857 35391 25891
rect 33149 25789 33183 25823
rect 34345 25789 34379 25823
rect 52377 25789 52411 25823
rect 53481 25789 53515 25823
rect 53757 25789 53791 25823
rect 1777 25721 1811 25755
rect 36461 25721 36495 25755
rect 25237 25653 25271 25687
rect 34713 25653 34747 25687
rect 35173 25653 35207 25687
rect 38853 25653 38887 25687
rect 52929 25653 52963 25687
rect 2237 25449 2271 25483
rect 25697 25449 25731 25483
rect 29009 25449 29043 25483
rect 31953 25449 31987 25483
rect 32413 25449 32447 25483
rect 35265 25449 35299 25483
rect 37657 25449 37691 25483
rect 52745 25449 52779 25483
rect 54217 25449 54251 25483
rect 39221 25381 39255 25415
rect 25697 25313 25731 25347
rect 26065 25313 26099 25347
rect 1593 25245 1627 25279
rect 2789 25245 2823 25279
rect 24869 25245 24903 25279
rect 26617 25245 26651 25279
rect 26985 25245 27019 25279
rect 27537 25245 27571 25279
rect 28181 25245 28215 25279
rect 28825 25245 28859 25279
rect 33149 25245 33183 25279
rect 33793 25245 33827 25279
rect 34069 25245 34103 25279
rect 34161 25245 34195 25279
rect 34989 25245 35023 25279
rect 35081 25245 35115 25279
rect 35909 25245 35943 25279
rect 36369 25245 36403 25279
rect 38393 25245 38427 25279
rect 39037 25245 39071 25279
rect 53297 25245 53331 25279
rect 54033 25245 54067 25279
rect 28641 25177 28675 25211
rect 31401 25177 31435 25211
rect 33977 25177 34011 25211
rect 40049 25177 40083 25211
rect 1777 25109 1811 25143
rect 25053 25109 25087 25143
rect 25881 25109 25915 25143
rect 26617 25109 26651 25143
rect 33333 25109 33367 25143
rect 34345 25109 34379 25143
rect 35725 25109 35759 25143
rect 36553 25109 36587 25143
rect 37105 25109 37139 25143
rect 38577 25109 38611 25143
rect 53481 25109 53515 25143
rect 26433 24905 26467 24939
rect 28549 24905 28583 24939
rect 31493 24905 31527 24939
rect 33149 24905 33183 24939
rect 34989 24905 35023 24939
rect 25298 24837 25332 24871
rect 33854 24837 33888 24871
rect 35716 24837 35750 24871
rect 1685 24769 1719 24803
rect 2329 24769 2363 24803
rect 24409 24769 24443 24803
rect 27425 24769 27459 24803
rect 29193 24769 29227 24803
rect 30757 24769 30791 24803
rect 32873 24769 32907 24803
rect 32965 24769 32999 24803
rect 37749 24769 37783 24803
rect 38660 24769 38694 24803
rect 40417 24769 40451 24803
rect 53297 24769 53331 24803
rect 54217 24769 54251 24803
rect 25053 24701 25087 24735
rect 27169 24701 27203 24735
rect 33609 24701 33643 24735
rect 35449 24701 35483 24735
rect 38393 24701 38427 24735
rect 24593 24633 24627 24667
rect 36829 24633 36863 24667
rect 54033 24633 54067 24667
rect 1777 24565 1811 24599
rect 23949 24565 23983 24599
rect 29101 24565 29135 24599
rect 30941 24565 30975 24599
rect 37933 24565 37967 24599
rect 39773 24565 39807 24599
rect 40601 24565 40635 24599
rect 53481 24565 53515 24599
rect 14657 24361 14691 24395
rect 15209 24361 15243 24395
rect 24041 24361 24075 24395
rect 26341 24361 26375 24395
rect 28273 24361 28307 24395
rect 30941 24361 30975 24395
rect 33701 24361 33735 24395
rect 36277 24361 36311 24395
rect 38577 24361 38611 24395
rect 41429 24361 41463 24395
rect 53573 24361 53607 24395
rect 38117 24293 38151 24327
rect 39405 24293 39439 24327
rect 23121 24225 23155 24259
rect 23857 24225 23891 24259
rect 30573 24225 30607 24259
rect 31401 24225 31435 24259
rect 32873 24225 32907 24259
rect 34897 24225 34931 24259
rect 40049 24225 40083 24259
rect 14749 24157 14783 24191
rect 23765 24157 23799 24191
rect 24961 24157 24995 24191
rect 26893 24157 26927 24191
rect 30757 24157 30791 24191
rect 31585 24157 31619 24191
rect 31769 24157 31803 24191
rect 32413 24157 32447 24191
rect 33057 24157 33091 24191
rect 33885 24157 33919 24191
rect 33977 24157 34011 24191
rect 34253 24157 34287 24191
rect 36737 24157 36771 24191
rect 36993 24157 37027 24191
rect 38761 24157 38795 24191
rect 38945 24157 38979 24191
rect 40305 24157 40339 24191
rect 53021 24157 53055 24191
rect 54217 24157 54251 24191
rect 1685 24089 1719 24123
rect 2329 24089 2363 24123
rect 24041 24089 24075 24123
rect 25228 24089 25262 24123
rect 27160 24089 27194 24123
rect 34069 24089 34103 24123
rect 35164 24089 35198 24123
rect 1777 24021 1811 24055
rect 14289 24021 14323 24055
rect 23581 24021 23615 24055
rect 30113 24021 30147 24055
rect 32229 24021 32263 24055
rect 33241 24021 33275 24055
rect 54125 24021 54159 24055
rect 24961 23817 24995 23851
rect 27537 23817 27571 23851
rect 31769 23817 31803 23851
rect 32597 23817 32631 23851
rect 34437 23817 34471 23851
rect 35725 23817 35759 23851
rect 37841 23817 37875 23851
rect 40233 23817 40267 23851
rect 24593 23749 24627 23783
rect 36461 23749 36495 23783
rect 36553 23749 36587 23783
rect 38546 23749 38580 23783
rect 40938 23749 40972 23783
rect 54217 23749 54251 23783
rect 1869 23681 1903 23715
rect 22753 23681 22787 23715
rect 23673 23681 23707 23715
rect 25697 23681 25731 23715
rect 26157 23681 26191 23715
rect 30021 23681 30055 23715
rect 31125 23681 31159 23715
rect 32689 23681 32723 23715
rect 33885 23681 33919 23715
rect 34069 23681 34103 23715
rect 34161 23681 34195 23715
rect 34253 23681 34287 23715
rect 35541 23681 35575 23715
rect 36369 23681 36403 23715
rect 36737 23681 36771 23715
rect 37657 23681 37691 23715
rect 38301 23681 38335 23715
rect 40693 23681 40727 23715
rect 53481 23681 53515 23715
rect 23213 23613 23247 23647
rect 24317 23613 24351 23647
rect 24501 23613 24535 23647
rect 26341 23613 26375 23647
rect 27629 23613 27663 23647
rect 27721 23613 27755 23647
rect 28365 23613 28399 23647
rect 32413 23613 32447 23647
rect 35357 23613 35391 23647
rect 37473 23613 37507 23647
rect 54033 23613 54067 23647
rect 2421 23545 2455 23579
rect 22569 23545 22603 23579
rect 25605 23545 25639 23579
rect 29469 23545 29503 23579
rect 36185 23545 36219 23579
rect 42073 23545 42107 23579
rect 53297 23545 53331 23579
rect 1685 23477 1719 23511
rect 14841 23477 14875 23511
rect 22109 23477 22143 23511
rect 23397 23477 23431 23511
rect 27169 23477 27203 23511
rect 29009 23477 29043 23511
rect 30205 23477 30239 23511
rect 30849 23477 30883 23511
rect 33057 23477 33091 23511
rect 39681 23477 39715 23511
rect 22569 23273 22603 23307
rect 24041 23273 24075 23307
rect 24777 23273 24811 23307
rect 25881 23273 25915 23307
rect 27077 23273 27111 23307
rect 29101 23273 29135 23307
rect 38117 23273 38151 23307
rect 40417 23273 40451 23307
rect 54217 23273 54251 23307
rect 35633 23205 35667 23239
rect 42349 23205 42383 23239
rect 53573 23205 53607 23239
rect 23949 23137 23983 23171
rect 24869 23137 24903 23171
rect 26433 23137 26467 23171
rect 28365 23137 28399 23171
rect 33793 23137 33827 23171
rect 34069 23137 34103 23171
rect 34989 23137 35023 23171
rect 40049 23137 40083 23171
rect 40969 23137 41003 23171
rect 1869 23069 1903 23103
rect 23213 23069 23247 23103
rect 24041 23069 24075 23103
rect 24961 23069 24995 23103
rect 26249 23069 26283 23103
rect 27261 23069 27295 23103
rect 29837 23069 29871 23103
rect 31677 23069 31711 23103
rect 34161 23069 34195 23103
rect 36461 23069 36495 23103
rect 37105 23069 37139 23103
rect 37565 23069 37599 23103
rect 37749 23069 37783 23103
rect 37933 23069 37967 23103
rect 38577 23069 38611 23103
rect 38761 23069 38795 23103
rect 38945 23069 38979 23103
rect 40233 23069 40267 23103
rect 42993 23069 43027 23103
rect 54033 23069 54067 23103
rect 30104 23001 30138 23035
rect 31922 23001 31956 23035
rect 37841 23001 37875 23035
rect 38853 23001 38887 23035
rect 41236 23001 41270 23035
rect 1685 22933 1719 22967
rect 14657 22933 14691 22967
rect 23029 22933 23063 22967
rect 23673 22933 23707 22967
rect 24593 22933 24627 22967
rect 26341 22933 26375 22967
rect 27813 22933 27847 22967
rect 31217 22933 31251 22967
rect 33057 22933 33091 22967
rect 35173 22933 35207 22967
rect 35265 22933 35299 22967
rect 39129 22933 39163 22967
rect 42809 22933 42843 22967
rect 2329 22729 2363 22763
rect 14933 22729 14967 22763
rect 22937 22729 22971 22763
rect 24777 22729 24811 22763
rect 25329 22729 25363 22763
rect 25697 22729 25731 22763
rect 29929 22729 29963 22763
rect 31769 22729 31803 22763
rect 32321 22729 32355 22763
rect 32689 22729 32723 22763
rect 33885 22729 33919 22763
rect 35541 22729 35575 22763
rect 36001 22729 36035 22763
rect 38025 22729 38059 22763
rect 39313 22729 39347 22763
rect 53481 22729 53515 22763
rect 54217 22729 54251 22763
rect 33793 22661 33827 22695
rect 35081 22661 35115 22695
rect 36369 22661 36403 22695
rect 37657 22661 37691 22695
rect 38945 22661 38979 22695
rect 39773 22661 39807 22695
rect 43269 22661 43303 22695
rect 1869 22593 1903 22627
rect 2513 22593 2547 22627
rect 14473 22593 14507 22627
rect 15393 22593 15427 22627
rect 15853 22593 15887 22627
rect 23489 22593 23523 22627
rect 27537 22593 27571 22627
rect 27721 22593 27755 22627
rect 28365 22593 28399 22627
rect 29101 22593 29135 22627
rect 29653 22593 29687 22627
rect 29745 22593 29779 22627
rect 30389 22593 30423 22627
rect 30656 22593 30690 22627
rect 35173 22593 35207 22627
rect 36461 22593 36495 22627
rect 37473 22593 37507 22627
rect 37749 22593 37783 22627
rect 37841 22593 37875 22627
rect 38761 22593 38795 22627
rect 39037 22593 39071 22627
rect 39129 22593 39163 22627
rect 39957 22593 39991 22627
rect 40693 22593 40727 22627
rect 40960 22593 40994 22627
rect 42809 22593 42843 22627
rect 54033 22593 54067 22627
rect 23765 22525 23799 22559
rect 25789 22525 25823 22559
rect 25881 22525 25915 22559
rect 27353 22525 27387 22559
rect 32781 22525 32815 22559
rect 32873 22525 32907 22559
rect 33609 22525 33643 22559
rect 34897 22525 34931 22559
rect 36553 22525 36587 22559
rect 40141 22525 40175 22559
rect 42625 22457 42659 22491
rect 1685 22389 1719 22423
rect 14013 22389 14047 22423
rect 14381 22389 14415 22423
rect 15301 22389 15335 22423
rect 22477 22389 22511 22423
rect 26525 22389 26559 22423
rect 28181 22389 28215 22423
rect 34253 22389 34287 22423
rect 42073 22389 42107 22423
rect 14749 22185 14783 22219
rect 22753 22185 22787 22219
rect 30941 22185 30975 22219
rect 40601 22185 40635 22219
rect 43361 22185 43395 22219
rect 2421 22117 2455 22151
rect 36737 22117 36771 22151
rect 15485 22049 15519 22083
rect 20729 22049 20763 22083
rect 21281 22049 21315 22083
rect 27445 22049 27479 22083
rect 29837 22049 29871 22083
rect 31493 22049 31527 22083
rect 32781 22049 32815 22083
rect 36277 22049 36311 22083
rect 37565 22049 37599 22083
rect 37749 22049 37783 22083
rect 41429 22049 41463 22083
rect 42809 22049 42843 22083
rect 1869 21981 1903 22015
rect 21925 21981 21959 22015
rect 22845 21981 22879 22015
rect 23765 21981 23799 22015
rect 24777 21981 24811 22015
rect 24961 21981 24995 22015
rect 25789 21981 25823 22015
rect 25973 21981 26007 22015
rect 27712 21981 27746 22015
rect 31309 21981 31343 22015
rect 32505 21981 32539 22015
rect 33885 21981 33919 22015
rect 36921 21981 36955 22015
rect 38669 21981 38703 22015
rect 38839 21981 38873 22015
rect 40049 21981 40083 22015
rect 40417 21981 40451 22015
rect 41061 21981 41095 22015
rect 41245 21981 41279 22015
rect 41889 21981 41923 22015
rect 42073 21981 42107 22015
rect 42257 21981 42291 22015
rect 54217 21981 54251 22015
rect 26433 21913 26467 21947
rect 26617 21913 26651 21947
rect 26801 21913 26835 21947
rect 30113 21913 30147 21947
rect 36032 21913 36066 21947
rect 40233 21913 40267 21947
rect 40325 21913 40359 21947
rect 53297 21913 53331 21947
rect 53481 21913 53515 21947
rect 54033 21913 54067 21947
rect 1685 21845 1719 21879
rect 22385 21845 22419 21879
rect 23581 21845 23615 21879
rect 24593 21845 24627 21879
rect 25605 21845 25639 21879
rect 28825 21845 28859 21879
rect 30021 21845 30055 21879
rect 30481 21845 30515 21879
rect 31401 21845 31435 21879
rect 32137 21845 32171 21879
rect 32597 21845 32631 21879
rect 33333 21845 33367 21879
rect 34897 21845 34931 21879
rect 37841 21845 37875 21879
rect 38209 21845 38243 21879
rect 39037 21845 39071 21879
rect 43821 21845 43855 21879
rect 52837 21845 52871 21879
rect 2421 21641 2455 21675
rect 25329 21641 25363 21675
rect 27169 21641 27203 21675
rect 33517 21641 33551 21675
rect 35449 21641 35483 21675
rect 35909 21641 35943 21675
rect 40049 21641 40083 21675
rect 53573 21641 53607 21675
rect 54217 21641 54251 21675
rect 20821 21573 20855 21607
rect 28733 21573 28767 21607
rect 39773 21573 39807 21607
rect 42625 21573 42659 21607
rect 1869 21505 1903 21539
rect 14105 21505 14139 21539
rect 21465 21505 21499 21539
rect 22477 21505 22511 21539
rect 23305 21505 23339 21539
rect 23949 21505 23983 21539
rect 24205 21505 24239 21539
rect 25881 21505 25915 21539
rect 27537 21505 27571 21539
rect 31401 21505 31435 21539
rect 32689 21505 32723 21539
rect 35541 21505 35575 21539
rect 36553 21505 36587 21539
rect 36645 21505 36679 21539
rect 36737 21505 36771 21539
rect 38586 21505 38620 21539
rect 38853 21505 38887 21539
rect 39497 21505 39531 21539
rect 39681 21505 39715 21539
rect 39865 21505 39899 21539
rect 40960 21505 40994 21539
rect 54033 21505 54067 21539
rect 22017 21437 22051 21471
rect 27629 21437 27663 21471
rect 27721 21437 27755 21471
rect 28549 21437 28583 21471
rect 28641 21437 28675 21471
rect 29653 21437 29687 21471
rect 32413 21437 32447 21471
rect 32597 21437 32631 21471
rect 34713 21437 34747 21471
rect 35265 21437 35299 21471
rect 40693 21437 40727 21471
rect 21281 21369 21315 21403
rect 23489 21369 23523 21403
rect 33057 21369 33091 21403
rect 34069 21369 34103 21403
rect 36921 21369 36955 21403
rect 42073 21369 42107 21403
rect 1685 21301 1719 21335
rect 13921 21301 13955 21335
rect 22385 21301 22419 21335
rect 26433 21301 26467 21335
rect 29101 21301 29135 21335
rect 30205 21301 30239 21335
rect 30849 21301 30883 21335
rect 36369 21301 36403 21335
rect 37473 21301 37507 21335
rect 2421 21097 2455 21131
rect 22017 21097 22051 21131
rect 23029 21097 23063 21131
rect 26617 21097 26651 21131
rect 34897 21097 34931 21131
rect 40049 21097 40083 21131
rect 44005 21097 44039 21131
rect 19901 21029 19935 21063
rect 27905 21029 27939 21063
rect 42165 21029 42199 21063
rect 54217 21029 54251 21063
rect 20453 20961 20487 20995
rect 22661 20961 22695 20995
rect 28549 20961 28583 20995
rect 32321 20961 32355 20995
rect 33793 20961 33827 20995
rect 35541 20961 35575 20995
rect 36461 20961 36495 20995
rect 1869 20893 1903 20927
rect 22201 20893 22235 20927
rect 23121 20893 23155 20927
rect 23857 20893 23891 20927
rect 24593 20893 24627 20927
rect 27169 20893 27203 20927
rect 30297 20893 30331 20927
rect 31861 20893 31895 20927
rect 38945 20893 38979 20927
rect 39221 20893 39255 20927
rect 39313 20893 39347 20927
rect 40233 20893 40267 20927
rect 40785 20893 40819 20927
rect 42809 20893 42843 20927
rect 43453 20893 43487 20927
rect 54033 20893 54067 20927
rect 21005 20825 21039 20859
rect 24838 20825 24872 20859
rect 28641 20825 28675 20859
rect 35265 20825 35299 20859
rect 38209 20825 38243 20859
rect 39129 20825 39163 20859
rect 41052 20825 41086 20859
rect 1685 20757 1719 20791
rect 21465 20757 21499 20791
rect 24041 20757 24075 20791
rect 25973 20757 26007 20791
rect 28733 20757 28767 20791
rect 29101 20757 29135 20791
rect 29745 20757 29779 20791
rect 31217 20757 31251 20791
rect 32965 20757 32999 20791
rect 34345 20757 34379 20791
rect 35357 20757 35391 20791
rect 39497 20757 39531 20791
rect 42625 20757 42659 20791
rect 43269 20757 43303 20791
rect 53573 20757 53607 20791
rect 22017 20553 22051 20587
rect 23581 20553 23615 20587
rect 24041 20553 24075 20587
rect 24501 20553 24535 20587
rect 26617 20553 26651 20587
rect 27169 20553 27203 20587
rect 27813 20553 27847 20587
rect 29745 20553 29779 20587
rect 36093 20553 36127 20587
rect 39497 20553 39531 20587
rect 43177 20553 43211 20587
rect 44281 20553 44315 20587
rect 20361 20485 20395 20519
rect 20913 20485 20947 20519
rect 40785 20485 40819 20519
rect 54033 20485 54067 20519
rect 54217 20485 54251 20519
rect 1869 20417 1903 20451
rect 2421 20417 2455 20451
rect 19441 20417 19475 20451
rect 22201 20417 22235 20451
rect 23397 20417 23431 20451
rect 24409 20417 24443 20451
rect 25237 20417 25271 20451
rect 25493 20417 25527 20451
rect 27169 20417 27203 20451
rect 27353 20417 27387 20451
rect 28937 20417 28971 20451
rect 29193 20417 29227 20451
rect 29929 20417 29963 20451
rect 30021 20417 30055 20451
rect 30205 20417 30239 20451
rect 34969 20417 35003 20451
rect 36737 20417 36771 20451
rect 41383 20417 41417 20451
rect 41521 20417 41555 20451
rect 41613 20417 41647 20451
rect 41797 20417 41831 20451
rect 43729 20417 43763 20451
rect 53297 20417 53331 20451
rect 53481 20417 53515 20451
rect 23213 20349 23247 20383
rect 24685 20349 24719 20383
rect 30113 20349 30147 20383
rect 31493 20349 31527 20383
rect 32321 20349 32355 20383
rect 33609 20349 33643 20383
rect 34713 20349 34747 20383
rect 36553 20349 36587 20383
rect 37565 20349 37599 20383
rect 21373 20281 21407 20315
rect 22753 20281 22787 20315
rect 32965 20281 32999 20315
rect 36921 20281 36955 20315
rect 1685 20213 1719 20247
rect 19257 20213 19291 20247
rect 30849 20213 30883 20247
rect 34253 20213 34287 20247
rect 38117 20213 38151 20247
rect 41245 20213 41279 20247
rect 42625 20213 42659 20247
rect 2421 20009 2455 20043
rect 19625 20009 19659 20043
rect 24593 20009 24627 20043
rect 27169 20009 27203 20043
rect 32689 20009 32723 20043
rect 34897 20009 34931 20043
rect 39313 20009 39347 20043
rect 42441 20009 42475 20043
rect 54217 20009 54251 20043
rect 22017 19941 22051 19975
rect 27997 19941 28031 19975
rect 32229 19941 32263 19975
rect 37473 19941 37507 19975
rect 53573 19941 53607 19975
rect 20269 19873 20303 19907
rect 22569 19873 22603 19907
rect 23489 19873 23523 19907
rect 24041 19873 24075 19907
rect 25145 19873 25179 19907
rect 25789 19873 25823 19907
rect 28089 19873 28123 19907
rect 28549 19873 28583 19907
rect 30113 19873 30147 19907
rect 30849 19873 30883 19907
rect 38853 19873 38887 19907
rect 42073 19873 42107 19907
rect 1869 19805 1903 19839
rect 14473 19805 14507 19839
rect 19993 19805 20027 19839
rect 21373 19805 21407 19839
rect 22385 19805 22419 19839
rect 27629 19805 27663 19839
rect 30021 19805 30055 19839
rect 31116 19805 31150 19839
rect 34069 19805 34103 19839
rect 36277 19805 36311 19839
rect 36921 19805 36955 19839
rect 39497 19805 39531 19839
rect 41613 19805 41647 19839
rect 42257 19805 42291 19839
rect 54033 19805 54067 19839
rect 18889 19737 18923 19771
rect 22477 19737 22511 19771
rect 24961 19737 24995 19771
rect 26056 19737 26090 19771
rect 33824 19737 33858 19771
rect 36032 19737 36066 19771
rect 38608 19737 38642 19771
rect 41368 19737 41402 19771
rect 43453 19737 43487 19771
rect 1685 19669 1719 19703
rect 14289 19669 14323 19703
rect 20085 19669 20119 19703
rect 20821 19669 20855 19703
rect 21557 19669 21591 19703
rect 25053 19669 25087 19703
rect 29193 19669 29227 19703
rect 30389 19669 30423 19703
rect 36737 19669 36771 19703
rect 40233 19669 40267 19703
rect 42901 19669 42935 19703
rect 20085 19465 20119 19499
rect 22017 19465 22051 19499
rect 23949 19465 23983 19499
rect 25973 19465 26007 19499
rect 27629 19465 27663 19499
rect 29377 19465 29411 19499
rect 30481 19465 30515 19499
rect 33425 19465 33459 19499
rect 35725 19465 35759 19499
rect 37657 19465 37691 19499
rect 38025 19465 38059 19499
rect 38117 19465 38151 19499
rect 38853 19465 38887 19499
rect 39773 19465 39807 19499
rect 40509 19465 40543 19499
rect 41521 19465 41555 19499
rect 54217 19465 54251 19499
rect 31585 19397 31619 19431
rect 34590 19397 34624 19431
rect 40785 19397 40819 19431
rect 1869 19329 1903 19363
rect 18705 19329 18739 19363
rect 18972 19329 19006 19363
rect 21097 19329 21131 19363
rect 23130 19329 23164 19363
rect 23397 19329 23431 19363
rect 24133 19329 24167 19363
rect 24225 19329 24259 19363
rect 27537 19329 27571 19363
rect 27721 19329 27755 19363
rect 27905 19329 27939 19363
rect 28549 19329 28583 19363
rect 28733 19329 28767 19363
rect 29561 19329 29595 19363
rect 30021 19329 30055 19363
rect 32321 19329 32355 19363
rect 33609 19329 33643 19363
rect 39313 19329 39347 19363
rect 39773 19329 39807 19363
rect 39957 19329 39991 19363
rect 40693 19329 40727 19363
rect 40877 19329 40911 19363
rect 41061 19329 41095 19363
rect 41705 19329 41739 19363
rect 54033 19329 54067 19363
rect 21189 19261 21223 19295
rect 21281 19261 21315 19295
rect 25329 19261 25363 19295
rect 26525 19261 26559 19295
rect 27353 19261 27387 19295
rect 28641 19261 28675 19295
rect 28825 19261 28859 19295
rect 31033 19261 31067 19295
rect 32873 19261 32907 19295
rect 33793 19261 33827 19295
rect 34345 19261 34379 19295
rect 36185 19261 36219 19295
rect 38301 19261 38335 19295
rect 30297 19193 30331 19227
rect 38945 19193 38979 19227
rect 1685 19125 1719 19159
rect 18245 19125 18279 19159
rect 20729 19125 20763 19159
rect 24777 19125 24811 19159
rect 28365 19125 28399 19159
rect 36829 19125 36863 19159
rect 42625 19125 42659 19159
rect 53573 19125 53607 19159
rect 2421 18921 2455 18955
rect 24869 18921 24903 18955
rect 26525 18921 26559 18955
rect 29745 18921 29779 18955
rect 33241 18921 33275 18955
rect 34345 18921 34379 18955
rect 36001 18921 36035 18955
rect 37013 18921 37047 18955
rect 40049 18921 40083 18955
rect 54125 18921 54159 18955
rect 21097 18853 21131 18887
rect 27721 18853 27755 18887
rect 32781 18853 32815 18887
rect 34897 18853 34931 18887
rect 42533 18853 42567 18887
rect 22477 18785 22511 18819
rect 23765 18785 23799 18819
rect 24041 18785 24075 18819
rect 25881 18785 25915 18819
rect 26893 18785 26927 18819
rect 28733 18785 28767 18819
rect 31401 18785 31435 18819
rect 33517 18785 33551 18819
rect 33701 18785 33735 18819
rect 36277 18785 36311 18819
rect 36461 18785 36495 18819
rect 37657 18785 37691 18819
rect 41429 18785 41463 18819
rect 1869 18717 1903 18751
rect 19441 18717 19475 18751
rect 20453 18717 20487 18751
rect 23673 18717 23707 18751
rect 24685 18717 24719 18751
rect 26801 18717 26835 18751
rect 27537 18717 27571 18751
rect 30297 18717 30331 18751
rect 31668 18717 31702 18751
rect 33425 18717 33459 18751
rect 33609 18717 33643 18751
rect 35449 18717 35483 18751
rect 36185 18717 36219 18751
rect 36369 18717 36403 18751
rect 38301 18717 38335 18751
rect 38761 18717 38795 18751
rect 39037 18717 39071 18751
rect 39175 18717 39209 18751
rect 42073 18717 42107 18751
rect 54217 18717 54251 18751
rect 18797 18649 18831 18683
rect 22210 18649 22244 18683
rect 23029 18649 23063 18683
rect 38945 18649 38979 18683
rect 41184 18649 41218 18683
rect 53297 18649 53331 18683
rect 53481 18649 53515 18683
rect 1685 18581 1719 18615
rect 18337 18581 18371 18615
rect 19625 18581 19659 18615
rect 20637 18581 20671 18615
rect 25329 18581 25363 18615
rect 28181 18581 28215 18615
rect 30849 18581 30883 18615
rect 38117 18581 38151 18615
rect 39313 18581 39347 18615
rect 41889 18581 41923 18615
rect 43177 18581 43211 18615
rect 52837 18581 52871 18615
rect 20637 18377 20671 18411
rect 31585 18377 31619 18411
rect 38577 18377 38611 18411
rect 41981 18377 42015 18411
rect 43269 18377 43303 18411
rect 54217 18377 54251 18411
rect 21005 18309 21039 18343
rect 28089 18309 28123 18343
rect 28273 18309 28307 18343
rect 28457 18309 28491 18343
rect 30757 18309 30791 18343
rect 30941 18309 30975 18343
rect 32597 18309 32631 18343
rect 34704 18309 34738 18343
rect 1777 18241 1811 18275
rect 18797 18241 18831 18275
rect 19053 18241 19087 18275
rect 22477 18241 22511 18275
rect 23121 18241 23155 18275
rect 23377 18241 23411 18275
rect 24961 18241 24995 18275
rect 25228 18241 25262 18275
rect 27261 18241 27295 18275
rect 28181 18241 28215 18275
rect 30030 18241 30064 18275
rect 31585 18241 31619 18275
rect 31769 18241 31803 18275
rect 32505 18241 32539 18275
rect 32689 18241 32723 18275
rect 32873 18241 32907 18275
rect 33793 18241 33827 18275
rect 34437 18241 34471 18275
rect 37657 18241 37691 18275
rect 38393 18241 38427 18275
rect 39221 18241 39255 18275
rect 39865 18241 39899 18275
rect 40693 18241 40727 18275
rect 41521 18241 41555 18275
rect 42717 18241 42751 18275
rect 54033 18241 54067 18275
rect 21097 18173 21131 18207
rect 21281 18173 21315 18207
rect 30297 18173 30331 18207
rect 33425 18173 33459 18207
rect 33701 18173 33735 18207
rect 36277 18173 36311 18207
rect 38209 18173 38243 18207
rect 39681 18173 39715 18207
rect 40509 18173 40543 18207
rect 17785 18105 17819 18139
rect 27445 18105 27479 18139
rect 27905 18105 27939 18139
rect 31125 18105 31159 18139
rect 35817 18105 35851 18139
rect 40049 18105 40083 18139
rect 40877 18105 40911 18139
rect 1593 18037 1627 18071
rect 2329 18037 2363 18071
rect 18337 18037 18371 18071
rect 20177 18037 20211 18071
rect 22661 18037 22695 18071
rect 24501 18037 24535 18071
rect 26341 18037 26375 18071
rect 28917 18037 28951 18071
rect 32321 18037 32355 18071
rect 36921 18037 36955 18071
rect 37565 18037 37599 18071
rect 39037 18037 39071 18071
rect 41337 18037 41371 18071
rect 53481 18037 53515 18071
rect 23121 17833 23155 17867
rect 24593 17833 24627 17867
rect 30941 17833 30975 17867
rect 21281 17765 21315 17799
rect 22661 17765 22695 17799
rect 33977 17765 34011 17799
rect 41521 17765 41555 17799
rect 42165 17765 42199 17799
rect 42809 17765 42843 17799
rect 54217 17765 54251 17799
rect 18245 17697 18279 17731
rect 19441 17697 19475 17731
rect 21925 17697 21959 17731
rect 25145 17697 25179 17731
rect 27537 17697 27571 17731
rect 27721 17697 27755 17731
rect 28549 17697 28583 17731
rect 29929 17697 29963 17731
rect 32505 17697 32539 17731
rect 33701 17697 33735 17731
rect 35541 17697 35575 17731
rect 1869 17629 1903 17663
rect 18705 17629 18739 17663
rect 21649 17629 21683 17663
rect 22477 17629 22511 17663
rect 23305 17629 23339 17663
rect 23397 17629 23431 17663
rect 25789 17629 25823 17663
rect 27445 17629 27479 17663
rect 27629 17629 27663 17663
rect 28825 17629 28859 17663
rect 31125 17629 31159 17663
rect 31309 17629 31343 17663
rect 32229 17629 32263 17663
rect 33609 17629 33643 17663
rect 35265 17629 35299 17663
rect 38025 17629 38059 17663
rect 38669 17629 38703 17663
rect 38853 17629 38887 17663
rect 39037 17629 39071 17663
rect 40325 17629 40359 17663
rect 40785 17629 40819 17663
rect 41705 17629 41739 17663
rect 54033 17629 54067 17663
rect 19686 17561 19720 17595
rect 30113 17561 30147 17595
rect 37780 17561 37814 17595
rect 38945 17561 38979 17595
rect 40141 17561 40175 17595
rect 1685 17493 1719 17527
rect 17141 17493 17175 17527
rect 17693 17493 17727 17527
rect 18889 17493 18923 17527
rect 20821 17493 20855 17527
rect 21741 17493 21775 17527
rect 24041 17493 24075 17527
rect 24961 17493 24995 17527
rect 25053 17493 25087 17527
rect 26433 17493 26467 17527
rect 27905 17493 27939 17527
rect 28733 17493 28767 17527
rect 29193 17493 29227 17527
rect 30021 17493 30055 17527
rect 30481 17493 30515 17527
rect 31861 17493 31895 17527
rect 32321 17493 32355 17527
rect 34897 17493 34931 17527
rect 35357 17493 35391 17527
rect 36093 17493 36127 17527
rect 36645 17493 36679 17527
rect 39221 17493 39255 17527
rect 40969 17493 41003 17527
rect 43269 17493 43303 17527
rect 53573 17493 53607 17527
rect 17233 17289 17267 17323
rect 24685 17289 24719 17323
rect 27169 17289 27203 17323
rect 36737 17289 36771 17323
rect 37565 17289 37599 17323
rect 38853 17289 38887 17323
rect 41521 17289 41555 17323
rect 54125 17289 54159 17323
rect 16313 17221 16347 17255
rect 20085 17221 20119 17255
rect 22998 17221 23032 17255
rect 26350 17221 26384 17255
rect 39988 17221 40022 17255
rect 54217 17221 54251 17255
rect 1869 17153 1903 17187
rect 21097 17153 21131 17187
rect 22109 17153 22143 17187
rect 24593 17153 24627 17187
rect 24777 17153 24811 17187
rect 26617 17153 26651 17187
rect 28365 17153 28399 17187
rect 28621 17153 28655 17187
rect 30205 17153 30239 17187
rect 30472 17153 30506 17187
rect 33445 17153 33479 17187
rect 33701 17153 33735 17187
rect 35561 17153 35595 17187
rect 35817 17153 35851 17187
rect 36461 17153 36495 17187
rect 38209 17153 38243 17187
rect 40233 17153 40267 17187
rect 40877 17153 40911 17187
rect 41705 17153 41739 17187
rect 53481 17153 53515 17187
rect 18337 17085 18371 17119
rect 20913 17085 20947 17119
rect 21005 17085 21039 17119
rect 22753 17085 22787 17119
rect 27721 17085 27755 17119
rect 38025 17085 38059 17119
rect 40693 17085 40727 17119
rect 29745 17017 29779 17051
rect 34437 17017 34471 17051
rect 38393 17017 38427 17051
rect 53297 17017 53331 17051
rect 1685 16949 1719 16983
rect 17785 16949 17819 16983
rect 21465 16949 21499 16983
rect 22293 16949 22327 16983
rect 24133 16949 24167 16983
rect 25237 16949 25271 16983
rect 31585 16949 31619 16983
rect 32321 16949 32355 16983
rect 41061 16949 41095 16983
rect 42717 16949 42751 16983
rect 43177 16949 43211 16983
rect 43821 16949 43855 16983
rect 44373 16949 44407 16983
rect 15669 16745 15703 16779
rect 22385 16745 22419 16779
rect 23029 16745 23063 16779
rect 23213 16745 23247 16779
rect 24041 16745 24075 16779
rect 24593 16745 24627 16779
rect 31033 16745 31067 16779
rect 33149 16745 33183 16779
rect 34161 16745 34195 16779
rect 35265 16745 35299 16779
rect 37657 16745 37691 16779
rect 38209 16745 38243 16779
rect 39405 16745 39439 16779
rect 44281 16745 44315 16779
rect 54217 16745 54251 16779
rect 26433 16677 26467 16711
rect 26893 16677 26927 16711
rect 27445 16677 27479 16711
rect 36185 16677 36219 16711
rect 41889 16677 41923 16711
rect 43085 16677 43119 16711
rect 53573 16677 53607 16711
rect 16129 16609 16163 16643
rect 16773 16609 16807 16643
rect 17877 16609 17911 16643
rect 21281 16609 21315 16643
rect 23673 16609 23707 16643
rect 25053 16609 25087 16643
rect 25145 16609 25179 16643
rect 28365 16609 28399 16643
rect 28457 16609 28491 16643
rect 30389 16609 30423 16643
rect 32505 16609 32539 16643
rect 34897 16609 34931 16643
rect 36829 16609 36863 16643
rect 41429 16609 41463 16643
rect 43637 16609 43671 16643
rect 1869 16541 1903 16575
rect 17233 16541 17267 16575
rect 18061 16541 18095 16575
rect 18245 16541 18279 16575
rect 18705 16541 18739 16575
rect 22201 16541 22235 16575
rect 22385 16541 22419 16575
rect 23857 16541 23891 16575
rect 24961 16541 24995 16575
rect 25789 16541 25823 16575
rect 27169 16541 27203 16575
rect 28549 16541 28583 16575
rect 28641 16541 28675 16575
rect 29745 16541 29779 16575
rect 33977 16541 34011 16575
rect 35081 16541 35115 16575
rect 36369 16541 36403 16575
rect 37289 16541 37323 16575
rect 37473 16541 37507 16575
rect 38853 16541 38887 16575
rect 39221 16541 39255 16575
rect 41173 16541 41207 16575
rect 42073 16541 42107 16575
rect 42533 16541 42567 16575
rect 54033 16541 54067 16575
rect 15117 16473 15151 16507
rect 21036 16473 21070 16507
rect 22845 16473 22879 16507
rect 23061 16473 23095 16507
rect 27261 16473 27295 16507
rect 33425 16473 33459 16507
rect 36461 16473 36495 16507
rect 36553 16473 36587 16507
rect 36691 16473 36725 16507
rect 38301 16473 38335 16507
rect 39037 16473 39071 16507
rect 39129 16473 39163 16507
rect 1685 16405 1719 16439
rect 17417 16405 17451 16439
rect 18889 16405 18923 16439
rect 19901 16405 19935 16439
rect 27077 16405 27111 16439
rect 28181 16405 28215 16439
rect 29929 16405 29963 16439
rect 31861 16405 31895 16439
rect 40049 16405 40083 16439
rect 14565 16201 14599 16235
rect 16865 16201 16899 16235
rect 20545 16201 20579 16235
rect 21005 16201 21039 16235
rect 22569 16201 22603 16235
rect 25605 16201 25639 16235
rect 28181 16201 28215 16235
rect 30297 16201 30331 16235
rect 33333 16201 33367 16235
rect 41981 16201 42015 16235
rect 44833 16201 44867 16235
rect 54217 16201 54251 16235
rect 15117 16133 15151 16167
rect 18245 16133 18279 16167
rect 23489 16133 23523 16167
rect 25145 16133 25179 16167
rect 34253 16133 34287 16167
rect 35173 16133 35207 16167
rect 39037 16133 39071 16167
rect 1869 16065 1903 16099
rect 16129 16065 16163 16099
rect 17325 16065 17359 16099
rect 20913 16065 20947 16099
rect 22753 16065 22787 16099
rect 27169 16065 27203 16099
rect 27353 16065 27387 16099
rect 27445 16065 27479 16099
rect 27537 16065 27571 16099
rect 28641 16065 28675 16099
rect 29101 16065 29135 16099
rect 29285 16065 29319 16099
rect 29929 16065 29963 16099
rect 31125 16065 31159 16099
rect 31217 16065 31251 16099
rect 32321 16065 32355 16099
rect 32505 16065 32539 16099
rect 32965 16065 32999 16099
rect 33149 16065 33183 16099
rect 36921 16065 36955 16099
rect 37657 16065 37691 16099
rect 38485 16065 38519 16099
rect 41245 16065 41279 16099
rect 54033 16065 54067 16099
rect 17049 15997 17083 16031
rect 17141 15997 17175 16031
rect 17233 15997 17267 16031
rect 19993 15997 20027 16031
rect 21189 15997 21223 16031
rect 22937 15997 22971 16031
rect 26249 15997 26283 16031
rect 29193 15997 29227 16031
rect 29837 15997 29871 16031
rect 31401 15997 31435 16031
rect 32413 15997 32447 16031
rect 40785 15997 40819 16031
rect 27721 15929 27755 15963
rect 28273 15929 28307 15963
rect 43729 15929 43763 15963
rect 1685 15861 1719 15895
rect 15577 15861 15611 15895
rect 16313 15861 16347 15895
rect 22109 15861 22143 15895
rect 33977 15861 34011 15895
rect 37473 15861 37507 15895
rect 38209 15861 38243 15895
rect 41429 15861 41463 15895
rect 42625 15861 42659 15895
rect 43177 15861 43211 15895
rect 44373 15861 44407 15895
rect 16773 15657 16807 15691
rect 21649 15657 21683 15691
rect 25973 15657 26007 15691
rect 29745 15657 29779 15691
rect 33885 15657 33919 15691
rect 36001 15657 36035 15691
rect 37933 15657 37967 15691
rect 40049 15657 40083 15691
rect 43821 15657 43855 15691
rect 20821 15589 20855 15623
rect 28549 15589 28583 15623
rect 53297 15589 53331 15623
rect 13737 15521 13771 15555
rect 17049 15521 17083 15555
rect 18797 15521 18831 15555
rect 22293 15521 22327 15555
rect 29101 15521 29135 15555
rect 32781 15521 32815 15555
rect 35265 15521 35299 15555
rect 41429 15521 41463 15555
rect 54033 15521 54067 15555
rect 1869 15453 1903 15487
rect 16129 15453 16163 15487
rect 16957 15453 16991 15487
rect 17141 15453 17175 15487
rect 17233 15453 17267 15487
rect 19441 15453 19475 15487
rect 19697 15453 19731 15487
rect 21833 15453 21867 15487
rect 24593 15453 24627 15487
rect 26525 15453 26559 15487
rect 28089 15453 28123 15487
rect 28365 15453 28399 15487
rect 29009 15453 29043 15487
rect 29929 15453 29963 15487
rect 30021 15453 30055 15487
rect 30757 15453 30791 15487
rect 33241 15453 33275 15487
rect 35081 15453 35115 15487
rect 35173 15453 35207 15487
rect 35357 15453 35391 15487
rect 36461 15453 36495 15487
rect 38945 15453 38979 15487
rect 39129 15453 39163 15487
rect 39221 15453 39255 15487
rect 39313 15453 39347 15487
rect 41889 15453 41923 15487
rect 42073 15453 42107 15487
rect 42533 15453 42567 15487
rect 42717 15453 42751 15487
rect 43361 15453 43395 15487
rect 54217 15453 54251 15487
rect 14565 15385 14599 15419
rect 15669 15385 15703 15419
rect 22538 15385 22572 15419
rect 24838 15385 24872 15419
rect 27077 15385 27111 15419
rect 30941 15385 30975 15419
rect 32536 15385 32570 15419
rect 41184 15385 41218 15419
rect 45201 15385 45235 15419
rect 52837 15385 52871 15419
rect 53481 15385 53515 15419
rect 1685 15317 1719 15351
rect 15025 15317 15059 15351
rect 16313 15317 16347 15351
rect 18153 15317 18187 15351
rect 18521 15317 18555 15351
rect 18613 15317 18647 15351
rect 23673 15317 23707 15351
rect 27537 15317 27571 15351
rect 28181 15317 28215 15351
rect 30573 15317 30607 15351
rect 31401 15317 31435 15351
rect 34897 15317 34931 15351
rect 39497 15317 39531 15351
rect 41981 15317 42015 15351
rect 42625 15317 42659 15351
rect 43177 15317 43211 15351
rect 44465 15317 44499 15351
rect 13737 15113 13771 15147
rect 19533 15113 19567 15147
rect 20821 15113 20855 15147
rect 23305 15113 23339 15147
rect 27169 15113 27203 15147
rect 29101 15113 29135 15147
rect 41321 15113 41355 15147
rect 43177 15113 43211 15147
rect 53573 15113 53607 15147
rect 54217 15113 54251 15147
rect 14289 15045 14323 15079
rect 15945 15045 15979 15079
rect 18245 15045 18279 15079
rect 23765 15045 23799 15079
rect 29561 15045 29595 15079
rect 36737 15045 36771 15079
rect 39681 15045 39715 15079
rect 41521 15045 41555 15079
rect 1869 14977 1903 15011
rect 14749 14977 14783 15011
rect 17141 14977 17175 15011
rect 22661 14977 22695 15011
rect 23673 14977 23707 15011
rect 24777 14977 24811 15011
rect 27537 14977 27571 15011
rect 28181 14977 28215 15011
rect 28365 14977 28399 15011
rect 28457 14977 28491 15011
rect 28554 14977 28588 15011
rect 30573 14977 30607 15011
rect 33445 14977 33479 15011
rect 34161 14977 34195 15011
rect 35633 14977 35667 15011
rect 36921 14977 36955 15011
rect 38597 14977 38631 15011
rect 38853 14977 38887 15011
rect 39497 14977 39531 15011
rect 39589 14977 39623 15011
rect 39865 14977 39899 15011
rect 40509 14977 40543 15011
rect 40693 14977 40727 15011
rect 54033 14977 54067 15011
rect 16865 14909 16899 14943
rect 17049 14909 17083 14943
rect 17233 14909 17267 14943
rect 17325 14909 17359 14943
rect 20913 14909 20947 14943
rect 21097 14909 21131 14943
rect 22845 14909 22879 14943
rect 23857 14909 23891 14943
rect 25329 14909 25363 14943
rect 25789 14909 25823 14943
rect 26341 14909 26375 14943
rect 27345 14909 27379 14943
rect 27445 14909 27479 14943
rect 27629 14909 27663 14943
rect 31677 14909 31711 14943
rect 33701 14909 33735 14943
rect 34713 14909 34747 14943
rect 35541 14909 35575 14943
rect 40325 14909 40359 14943
rect 20453 14841 20487 14875
rect 29193 14841 29227 14875
rect 30297 14841 30331 14875
rect 31033 14841 31067 14875
rect 37473 14841 37507 14875
rect 1685 14773 1719 14807
rect 13185 14773 13219 14807
rect 15393 14773 15427 14807
rect 16037 14773 16071 14807
rect 22477 14773 22511 14807
rect 28181 14773 28215 14807
rect 30113 14773 30147 14807
rect 32321 14773 32355 14807
rect 35357 14773 35391 14807
rect 36553 14773 36587 14807
rect 39313 14773 39347 14807
rect 41153 14773 41187 14807
rect 41337 14773 41371 14807
rect 41981 14773 42015 14807
rect 42625 14773 42659 14807
rect 43729 14773 43763 14807
rect 44281 14773 44315 14807
rect 44925 14773 44959 14807
rect 15117 14569 15151 14603
rect 15577 14569 15611 14603
rect 16589 14569 16623 14603
rect 17693 14569 17727 14603
rect 23949 14569 23983 14603
rect 25237 14569 25271 14603
rect 31677 14569 31711 14603
rect 33149 14569 33183 14603
rect 37013 14569 37047 14603
rect 37565 14569 37599 14603
rect 43085 14569 43119 14603
rect 13737 14501 13771 14535
rect 28089 14501 28123 14535
rect 54217 14501 54251 14535
rect 14565 14433 14599 14467
rect 15853 14433 15887 14467
rect 15945 14433 15979 14467
rect 16773 14433 16807 14467
rect 18797 14433 18831 14467
rect 21833 14433 21867 14467
rect 22569 14433 22603 14467
rect 26617 14433 26651 14467
rect 29837 14433 29871 14467
rect 31953 14433 31987 14467
rect 32045 14433 32079 14467
rect 32965 14433 32999 14467
rect 33793 14433 33827 14467
rect 1869 14365 1903 14399
rect 15761 14365 15795 14399
rect 16037 14365 16071 14399
rect 16865 14365 16899 14399
rect 16957 14365 16991 14399
rect 17049 14365 17083 14399
rect 19441 14365 19475 14399
rect 21649 14365 21683 14399
rect 24593 14365 24627 14399
rect 24777 14365 24811 14399
rect 27537 14365 27571 14399
rect 27721 14365 27755 14399
rect 27905 14365 27939 14399
rect 28917 14365 28951 14399
rect 31861 14365 31895 14399
rect 32137 14365 32171 14399
rect 32873 14365 32907 14399
rect 36277 14365 36311 14399
rect 36921 14365 36955 14399
rect 37440 14365 37474 14399
rect 38209 14365 38243 14399
rect 38301 14365 38335 14399
rect 39129 14365 39163 14399
rect 39333 14365 39367 14399
rect 41429 14365 41463 14399
rect 43545 14365 43579 14399
rect 54033 14365 54067 14399
rect 18613 14297 18647 14331
rect 19686 14297 19720 14331
rect 22814 14297 22848 14331
rect 24685 14297 24719 14331
rect 26350 14297 26384 14331
rect 27813 14297 27847 14331
rect 30082 14297 30116 14331
rect 36010 14297 36044 14331
rect 39497 14297 39531 14331
rect 41162 14297 41196 14331
rect 41889 14297 41923 14331
rect 42441 14297 42475 14331
rect 1685 14229 1719 14263
rect 12633 14229 12667 14263
rect 13185 14229 13219 14263
rect 18153 14229 18187 14263
rect 18521 14229 18555 14263
rect 20821 14229 20855 14263
rect 21281 14229 21315 14263
rect 21741 14229 21775 14263
rect 29101 14229 29135 14263
rect 31217 14229 31251 14263
rect 34345 14229 34379 14263
rect 34897 14229 34931 14263
rect 37381 14229 37415 14263
rect 38301 14229 38335 14263
rect 40049 14229 40083 14263
rect 44189 14229 44223 14263
rect 53573 14229 53607 14263
rect 13921 14025 13955 14059
rect 18337 14025 18371 14059
rect 20269 14025 20303 14059
rect 23397 14025 23431 14059
rect 23765 14025 23799 14059
rect 23857 14025 23891 14059
rect 29377 14025 29411 14059
rect 31309 14025 31343 14059
rect 31401 14025 31435 14059
rect 35541 14025 35575 14059
rect 43269 14025 43303 14059
rect 43821 14025 43855 14059
rect 13369 13957 13403 13991
rect 15117 13957 15151 13991
rect 22477 13957 22511 13991
rect 22845 13957 22879 13991
rect 32321 13957 32355 13991
rect 38597 13957 38631 13991
rect 54217 13957 54251 13991
rect 1869 13889 1903 13923
rect 12265 13889 12299 13923
rect 14933 13889 14967 13923
rect 16129 13889 16163 13923
rect 17224 13889 17258 13923
rect 19450 13889 19484 13923
rect 21097 13889 21131 13923
rect 21189 13889 21223 13923
rect 24593 13889 24627 13923
rect 24777 13889 24811 13923
rect 25237 13889 25271 13923
rect 25504 13889 25538 13923
rect 28282 13889 28316 13923
rect 28549 13889 28583 13923
rect 29561 13889 29595 13923
rect 30021 13889 30055 13923
rect 31217 13889 31251 13923
rect 31585 13889 31619 13923
rect 33517 13889 33551 13923
rect 34161 13889 34195 13923
rect 34428 13889 34462 13923
rect 38853 13889 38887 13923
rect 39405 13889 39439 13923
rect 40141 13889 40175 13923
rect 41061 13889 41095 13923
rect 53481 13889 53515 13923
rect 14473 13821 14507 13855
rect 15945 13821 15979 13855
rect 16037 13821 16071 13855
rect 16221 13821 16255 13855
rect 17049 13821 17083 13855
rect 17141 13821 17175 13855
rect 17325 13821 17359 13855
rect 19717 13821 19751 13855
rect 21281 13821 21315 13855
rect 23949 13821 23983 13855
rect 29745 13821 29779 13855
rect 31033 13821 31067 13855
rect 32965 13821 32999 13855
rect 33701 13821 33735 13855
rect 36553 13821 36587 13855
rect 42625 13821 42659 13855
rect 54033 13821 54067 13855
rect 24777 13753 24811 13787
rect 26617 13753 26651 13787
rect 30481 13753 30515 13787
rect 53297 13753 53331 13787
rect 1685 13685 1719 13719
rect 12817 13685 12851 13719
rect 15301 13685 15335 13719
rect 15761 13685 15795 13719
rect 16865 13685 16899 13719
rect 20729 13685 20763 13719
rect 27169 13685 27203 13719
rect 29929 13685 29963 13719
rect 36001 13685 36035 13719
rect 37473 13685 37507 13719
rect 39497 13685 39531 13719
rect 40141 13685 40175 13719
rect 40877 13685 40911 13719
rect 41521 13685 41555 13719
rect 14841 13481 14875 13515
rect 16037 13481 16071 13515
rect 22293 13481 22327 13515
rect 23397 13481 23431 13515
rect 24593 13481 24627 13515
rect 26065 13481 26099 13515
rect 26893 13481 26927 13515
rect 29101 13481 29135 13515
rect 30297 13481 30331 13515
rect 32321 13481 32355 13515
rect 32965 13481 32999 13515
rect 37197 13481 37231 13515
rect 38393 13481 38427 13515
rect 40785 13481 40819 13515
rect 41521 13481 41555 13515
rect 41981 13481 42015 13515
rect 42533 13481 42567 13515
rect 54217 13481 54251 13515
rect 20361 13413 20395 13447
rect 27445 13413 27479 13447
rect 53573 13413 53607 13447
rect 13645 13345 13679 13379
rect 16313 13345 16347 13379
rect 18889 13345 18923 13379
rect 23949 13345 23983 13379
rect 24961 13345 24995 13379
rect 26801 13345 26835 13379
rect 29929 13345 29963 13379
rect 31677 13345 31711 13379
rect 33517 13345 33551 13379
rect 36277 13345 36311 13379
rect 1869 13277 1903 13311
rect 14657 13277 14691 13311
rect 15301 13277 15335 13311
rect 16221 13277 16255 13311
rect 16405 13277 16439 13311
rect 16497 13277 16531 13311
rect 19441 13277 19475 13311
rect 20085 13277 20119 13311
rect 20821 13277 20855 13311
rect 24777 13277 24811 13311
rect 25421 13277 25455 13311
rect 27320 13277 27354 13311
rect 27997 13277 28031 13311
rect 29193 13277 29227 13311
rect 30113 13277 30147 13311
rect 30757 13277 30791 13311
rect 30849 13277 30883 13311
rect 31033 13277 31067 13311
rect 37105 13277 37139 13311
rect 37568 13277 37602 13311
rect 38209 13277 38243 13311
rect 39221 13277 39255 13311
rect 39405 13277 39439 13311
rect 40049 13277 40083 13311
rect 40969 13277 41003 13311
rect 54033 13277 54067 13311
rect 18622 13209 18656 13243
rect 20361 13209 20395 13243
rect 34253 13209 34287 13243
rect 36010 13209 36044 13243
rect 1685 13141 1719 13175
rect 12633 13141 12667 13175
rect 13185 13141 13219 13175
rect 15485 13141 15519 13175
rect 17509 13141 17543 13175
rect 19625 13141 19659 13175
rect 20177 13141 20211 13175
rect 27261 13141 27295 13175
rect 28549 13141 28583 13175
rect 31217 13141 31251 13175
rect 34161 13141 34195 13175
rect 34897 13141 34931 13175
rect 37565 13141 37599 13175
rect 37749 13141 37783 13175
rect 39037 13141 39071 13175
rect 40233 13141 40267 13175
rect 12449 12937 12483 12971
rect 14473 12937 14507 12971
rect 17049 12937 17083 12971
rect 17693 12937 17727 12971
rect 18245 12937 18279 12971
rect 24961 12937 24995 12971
rect 27997 12937 28031 12971
rect 30757 12937 30791 12971
rect 36001 12937 36035 12971
rect 40233 12937 40267 12971
rect 41889 12937 41923 12971
rect 54217 12937 54251 12971
rect 11897 12869 11931 12903
rect 15117 12869 15151 12903
rect 15301 12869 15335 12903
rect 23029 12869 23063 12903
rect 26157 12869 26191 12903
rect 29929 12869 29963 12903
rect 34094 12869 34128 12903
rect 34713 12869 34747 12903
rect 37641 12869 37675 12903
rect 37841 12869 37875 12903
rect 1869 12801 1903 12835
rect 13001 12801 13035 12835
rect 13461 12801 13495 12835
rect 13553 12801 13587 12835
rect 13737 12801 13771 12835
rect 14933 12801 14967 12835
rect 16129 12801 16163 12835
rect 16865 12801 16899 12835
rect 17509 12801 17543 12835
rect 19369 12801 19403 12835
rect 20085 12801 20119 12835
rect 20352 12801 20386 12835
rect 22385 12801 22419 12835
rect 24041 12801 24075 12835
rect 25053 12801 25087 12835
rect 28825 12801 28859 12835
rect 29653 12801 29687 12835
rect 29746 12801 29780 12835
rect 30021 12801 30055 12835
rect 30159 12801 30193 12835
rect 30941 12801 30975 12835
rect 31033 12801 31067 12835
rect 31217 12801 31251 12835
rect 32597 12801 32631 12835
rect 32689 12801 32723 12835
rect 33609 12801 33643 12835
rect 35357 12801 35391 12835
rect 36369 12801 36403 12835
rect 38557 12801 38591 12835
rect 40141 12801 40175 12835
rect 40325 12801 40359 12835
rect 54033 12801 54067 12835
rect 15761 12733 15795 12767
rect 15945 12733 15979 12767
rect 16037 12733 16071 12767
rect 16221 12733 16255 12767
rect 19625 12733 19659 12767
rect 23489 12733 23523 12767
rect 25145 12733 25179 12767
rect 26249 12733 26283 12767
rect 26341 12733 26375 12767
rect 27445 12733 27479 12767
rect 28733 12733 28767 12767
rect 31125 12733 31159 12767
rect 32505 12733 32539 12767
rect 32781 12733 32815 12767
rect 33885 12733 33919 12767
rect 33977 12733 34011 12767
rect 36277 12733 36311 12767
rect 38301 12733 38335 12767
rect 21465 12665 21499 12699
rect 28457 12665 28491 12699
rect 39681 12665 39715 12699
rect 1685 12597 1719 12631
rect 13921 12597 13955 12631
rect 22109 12597 22143 12631
rect 24593 12597 24627 12631
rect 25789 12597 25823 12631
rect 30297 12597 30331 12631
rect 32321 12597 32355 12631
rect 34253 12597 34287 12631
rect 37473 12597 37507 12631
rect 37657 12597 37691 12631
rect 40785 12597 40819 12631
rect 41429 12597 41463 12631
rect 12081 12393 12115 12427
rect 15853 12393 15887 12427
rect 17325 12393 17359 12427
rect 25973 12393 26007 12427
rect 31125 12393 31159 12427
rect 36185 12393 36219 12427
rect 37657 12393 37691 12427
rect 38301 12393 38335 12427
rect 40049 12393 40083 12427
rect 13185 12325 13219 12359
rect 13737 12325 13771 12359
rect 17141 12325 17175 12359
rect 22753 12325 22787 12359
rect 29193 12325 29227 12359
rect 34989 12325 35023 12359
rect 38669 12325 38703 12359
rect 40601 12325 40635 12359
rect 41153 12325 41187 12359
rect 16129 12257 16163 12291
rect 18797 12257 18831 12291
rect 21189 12257 21223 12291
rect 23765 12257 23799 12291
rect 24041 12257 24075 12291
rect 24593 12257 24627 12291
rect 27261 12257 27295 12291
rect 29745 12257 29779 12291
rect 32137 12257 32171 12291
rect 37749 12257 37783 12291
rect 38761 12257 38795 12291
rect 1869 12189 1903 12223
rect 14381 12189 14415 12223
rect 16037 12189 16071 12223
rect 16221 12189 16255 12223
rect 16313 12189 16347 12223
rect 16865 12189 16899 12223
rect 18613 12189 18647 12223
rect 19901 12189 19935 12223
rect 20085 12189 20119 12223
rect 23673 12189 23707 12223
rect 26433 12189 26467 12223
rect 26617 12189 26651 12223
rect 28825 12189 28859 12223
rect 29009 12189 29043 12223
rect 33839 12189 33873 12223
rect 34069 12189 34103 12223
rect 34252 12189 34286 12223
rect 34345 12189 34379 12223
rect 36829 12189 36863 12223
rect 37473 12189 37507 12223
rect 38485 12189 38519 12223
rect 39221 12189 39255 12223
rect 54033 12189 54067 12223
rect 54217 12189 54251 12223
rect 22201 12121 22235 12155
rect 22477 12121 22511 12155
rect 24838 12121 24872 12155
rect 29990 12121 30024 12155
rect 33977 12121 34011 12155
rect 35357 12121 35391 12155
rect 53297 12121 53331 12155
rect 53481 12121 53515 12155
rect 1685 12053 1719 12087
rect 12633 12053 12667 12087
rect 14473 12053 14507 12087
rect 15301 12053 15335 12087
rect 18153 12053 18187 12087
rect 18521 12053 18555 12087
rect 19993 12053 20027 12087
rect 20545 12053 20579 12087
rect 20913 12053 20947 12087
rect 21005 12053 21039 12087
rect 22293 12053 22327 12087
rect 26801 12053 26835 12087
rect 27905 12053 27939 12087
rect 31585 12053 31619 12087
rect 32781 12053 32815 12087
rect 33701 12053 33735 12087
rect 34897 12053 34931 12087
rect 37289 12053 37323 12087
rect 39313 12053 39347 12087
rect 41797 12053 41831 12087
rect 52837 12053 52871 12087
rect 12633 11849 12667 11883
rect 15761 11849 15795 11883
rect 26157 11849 26191 11883
rect 29653 11849 29687 11883
rect 30021 11849 30055 11883
rect 31493 11849 31527 11883
rect 32321 11849 32355 11883
rect 32873 11849 32907 11883
rect 34989 11849 35023 11883
rect 36829 11849 36863 11883
rect 41153 11849 41187 11883
rect 41705 11849 41739 11883
rect 53573 11849 53607 11883
rect 54217 11849 54251 11883
rect 13737 11781 13771 11815
rect 17049 11781 17083 11815
rect 20146 11781 20180 11815
rect 22845 11781 22879 11815
rect 25022 11781 25056 11815
rect 29101 11781 29135 11815
rect 30113 11781 30147 11815
rect 34008 11781 34042 11815
rect 1869 11713 1903 11747
rect 15025 11713 15059 11747
rect 16037 11713 16071 11747
rect 17877 11713 17911 11747
rect 18133 11713 18167 11747
rect 24133 11713 24167 11747
rect 28293 11713 28327 11747
rect 29009 11713 29043 11747
rect 29193 11713 29227 11747
rect 30849 11713 30883 11747
rect 31033 11713 31067 11747
rect 31125 11713 31159 11747
rect 31217 11713 31251 11747
rect 34805 11713 34839 11747
rect 35716 11713 35750 11747
rect 37565 11713 37599 11747
rect 37657 11713 37691 11747
rect 38485 11713 38519 11747
rect 38752 11713 38786 11747
rect 40509 11713 40543 11747
rect 54033 11713 54067 11747
rect 14749 11645 14783 11679
rect 14933 11645 14967 11679
rect 15117 11645 15151 11679
rect 15209 11645 15243 11679
rect 15945 11645 15979 11679
rect 16129 11645 16163 11679
rect 16221 11645 16255 11679
rect 19901 11645 19935 11679
rect 22845 11645 22879 11679
rect 22937 11645 22971 11679
rect 24317 11645 24351 11679
rect 24777 11645 24811 11679
rect 28549 11645 28583 11679
rect 30205 11645 30239 11679
rect 34253 11645 34287 11679
rect 35449 11645 35483 11679
rect 40693 11645 40727 11679
rect 21281 11577 21315 11611
rect 22385 11577 22419 11611
rect 39865 11577 39899 11611
rect 1685 11509 1719 11543
rect 13185 11509 13219 11543
rect 14289 11509 14323 11543
rect 16957 11509 16991 11543
rect 19257 11509 19291 11543
rect 23949 11509 23983 11543
rect 27169 11509 27203 11543
rect 37841 11509 37875 11543
rect 40325 11509 40359 11543
rect 15209 11305 15243 11339
rect 16129 11305 16163 11339
rect 25053 11305 25087 11339
rect 36001 11305 36035 11339
rect 39129 11305 39163 11339
rect 40049 11305 40083 11339
rect 40969 11305 41003 11339
rect 15025 11237 15059 11271
rect 15945 11237 15979 11271
rect 16865 11237 16899 11271
rect 26157 11237 26191 11271
rect 29837 11237 29871 11271
rect 31217 11237 31251 11271
rect 32321 11237 32355 11271
rect 33701 11237 33735 11271
rect 36277 11237 36311 11271
rect 40417 11237 40451 11271
rect 54217 11237 54251 11271
rect 25697 11169 25731 11203
rect 27721 11169 27755 11203
rect 27905 11169 27939 11203
rect 33149 11169 33183 11203
rect 36369 11169 36403 11203
rect 40509 11169 40543 11203
rect 1869 11101 1903 11135
rect 17049 11101 17083 11135
rect 17509 11101 17543 11135
rect 19533 11101 19567 11135
rect 21373 11101 21407 11135
rect 22293 11101 22327 11135
rect 26341 11101 26375 11135
rect 26525 11101 26559 11135
rect 27629 11101 27663 11135
rect 28825 11101 28859 11135
rect 29745 11101 29779 11135
rect 30021 11101 30055 11135
rect 30573 11101 30607 11135
rect 30752 11101 30786 11135
rect 30849 11101 30883 11135
rect 30987 11101 31021 11135
rect 31677 11101 31711 11135
rect 31861 11101 31895 11135
rect 31953 11101 31987 11135
rect 32045 11101 32079 11135
rect 33333 11101 33367 11135
rect 34161 11101 34195 11135
rect 34345 11101 34379 11135
rect 34989 11101 35023 11135
rect 36185 11101 36219 11135
rect 36461 11101 36495 11135
rect 36645 11101 36679 11135
rect 37243 11101 37277 11135
rect 37473 11101 37507 11135
rect 37601 11101 37635 11135
rect 37749 11101 37783 11135
rect 38393 11101 38427 11135
rect 38577 11101 38611 11135
rect 38669 11101 38703 11135
rect 39313 11101 39347 11135
rect 40233 11101 40267 11135
rect 54033 11101 54067 11135
rect 13185 11033 13219 11067
rect 14749 11033 14783 11067
rect 15669 11033 15703 11067
rect 17776 11033 17810 11067
rect 21106 11033 21140 11067
rect 22538 11033 22572 11067
rect 28733 11033 28767 11067
rect 34253 11033 34287 11067
rect 37381 11033 37415 11067
rect 38209 11033 38243 11067
rect 53573 11033 53607 11067
rect 1685 10965 1719 10999
rect 13737 10965 13771 10999
rect 18889 10965 18923 10999
rect 19993 10965 20027 10999
rect 23673 10965 23707 10999
rect 27261 10965 27295 10999
rect 33241 10965 33275 10999
rect 35541 10965 35575 10999
rect 37105 10965 37139 10999
rect 14933 10761 14967 10795
rect 16313 10761 16347 10795
rect 16865 10761 16899 10795
rect 24685 10761 24719 10795
rect 26617 10761 26651 10795
rect 29193 10761 29227 10795
rect 30205 10761 30239 10795
rect 32597 10761 32631 10795
rect 33977 10761 34011 10795
rect 37565 10761 37599 10795
rect 40049 10761 40083 10795
rect 40417 10761 40451 10795
rect 40969 10761 41003 10795
rect 41981 10761 42015 10795
rect 14013 10693 14047 10727
rect 26157 10693 26191 10727
rect 31309 10693 31343 10727
rect 54217 10693 54251 10727
rect 1869 10625 1903 10659
rect 15209 10625 15243 10659
rect 16129 10625 16163 10659
rect 18409 10625 18443 10659
rect 19993 10625 20027 10659
rect 21005 10625 21039 10659
rect 22753 10625 22787 10659
rect 23397 10625 23431 10659
rect 26249 10625 26283 10659
rect 27353 10625 27387 10659
rect 28181 10625 28215 10659
rect 29009 10625 29043 10659
rect 29837 10625 29871 10659
rect 30021 10625 30055 10659
rect 30665 10625 30699 10659
rect 30849 10625 30883 10659
rect 30941 10625 30975 10659
rect 31079 10625 31113 10659
rect 32781 10625 32815 10659
rect 32965 10625 32999 10659
rect 33057 10625 33091 10659
rect 35101 10625 35135 10659
rect 36185 10625 36219 10659
rect 36369 10625 36403 10659
rect 36461 10625 36495 10659
rect 36737 10625 36771 10659
rect 37749 10625 37783 10659
rect 38476 10625 38510 10659
rect 40233 10625 40267 10659
rect 40509 10625 40543 10659
rect 41429 10625 41463 10659
rect 53481 10625 53515 10659
rect 13553 10557 13587 10591
rect 15117 10557 15151 10591
rect 15301 10557 15335 10591
rect 15393 10557 15427 10591
rect 17325 10557 17359 10591
rect 18153 10557 18187 10591
rect 21097 10557 21131 10591
rect 21189 10557 21223 10591
rect 22569 10557 22603 10591
rect 26065 10557 26099 10591
rect 27169 10557 27203 10591
rect 28365 10557 28399 10591
rect 29745 10557 29779 10591
rect 29929 10557 29963 10591
rect 35357 10557 35391 10591
rect 36553 10557 36587 10591
rect 38209 10557 38243 10591
rect 14289 10489 14323 10523
rect 16957 10489 16991 10523
rect 19533 10489 19567 10523
rect 20177 10489 20211 10523
rect 54033 10489 54067 10523
rect 1685 10421 1719 10455
rect 14473 10421 14507 10455
rect 20637 10421 20671 10455
rect 22109 10421 22143 10455
rect 22937 10421 22971 10455
rect 27537 10421 27571 10455
rect 27997 10421 28031 10455
rect 36921 10421 36955 10455
rect 39589 10421 39623 10455
rect 41337 10421 41371 10455
rect 53389 10421 53423 10455
rect 13737 10217 13771 10251
rect 15025 10217 15059 10251
rect 16589 10217 16623 10251
rect 17693 10217 17727 10251
rect 18153 10217 18187 10251
rect 20637 10217 20671 10251
rect 23581 10217 23615 10251
rect 28365 10217 28399 10251
rect 29193 10217 29227 10251
rect 32689 10217 32723 10251
rect 35817 10217 35851 10251
rect 38393 10217 38427 10251
rect 54217 10217 54251 10251
rect 13553 10149 13587 10183
rect 16773 10149 16807 10183
rect 30205 10149 30239 10183
rect 31217 10149 31251 10183
rect 33609 10149 33643 10183
rect 38761 10149 38795 10183
rect 53481 10149 53515 10183
rect 13277 10081 13311 10115
rect 15393 10081 15427 10115
rect 16129 10081 16163 10115
rect 18797 10081 18831 10115
rect 19993 10081 20027 10115
rect 25237 10081 25271 10115
rect 31861 10081 31895 10115
rect 34161 10081 34195 10115
rect 40417 10081 40451 10115
rect 53021 10081 53055 10115
rect 1869 10013 1903 10047
rect 15209 10013 15243 10047
rect 15301 10013 15335 10047
rect 15485 10013 15519 10047
rect 17049 10013 17083 10047
rect 17509 10013 17543 10047
rect 20821 10013 20855 10047
rect 21649 10013 21683 10047
rect 22201 10013 22235 10047
rect 22468 10013 22502 10047
rect 24961 10013 24995 10047
rect 26065 10013 26099 10047
rect 28273 10013 28307 10047
rect 29009 10013 29043 10047
rect 30389 10013 30423 10047
rect 31401 10013 31435 10047
rect 32045 10013 32079 10047
rect 32873 10013 32907 10047
rect 33149 10013 33183 10047
rect 33977 10013 34011 10047
rect 34989 10013 35023 10047
rect 35081 10013 35115 10047
rect 35725 10013 35759 10047
rect 35909 10013 35943 10047
rect 36553 10013 36587 10047
rect 38577 10013 38611 10047
rect 38853 10013 38887 10047
rect 40049 10013 40083 10047
rect 40233 10013 40267 10047
rect 54033 10013 54067 10047
rect 19901 9945 19935 9979
rect 30481 9945 30515 9979
rect 30757 9945 30791 9979
rect 33057 9945 33091 9979
rect 36820 9945 36854 9979
rect 39313 9945 39347 9979
rect 1685 9877 1719 9911
rect 14565 9877 14599 9911
rect 18521 9877 18555 9911
rect 18613 9877 18647 9911
rect 19441 9877 19475 9911
rect 19809 9877 19843 9911
rect 21557 9877 21591 9911
rect 24593 9877 24627 9911
rect 25053 9877 25087 9911
rect 27537 9877 27571 9911
rect 30573 9877 30607 9911
rect 32229 9877 32263 9911
rect 34069 9877 34103 9911
rect 35265 9877 35299 9911
rect 37933 9877 37967 9911
rect 17969 9673 18003 9707
rect 19625 9673 19659 9707
rect 22845 9673 22879 9707
rect 13093 9605 13127 9639
rect 16313 9605 16347 9639
rect 17325 9605 17359 9639
rect 23213 9605 23247 9639
rect 30849 9605 30883 9639
rect 36553 9605 36587 9639
rect 39865 9605 39899 9639
rect 48329 9605 48363 9639
rect 1869 9537 1903 9571
rect 14289 9537 14323 9571
rect 14473 9537 14507 9571
rect 15117 9537 15151 9571
rect 15323 9537 15357 9571
rect 17785 9537 17819 9571
rect 18613 9537 18647 9571
rect 19717 9537 19751 9571
rect 20637 9537 20671 9571
rect 21281 9537 21315 9571
rect 22201 9537 22235 9571
rect 24133 9537 24167 9571
rect 24593 9537 24627 9571
rect 24777 9537 24811 9571
rect 26065 9537 26099 9571
rect 26157 9537 26191 9571
rect 27537 9537 27571 9571
rect 27629 9537 27663 9571
rect 28549 9537 28583 9571
rect 28673 9537 28707 9571
rect 29653 9537 29687 9571
rect 29745 9537 29779 9571
rect 30573 9537 30607 9571
rect 30665 9537 30699 9571
rect 31493 9537 31527 9571
rect 31585 9537 31619 9571
rect 33434 9537 33468 9571
rect 34877 9537 34911 9571
rect 36461 9537 36495 9571
rect 36645 9537 36679 9571
rect 38025 9537 38059 9571
rect 38281 9537 38315 9571
rect 48789 9537 48823 9571
rect 49056 9537 49090 9571
rect 50813 9537 50847 9571
rect 53297 9537 53331 9571
rect 53481 9537 53515 9571
rect 54033 9537 54067 9571
rect 14013 9469 14047 9503
rect 14197 9469 14231 9503
rect 14381 9469 14415 9503
rect 15209 9469 15243 9503
rect 15401 9469 15435 9503
rect 16865 9469 16899 9503
rect 19809 9469 19843 9503
rect 23305 9469 23339 9503
rect 23397 9469 23431 9503
rect 24869 9469 24903 9503
rect 26341 9469 26375 9503
rect 27813 9469 27847 9503
rect 28457 9469 28491 9503
rect 29469 9469 29503 9503
rect 33701 9469 33735 9503
rect 34621 9469 34655 9503
rect 50629 9469 50663 9503
rect 13369 9401 13403 9435
rect 13553 9401 13587 9435
rect 16957 9401 16991 9435
rect 18797 9401 18831 9435
rect 20821 9401 20855 9435
rect 21465 9401 21499 9435
rect 22385 9401 22419 9435
rect 25697 9401 25731 9435
rect 27169 9401 27203 9435
rect 30849 9401 30883 9435
rect 32321 9401 32355 9435
rect 50169 9401 50203 9435
rect 54217 9401 54251 9435
rect 1685 9333 1719 9367
rect 15577 9333 15611 9367
rect 19257 9333 19291 9367
rect 28917 9333 28951 9367
rect 30113 9333 30147 9367
rect 31769 9333 31803 9367
rect 36001 9333 36035 9367
rect 37565 9333 37599 9367
rect 39405 9333 39439 9367
rect 50997 9333 51031 9367
rect 52285 9333 52319 9367
rect 13737 9129 13771 9163
rect 15485 9129 15519 9163
rect 16405 9129 16439 9163
rect 16957 9129 16991 9163
rect 18245 9129 18279 9163
rect 23029 9129 23063 9163
rect 24041 9129 24075 9163
rect 27997 9129 28031 9163
rect 31125 9129 31159 9163
rect 31677 9129 31711 9163
rect 34345 9129 34379 9163
rect 36093 9129 36127 9163
rect 38761 9129 38795 9163
rect 48973 9129 49007 9163
rect 53573 9129 53607 9163
rect 13553 9061 13587 9095
rect 16221 9061 16255 9095
rect 53757 9061 53791 9095
rect 14289 8993 14323 9027
rect 14565 8993 14599 9027
rect 19993 8993 20027 9027
rect 21557 8993 21591 9027
rect 25053 8993 25087 9027
rect 25145 8993 25179 9027
rect 28457 8993 28491 9027
rect 28641 8993 28675 9027
rect 32137 8993 32171 9027
rect 32321 8993 32355 9027
rect 33701 8993 33735 9027
rect 35449 8993 35483 9027
rect 37933 8993 37967 9027
rect 1869 8925 1903 8959
rect 14473 8925 14507 8959
rect 14657 8925 14691 8959
rect 14749 8925 14783 8959
rect 15301 8925 15335 8959
rect 18061 8925 18095 8959
rect 18705 8925 18739 8959
rect 21373 8925 21407 8959
rect 22385 8925 22419 8959
rect 23213 8925 23247 8959
rect 23857 8925 23891 8959
rect 27537 8925 27571 8959
rect 29745 8925 29779 8959
rect 30001 8925 30035 8959
rect 32873 8925 32907 8959
rect 36277 8925 36311 8959
rect 36737 8925 36771 8959
rect 38945 8925 38979 8959
rect 39129 8925 39163 8959
rect 48789 8925 48823 8959
rect 48973 8925 49007 8959
rect 51641 8925 51675 8959
rect 52745 8925 52779 8959
rect 52929 8925 52963 8959
rect 13277 8857 13311 8891
rect 15945 8857 15979 8891
rect 17049 8857 17083 8891
rect 19809 8857 19843 8891
rect 27270 8857 27304 8891
rect 37289 8857 37323 8891
rect 50445 8857 50479 8891
rect 52837 8857 52871 8891
rect 53389 8857 53423 8891
rect 1685 8789 1719 8823
rect 18889 8789 18923 8823
rect 19441 8789 19475 8823
rect 19901 8789 19935 8823
rect 21005 8789 21039 8823
rect 21465 8789 21499 8823
rect 22569 8789 22603 8823
rect 24593 8789 24627 8823
rect 24961 8789 24995 8823
rect 26157 8789 26191 8823
rect 28365 8789 28399 8823
rect 32045 8789 32079 8823
rect 33057 8789 33091 8823
rect 33885 8789 33919 8823
rect 33977 8789 34011 8823
rect 34897 8789 34931 8823
rect 35265 8789 35299 8823
rect 35357 8789 35391 8823
rect 49525 8789 49559 8823
rect 51825 8789 51859 8823
rect 53573 8789 53607 8823
rect 14841 8585 14875 8619
rect 17325 8585 17359 8619
rect 22017 8585 22051 8619
rect 22385 8585 22419 8619
rect 25789 8585 25823 8619
rect 28549 8585 28583 8619
rect 32505 8585 32539 8619
rect 35265 8585 35299 8619
rect 36553 8585 36587 8619
rect 38117 8585 38151 8619
rect 38577 8585 38611 8619
rect 53389 8585 53423 8619
rect 54217 8585 54251 8619
rect 14381 8517 14415 8551
rect 16313 8517 16347 8551
rect 16865 8517 16899 8551
rect 20330 8517 20364 8551
rect 26249 8517 26283 8551
rect 1869 8449 1903 8483
rect 13921 8449 13955 8483
rect 15485 8449 15519 8483
rect 18245 8449 18279 8483
rect 18512 8449 18546 8483
rect 23305 8449 23339 8483
rect 23572 8449 23606 8483
rect 25145 8449 25179 8483
rect 26157 8449 26191 8483
rect 27169 8449 27203 8483
rect 27425 8449 27459 8483
rect 29377 8449 29411 8483
rect 29633 8449 29667 8483
rect 31401 8449 31435 8483
rect 32321 8449 32355 8483
rect 33425 8449 33459 8483
rect 33681 8449 33715 8483
rect 35449 8449 35483 8483
rect 51733 8449 51767 8483
rect 52193 8449 52227 8483
rect 53481 8449 53515 8483
rect 54033 8449 54067 8483
rect 20085 8381 20119 8415
rect 22477 8381 22511 8415
rect 22569 8381 22603 8415
rect 26433 8381 26467 8415
rect 31585 8381 31619 8415
rect 51181 8381 51215 8415
rect 1685 8313 1719 8347
rect 14657 8313 14691 8347
rect 15669 8313 15703 8347
rect 17233 8313 17267 8347
rect 19625 8313 19659 8347
rect 21465 8313 21499 8347
rect 24685 8313 24719 8347
rect 25329 8313 25363 8347
rect 30757 8313 30791 8347
rect 34805 8313 34839 8347
rect 37565 8313 37599 8347
rect 52377 8313 52411 8347
rect 31217 8245 31251 8279
rect 35909 8245 35943 8279
rect 14657 8041 14691 8075
rect 15669 8041 15703 8075
rect 16773 8041 16807 8075
rect 17233 8041 17267 8075
rect 22201 8041 22235 8075
rect 24685 8041 24719 8075
rect 25145 8041 25179 8075
rect 28181 8041 28215 8075
rect 31125 8041 31159 8075
rect 32229 8041 32263 8075
rect 32689 8041 32723 8075
rect 33333 8041 33367 8075
rect 35541 8041 35575 8075
rect 36001 8041 36035 8075
rect 36645 8041 36679 8075
rect 52469 8041 52503 8075
rect 17417 7973 17451 8007
rect 12449 7905 12483 7939
rect 12633 7905 12667 7939
rect 12817 7905 12851 7939
rect 13553 7905 13587 7939
rect 18337 7905 18371 7939
rect 22661 7905 22695 7939
rect 25697 7905 25731 7939
rect 27353 7905 27387 7939
rect 27537 7905 27571 7939
rect 29193 7905 29227 7939
rect 29745 7905 29779 7939
rect 34989 7905 35023 7939
rect 1869 7837 1903 7871
rect 12725 7837 12759 7871
rect 12909 7837 12943 7871
rect 19901 7837 19935 7871
rect 22017 7837 22051 7871
rect 22917 7837 22951 7871
rect 27261 7837 27295 7871
rect 28181 7837 28215 7871
rect 28365 7837 28399 7871
rect 29009 7837 29043 7871
rect 33517 7837 33551 7871
rect 33701 7837 33735 7871
rect 51825 7837 51859 7871
rect 52285 7837 52319 7871
rect 52929 7837 52963 7871
rect 17693 7769 17727 7803
rect 18429 7769 18463 7803
rect 20146 7769 20180 7803
rect 25605 7769 25639 7803
rect 30012 7769 30046 7803
rect 53174 7769 53208 7803
rect 1685 7701 1719 7735
rect 15209 7701 15243 7735
rect 18521 7701 18555 7735
rect 18889 7701 18923 7735
rect 21281 7701 21315 7735
rect 24041 7701 24075 7735
rect 25513 7701 25547 7735
rect 26433 7701 26467 7735
rect 26893 7701 26927 7735
rect 28825 7701 28859 7735
rect 31585 7701 31619 7735
rect 34161 7701 34195 7735
rect 54309 7701 54343 7735
rect 12633 7497 12667 7531
rect 13737 7497 13771 7531
rect 15761 7497 15795 7531
rect 17233 7497 17267 7531
rect 22385 7497 22419 7531
rect 27353 7497 27387 7531
rect 29193 7497 29227 7531
rect 30389 7497 30423 7531
rect 31033 7497 31067 7531
rect 33425 7497 33459 7531
rect 33977 7497 34011 7531
rect 34529 7497 34563 7531
rect 35081 7497 35115 7531
rect 52377 7497 52411 7531
rect 53205 7497 53239 7531
rect 17693 7429 17727 7463
rect 28641 7429 28675 7463
rect 32321 7429 32355 7463
rect 53849 7429 53883 7463
rect 1869 7361 1903 7395
rect 13093 7361 13127 7395
rect 16313 7361 16347 7395
rect 18245 7361 18279 7395
rect 18501 7361 18535 7395
rect 21209 7361 21243 7395
rect 24797 7361 24831 7395
rect 25053 7361 25087 7395
rect 26249 7361 26283 7395
rect 26433 7361 26467 7395
rect 27169 7361 27203 7395
rect 27905 7361 27939 7395
rect 28549 7361 28583 7395
rect 29561 7361 29595 7395
rect 29653 7361 29687 7395
rect 30573 7361 30607 7395
rect 53389 7361 53423 7395
rect 54217 7361 54251 7395
rect 12817 7293 12851 7327
rect 12909 7293 12943 7327
rect 13001 7293 13035 7327
rect 21465 7293 21499 7327
rect 22477 7293 22511 7327
rect 22569 7293 22603 7327
rect 26065 7293 26099 7327
rect 29745 7293 29779 7327
rect 32873 7293 32907 7327
rect 17417 7225 17451 7259
rect 20085 7225 20119 7259
rect 25605 7225 25639 7259
rect 28089 7225 28123 7259
rect 1685 7157 1719 7191
rect 19625 7157 19659 7191
rect 22017 7157 22051 7191
rect 23673 7157 23707 7191
rect 31585 7157 31619 7191
rect 18245 6953 18279 6987
rect 21465 6953 21499 6987
rect 25789 6953 25823 6987
rect 33885 6953 33919 6987
rect 53481 6953 53515 6987
rect 54125 6953 54159 6987
rect 17233 6885 17267 6919
rect 13093 6817 13127 6851
rect 13369 6817 13403 6851
rect 17509 6817 17543 6851
rect 20821 6817 20855 6851
rect 24777 6817 24811 6851
rect 26525 6817 26559 6851
rect 27721 6817 27755 6851
rect 29745 6817 29779 6851
rect 30849 6817 30883 6851
rect 31953 6817 31987 6851
rect 33057 6817 33091 6851
rect 1869 6749 1903 6783
rect 13277 6749 13311 6783
rect 13461 6749 13495 6783
rect 13553 6749 13587 6783
rect 14565 6749 14599 6783
rect 15209 6749 15243 6783
rect 18705 6749 18739 6783
rect 21649 6749 21683 6783
rect 24041 6749 24075 6783
rect 24961 6749 24995 6783
rect 25973 6749 26007 6783
rect 30389 6749 30423 6783
rect 54309 6749 54343 6783
rect 14381 6681 14415 6715
rect 20554 6681 20588 6715
rect 23774 6681 23808 6715
rect 26985 6681 27019 6715
rect 29101 6681 29135 6715
rect 31401 6681 31435 6715
rect 32505 6681 32539 6715
rect 1685 6613 1719 6647
rect 17049 6613 17083 6647
rect 18889 6613 18923 6647
rect 19441 6613 19475 6647
rect 22201 6613 22235 6647
rect 22661 6613 22695 6647
rect 24869 6613 24903 6647
rect 25329 6613 25363 6647
rect 28641 6613 28675 6647
rect 12541 6409 12575 6443
rect 13001 6409 13035 6443
rect 14105 6409 14139 6443
rect 14565 6409 14599 6443
rect 17325 6409 17359 6443
rect 17785 6409 17819 6443
rect 18705 6409 18739 6443
rect 19533 6409 19567 6443
rect 20177 6409 20211 6443
rect 20729 6409 20763 6443
rect 21465 6409 21499 6443
rect 22477 6409 22511 6443
rect 23673 6409 23707 6443
rect 24961 6409 24995 6443
rect 25789 6409 25823 6443
rect 26617 6409 26651 6443
rect 27629 6409 27663 6443
rect 28641 6409 28675 6443
rect 29929 6409 29963 6443
rect 31493 6409 31527 6443
rect 32413 6409 32447 6443
rect 54309 6409 54343 6443
rect 28089 6341 28123 6375
rect 31033 6341 31067 6375
rect 1869 6273 1903 6307
rect 13185 6273 13219 6307
rect 13277 6273 13311 6307
rect 18889 6273 18923 6307
rect 19349 6273 19383 6307
rect 23489 6273 23523 6307
rect 30481 6273 30515 6307
rect 12081 6205 12115 6239
rect 13369 6205 13403 6239
rect 13461 6205 13495 6239
rect 25053 6205 25087 6239
rect 25145 6205 25179 6239
rect 29377 6205 29411 6239
rect 12357 6137 12391 6171
rect 24593 6137 24627 6171
rect 1685 6069 1719 6103
rect 23029 6069 23063 6103
rect 12633 5865 12667 5899
rect 13093 5865 13127 5899
rect 22937 5865 22971 5899
rect 24041 5865 24075 5899
rect 24685 5865 24719 5899
rect 25237 5865 25271 5899
rect 27905 5865 27939 5899
rect 28549 5865 28583 5899
rect 30757 5865 30791 5899
rect 11529 5797 11563 5831
rect 12541 5797 12575 5831
rect 26249 5797 26283 5831
rect 11713 5729 11747 5763
rect 13461 5729 13495 5763
rect 26985 5729 27019 5763
rect 1869 5661 1903 5695
rect 13277 5661 13311 5695
rect 13369 5661 13403 5695
rect 13553 5661 13587 5695
rect 23397 5661 23431 5695
rect 25789 5661 25823 5695
rect 30297 5661 30331 5695
rect 11253 5593 11287 5627
rect 12173 5593 12207 5627
rect 30021 5593 30055 5627
rect 1685 5525 1719 5559
rect 10701 5525 10735 5559
rect 14381 5525 14415 5559
rect 29009 5525 29043 5559
rect 12449 5321 12483 5355
rect 24501 5321 24535 5355
rect 25605 5321 25639 5355
rect 26065 5321 26099 5355
rect 27721 5321 27755 5355
rect 28549 5321 28583 5355
rect 30021 5321 30055 5355
rect 30573 5321 30607 5355
rect 14473 5253 14507 5287
rect 1869 5185 1903 5219
rect 12629 5185 12663 5219
rect 12910 5185 12944 5219
rect 14933 5185 14967 5219
rect 27261 5185 27295 5219
rect 29285 5185 29319 5219
rect 12726 5117 12760 5151
rect 12817 5117 12851 5151
rect 13461 5117 13495 5151
rect 10609 5049 10643 5083
rect 13737 5049 13771 5083
rect 13921 5049 13955 5083
rect 1685 4981 1719 5015
rect 9321 4981 9355 5015
rect 9873 4981 9907 5015
rect 11161 4981 11195 5015
rect 11713 4981 11747 5015
rect 24961 4981 24995 5015
rect 10517 4777 10551 4811
rect 12541 4777 12575 4811
rect 13001 4777 13035 4811
rect 25145 4777 25179 4811
rect 26249 4777 26283 4811
rect 38393 4777 38427 4811
rect 41429 4777 41463 4811
rect 42441 4777 42475 4811
rect 42993 4777 43027 4811
rect 12357 4709 12391 4743
rect 13093 4709 13127 4743
rect 10793 4641 10827 4675
rect 1869 4573 1903 4607
rect 10701 4573 10735 4607
rect 10885 4573 10919 4607
rect 10977 4573 11011 4607
rect 14565 4573 14599 4607
rect 45569 4573 45603 4607
rect 7389 4505 7423 4539
rect 10057 4505 10091 4539
rect 12081 4505 12115 4539
rect 13461 4505 13495 4539
rect 15301 4505 15335 4539
rect 22753 4505 22787 4539
rect 1685 4437 1719 4471
rect 8033 4437 8067 4471
rect 9505 4437 9539 4471
rect 11621 4437 11655 4471
rect 14749 4437 14783 4471
rect 23305 4437 23339 4471
rect 23765 4437 23799 4471
rect 25605 4437 25639 4471
rect 38945 4437 38979 4471
rect 43637 4437 43671 4471
rect 45753 4437 45787 4471
rect 10057 4233 10091 4267
rect 25421 4233 25455 4267
rect 9137 4165 9171 4199
rect 32781 4165 32815 4199
rect 36737 4165 36771 4199
rect 1869 4097 1903 4131
rect 10793 4097 10827 4131
rect 22661 4097 22695 4131
rect 26065 4097 26099 4131
rect 39865 4097 39899 4131
rect 40969 4097 41003 4131
rect 42717 4097 42751 4131
rect 43913 4097 43947 4131
rect 44557 4097 44591 4131
rect 45201 4097 45235 4131
rect 45845 4097 45879 4131
rect 46489 4097 46523 4131
rect 9597 4029 9631 4063
rect 10517 4029 10551 4063
rect 10701 4029 10735 4063
rect 10885 4029 10919 4063
rect 10977 4029 11011 4063
rect 11989 4029 12023 4063
rect 12449 4029 12483 4063
rect 15209 4029 15243 4063
rect 24317 4029 24351 4063
rect 26525 4029 26559 4063
rect 9873 3961 9907 3995
rect 12265 3961 12299 3995
rect 37473 3961 37507 3995
rect 38025 3961 38059 3995
rect 40417 3961 40451 3995
rect 42901 3961 42935 3995
rect 44741 3961 44775 3995
rect 1685 3893 1719 3927
rect 6837 3893 6871 3927
rect 7481 3893 7515 3927
rect 8033 3893 8067 3927
rect 8493 3893 8527 3927
rect 13461 3893 13495 3927
rect 14105 3893 14139 3927
rect 14657 3893 14691 3927
rect 15669 3893 15703 3927
rect 17785 3893 17819 3927
rect 23213 3893 23247 3927
rect 23765 3893 23799 3927
rect 24869 3893 24903 3927
rect 30941 3893 30975 3927
rect 38853 3893 38887 3927
rect 39313 3893 39347 3927
rect 41797 3893 41831 3927
rect 43361 3893 43395 3927
rect 44097 3893 44131 3927
rect 45385 3893 45419 3927
rect 46029 3893 46063 3927
rect 46673 3893 46707 3927
rect 49065 3893 49099 3927
rect 50169 3893 50203 3927
rect 50997 3893 51031 3927
rect 7113 3689 7147 3723
rect 7941 3689 7975 3723
rect 10425 3689 10459 3723
rect 12449 3689 12483 3723
rect 13553 3689 13587 3723
rect 26801 3689 26835 3723
rect 27445 3689 27479 3723
rect 27997 3689 28031 3723
rect 28641 3689 28675 3723
rect 31309 3689 31343 3723
rect 32781 3689 32815 3723
rect 33333 3689 33367 3723
rect 33885 3689 33919 3723
rect 34897 3689 34931 3723
rect 41429 3689 41463 3723
rect 42993 3689 43027 3723
rect 51181 3689 51215 3723
rect 9781 3621 9815 3655
rect 11621 3621 11655 3655
rect 23167 3621 23201 3655
rect 30573 3621 30607 3655
rect 31861 3621 31895 3655
rect 40877 3621 40911 3655
rect 10609 3553 10643 3587
rect 10793 3553 10827 3587
rect 14473 3553 14507 3587
rect 14657 3553 14691 3587
rect 14749 3553 14783 3587
rect 1869 3485 1903 3519
rect 6929 3485 6963 3519
rect 7757 3485 7791 3519
rect 8401 3485 8435 3519
rect 10690 3485 10724 3519
rect 10886 3485 10920 3519
rect 11437 3485 11471 3519
rect 12633 3485 12667 3519
rect 13737 3485 13771 3519
rect 14841 3485 14875 3519
rect 14933 3485 14967 3519
rect 19809 3485 19843 3519
rect 21649 3485 21683 3519
rect 22477 3485 22511 3519
rect 22937 3485 22971 3519
rect 25237 3485 25271 3519
rect 37289 3485 37323 3519
rect 37933 3485 37967 3519
rect 38945 3485 38979 3519
rect 40049 3485 40083 3519
rect 40693 3485 40727 3519
rect 41889 3485 41923 3519
rect 43085 3485 43119 3519
rect 43637 3485 43671 3519
rect 44281 3485 44315 3519
rect 45201 3485 45235 3519
rect 45937 3485 45971 3519
rect 46949 3485 46983 3519
rect 47409 3485 47443 3519
rect 9505 3417 9539 3451
rect 22109 3417 22143 3451
rect 22293 3417 22327 3451
rect 26249 3417 26283 3451
rect 51273 3417 51307 3451
rect 1685 3349 1719 3383
rect 6469 3349 6503 3383
rect 8585 3349 8619 3383
rect 9965 3349 9999 3383
rect 15945 3349 15979 3383
rect 16405 3349 16439 3383
rect 17509 3349 17543 3383
rect 18245 3349 18279 3383
rect 25053 3349 25087 3383
rect 36001 3349 36035 3383
rect 36645 3349 36679 3383
rect 37473 3349 37507 3383
rect 38117 3349 38151 3383
rect 39129 3349 39163 3383
rect 40233 3349 40267 3383
rect 42073 3349 42107 3383
rect 43821 3349 43855 3383
rect 44465 3349 44499 3383
rect 45385 3349 45419 3383
rect 46121 3349 46155 3383
rect 46765 3349 46799 3383
rect 48329 3349 48363 3383
rect 48881 3349 48915 3383
rect 49433 3349 49467 3383
rect 50353 3349 50387 3383
rect 51825 3349 51859 3383
rect 52469 3349 52503 3383
rect 8493 3145 8527 3179
rect 9781 3145 9815 3179
rect 10701 3145 10735 3179
rect 11989 3145 12023 3179
rect 13277 3145 13311 3179
rect 13921 3145 13955 3179
rect 14841 3145 14875 3179
rect 15577 3145 15611 3179
rect 16313 3145 16347 3179
rect 16957 3145 16991 3179
rect 17601 3145 17635 3179
rect 18337 3145 18371 3179
rect 29009 3145 29043 3179
rect 29653 3145 29687 3179
rect 31585 3145 31619 3179
rect 47869 3145 47903 3179
rect 48605 3145 48639 3179
rect 49341 3145 49375 3179
rect 50077 3145 50111 3179
rect 50813 3145 50847 3179
rect 51549 3145 51583 3179
rect 6009 3077 6043 3111
rect 35081 3077 35115 3111
rect 48697 3077 48731 3111
rect 51641 3077 51675 3111
rect 7021 3009 7055 3043
rect 7665 3009 7699 3043
rect 8309 3009 8343 3043
rect 8953 3009 8987 3043
rect 9597 3009 9631 3043
rect 10241 3009 10275 3043
rect 11805 3009 11839 3043
rect 12449 3009 12483 3043
rect 13093 3009 13127 3043
rect 13737 3009 13771 3043
rect 15393 3009 15427 3043
rect 16129 3009 16163 3043
rect 17141 3009 17175 3043
rect 17785 3009 17819 3043
rect 18521 3009 18555 3043
rect 23673 3009 23707 3043
rect 24409 3009 24443 3043
rect 24869 3009 24903 3043
rect 25605 3009 25639 3043
rect 26341 3009 26375 3043
rect 27813 3009 27847 3043
rect 28549 3009 28583 3043
rect 30389 3009 30423 3043
rect 31125 3009 31159 3043
rect 32597 3009 32631 3043
rect 33333 3009 33367 3043
rect 36369 3009 36403 3043
rect 38117 3009 38151 3043
rect 38577 3009 38611 3043
rect 39313 3009 39347 3043
rect 40325 3009 40359 3043
rect 41061 3009 41095 3043
rect 41797 3009 41831 3043
rect 42625 3009 42659 3043
rect 43637 3009 43671 3043
rect 44097 3009 44131 3043
rect 44833 3009 44867 3043
rect 45569 3009 45603 3043
rect 46305 3009 46339 3043
rect 47225 3009 47259 3043
rect 47961 3009 47995 3043
rect 49433 3009 49467 3043
rect 50261 3009 50295 3043
rect 50997 3009 51031 3043
rect 14381 2941 14415 2975
rect 33793 2941 33827 2975
rect 34437 2941 34471 2975
rect 35725 2941 35759 2975
rect 7205 2873 7239 2907
rect 7849 2873 7883 2907
rect 9137 2873 9171 2907
rect 10517 2873 10551 2907
rect 12633 2873 12667 2907
rect 14657 2873 14691 2907
rect 32413 2873 32447 2907
rect 45017 2873 45051 2907
rect 46489 2873 46523 2907
rect 52193 2873 52227 2907
rect 19073 2805 19107 2839
rect 20085 2805 20119 2839
rect 20545 2805 20579 2839
rect 21465 2805 21499 2839
rect 22293 2805 22327 2839
rect 22753 2805 22787 2839
rect 23489 2805 23523 2839
rect 24225 2805 24259 2839
rect 25053 2805 25087 2839
rect 25789 2805 25823 2839
rect 26525 2805 26559 2839
rect 27629 2805 27663 2839
rect 28365 2805 28399 2839
rect 30205 2805 30239 2839
rect 30941 2805 30975 2839
rect 33149 2805 33183 2839
rect 37933 2805 37967 2839
rect 38761 2805 38795 2839
rect 39497 2805 39531 2839
rect 40141 2805 40175 2839
rect 40877 2805 40911 2839
rect 41613 2805 41647 2839
rect 42809 2805 42843 2839
rect 43453 2805 43487 2839
rect 44281 2805 44315 2839
rect 45753 2805 45787 2839
rect 9873 2601 9907 2635
rect 11161 2601 11195 2635
rect 11805 2601 11839 2635
rect 13093 2601 13127 2635
rect 13737 2601 13771 2635
rect 15669 2601 15703 2635
rect 16313 2601 16347 2635
rect 17417 2601 17451 2635
rect 18061 2601 18095 2635
rect 36829 2601 36863 2635
rect 49433 2601 49467 2635
rect 7205 2533 7239 2567
rect 9229 2533 9263 2567
rect 10517 2533 10551 2567
rect 15025 2533 15059 2567
rect 20177 2533 20211 2567
rect 29837 2533 29871 2567
rect 31309 2533 31343 2567
rect 33149 2533 33183 2567
rect 38393 2533 38427 2567
rect 40969 2533 41003 2567
rect 42717 2533 42751 2567
rect 44281 2533 44315 2567
rect 46121 2533 46155 2567
rect 47961 2533 47995 2567
rect 48513 2533 48547 2567
rect 50353 2533 50387 2567
rect 51089 2533 51123 2567
rect 4905 2465 4939 2499
rect 7941 2465 7975 2499
rect 34897 2465 34931 2499
rect 7021 2397 7055 2431
rect 7665 2397 7699 2431
rect 9689 2397 9723 2431
rect 10333 2397 10367 2431
rect 10977 2397 11011 2431
rect 12265 2397 12299 2431
rect 12909 2397 12943 2431
rect 13553 2397 13587 2431
rect 14841 2397 14875 2431
rect 15485 2397 15519 2431
rect 16129 2397 16163 2431
rect 17601 2397 17635 2431
rect 18245 2397 18279 2431
rect 18889 2397 18923 2431
rect 20821 2397 20855 2431
rect 21465 2397 21499 2431
rect 22569 2397 22603 2431
rect 23305 2397 23339 2431
rect 23765 2397 23799 2431
rect 24869 2397 24903 2431
rect 25605 2397 25639 2431
rect 26341 2397 26375 2431
rect 27445 2397 27479 2431
rect 28181 2397 28215 2431
rect 29193 2397 29227 2431
rect 30021 2397 30055 2431
rect 30757 2397 30791 2431
rect 31493 2397 31527 2431
rect 32597 2397 32631 2431
rect 33333 2397 33367 2431
rect 34069 2397 34103 2431
rect 35541 2397 35575 2431
rect 37473 2397 37507 2431
rect 38209 2397 38243 2431
rect 38945 2397 38979 2431
rect 40049 2397 40083 2431
rect 40785 2397 40819 2431
rect 41521 2397 41555 2431
rect 42901 2397 42935 2431
rect 43361 2397 43395 2431
rect 44097 2397 44131 2431
rect 45201 2397 45235 2431
rect 45937 2397 45971 2431
rect 46673 2397 46707 2431
rect 47777 2397 47811 2431
rect 49249 2397 49283 2431
rect 51273 2397 51307 2431
rect 52929 2397 52963 2431
rect 14381 2329 14415 2363
rect 19441 2329 19475 2363
rect 36185 2329 36219 2363
rect 48697 2329 48731 2363
rect 50537 2329 50571 2363
rect 51825 2329 51859 2363
rect 52009 2329 52043 2363
rect 5457 2261 5491 2295
rect 6009 2261 6043 2295
rect 12449 2261 12483 2295
rect 16957 2261 16991 2295
rect 22385 2261 22419 2295
rect 23121 2261 23155 2295
rect 23949 2261 23983 2295
rect 25053 2261 25087 2295
rect 25789 2261 25823 2295
rect 26525 2261 26559 2295
rect 27629 2261 27663 2295
rect 28365 2261 28399 2295
rect 29009 2261 29043 2295
rect 30573 2261 30607 2295
rect 32413 2261 32447 2295
rect 33885 2261 33919 2295
rect 37657 2261 37691 2295
rect 39129 2261 39163 2295
rect 40233 2261 40267 2295
rect 41705 2261 41739 2295
rect 43545 2261 43579 2295
rect 45385 2261 45419 2295
rect 46857 2261 46891 2295
<< metal1 >>
rect 1104 53338 54832 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 54832 53338
rect 1104 53264 54832 53286
rect 8570 53224 8576 53236
rect 8531 53196 8576 53224
rect 8570 53184 8576 53196
rect 8628 53184 8634 53236
rect 9306 53224 9312 53236
rect 9267 53196 9312 53224
rect 9306 53184 9312 53196
rect 9364 53184 9370 53236
rect 21085 53227 21143 53233
rect 21085 53193 21097 53227
rect 21131 53224 21143 53227
rect 25590 53224 25596 53236
rect 21131 53196 25596 53224
rect 21131 53193 21143 53196
rect 21085 53187 21143 53193
rect 25590 53184 25596 53196
rect 25648 53184 25654 53236
rect 26602 53224 26608 53236
rect 26563 53196 26608 53224
rect 26602 53184 26608 53196
rect 26660 53184 26666 53236
rect 29178 53224 29184 53236
rect 29139 53196 29184 53224
rect 29178 53184 29184 53196
rect 29236 53184 29242 53236
rect 31754 53224 31760 53236
rect 31715 53196 31760 53224
rect 31754 53184 31760 53196
rect 31812 53184 31818 53236
rect 47118 53224 47124 53236
rect 47079 53196 47124 53224
rect 47118 53184 47124 53196
rect 47176 53184 47182 53236
rect 49694 53224 49700 53236
rect 49655 53196 49700 53224
rect 49694 53184 49700 53196
rect 49752 53184 49758 53236
rect 3142 53156 3148 53168
rect 3103 53128 3148 53156
rect 3142 53116 3148 53128
rect 3200 53116 3206 53168
rect 4893 53159 4951 53165
rect 4893 53125 4905 53159
rect 4939 53156 4951 53159
rect 5442 53156 5448 53168
rect 4939 53128 5448 53156
rect 4939 53125 4951 53128
rect 4893 53119 4951 53125
rect 5442 53116 5448 53128
rect 5500 53116 5506 53168
rect 6638 53156 6644 53168
rect 6599 53128 6644 53156
rect 6638 53116 6644 53128
rect 6696 53116 6702 53168
rect 2317 53091 2375 53097
rect 2317 53057 2329 53091
rect 2363 53088 2375 53091
rect 2363 53060 3096 53088
rect 2363 53057 2375 53060
rect 2317 53051 2375 53057
rect 1670 52980 1676 53032
rect 1728 53020 1734 53032
rect 2590 53020 2596 53032
rect 1728 52992 2596 53020
rect 1728 52980 1734 52992
rect 2590 52980 2596 52992
rect 2648 52980 2654 53032
rect 3068 53020 3096 53060
rect 4062 53048 4068 53100
rect 4120 53088 4126 53100
rect 4157 53091 4215 53097
rect 4157 53088 4169 53091
rect 4120 53060 4169 53088
rect 4120 53048 4126 53060
rect 4157 53057 4169 53060
rect 4203 53057 4215 53091
rect 7742 53088 7748 53100
rect 7703 53060 7748 53088
rect 4157 53051 4215 53057
rect 7742 53048 7748 53060
rect 7800 53048 7806 53100
rect 8588 53088 8616 53184
rect 24486 53156 24492 53168
rect 18340 53128 24492 53156
rect 9125 53091 9183 53097
rect 9125 53088 9137 53091
rect 8588 53060 9137 53088
rect 9125 53057 9137 53060
rect 9171 53057 9183 53091
rect 10134 53088 10140 53100
rect 10095 53060 10140 53088
rect 9125 53051 9183 53057
rect 10134 53048 10140 53060
rect 10192 53048 10198 53100
rect 12069 53091 12127 53097
rect 12069 53057 12081 53091
rect 12115 53088 12127 53091
rect 12526 53088 12532 53100
rect 12115 53060 12532 53088
rect 12115 53057 12127 53060
rect 12069 53051 12127 53057
rect 12526 53048 12532 53060
rect 12584 53048 12590 53100
rect 14826 53088 14832 53100
rect 14787 53060 14832 53088
rect 14826 53048 14832 53060
rect 14884 53048 14890 53100
rect 16298 53088 16304 53100
rect 16259 53060 16304 53088
rect 16298 53048 16304 53060
rect 16356 53088 16362 53100
rect 16853 53091 16911 53097
rect 16853 53088 16865 53091
rect 16356 53060 16865 53088
rect 16356 53048 16362 53060
rect 16853 53057 16865 53060
rect 16899 53057 16911 53091
rect 16853 53051 16911 53057
rect 8202 53020 8208 53032
rect 3068 52992 8208 53020
rect 8202 52980 8208 52992
rect 8260 52980 8266 53032
rect 10410 53020 10416 53032
rect 10371 52992 10416 53020
rect 10410 52980 10416 52992
rect 10468 52980 10474 53032
rect 12802 53020 12808 53032
rect 12763 52992 12808 53020
rect 12802 52980 12808 52992
rect 12860 52980 12866 53032
rect 16022 53020 16028 53032
rect 15983 52992 16028 53020
rect 16022 52980 16028 52992
rect 16080 52980 16086 53032
rect 18340 53020 18368 53128
rect 24486 53116 24492 53128
rect 24544 53116 24550 53168
rect 18414 53048 18420 53100
rect 18472 53088 18478 53100
rect 18782 53088 18788 53100
rect 18472 53060 18788 53088
rect 18472 53048 18478 53060
rect 18782 53048 18788 53060
rect 18840 53088 18846 53100
rect 18877 53091 18935 53097
rect 18877 53088 18889 53091
rect 18840 53060 18889 53088
rect 18840 53048 18846 53060
rect 18877 53057 18889 53060
rect 18923 53057 18935 53091
rect 18877 53051 18935 53057
rect 19426 53048 19432 53100
rect 19484 53088 19490 53100
rect 19705 53091 19763 53097
rect 19705 53088 19717 53091
rect 19484 53060 19717 53088
rect 19484 53048 19490 53060
rect 19705 53057 19717 53060
rect 19751 53057 19763 53091
rect 19705 53051 19763 53057
rect 20441 53091 20499 53097
rect 20441 53057 20453 53091
rect 20487 53088 20499 53091
rect 20898 53088 20904 53100
rect 20487 53060 20904 53088
rect 20487 53057 20499 53060
rect 20441 53051 20499 53057
rect 20898 53048 20904 53060
rect 20956 53048 20962 53100
rect 22002 53048 22008 53100
rect 22060 53088 22066 53100
rect 22097 53091 22155 53097
rect 22097 53088 22109 53091
rect 22060 53060 22109 53088
rect 22060 53048 22066 53060
rect 22097 53057 22109 53060
rect 22143 53057 22155 53091
rect 22097 53051 22155 53057
rect 22833 53091 22891 53097
rect 22833 53057 22845 53091
rect 22879 53088 22891 53091
rect 23290 53088 23296 53100
rect 22879 53060 23296 53088
rect 22879 53057 22891 53060
rect 22833 53051 22891 53057
rect 23290 53048 23296 53060
rect 23348 53048 23354 53100
rect 24029 53091 24087 53097
rect 24029 53057 24041 53091
rect 24075 53088 24087 53091
rect 24578 53088 24584 53100
rect 24075 53060 24584 53088
rect 24075 53057 24087 53060
rect 24029 53051 24087 53057
rect 24578 53048 24584 53060
rect 24636 53048 24642 53100
rect 25682 53088 25688 53100
rect 25643 53060 25688 53088
rect 25682 53048 25688 53060
rect 25740 53048 25746 53100
rect 26620 53088 26648 53184
rect 27157 53091 27215 53097
rect 27157 53088 27169 53091
rect 26620 53060 27169 53088
rect 27157 53057 27169 53060
rect 27203 53057 27215 53091
rect 28258 53088 28264 53100
rect 28219 53060 28264 53088
rect 27157 53051 27215 53057
rect 28258 53048 28264 53060
rect 28316 53048 28322 53100
rect 29196 53088 29224 53184
rect 29917 53091 29975 53097
rect 29917 53088 29929 53091
rect 29196 53060 29929 53088
rect 29917 53057 29929 53060
rect 29963 53057 29975 53091
rect 30650 53088 30656 53100
rect 30611 53060 30656 53088
rect 29917 53051 29975 53057
rect 30650 53048 30656 53060
rect 30708 53088 30714 53100
rect 31113 53091 31171 53097
rect 31113 53088 31125 53091
rect 30708 53060 31125 53088
rect 30708 53048 30714 53060
rect 31113 53057 31125 53060
rect 31159 53057 31171 53091
rect 31772 53088 31800 53184
rect 32214 53116 32220 53168
rect 32272 53156 32278 53168
rect 47026 53156 47032 53168
rect 32272 53128 47032 53156
rect 32272 53116 32278 53128
rect 47026 53116 47032 53128
rect 47084 53116 47090 53168
rect 32493 53091 32551 53097
rect 32493 53088 32505 53091
rect 31772 53060 32505 53088
rect 31113 53051 31171 53057
rect 32493 53057 32505 53060
rect 32539 53057 32551 53091
rect 32493 53051 32551 53057
rect 32766 53048 32772 53100
rect 32824 53088 32830 53100
rect 33137 53091 33195 53097
rect 33137 53088 33149 53091
rect 32824 53060 33149 53088
rect 32824 53048 32830 53060
rect 33137 53057 33149 53060
rect 33183 53057 33195 53091
rect 34238 53088 34244 53100
rect 34199 53060 34244 53088
rect 33137 53051 33195 53057
rect 34238 53048 34244 53060
rect 34296 53048 34302 53100
rect 35434 53088 35440 53100
rect 35395 53060 35440 53088
rect 35434 53048 35440 53060
rect 35492 53088 35498 53100
rect 35897 53091 35955 53097
rect 35897 53088 35909 53091
rect 35492 53060 35909 53088
rect 35492 53048 35498 53060
rect 35897 53057 35909 53060
rect 35943 53057 35955 53091
rect 36630 53088 36636 53100
rect 36591 53060 36636 53088
rect 35897 53051 35955 53057
rect 36630 53048 36636 53060
rect 36688 53048 36694 53100
rect 37826 53088 37832 53100
rect 37787 53060 37832 53088
rect 37826 53048 37832 53060
rect 37884 53088 37890 53100
rect 38289 53091 38347 53097
rect 38289 53088 38301 53091
rect 37884 53060 38301 53088
rect 37884 53048 37890 53060
rect 38289 53057 38301 53060
rect 38335 53057 38347 53091
rect 39022 53088 39028 53100
rect 38983 53060 39028 53088
rect 38289 53051 38347 53057
rect 39022 53048 39028 53060
rect 39080 53048 39086 53100
rect 40034 53048 40040 53100
rect 40092 53088 40098 53100
rect 40221 53091 40279 53097
rect 40221 53088 40233 53091
rect 40092 53060 40233 53088
rect 40092 53048 40098 53060
rect 40221 53057 40233 53060
rect 40267 53088 40279 53091
rect 40681 53091 40739 53097
rect 40681 53088 40693 53091
rect 40267 53060 40693 53088
rect 40267 53057 40279 53060
rect 40221 53051 40279 53057
rect 40681 53057 40693 53060
rect 40727 53057 40739 53091
rect 41414 53088 41420 53100
rect 41375 53060 41420 53088
rect 40681 53051 40739 53057
rect 41414 53048 41420 53060
rect 41472 53088 41478 53100
rect 41877 53091 41935 53097
rect 41877 53088 41889 53091
rect 41472 53060 41889 53088
rect 41472 53048 41478 53060
rect 41877 53057 41889 53060
rect 41923 53057 41935 53091
rect 41877 53051 41935 53057
rect 42334 53048 42340 53100
rect 42392 53088 42398 53100
rect 42797 53091 42855 53097
rect 42797 53088 42809 53091
rect 42392 53060 42809 53088
rect 42392 53048 42398 53060
rect 42797 53057 42809 53060
rect 42843 53057 42855 53091
rect 43622 53088 43628 53100
rect 43583 53060 43628 53088
rect 42797 53051 42855 53057
rect 43622 53048 43628 53060
rect 43680 53048 43686 53100
rect 44726 53048 44732 53100
rect 44784 53088 44790 53100
rect 45186 53088 45192 53100
rect 44784 53060 45192 53088
rect 44784 53048 44790 53060
rect 45186 53048 45192 53060
rect 45244 53048 45250 53100
rect 47136 53088 47164 53184
rect 47765 53091 47823 53097
rect 47765 53088 47777 53091
rect 47136 53060 47777 53088
rect 47765 53057 47777 53060
rect 47811 53057 47823 53091
rect 49712 53088 49740 53184
rect 51074 53116 51080 53168
rect 51132 53156 51138 53168
rect 51442 53156 51448 53168
rect 51132 53128 51448 53156
rect 51132 53116 51138 53128
rect 51442 53116 51448 53128
rect 51500 53156 51506 53168
rect 51813 53159 51871 53165
rect 51813 53156 51825 53159
rect 51500 53128 51825 53156
rect 51500 53116 51506 53128
rect 51813 53125 51825 53128
rect 51859 53125 51871 53159
rect 51813 53119 51871 53125
rect 50341 53091 50399 53097
rect 50341 53088 50353 53091
rect 49712 53060 50353 53088
rect 47765 53051 47823 53057
rect 50341 53057 50353 53060
rect 50387 53057 50399 53091
rect 53190 53088 53196 53100
rect 53151 53060 53196 53088
rect 50341 53051 50399 53057
rect 53190 53048 53196 53060
rect 53248 53048 53254 53100
rect 16546 52992 18368 53020
rect 18601 53023 18659 53029
rect 4341 52955 4399 52961
rect 4341 52921 4353 52955
rect 4387 52952 4399 52955
rect 16546 52952 16574 52992
rect 18601 52989 18613 53023
rect 18647 53020 18659 53023
rect 21450 53020 21456 53032
rect 18647 52992 21456 53020
rect 18647 52989 18659 52992
rect 18601 52983 18659 52989
rect 21450 52980 21456 52992
rect 21508 52980 21514 53032
rect 34790 52980 34796 53032
rect 34848 53020 34854 53032
rect 43898 53020 43904 53032
rect 34848 52992 40724 53020
rect 43859 52992 43904 53020
rect 34848 52980 34854 52992
rect 4387 52924 16574 52952
rect 19889 52955 19947 52961
rect 4387 52921 4399 52924
rect 4341 52915 4399 52921
rect 19889 52921 19901 52955
rect 19935 52952 19947 52955
rect 24026 52952 24032 52964
rect 19935 52924 24032 52952
rect 19935 52921 19947 52924
rect 19889 52915 19947 52921
rect 24026 52912 24032 52924
rect 24084 52912 24090 52964
rect 24765 52955 24823 52961
rect 24765 52921 24777 52955
rect 24811 52952 24823 52955
rect 26694 52952 26700 52964
rect 24811 52924 26700 52952
rect 24811 52921 24823 52924
rect 24765 52915 24823 52921
rect 26694 52912 26700 52924
rect 26752 52912 26758 52964
rect 32122 52912 32128 52964
rect 32180 52952 32186 52964
rect 32953 52955 33011 52961
rect 32953 52952 32965 52955
rect 32180 52924 32965 52952
rect 32180 52912 32186 52924
rect 32953 52921 32965 52924
rect 32999 52921 33011 52955
rect 32953 52915 33011 52921
rect 34698 52912 34704 52964
rect 34756 52952 34762 52964
rect 37645 52955 37703 52961
rect 37645 52952 37657 52955
rect 34756 52924 37657 52952
rect 34756 52912 34762 52924
rect 37645 52921 37657 52924
rect 37691 52921 37703 52955
rect 40696 52952 40724 52992
rect 43898 52980 43904 52992
rect 43956 52980 43962 53032
rect 45462 53020 45468 53032
rect 45423 52992 45468 53020
rect 45462 52980 45468 52992
rect 45520 52980 45526 53032
rect 48038 53020 48044 53032
rect 47999 52992 48044 53020
rect 48038 52980 48044 52992
rect 48096 52980 48102 53032
rect 50154 52980 50160 53032
rect 50212 53020 50218 53032
rect 50617 53023 50675 53029
rect 50617 53020 50629 53023
rect 50212 52992 50629 53020
rect 50212 52980 50218 52992
rect 50617 52989 50629 52992
rect 50663 52989 50675 53023
rect 50617 52983 50675 52989
rect 53469 53023 53527 53029
rect 53469 52989 53481 53023
rect 53515 52989 53527 53023
rect 53469 52983 53527 52989
rect 51629 52955 51687 52961
rect 51629 52952 51641 52955
rect 40696 52924 51641 52952
rect 37645 52915 37703 52921
rect 51629 52921 51641 52924
rect 51675 52921 51687 52955
rect 51629 52915 51687 52921
rect 3234 52884 3240 52896
rect 3195 52856 3240 52884
rect 3234 52844 3240 52856
rect 3292 52844 3298 52896
rect 5534 52884 5540 52896
rect 5495 52856 5540 52884
rect 5534 52844 5540 52856
rect 5592 52844 5598 52896
rect 6730 52884 6736 52896
rect 6691 52856 6736 52884
rect 6730 52844 6736 52856
rect 6788 52844 6794 52896
rect 7929 52887 7987 52893
rect 7929 52853 7941 52887
rect 7975 52884 7987 52887
rect 11698 52884 11704 52896
rect 7975 52856 11704 52884
rect 7975 52853 7987 52856
rect 7929 52847 7987 52853
rect 11698 52844 11704 52856
rect 11756 52844 11762 52896
rect 15010 52884 15016 52896
rect 14971 52856 15016 52884
rect 15010 52844 15016 52856
rect 15068 52844 15074 52896
rect 22278 52884 22284 52896
rect 22239 52856 22284 52884
rect 22278 52844 22284 52856
rect 22336 52844 22342 52896
rect 23477 52887 23535 52893
rect 23477 52853 23489 52887
rect 23523 52884 23535 52887
rect 25406 52884 25412 52896
rect 23523 52856 25412 52884
rect 23523 52853 23535 52856
rect 23477 52847 23535 52853
rect 25406 52844 25412 52856
rect 25464 52844 25470 52896
rect 25869 52887 25927 52893
rect 25869 52853 25881 52887
rect 25915 52884 25927 52887
rect 25958 52884 25964 52896
rect 25915 52856 25964 52884
rect 25915 52853 25927 52856
rect 25869 52847 25927 52853
rect 25958 52844 25964 52856
rect 26016 52844 26022 52896
rect 26970 52844 26976 52896
rect 27028 52884 27034 52896
rect 27341 52887 27399 52893
rect 27341 52884 27353 52887
rect 27028 52856 27353 52884
rect 27028 52844 27034 52856
rect 27341 52853 27353 52856
rect 27387 52853 27399 52887
rect 28074 52884 28080 52896
rect 28035 52856 28080 52884
rect 27341 52847 27399 52853
rect 28074 52844 28080 52856
rect 28132 52844 28138 52896
rect 28718 52844 28724 52896
rect 28776 52884 28782 52896
rect 29733 52887 29791 52893
rect 29733 52884 29745 52887
rect 28776 52856 29745 52884
rect 28776 52844 28782 52856
rect 29733 52853 29745 52856
rect 29779 52853 29791 52887
rect 29733 52847 29791 52853
rect 30098 52844 30104 52896
rect 30156 52884 30162 52896
rect 30469 52887 30527 52893
rect 30469 52884 30481 52887
rect 30156 52856 30481 52884
rect 30156 52844 30162 52856
rect 30469 52853 30481 52856
rect 30515 52853 30527 52887
rect 30469 52847 30527 52853
rect 31202 52844 31208 52896
rect 31260 52884 31266 52896
rect 32309 52887 32367 52893
rect 32309 52884 32321 52887
rect 31260 52856 32321 52884
rect 31260 52844 31266 52856
rect 32309 52853 32321 52856
rect 32355 52853 32367 52887
rect 32309 52847 32367 52853
rect 32582 52844 32588 52896
rect 32640 52884 32646 52896
rect 34057 52887 34115 52893
rect 34057 52884 34069 52887
rect 32640 52856 34069 52884
rect 32640 52844 32646 52856
rect 34057 52853 34069 52856
rect 34103 52853 34115 52887
rect 34057 52847 34115 52853
rect 34330 52844 34336 52896
rect 34388 52884 34394 52896
rect 35253 52887 35311 52893
rect 35253 52884 35265 52887
rect 34388 52856 35265 52884
rect 34388 52844 34394 52856
rect 35253 52853 35265 52856
rect 35299 52853 35311 52887
rect 35253 52847 35311 52853
rect 35342 52844 35348 52896
rect 35400 52884 35406 52896
rect 36449 52887 36507 52893
rect 36449 52884 36461 52887
rect 35400 52856 36461 52884
rect 35400 52844 35406 52856
rect 36449 52853 36461 52856
rect 36495 52853 36507 52887
rect 38838 52884 38844 52896
rect 38799 52856 38844 52884
rect 36449 52847 36507 52853
rect 38838 52844 38844 52856
rect 38896 52844 38902 52896
rect 38930 52844 38936 52896
rect 38988 52884 38994 52896
rect 40037 52887 40095 52893
rect 40037 52884 40049 52887
rect 38988 52856 40049 52884
rect 38988 52844 38994 52856
rect 40037 52853 40049 52856
rect 40083 52853 40095 52887
rect 41230 52884 41236 52896
rect 41191 52856 41236 52884
rect 40037 52847 40095 52853
rect 41230 52844 41236 52856
rect 41288 52844 41294 52896
rect 42610 52884 42616 52896
rect 42571 52856 42616 52884
rect 42610 52844 42616 52856
rect 42668 52844 42674 52896
rect 49510 52844 49516 52896
rect 49568 52884 49574 52896
rect 53484 52884 53512 52983
rect 49568 52856 53512 52884
rect 49568 52844 49574 52856
rect 1104 52794 54832 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 54832 52794
rect 1104 52720 54832 52742
rect 3142 52680 3148 52692
rect 3103 52652 3148 52680
rect 3142 52640 3148 52652
rect 3200 52640 3206 52692
rect 4062 52680 4068 52692
rect 4023 52652 4068 52680
rect 4062 52640 4068 52652
rect 4120 52640 4126 52692
rect 6457 52683 6515 52689
rect 6457 52649 6469 52683
rect 6503 52680 6515 52683
rect 6638 52680 6644 52692
rect 6503 52652 6644 52680
rect 6503 52649 6515 52652
rect 6457 52643 6515 52649
rect 6638 52640 6644 52652
rect 6696 52640 6702 52692
rect 7653 52683 7711 52689
rect 7653 52649 7665 52683
rect 7699 52680 7711 52683
rect 7742 52680 7748 52692
rect 7699 52652 7748 52680
rect 7699 52649 7711 52652
rect 7653 52643 7711 52649
rect 7742 52640 7748 52652
rect 7800 52640 7806 52692
rect 10045 52683 10103 52689
rect 10045 52649 10057 52683
rect 10091 52680 10103 52683
rect 10134 52680 10140 52692
rect 10091 52652 10140 52680
rect 10091 52649 10103 52652
rect 10045 52643 10103 52649
rect 10134 52640 10140 52652
rect 10192 52640 10198 52692
rect 13630 52680 13636 52692
rect 13591 52652 13636 52680
rect 13630 52640 13636 52652
rect 13688 52640 13694 52692
rect 14826 52640 14832 52692
rect 14884 52680 14890 52692
rect 15105 52683 15163 52689
rect 15105 52680 15117 52683
rect 14884 52652 15117 52680
rect 14884 52640 14890 52652
rect 15105 52649 15117 52652
rect 15151 52649 15163 52683
rect 18782 52680 18788 52692
rect 18743 52652 18788 52680
rect 15105 52643 15163 52649
rect 18782 52640 18788 52652
rect 18840 52640 18846 52692
rect 19426 52640 19432 52692
rect 19484 52680 19490 52692
rect 19521 52683 19579 52689
rect 19521 52680 19533 52683
rect 19484 52652 19533 52680
rect 19484 52640 19490 52652
rect 19521 52649 19533 52652
rect 19567 52649 19579 52683
rect 22002 52680 22008 52692
rect 21963 52652 22008 52680
rect 19521 52643 19579 52649
rect 22002 52640 22008 52652
rect 22060 52640 22066 52692
rect 25682 52640 25688 52692
rect 25740 52680 25746 52692
rect 26329 52683 26387 52689
rect 26329 52680 26341 52683
rect 25740 52652 26341 52680
rect 25740 52640 25746 52652
rect 26329 52649 26341 52652
rect 26375 52649 26387 52683
rect 26329 52643 26387 52649
rect 27985 52683 28043 52689
rect 27985 52649 27997 52683
rect 28031 52680 28043 52683
rect 28258 52680 28264 52692
rect 28031 52652 28264 52680
rect 28031 52649 28043 52652
rect 27985 52643 28043 52649
rect 28258 52640 28264 52652
rect 28316 52640 28322 52692
rect 32766 52680 32772 52692
rect 32727 52652 32772 52680
rect 32766 52640 32772 52652
rect 32824 52640 32830 52692
rect 33965 52683 34023 52689
rect 33965 52649 33977 52683
rect 34011 52680 34023 52683
rect 34238 52680 34244 52692
rect 34011 52652 34244 52680
rect 34011 52649 34023 52652
rect 33965 52643 34023 52649
rect 34238 52640 34244 52652
rect 34296 52640 34302 52692
rect 36357 52683 36415 52689
rect 36357 52649 36369 52683
rect 36403 52680 36415 52683
rect 36630 52680 36636 52692
rect 36403 52652 36636 52680
rect 36403 52649 36415 52652
rect 36357 52643 36415 52649
rect 36630 52640 36636 52652
rect 36688 52640 36694 52692
rect 38749 52683 38807 52689
rect 38749 52649 38761 52683
rect 38795 52680 38807 52683
rect 39022 52680 39028 52692
rect 38795 52652 39028 52680
rect 38795 52649 38807 52652
rect 38749 52643 38807 52649
rect 39022 52640 39028 52652
rect 39080 52640 39086 52692
rect 42334 52640 42340 52692
rect 42392 52680 42398 52692
rect 42429 52683 42487 52689
rect 42429 52680 42441 52683
rect 42392 52652 42441 52680
rect 42392 52640 42398 52652
rect 42429 52649 42441 52652
rect 42475 52649 42487 52683
rect 42429 52643 42487 52649
rect 43533 52683 43591 52689
rect 43533 52649 43545 52683
rect 43579 52680 43591 52683
rect 43622 52680 43628 52692
rect 43579 52652 43628 52680
rect 43579 52649 43591 52652
rect 43533 52643 43591 52649
rect 43622 52640 43628 52652
rect 43680 52640 43686 52692
rect 45186 52680 45192 52692
rect 45147 52652 45192 52680
rect 45186 52640 45192 52652
rect 45244 52640 45250 52692
rect 51537 52683 51595 52689
rect 51537 52649 51549 52683
rect 51583 52680 51595 52683
rect 51902 52680 51908 52692
rect 51583 52652 51908 52680
rect 51583 52649 51595 52652
rect 51537 52643 51595 52649
rect 51902 52640 51908 52652
rect 51960 52640 51966 52692
rect 53101 52683 53159 52689
rect 53101 52649 53113 52683
rect 53147 52680 53159 52683
rect 53190 52680 53196 52692
rect 53147 52652 53196 52680
rect 53147 52649 53159 52652
rect 53101 52643 53159 52649
rect 53190 52640 53196 52652
rect 53248 52640 53254 52692
rect 34514 52572 34520 52624
rect 34572 52612 34578 52624
rect 41230 52612 41236 52624
rect 34572 52584 41236 52612
rect 34572 52572 34578 52584
rect 41230 52572 41236 52584
rect 41288 52572 41294 52624
rect 47026 52572 47032 52624
rect 47084 52612 47090 52624
rect 47084 52584 48728 52612
rect 47084 52572 47090 52584
rect 10873 52547 10931 52553
rect 10873 52513 10885 52547
rect 10919 52544 10931 52547
rect 11330 52544 11336 52556
rect 10919 52516 11336 52544
rect 10919 52513 10931 52516
rect 10873 52507 10931 52513
rect 11330 52504 11336 52516
rect 11388 52504 11394 52556
rect 16853 52547 16911 52553
rect 16853 52513 16865 52547
rect 16899 52544 16911 52547
rect 17310 52544 17316 52556
rect 16899 52516 17316 52544
rect 16899 52513 16911 52516
rect 16853 52507 16911 52513
rect 17310 52504 17316 52516
rect 17368 52504 17374 52556
rect 33042 52504 33048 52556
rect 33100 52544 33106 52556
rect 42610 52544 42616 52556
rect 33100 52516 42616 52544
rect 33100 52504 33106 52516
rect 42610 52504 42616 52516
rect 42668 52504 42674 52556
rect 46014 52544 46020 52556
rect 45975 52516 46020 52544
rect 46014 52504 46020 52516
rect 46072 52504 46078 52556
rect 47949 52547 48007 52553
rect 47949 52513 47961 52547
rect 47995 52544 48007 52547
rect 48406 52544 48412 52556
rect 47995 52516 48412 52544
rect 47995 52513 48007 52516
rect 47949 52507 48007 52513
rect 48406 52504 48412 52516
rect 48464 52504 48470 52556
rect 48700 52553 48728 52584
rect 48685 52547 48743 52553
rect 48685 52513 48697 52547
rect 48731 52513 48743 52547
rect 51994 52544 52000 52556
rect 51955 52516 52000 52544
rect 48685 52507 48743 52513
rect 51994 52504 52000 52516
rect 52052 52504 52058 52556
rect 1762 52436 1768 52488
rect 1820 52476 1826 52488
rect 1857 52479 1915 52485
rect 1857 52476 1869 52479
rect 1820 52448 1869 52476
rect 1820 52436 1826 52448
rect 1857 52445 1869 52448
rect 1903 52445 1915 52479
rect 1857 52439 1915 52445
rect 2498 52436 2504 52488
rect 2556 52476 2562 52488
rect 2593 52479 2651 52485
rect 2593 52476 2605 52479
rect 2556 52448 2605 52476
rect 2556 52436 2562 52448
rect 2593 52445 2605 52448
rect 2639 52445 2651 52479
rect 11606 52476 11612 52488
rect 11567 52448 11612 52476
rect 2593 52439 2651 52445
rect 11606 52436 11612 52448
rect 11664 52436 11670 52488
rect 13630 52436 13636 52488
rect 13688 52476 13694 52488
rect 14461 52479 14519 52485
rect 14461 52476 14473 52479
rect 13688 52448 14473 52476
rect 13688 52436 13694 52448
rect 14461 52445 14473 52448
rect 14507 52445 14519 52479
rect 14461 52439 14519 52445
rect 17589 52479 17647 52485
rect 17589 52445 17601 52479
rect 17635 52476 17647 52479
rect 22830 52476 22836 52488
rect 17635 52448 22836 52476
rect 17635 52445 17647 52448
rect 17589 52439 17647 52445
rect 22830 52436 22836 52448
rect 22888 52436 22894 52488
rect 26050 52436 26056 52488
rect 26108 52476 26114 52488
rect 27154 52476 27160 52488
rect 26108 52448 27160 52476
rect 26108 52436 26114 52448
rect 27154 52436 27160 52448
rect 27212 52436 27218 52488
rect 46290 52476 46296 52488
rect 46251 52448 46296 52476
rect 46290 52436 46296 52448
rect 46348 52436 46354 52488
rect 51902 52436 51908 52488
rect 51960 52476 51966 52488
rect 52181 52479 52239 52485
rect 52181 52476 52193 52479
rect 51960 52448 52193 52476
rect 51960 52436 51966 52448
rect 52181 52445 52193 52448
rect 52227 52445 52239 52479
rect 54018 52476 54024 52488
rect 53979 52448 54024 52476
rect 52181 52439 52239 52445
rect 54018 52436 54024 52448
rect 54076 52436 54082 52488
rect 1673 52411 1731 52417
rect 1673 52377 1685 52411
rect 1719 52408 1731 52411
rect 2409 52411 2467 52417
rect 1719 52380 1808 52408
rect 1719 52377 1731 52380
rect 1673 52371 1731 52377
rect 1486 52300 1492 52352
rect 1544 52340 1550 52352
rect 1780 52340 1808 52380
rect 2409 52377 2421 52411
rect 2455 52408 2467 52411
rect 2774 52408 2780 52420
rect 2455 52380 2780 52408
rect 2455 52377 2467 52380
rect 2409 52371 2467 52377
rect 2774 52368 2780 52380
rect 2832 52368 2838 52420
rect 54205 52411 54263 52417
rect 54205 52377 54217 52411
rect 54251 52408 54263 52411
rect 54294 52408 54300 52420
rect 54251 52380 54300 52408
rect 54251 52377 54263 52380
rect 54205 52371 54263 52377
rect 54294 52368 54300 52380
rect 54352 52368 54358 52420
rect 2866 52340 2872 52352
rect 1544 52312 2872 52340
rect 1544 52300 1550 52312
rect 2866 52300 2872 52312
rect 2924 52300 2930 52352
rect 14274 52340 14280 52352
rect 14235 52312 14280 52340
rect 14274 52300 14280 52312
rect 14332 52300 14338 52352
rect 25498 52300 25504 52352
rect 25556 52340 25562 52352
rect 25777 52343 25835 52349
rect 25777 52340 25789 52343
rect 25556 52312 25789 52340
rect 25556 52300 25562 52312
rect 25777 52309 25789 52312
rect 25823 52309 25835 52343
rect 25777 52303 25835 52309
rect 1104 52250 54832 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 54832 52250
rect 1104 52176 54832 52198
rect 2409 52139 2467 52145
rect 2409 52105 2421 52139
rect 2455 52136 2467 52139
rect 2774 52136 2780 52148
rect 2455 52108 2780 52136
rect 2455 52105 2467 52108
rect 2409 52099 2467 52105
rect 2774 52096 2780 52108
rect 2832 52096 2838 52148
rect 24486 52096 24492 52148
rect 24544 52136 24550 52148
rect 24581 52139 24639 52145
rect 24581 52136 24593 52139
rect 24544 52108 24593 52136
rect 24544 52096 24550 52108
rect 24581 52105 24593 52108
rect 24627 52105 24639 52139
rect 26050 52136 26056 52148
rect 24581 52099 24639 52105
rect 25240 52108 26056 52136
rect 2590 52028 2596 52080
rect 2648 52068 2654 52080
rect 3421 52071 3479 52077
rect 3421 52068 3433 52071
rect 2648 52040 3433 52068
rect 2648 52028 2654 52040
rect 3421 52037 3433 52040
rect 3467 52037 3479 52071
rect 3421 52031 3479 52037
rect 1670 52000 1676 52012
rect 1631 51972 1676 52000
rect 1670 51960 1676 51972
rect 1728 52000 1734 52012
rect 2869 52003 2927 52009
rect 2869 52000 2881 52003
rect 1728 51972 2881 52000
rect 1728 51960 1734 51972
rect 2869 51969 2881 51972
rect 2915 51969 2927 52003
rect 24596 52000 24624 52099
rect 25133 52003 25191 52009
rect 25133 52000 25145 52003
rect 24596 51972 25145 52000
rect 2869 51963 2927 51969
rect 25133 51969 25145 51972
rect 25179 51969 25191 52003
rect 25240 52000 25268 52108
rect 26050 52096 26056 52108
rect 26108 52096 26114 52148
rect 45925 52139 45983 52145
rect 45925 52105 45937 52139
rect 45971 52136 45983 52139
rect 46014 52136 46020 52148
rect 45971 52108 46020 52136
rect 45971 52105 45983 52108
rect 45925 52099 45983 52105
rect 46014 52096 46020 52108
rect 46072 52096 46078 52148
rect 51442 52136 51448 52148
rect 51403 52108 51448 52136
rect 51442 52096 51448 52108
rect 51500 52096 51506 52148
rect 54294 52136 54300 52148
rect 54255 52108 54300 52136
rect 54294 52096 54300 52108
rect 54352 52096 54358 52148
rect 25406 52068 25412 52080
rect 25367 52040 25412 52068
rect 25406 52028 25412 52040
rect 25464 52028 25470 52080
rect 27154 52028 27160 52080
rect 27212 52068 27218 52080
rect 27709 52071 27767 52077
rect 27709 52068 27721 52071
rect 27212 52040 27721 52068
rect 27212 52028 27218 52040
rect 27709 52037 27721 52040
rect 27755 52037 27767 52071
rect 27709 52031 27767 52037
rect 27801 52071 27859 52077
rect 27801 52037 27813 52071
rect 27847 52068 27859 52071
rect 28074 52068 28080 52080
rect 27847 52040 28080 52068
rect 27847 52037 27859 52040
rect 27801 52031 27859 52037
rect 28074 52028 28080 52040
rect 28132 52028 28138 52080
rect 25317 52003 25375 52009
rect 25317 52000 25329 52003
rect 25240 51972 25329 52000
rect 25133 51963 25191 51969
rect 25317 51969 25329 51972
rect 25363 51969 25375 52003
rect 25317 51963 25375 51969
rect 25498 51960 25504 52012
rect 25556 52000 25562 52012
rect 26605 52003 26663 52009
rect 26605 52000 26617 52003
rect 25556 51972 25601 52000
rect 26206 51972 26617 52000
rect 25556 51960 25562 51972
rect 9306 51892 9312 51944
rect 9364 51932 9370 51944
rect 26206 51932 26234 51972
rect 26605 51969 26617 51972
rect 26651 52000 26663 52003
rect 27525 52003 27583 52009
rect 27525 52000 27537 52003
rect 26651 51972 27537 52000
rect 26651 51969 26663 51972
rect 26605 51963 26663 51969
rect 27525 51969 27537 51972
rect 27571 51969 27583 52003
rect 27890 52000 27896 52012
rect 27851 51972 27896 52000
rect 27525 51963 27583 51969
rect 27890 51960 27896 51972
rect 27948 51960 27954 52012
rect 9364 51904 26234 51932
rect 9364 51892 9370 51904
rect 1854 51864 1860 51876
rect 1815 51836 1860 51864
rect 1854 51824 1860 51836
rect 1912 51824 1918 51876
rect 32674 51824 32680 51876
rect 32732 51864 32738 51876
rect 49510 51864 49516 51876
rect 32732 51836 49516 51864
rect 32732 51824 32738 51836
rect 49510 51824 49516 51836
rect 49568 51824 49574 51876
rect 25685 51799 25743 51805
rect 25685 51765 25697 51799
rect 25731 51796 25743 51799
rect 27614 51796 27620 51808
rect 25731 51768 27620 51796
rect 25731 51765 25743 51768
rect 25685 51759 25743 51765
rect 27614 51756 27620 51768
rect 27672 51756 27678 51808
rect 28077 51799 28135 51805
rect 28077 51765 28089 51799
rect 28123 51796 28135 51799
rect 29822 51796 29828 51808
rect 28123 51768 29828 51796
rect 28123 51765 28135 51768
rect 28077 51759 28135 51765
rect 29822 51756 29828 51768
rect 29880 51756 29886 51808
rect 1104 51706 54832 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 54832 51706
rect 1104 51632 54832 51654
rect 2866 51592 2872 51604
rect 2827 51564 2872 51592
rect 2866 51552 2872 51564
rect 2924 51552 2930 51604
rect 25498 51552 25504 51604
rect 25556 51592 25562 51604
rect 27341 51595 27399 51601
rect 27341 51592 27353 51595
rect 25556 51564 27353 51592
rect 25556 51552 25562 51564
rect 27341 51561 27353 51564
rect 27387 51592 27399 51595
rect 27890 51592 27896 51604
rect 27387 51564 27896 51592
rect 27387 51561 27399 51564
rect 27341 51555 27399 51561
rect 27890 51552 27896 51564
rect 27948 51592 27954 51604
rect 29638 51592 29644 51604
rect 27948 51564 29644 51592
rect 27948 51552 27954 51564
rect 29638 51552 29644 51564
rect 29696 51552 29702 51604
rect 1670 51320 1676 51332
rect 1631 51292 1676 51320
rect 1670 51280 1676 51292
rect 1728 51320 1734 51332
rect 2317 51323 2375 51329
rect 2317 51320 2329 51323
rect 1728 51292 2329 51320
rect 1728 51280 1734 51292
rect 2317 51289 2329 51292
rect 2363 51289 2375 51323
rect 2317 51283 2375 51289
rect 53745 51323 53803 51329
rect 53745 51289 53757 51323
rect 53791 51320 53803 51323
rect 54386 51320 54392 51332
rect 53791 51292 54392 51320
rect 53791 51289 53803 51292
rect 53745 51283 53803 51289
rect 54386 51280 54392 51292
rect 54444 51280 54450 51332
rect 1765 51255 1823 51261
rect 1765 51221 1777 51255
rect 1811 51252 1823 51255
rect 2682 51252 2688 51264
rect 1811 51224 2688 51252
rect 1811 51221 1823 51224
rect 1765 51215 1823 51221
rect 2682 51212 2688 51224
rect 2740 51212 2746 51264
rect 26050 51252 26056 51264
rect 26011 51224 26056 51252
rect 26050 51212 26056 51224
rect 26108 51212 26114 51264
rect 54294 51252 54300 51264
rect 54255 51224 54300 51252
rect 54294 51212 54300 51224
rect 54352 51212 54358 51264
rect 1104 51162 54832 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 54832 51162
rect 1104 51088 54832 51110
rect 54297 50915 54355 50921
rect 54297 50881 54309 50915
rect 54343 50912 54355 50915
rect 54386 50912 54392 50924
rect 54343 50884 54392 50912
rect 54343 50881 54355 50884
rect 54297 50875 54355 50881
rect 54386 50872 54392 50884
rect 54444 50872 54450 50924
rect 2133 50847 2191 50853
rect 2133 50813 2145 50847
rect 2179 50844 2191 50847
rect 2314 50844 2320 50856
rect 2179 50816 2320 50844
rect 2179 50813 2191 50816
rect 2133 50807 2191 50813
rect 2314 50804 2320 50816
rect 2372 50804 2378 50856
rect 2409 50847 2467 50853
rect 2409 50813 2421 50847
rect 2455 50844 2467 50847
rect 2774 50844 2780 50856
rect 2455 50816 2780 50844
rect 2455 50813 2467 50816
rect 2409 50807 2467 50813
rect 2774 50804 2780 50816
rect 2832 50844 2838 50856
rect 2869 50847 2927 50853
rect 2869 50844 2881 50847
rect 2832 50816 2881 50844
rect 2832 50804 2838 50816
rect 2869 50813 2881 50816
rect 2915 50813 2927 50847
rect 2869 50807 2927 50813
rect 53558 50708 53564 50720
rect 53519 50680 53564 50708
rect 53558 50668 53564 50680
rect 53616 50668 53622 50720
rect 53926 50668 53932 50720
rect 53984 50708 53990 50720
rect 54113 50711 54171 50717
rect 54113 50708 54125 50711
rect 53984 50680 54125 50708
rect 53984 50668 53990 50680
rect 54113 50677 54125 50680
rect 54159 50677 54171 50711
rect 54113 50671 54171 50677
rect 1104 50618 54832 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 54832 50618
rect 1104 50544 54832 50566
rect 16022 50396 16028 50448
rect 16080 50436 16086 50448
rect 25130 50436 25136 50448
rect 16080 50408 25136 50436
rect 16080 50396 16086 50408
rect 25130 50396 25136 50408
rect 25188 50396 25194 50448
rect 52270 50396 52276 50448
rect 52328 50436 52334 50448
rect 54113 50439 54171 50445
rect 54113 50436 54125 50439
rect 52328 50408 54125 50436
rect 52328 50396 52334 50408
rect 54113 50405 54125 50408
rect 54159 50405 54171 50439
rect 54113 50399 54171 50405
rect 8202 50328 8208 50380
rect 8260 50368 8266 50380
rect 25406 50368 25412 50380
rect 8260 50340 25412 50368
rect 8260 50328 8266 50340
rect 25406 50328 25412 50340
rect 25464 50328 25470 50380
rect 29914 50328 29920 50380
rect 29972 50368 29978 50380
rect 45462 50368 45468 50380
rect 29972 50340 45468 50368
rect 29972 50328 29978 50340
rect 45462 50328 45468 50340
rect 45520 50328 45526 50380
rect 2130 50300 2136 50312
rect 2091 50272 2136 50300
rect 2130 50260 2136 50272
rect 2188 50260 2194 50312
rect 2409 50303 2467 50309
rect 2409 50269 2421 50303
rect 2455 50300 2467 50303
rect 2774 50300 2780 50312
rect 2455 50272 2780 50300
rect 2455 50269 2467 50272
rect 2409 50263 2467 50269
rect 2774 50260 2780 50272
rect 2832 50300 2838 50312
rect 2869 50303 2927 50309
rect 2869 50300 2881 50303
rect 2832 50272 2881 50300
rect 2832 50260 2838 50272
rect 2869 50269 2881 50272
rect 2915 50269 2927 50303
rect 54294 50300 54300 50312
rect 54255 50272 54300 50300
rect 2869 50263 2927 50269
rect 54294 50260 54300 50272
rect 54352 50260 54358 50312
rect 52641 50235 52699 50241
rect 52641 50201 52653 50235
rect 52687 50232 52699 50235
rect 54478 50232 54484 50244
rect 52687 50204 54484 50232
rect 52687 50201 52699 50204
rect 52641 50195 52699 50201
rect 54478 50192 54484 50204
rect 54536 50192 54542 50244
rect 53098 50164 53104 50176
rect 53059 50136 53104 50164
rect 53098 50124 53104 50136
rect 53156 50124 53162 50176
rect 1104 50074 54832 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 54832 50074
rect 1104 50000 54832 50022
rect 54113 49963 54171 49969
rect 54113 49960 54125 49963
rect 51046 49932 54125 49960
rect 48130 49852 48136 49904
rect 48188 49892 48194 49904
rect 51046 49892 51074 49932
rect 54113 49929 54125 49932
rect 54159 49929 54171 49963
rect 54113 49923 54171 49929
rect 48188 49864 51074 49892
rect 48188 49852 48194 49864
rect 1670 49824 1676 49836
rect 1631 49796 1676 49824
rect 1670 49784 1676 49796
rect 1728 49824 1734 49836
rect 2317 49827 2375 49833
rect 2317 49824 2329 49827
rect 1728 49796 2329 49824
rect 1728 49784 1734 49796
rect 2317 49793 2329 49796
rect 2363 49793 2375 49827
rect 2317 49787 2375 49793
rect 52365 49827 52423 49833
rect 52365 49793 52377 49827
rect 52411 49824 52423 49827
rect 53650 49824 53656 49836
rect 52411 49796 53656 49824
rect 52411 49793 52423 49796
rect 52365 49787 52423 49793
rect 53650 49784 53656 49796
rect 53708 49784 53714 49836
rect 54297 49827 54355 49833
rect 54297 49793 54309 49827
rect 54343 49824 54355 49827
rect 54478 49824 54484 49836
rect 54343 49796 54484 49824
rect 54343 49793 54355 49796
rect 54297 49787 54355 49793
rect 54478 49784 54484 49796
rect 54536 49784 54542 49836
rect 1857 49759 1915 49765
rect 1857 49725 1869 49759
rect 1903 49756 1915 49759
rect 2038 49756 2044 49768
rect 1903 49728 2044 49756
rect 1903 49725 1915 49728
rect 1857 49719 1915 49725
rect 2038 49716 2044 49728
rect 2096 49716 2102 49768
rect 51166 49716 51172 49768
rect 51224 49756 51230 49768
rect 51224 49728 53512 49756
rect 51224 49716 51230 49728
rect 53484 49697 53512 49728
rect 53469 49691 53527 49697
rect 53469 49657 53481 49691
rect 53515 49657 53527 49691
rect 53469 49651 53527 49657
rect 52914 49620 52920 49632
rect 52875 49592 52920 49620
rect 52914 49580 52920 49592
rect 52972 49580 52978 49632
rect 1104 49530 54832 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 54832 49530
rect 1104 49456 54832 49478
rect 53745 49283 53803 49289
rect 53745 49280 53757 49283
rect 45526 49252 53757 49280
rect 2133 49215 2191 49221
rect 2133 49181 2145 49215
rect 2179 49212 2191 49215
rect 2314 49212 2320 49224
rect 2179 49184 2320 49212
rect 2179 49181 2191 49184
rect 2133 49175 2191 49181
rect 2314 49172 2320 49184
rect 2372 49172 2378 49224
rect 2409 49215 2467 49221
rect 2409 49181 2421 49215
rect 2455 49212 2467 49215
rect 2774 49212 2780 49224
rect 2455 49184 2780 49212
rect 2455 49181 2467 49184
rect 2409 49175 2467 49181
rect 2774 49172 2780 49184
rect 2832 49212 2838 49224
rect 2869 49215 2927 49221
rect 2869 49212 2881 49215
rect 2832 49184 2881 49212
rect 2832 49172 2838 49184
rect 2869 49181 2881 49184
rect 2915 49181 2927 49215
rect 2869 49175 2927 49181
rect 38654 49172 38660 49224
rect 38712 49212 38718 49224
rect 45526 49212 45554 49252
rect 53745 49249 53757 49252
rect 53791 49249 53803 49283
rect 53745 49243 53803 49249
rect 38712 49184 45554 49212
rect 52273 49215 52331 49221
rect 38712 49172 38718 49184
rect 52273 49181 52285 49215
rect 52319 49212 52331 49215
rect 52638 49212 52644 49224
rect 52319 49184 52644 49212
rect 52319 49181 52331 49184
rect 52273 49175 52331 49181
rect 52638 49172 52644 49184
rect 52696 49172 52702 49224
rect 53009 49215 53067 49221
rect 53009 49181 53021 49215
rect 53055 49212 53067 49215
rect 53098 49212 53104 49224
rect 53055 49184 53104 49212
rect 53055 49181 53067 49184
rect 53009 49175 53067 49181
rect 53098 49172 53104 49184
rect 53156 49172 53162 49224
rect 53469 49215 53527 49221
rect 53469 49181 53481 49215
rect 53515 49212 53527 49215
rect 53558 49212 53564 49224
rect 53515 49184 53564 49212
rect 53515 49181 53527 49184
rect 53469 49175 53527 49181
rect 53558 49172 53564 49184
rect 53616 49172 53622 49224
rect 51813 49147 51871 49153
rect 51813 49113 51825 49147
rect 51859 49144 51871 49147
rect 52362 49144 52368 49156
rect 51859 49116 52368 49144
rect 51859 49113 51871 49116
rect 51813 49107 51871 49113
rect 52362 49104 52368 49116
rect 52420 49104 52426 49156
rect 32769 49079 32827 49085
rect 32769 49045 32781 49079
rect 32815 49076 32827 49079
rect 32858 49076 32864 49088
rect 32815 49048 32864 49076
rect 32815 49045 32827 49048
rect 32769 49039 32827 49045
rect 32858 49036 32864 49048
rect 32916 49036 32922 49088
rect 33321 49079 33379 49085
rect 33321 49045 33333 49079
rect 33367 49076 33379 49079
rect 33502 49076 33508 49088
rect 33367 49048 33508 49076
rect 33367 49045 33379 49048
rect 33321 49039 33379 49045
rect 33502 49036 33508 49048
rect 33560 49036 33566 49088
rect 52454 49036 52460 49088
rect 52512 49076 52518 49088
rect 52825 49079 52883 49085
rect 52825 49076 52837 49079
rect 52512 49048 52837 49076
rect 52512 49036 52518 49048
rect 52825 49045 52837 49048
rect 52871 49045 52883 49079
rect 52825 49039 52883 49045
rect 1104 48986 54832 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 54832 48986
rect 1104 48912 54832 48934
rect 52178 48832 52184 48884
rect 52236 48872 52242 48884
rect 52917 48875 52975 48881
rect 52917 48872 52929 48875
rect 52236 48844 52929 48872
rect 52236 48832 52242 48844
rect 52917 48841 52929 48844
rect 52963 48841 52975 48875
rect 52917 48835 52975 48841
rect 51169 48807 51227 48813
rect 51169 48773 51181 48807
rect 51215 48804 51227 48807
rect 53466 48804 53472 48816
rect 51215 48776 53472 48804
rect 51215 48773 51227 48776
rect 51169 48767 51227 48773
rect 53466 48764 53472 48776
rect 53524 48764 53530 48816
rect 52362 48736 52368 48748
rect 52323 48708 52368 48736
rect 52362 48696 52368 48708
rect 52420 48696 52426 48748
rect 53745 48739 53803 48745
rect 53745 48736 53757 48739
rect 52472 48708 53757 48736
rect 2133 48671 2191 48677
rect 2133 48637 2145 48671
rect 2179 48668 2191 48671
rect 2222 48668 2228 48680
rect 2179 48640 2228 48668
rect 2179 48637 2191 48640
rect 2133 48631 2191 48637
rect 2222 48628 2228 48640
rect 2280 48628 2286 48680
rect 2409 48671 2467 48677
rect 2409 48637 2421 48671
rect 2455 48668 2467 48671
rect 2774 48668 2780 48680
rect 2455 48640 2780 48668
rect 2455 48637 2467 48640
rect 2409 48631 2467 48637
rect 2774 48628 2780 48640
rect 2832 48668 2838 48680
rect 2869 48671 2927 48677
rect 2869 48668 2881 48671
rect 2832 48640 2881 48668
rect 2832 48628 2838 48640
rect 2869 48637 2881 48640
rect 2915 48637 2927 48671
rect 2869 48631 2927 48637
rect 38746 48628 38752 48680
rect 38804 48668 38810 48680
rect 52472 48668 52500 48708
rect 53745 48705 53757 48708
rect 53791 48705 53803 48739
rect 53745 48699 53803 48705
rect 53466 48668 53472 48680
rect 38804 48640 52500 48668
rect 53427 48640 53472 48668
rect 38804 48628 38810 48640
rect 53466 48628 53472 48640
rect 53524 48628 53530 48680
rect 32858 48560 32864 48612
rect 32916 48600 32922 48612
rect 52181 48603 52239 48609
rect 52181 48600 52193 48603
rect 32916 48572 33272 48600
rect 32916 48560 32922 48572
rect 33244 48544 33272 48572
rect 45526 48572 52193 48600
rect 2130 48492 2136 48544
rect 2188 48532 2194 48544
rect 32769 48535 32827 48541
rect 32769 48532 32781 48535
rect 2188 48504 32781 48532
rect 2188 48492 2194 48504
rect 32769 48501 32781 48504
rect 32815 48532 32827 48535
rect 33134 48532 33140 48544
rect 32815 48504 33140 48532
rect 32815 48501 32827 48504
rect 32769 48495 32827 48501
rect 33134 48492 33140 48504
rect 33192 48492 33198 48544
rect 33226 48492 33232 48544
rect 33284 48532 33290 48544
rect 33873 48535 33931 48541
rect 33284 48504 33329 48532
rect 33284 48492 33290 48504
rect 33873 48501 33885 48535
rect 33919 48532 33931 48535
rect 34054 48532 34060 48544
rect 33919 48504 34060 48532
rect 33919 48501 33931 48504
rect 33873 48495 33931 48501
rect 34054 48492 34060 48504
rect 34112 48492 34118 48544
rect 34422 48532 34428 48544
rect 34383 48504 34428 48532
rect 34422 48492 34428 48504
rect 34480 48492 34486 48544
rect 35618 48492 35624 48544
rect 35676 48532 35682 48544
rect 45526 48532 45554 48572
rect 52181 48569 52193 48572
rect 52227 48569 52239 48603
rect 52181 48563 52239 48569
rect 35676 48504 45554 48532
rect 35676 48492 35682 48504
rect 51258 48492 51264 48544
rect 51316 48532 51322 48544
rect 51629 48535 51687 48541
rect 51629 48532 51641 48535
rect 51316 48504 51641 48532
rect 51316 48492 51322 48504
rect 51629 48501 51641 48504
rect 51675 48501 51687 48535
rect 51629 48495 51687 48501
rect 1104 48442 54832 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 54832 48442
rect 1104 48368 54832 48390
rect 31110 48220 31116 48272
rect 31168 48260 31174 48272
rect 32309 48263 32367 48269
rect 32309 48260 32321 48263
rect 31168 48232 32321 48260
rect 31168 48220 31174 48232
rect 32309 48229 32321 48232
rect 32355 48229 32367 48263
rect 32309 48223 32367 48229
rect 33410 48220 33416 48272
rect 33468 48260 33474 48272
rect 38838 48260 38844 48272
rect 33468 48232 38844 48260
rect 33468 48220 33474 48232
rect 38838 48220 38844 48232
rect 38896 48220 38902 48272
rect 51258 48220 51264 48272
rect 51316 48260 51322 48272
rect 51316 48232 53696 48260
rect 51316 48220 51322 48232
rect 34149 48195 34207 48201
rect 34149 48192 34161 48195
rect 31726 48164 34161 48192
rect 2133 48127 2191 48133
rect 2133 48093 2145 48127
rect 2179 48093 2191 48127
rect 2133 48087 2191 48093
rect 2409 48127 2467 48133
rect 2409 48093 2421 48127
rect 2455 48124 2467 48127
rect 2774 48124 2780 48136
rect 2455 48096 2780 48124
rect 2455 48093 2467 48096
rect 2409 48087 2467 48093
rect 2148 48056 2176 48087
rect 2774 48084 2780 48096
rect 2832 48124 2838 48136
rect 2869 48127 2927 48133
rect 2869 48124 2881 48127
rect 2832 48096 2881 48124
rect 2832 48084 2838 48096
rect 2869 48093 2881 48096
rect 2915 48093 2927 48127
rect 2869 48087 2927 48093
rect 30466 48056 30472 48068
rect 2148 48028 30472 48056
rect 30466 48016 30472 48028
rect 30524 48016 30530 48068
rect 2682 47948 2688 48000
rect 2740 47988 2746 48000
rect 31726 47988 31754 48164
rect 33152 48133 33180 48164
rect 34149 48161 34161 48164
rect 34195 48161 34207 48195
rect 34149 48155 34207 48161
rect 52822 48152 52828 48204
rect 52880 48192 52886 48204
rect 52880 48164 53512 48192
rect 52880 48152 52886 48164
rect 33045 48127 33103 48133
rect 33045 48093 33057 48127
rect 33091 48093 33103 48127
rect 33045 48087 33103 48093
rect 33138 48127 33196 48133
rect 33138 48093 33150 48127
rect 33184 48093 33196 48127
rect 33410 48124 33416 48136
rect 33371 48096 33416 48124
rect 33138 48087 33196 48093
rect 31846 47988 31852 48000
rect 2740 47960 31754 47988
rect 31807 47960 31852 47988
rect 2740 47948 2746 47960
rect 31846 47948 31852 47960
rect 31904 47948 31910 48000
rect 33060 47988 33088 48087
rect 33410 48084 33416 48096
rect 33468 48084 33474 48136
rect 33502 48084 33508 48136
rect 33560 48133 33566 48136
rect 33560 48127 33609 48133
rect 33560 48093 33563 48127
rect 33597 48124 33609 48127
rect 33962 48124 33968 48136
rect 33597 48096 33968 48124
rect 33597 48093 33609 48096
rect 33560 48087 33609 48093
rect 33560 48084 33566 48087
rect 33962 48084 33968 48096
rect 34020 48084 34026 48136
rect 35529 48127 35587 48133
rect 35529 48093 35541 48127
rect 35575 48124 35587 48127
rect 51810 48124 51816 48136
rect 35575 48096 51816 48124
rect 35575 48093 35587 48096
rect 35529 48087 35587 48093
rect 33226 48016 33232 48068
rect 33284 48056 33290 48068
rect 33321 48059 33379 48065
rect 33321 48056 33333 48059
rect 33284 48028 33333 48056
rect 33284 48016 33290 48028
rect 33321 48025 33333 48028
rect 33367 48025 33379 48059
rect 35544 48056 35572 48087
rect 51810 48084 51816 48096
rect 51868 48084 51874 48136
rect 52178 48124 52184 48136
rect 52139 48096 52184 48124
rect 52178 48084 52184 48096
rect 52236 48084 52242 48136
rect 52638 48124 52644 48136
rect 52599 48096 52644 48124
rect 52638 48084 52644 48096
rect 52696 48084 52702 48136
rect 53484 48133 53512 48164
rect 53668 48133 53696 48232
rect 53285 48127 53343 48133
rect 53285 48093 53297 48127
rect 53331 48093 53343 48127
rect 53285 48087 53343 48093
rect 53469 48127 53527 48133
rect 53469 48093 53481 48127
rect 53515 48093 53527 48127
rect 53469 48087 53527 48093
rect 53653 48127 53711 48133
rect 53653 48093 53665 48127
rect 53699 48093 53711 48127
rect 53653 48087 53711 48093
rect 33321 48019 33379 48025
rect 33520 48028 35572 48056
rect 33520 47988 33548 48028
rect 51350 48016 51356 48068
rect 51408 48056 51414 48068
rect 53300 48056 53328 48087
rect 51408 48028 53328 48056
rect 53561 48059 53619 48065
rect 51408 48016 51414 48028
rect 53561 48025 53573 48059
rect 53607 48025 53619 48059
rect 53561 48019 53619 48025
rect 33060 47960 33548 47988
rect 33689 47991 33747 47997
rect 33689 47957 33701 47991
rect 33735 47988 33747 47991
rect 34146 47988 34152 48000
rect 33735 47960 34152 47988
rect 33735 47957 33747 47960
rect 33689 47951 33747 47957
rect 34146 47948 34152 47960
rect 34204 47948 34210 48000
rect 34882 47988 34888 48000
rect 34843 47960 34888 47988
rect 34882 47948 34888 47960
rect 34940 47948 34946 48000
rect 50985 47991 51043 47997
rect 50985 47957 50997 47991
rect 51031 47988 51043 47991
rect 51258 47988 51264 48000
rect 51031 47960 51264 47988
rect 51031 47957 51043 47960
rect 50985 47951 51043 47957
rect 51258 47948 51264 47960
rect 51316 47948 51322 48000
rect 51537 47991 51595 47997
rect 51537 47957 51549 47991
rect 51583 47988 51595 47991
rect 51626 47988 51632 48000
rect 51583 47960 51632 47988
rect 51583 47957 51595 47960
rect 51537 47951 51595 47957
rect 51626 47948 51632 47960
rect 51684 47948 51690 48000
rect 51994 47988 52000 48000
rect 51955 47960 52000 47988
rect 51994 47948 52000 47960
rect 52052 47948 52058 48000
rect 52825 47991 52883 47997
rect 52825 47957 52837 47991
rect 52871 47988 52883 47991
rect 53006 47988 53012 48000
rect 52871 47960 53012 47988
rect 52871 47957 52883 47960
rect 52825 47951 52883 47957
rect 53006 47948 53012 47960
rect 53064 47948 53070 48000
rect 53190 47948 53196 48000
rect 53248 47988 53254 48000
rect 53576 47988 53604 48019
rect 53834 47988 53840 48000
rect 53248 47960 53604 47988
rect 53795 47960 53840 47988
rect 53248 47948 53254 47960
rect 53834 47948 53840 47960
rect 53892 47948 53898 48000
rect 1104 47898 54832 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 54832 47898
rect 1104 47824 54832 47846
rect 29638 47784 29644 47796
rect 29599 47756 29644 47784
rect 29638 47744 29644 47756
rect 29696 47784 29702 47796
rect 33318 47784 33324 47796
rect 29696 47756 33324 47784
rect 29696 47744 29702 47756
rect 33318 47744 33324 47756
rect 33376 47744 33382 47796
rect 35342 47784 35348 47796
rect 33428 47756 35348 47784
rect 32766 47676 32772 47728
rect 32824 47716 32830 47728
rect 33226 47716 33232 47728
rect 32824 47688 33232 47716
rect 32824 47676 32830 47688
rect 33226 47676 33232 47688
rect 33284 47716 33290 47728
rect 33428 47725 33456 47756
rect 35342 47744 35348 47756
rect 35400 47744 35406 47796
rect 35434 47744 35440 47796
rect 35492 47784 35498 47796
rect 51994 47784 52000 47796
rect 35492 47756 52000 47784
rect 35492 47744 35498 47756
rect 51994 47744 52000 47756
rect 52052 47744 52058 47796
rect 52086 47744 52092 47796
rect 52144 47784 52150 47796
rect 52144 47756 52224 47784
rect 52144 47744 52150 47756
rect 33413 47719 33471 47725
rect 33284 47688 33364 47716
rect 33284 47676 33290 47688
rect 2133 47651 2191 47657
rect 2133 47617 2145 47651
rect 2179 47648 2191 47651
rect 29086 47648 29092 47660
rect 2179 47620 29092 47648
rect 2179 47617 2191 47620
rect 2133 47611 2191 47617
rect 29086 47608 29092 47620
rect 29144 47608 29150 47660
rect 33045 47651 33103 47657
rect 33045 47617 33057 47651
rect 33091 47617 33103 47651
rect 33045 47611 33103 47617
rect 2409 47583 2467 47589
rect 2409 47549 2421 47583
rect 2455 47580 2467 47583
rect 2774 47580 2780 47592
rect 2455 47552 2780 47580
rect 2455 47549 2467 47552
rect 2409 47543 2467 47549
rect 2774 47540 2780 47552
rect 2832 47580 2838 47592
rect 2869 47583 2927 47589
rect 2869 47580 2881 47583
rect 2832 47552 2881 47580
rect 2832 47540 2838 47552
rect 2869 47549 2881 47552
rect 2915 47549 2927 47583
rect 33060 47580 33088 47611
rect 33134 47608 33140 47660
rect 33192 47648 33198 47660
rect 33336 47657 33364 47688
rect 33413 47685 33425 47719
rect 33459 47685 33471 47719
rect 33413 47679 33471 47685
rect 34425 47719 34483 47725
rect 34425 47685 34437 47719
rect 34471 47716 34483 47719
rect 38930 47716 38936 47728
rect 34471 47688 38936 47716
rect 34471 47685 34483 47688
rect 34425 47679 34483 47685
rect 38930 47676 38936 47688
rect 38988 47676 38994 47728
rect 50157 47719 50215 47725
rect 50157 47685 50169 47719
rect 50203 47716 50215 47719
rect 51718 47716 51724 47728
rect 50203 47688 51724 47716
rect 50203 47685 50215 47688
rect 50157 47679 50215 47685
rect 51718 47676 51724 47688
rect 51776 47676 51782 47728
rect 52196 47725 52224 47756
rect 52181 47719 52239 47725
rect 52181 47685 52193 47719
rect 52227 47716 52239 47719
rect 52822 47716 52828 47728
rect 52227 47688 52828 47716
rect 52227 47685 52239 47688
rect 52181 47679 52239 47685
rect 52822 47676 52828 47688
rect 52880 47716 52886 47728
rect 52917 47719 52975 47725
rect 52917 47716 52929 47719
rect 52880 47688 52929 47716
rect 52880 47676 52886 47688
rect 52917 47685 52929 47688
rect 52963 47685 52975 47719
rect 52917 47679 52975 47685
rect 33321 47651 33379 47657
rect 33192 47620 33237 47648
rect 33192 47608 33198 47620
rect 33321 47617 33333 47651
rect 33367 47617 33379 47651
rect 33502 47648 33508 47660
rect 33461 47620 33508 47648
rect 33321 47611 33379 47617
rect 33502 47608 33508 47620
rect 33560 47657 33566 47660
rect 33560 47651 33609 47657
rect 33560 47617 33563 47651
rect 33597 47648 33609 47651
rect 34054 47648 34060 47660
rect 33597 47620 34060 47648
rect 33597 47617 33609 47620
rect 33560 47611 33609 47617
rect 33560 47608 33566 47611
rect 34054 47608 34060 47620
rect 34112 47648 34118 47660
rect 34333 47651 34391 47657
rect 34333 47648 34345 47651
rect 34112 47620 34345 47648
rect 34112 47608 34118 47620
rect 34333 47617 34345 47620
rect 34379 47617 34391 47651
rect 34514 47648 34520 47660
rect 34475 47620 34520 47648
rect 34333 47611 34391 47617
rect 34514 47608 34520 47620
rect 34572 47608 34578 47660
rect 34701 47651 34759 47657
rect 34701 47617 34713 47651
rect 34747 47648 34759 47651
rect 50709 47651 50767 47657
rect 34747 47620 36400 47648
rect 34747 47617 34759 47620
rect 34701 47611 34759 47617
rect 33060 47552 33180 47580
rect 2869 47543 2927 47549
rect 2314 47472 2320 47524
rect 2372 47512 2378 47524
rect 32030 47512 32036 47524
rect 2372 47484 32036 47512
rect 2372 47472 2378 47484
rect 32030 47472 32036 47484
rect 32088 47512 32094 47524
rect 32309 47515 32367 47521
rect 32309 47512 32321 47515
rect 32088 47484 32321 47512
rect 32088 47472 32094 47484
rect 32309 47481 32321 47484
rect 32355 47481 32367 47515
rect 33152 47512 33180 47552
rect 33612 47552 35848 47580
rect 33612 47512 33640 47552
rect 33152 47484 33640 47512
rect 32309 47475 32367 47481
rect 33870 47472 33876 47524
rect 33928 47512 33934 47524
rect 34149 47515 34207 47521
rect 34149 47512 34161 47515
rect 33928 47484 34161 47512
rect 33928 47472 33934 47484
rect 34149 47481 34161 47484
rect 34195 47481 34207 47515
rect 34149 47475 34207 47481
rect 34238 47472 34244 47524
rect 34296 47512 34302 47524
rect 35434 47512 35440 47524
rect 34296 47484 35440 47512
rect 34296 47472 34302 47484
rect 35434 47472 35440 47484
rect 35492 47472 35498 47524
rect 35820 47456 35848 47552
rect 36372 47521 36400 47620
rect 50709 47617 50721 47651
rect 50755 47648 50767 47651
rect 51169 47651 51227 47657
rect 51169 47648 51181 47651
rect 50755 47620 51181 47648
rect 50755 47617 50767 47620
rect 50709 47611 50767 47617
rect 51169 47617 51181 47620
rect 51215 47648 51227 47651
rect 51442 47648 51448 47660
rect 51215 47620 51448 47648
rect 51215 47617 51227 47620
rect 51169 47611 51227 47617
rect 51442 47608 51448 47620
rect 51500 47608 51506 47660
rect 51973 47651 52031 47657
rect 51973 47617 51985 47651
rect 52019 47648 52031 47651
rect 52097 47651 52155 47657
rect 52019 47617 52040 47648
rect 51973 47611 52040 47617
rect 52097 47617 52109 47651
rect 52143 47648 52155 47651
rect 52143 47620 52224 47648
rect 52143 47617 52155 47620
rect 52097 47611 52155 47617
rect 51258 47540 51264 47592
rect 51316 47580 51322 47592
rect 52012 47580 52040 47611
rect 51316 47552 52040 47580
rect 52196 47580 52224 47620
rect 52270 47608 52276 47660
rect 52328 47648 52334 47660
rect 52365 47651 52423 47657
rect 52365 47648 52377 47651
rect 52328 47620 52377 47648
rect 52328 47608 52334 47620
rect 52365 47617 52377 47620
rect 52411 47617 52423 47651
rect 52365 47611 52423 47617
rect 53282 47580 53288 47592
rect 52196 47552 53288 47580
rect 51316 47540 51322 47552
rect 53282 47540 53288 47552
rect 53340 47540 53346 47592
rect 53469 47583 53527 47589
rect 53469 47549 53481 47583
rect 53515 47580 53527 47583
rect 53558 47580 53564 47592
rect 53515 47552 53564 47580
rect 53515 47549 53527 47552
rect 53469 47543 53527 47549
rect 53558 47540 53564 47552
rect 53616 47540 53622 47592
rect 53745 47583 53803 47589
rect 53745 47549 53757 47583
rect 53791 47549 53803 47583
rect 53745 47543 53803 47549
rect 36357 47515 36415 47521
rect 36357 47481 36369 47515
rect 36403 47512 36415 47515
rect 51166 47512 51172 47524
rect 36403 47484 51172 47512
rect 36403 47481 36415 47484
rect 36357 47475 36415 47481
rect 51166 47472 51172 47484
rect 51224 47472 51230 47524
rect 51350 47512 51356 47524
rect 51311 47484 51356 47512
rect 51350 47472 51356 47484
rect 51408 47472 51414 47524
rect 51810 47512 51816 47524
rect 51771 47484 51816 47512
rect 51810 47472 51816 47484
rect 51868 47472 51874 47524
rect 52730 47472 52736 47524
rect 52788 47512 52794 47524
rect 53760 47512 53788 47543
rect 52788 47484 53788 47512
rect 52788 47472 52794 47484
rect 28258 47404 28264 47456
rect 28316 47444 28322 47456
rect 30653 47447 30711 47453
rect 30653 47444 30665 47447
rect 28316 47416 30665 47444
rect 28316 47404 28322 47416
rect 30653 47413 30665 47416
rect 30699 47444 30711 47447
rect 31110 47444 31116 47456
rect 30699 47416 31116 47444
rect 30699 47413 30711 47416
rect 30653 47407 30711 47413
rect 31110 47404 31116 47416
rect 31168 47404 31174 47456
rect 31662 47444 31668 47456
rect 31575 47416 31668 47444
rect 31662 47404 31668 47416
rect 31720 47444 31726 47456
rect 32398 47444 32404 47456
rect 31720 47416 32404 47444
rect 31720 47404 31726 47416
rect 32398 47404 32404 47416
rect 32456 47404 32462 47456
rect 33686 47444 33692 47456
rect 33647 47416 33692 47444
rect 33686 47404 33692 47416
rect 33744 47404 33750 47456
rect 34054 47404 34060 47456
rect 34112 47444 34118 47456
rect 34882 47444 34888 47456
rect 34112 47416 34888 47444
rect 34112 47404 34118 47416
rect 34882 47404 34888 47416
rect 34940 47444 34946 47456
rect 35161 47447 35219 47453
rect 35161 47444 35173 47447
rect 34940 47416 35173 47444
rect 34940 47404 34946 47416
rect 35161 47413 35173 47416
rect 35207 47413 35219 47447
rect 35802 47444 35808 47456
rect 35763 47416 35808 47444
rect 35161 47407 35219 47413
rect 35802 47404 35808 47416
rect 35860 47404 35866 47456
rect 51718 47404 51724 47456
rect 51776 47444 51782 47456
rect 53558 47444 53564 47456
rect 51776 47416 53564 47444
rect 51776 47404 51782 47416
rect 53558 47404 53564 47416
rect 53616 47404 53622 47456
rect 1104 47354 54832 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 54832 47354
rect 1104 47280 54832 47302
rect 29086 47240 29092 47252
rect 29047 47212 29092 47240
rect 29086 47200 29092 47212
rect 29144 47200 29150 47252
rect 31846 47200 31852 47252
rect 31904 47240 31910 47252
rect 52457 47243 52515 47249
rect 52457 47240 52469 47243
rect 31904 47212 52469 47240
rect 31904 47200 31910 47212
rect 52457 47209 52469 47212
rect 52503 47209 52515 47243
rect 52457 47203 52515 47209
rect 2133 47107 2191 47113
rect 2133 47073 2145 47107
rect 2179 47104 2191 47107
rect 2682 47104 2688 47116
rect 2179 47076 2688 47104
rect 2179 47073 2191 47076
rect 2133 47067 2191 47073
rect 2682 47064 2688 47076
rect 2740 47064 2746 47116
rect 2409 47039 2467 47045
rect 2409 47005 2421 47039
rect 2455 47036 2467 47039
rect 2774 47036 2780 47048
rect 2455 47008 2780 47036
rect 2455 47005 2467 47008
rect 2409 46999 2467 47005
rect 2774 46996 2780 47008
rect 2832 47036 2838 47048
rect 2869 47039 2927 47045
rect 2869 47036 2881 47039
rect 2832 47008 2881 47036
rect 2832 46996 2838 47008
rect 2869 47005 2881 47008
rect 2915 47005 2927 47039
rect 29104 47036 29132 47200
rect 31294 47132 31300 47184
rect 31352 47172 31358 47184
rect 31481 47175 31539 47181
rect 31481 47172 31493 47175
rect 31352 47144 31493 47172
rect 31352 47132 31358 47144
rect 31481 47141 31493 47144
rect 31527 47141 31539 47175
rect 31481 47135 31539 47141
rect 29638 47064 29644 47116
rect 29696 47104 29702 47116
rect 31864 47104 31892 47200
rect 29696 47076 30236 47104
rect 29696 47064 29702 47076
rect 29825 47039 29883 47045
rect 29825 47036 29837 47039
rect 29104 47008 29837 47036
rect 2869 46999 2927 47005
rect 29825 47005 29837 47008
rect 29871 47005 29883 47039
rect 30098 47036 30104 47048
rect 30059 47008 30104 47036
rect 29825 46999 29883 47005
rect 30098 46996 30104 47008
rect 30156 46996 30162 47048
rect 30208 47045 30236 47076
rect 30852 47076 31892 47104
rect 31956 47144 33645 47172
rect 30852 47045 30880 47076
rect 30193 47039 30251 47045
rect 30193 47005 30205 47039
rect 30239 47005 30251 47039
rect 30193 46999 30251 47005
rect 30837 47039 30895 47045
rect 30837 47005 30849 47039
rect 30883 47005 30895 47039
rect 30837 46999 30895 47005
rect 30930 47039 30988 47045
rect 30930 47005 30942 47039
rect 30976 47005 30988 47039
rect 31202 47036 31208 47048
rect 31163 47008 31208 47036
rect 30930 46999 30988 47005
rect 30006 46968 30012 46980
rect 29967 46940 30012 46968
rect 30006 46928 30012 46940
rect 30064 46928 30070 46980
rect 30466 46928 30472 46980
rect 30524 46968 30530 46980
rect 30944 46968 30972 46999
rect 31202 46996 31208 47008
rect 31260 46996 31266 47048
rect 31343 47039 31401 47045
rect 31343 47005 31355 47039
rect 31389 47036 31401 47039
rect 31662 47036 31668 47048
rect 31389 47008 31668 47036
rect 31389 47005 31401 47008
rect 31343 46999 31401 47005
rect 31662 46996 31668 47008
rect 31720 46996 31726 47048
rect 31956 47045 31984 47144
rect 32582 47104 32588 47116
rect 32324 47076 32588 47104
rect 31941 47039 31999 47045
rect 31941 47005 31953 47039
rect 31987 47005 31999 47039
rect 31941 46999 31999 47005
rect 32030 46996 32036 47048
rect 32088 47036 32094 47048
rect 32324 47045 32352 47076
rect 32582 47064 32588 47076
rect 32640 47064 32646 47116
rect 33502 47104 33508 47116
rect 32973 47076 33508 47104
rect 32309 47039 32367 47045
rect 32088 47008 32133 47036
rect 32088 46996 32094 47008
rect 32309 47005 32321 47039
rect 32355 47005 32367 47039
rect 32309 46999 32367 47005
rect 32398 46996 32404 47048
rect 32456 47045 32462 47048
rect 32456 47039 32505 47045
rect 32456 47005 32459 47039
rect 32493 47036 32505 47039
rect 32973 47036 33001 47076
rect 33502 47064 33508 47076
rect 33560 47064 33566 47116
rect 33617 47104 33645 47144
rect 33778 47132 33784 47184
rect 33836 47172 33842 47184
rect 33836 47144 33881 47172
rect 33836 47132 33842 47144
rect 35802 47132 35808 47184
rect 35860 47172 35866 47184
rect 51445 47175 51503 47181
rect 51445 47172 51457 47175
rect 35860 47144 51457 47172
rect 35860 47132 35866 47144
rect 51445 47141 51457 47144
rect 51491 47141 51503 47175
rect 51445 47135 51503 47141
rect 51534 47132 51540 47184
rect 51592 47172 51598 47184
rect 53650 47172 53656 47184
rect 51592 47144 53656 47172
rect 51592 47132 51598 47144
rect 53650 47132 53656 47144
rect 53708 47132 53714 47184
rect 34977 47107 35035 47113
rect 34977 47104 34989 47107
rect 33617 47076 34989 47104
rect 34977 47073 34989 47076
rect 35023 47104 35035 47107
rect 53834 47104 53840 47116
rect 35023 47076 53840 47104
rect 35023 47073 35035 47076
rect 34977 47067 35035 47073
rect 53834 47064 53840 47076
rect 53892 47064 53898 47116
rect 33134 47036 33140 47048
rect 32493 47008 33001 47036
rect 33095 47008 33140 47036
rect 32493 47005 32505 47008
rect 32456 46999 32505 47005
rect 32456 46996 32462 46999
rect 33134 46996 33140 47008
rect 33192 46996 33198 47048
rect 33318 47045 33324 47048
rect 33285 47039 33324 47045
rect 33285 47005 33297 47039
rect 33285 46999 33324 47005
rect 33318 46996 33324 46999
rect 33376 46996 33382 47048
rect 33643 47039 33701 47045
rect 33643 47005 33655 47039
rect 33689 47036 33701 47039
rect 34054 47036 34060 47048
rect 33689 47008 34060 47036
rect 33689 47005 33701 47008
rect 33643 46999 33701 47005
rect 34054 46996 34060 47008
rect 34112 47036 34118 47048
rect 34333 47039 34391 47045
rect 34333 47036 34345 47039
rect 34112 47008 34345 47036
rect 34112 46996 34118 47008
rect 34333 47005 34345 47008
rect 34379 47036 34391 47039
rect 34422 47036 34428 47048
rect 34379 47008 34428 47036
rect 34379 47005 34391 47008
rect 34333 46999 34391 47005
rect 34422 46996 34428 47008
rect 34480 46996 34486 47048
rect 48222 46996 48228 47048
rect 48280 47036 48286 47048
rect 50890 47036 50896 47048
rect 48280 47008 50896 47036
rect 48280 46996 48286 47008
rect 50890 46996 50896 47008
rect 50948 46996 50954 47048
rect 51605 47039 51663 47045
rect 51605 47005 51617 47039
rect 51651 47036 51663 47039
rect 51902 47036 51908 47048
rect 51651 47005 51672 47036
rect 51605 46999 51672 47005
rect 31110 46968 31116 46980
rect 30524 46940 30972 46968
rect 31071 46940 31116 46968
rect 30524 46928 30530 46940
rect 31110 46928 31116 46940
rect 31168 46968 31174 46980
rect 32217 46971 32275 46977
rect 32217 46968 32229 46971
rect 31168 46940 32229 46968
rect 31168 46928 31174 46940
rect 32217 46937 32229 46940
rect 32263 46937 32275 46971
rect 33413 46971 33471 46977
rect 32217 46931 32275 46937
rect 32600 46940 33272 46968
rect 30377 46903 30435 46909
rect 30377 46869 30389 46903
rect 30423 46900 30435 46903
rect 30926 46900 30932 46912
rect 30423 46872 30932 46900
rect 30423 46869 30435 46872
rect 30377 46863 30435 46869
rect 30926 46860 30932 46872
rect 30984 46860 30990 46912
rect 32600 46909 32628 46940
rect 33244 46912 33272 46940
rect 33413 46937 33425 46971
rect 33459 46937 33471 46971
rect 33413 46931 33471 46937
rect 33505 46971 33563 46977
rect 33505 46937 33517 46971
rect 33551 46968 33563 46971
rect 34698 46968 34704 46980
rect 33551 46940 34704 46968
rect 33551 46937 33563 46940
rect 33505 46931 33563 46937
rect 32585 46903 32643 46909
rect 32585 46869 32597 46903
rect 32631 46869 32643 46903
rect 32585 46863 32643 46869
rect 33226 46860 33232 46912
rect 33284 46860 33290 46912
rect 33428 46900 33456 46931
rect 34698 46928 34704 46940
rect 34756 46928 34762 46980
rect 49789 46971 49847 46977
rect 49789 46937 49801 46971
rect 49835 46968 49847 46971
rect 51442 46968 51448 46980
rect 49835 46940 51448 46968
rect 49835 46937 49847 46940
rect 49789 46931 49847 46937
rect 51442 46928 51448 46940
rect 51500 46928 51506 46980
rect 33594 46900 33600 46912
rect 33428 46872 33600 46900
rect 33594 46860 33600 46872
rect 33652 46900 33658 46912
rect 34514 46900 34520 46912
rect 33652 46872 34520 46900
rect 33652 46860 33658 46872
rect 34514 46860 34520 46872
rect 34572 46900 34578 46912
rect 35437 46903 35495 46909
rect 35437 46900 35449 46903
rect 34572 46872 35449 46900
rect 34572 46860 34578 46872
rect 35437 46869 35449 46872
rect 35483 46869 35495 46903
rect 35437 46863 35495 46869
rect 50433 46903 50491 46909
rect 50433 46869 50445 46903
rect 50479 46900 50491 46903
rect 51258 46900 51264 46912
rect 50479 46872 51264 46900
rect 50479 46869 50491 46872
rect 50433 46863 50491 46869
rect 51258 46860 51264 46872
rect 51316 46900 51322 46912
rect 51644 46900 51672 46999
rect 51736 47008 51908 47036
rect 51736 46977 51764 47008
rect 51902 46996 51908 47008
rect 51960 46996 51966 47048
rect 51997 47039 52055 47045
rect 51997 47005 52009 47039
rect 52043 47036 52055 47039
rect 52454 47036 52460 47048
rect 52043 47008 52460 47036
rect 52043 47005 52055 47008
rect 51997 46999 52055 47005
rect 52454 46996 52460 47008
rect 52512 46996 52518 47048
rect 52641 47039 52699 47045
rect 52641 47005 52653 47039
rect 52687 47005 52699 47039
rect 52822 47036 52828 47048
rect 52783 47008 52828 47036
rect 52641 46999 52699 47005
rect 51721 46971 51779 46977
rect 51721 46937 51733 46971
rect 51767 46937 51779 46971
rect 51721 46931 51779 46937
rect 51810 46928 51816 46980
rect 51868 46968 51874 46980
rect 52086 46968 52092 46980
rect 51868 46940 52092 46968
rect 51868 46928 51874 46940
rect 52086 46928 52092 46940
rect 52144 46928 52150 46980
rect 52656 46900 52684 46999
rect 52822 46996 52828 47008
rect 52880 46996 52886 47048
rect 53006 47036 53012 47048
rect 52967 47008 53012 47036
rect 53006 46996 53012 47008
rect 53064 46996 53070 47048
rect 53469 47039 53527 47045
rect 53469 47005 53481 47039
rect 53515 47036 53527 47039
rect 53650 47036 53656 47048
rect 53515 47008 53656 47036
rect 53515 47005 53527 47008
rect 53469 46999 53527 47005
rect 53650 46996 53656 47008
rect 53708 46996 53714 47048
rect 53745 47039 53803 47045
rect 53745 47005 53757 47039
rect 53791 47005 53803 47039
rect 53745 46999 53803 47005
rect 52733 46971 52791 46977
rect 52733 46937 52745 46971
rect 52779 46937 52791 46971
rect 52733 46931 52791 46937
rect 51316 46872 52684 46900
rect 52748 46900 52776 46931
rect 52914 46928 52920 46980
rect 52972 46968 52978 46980
rect 53760 46968 53788 46999
rect 54110 46968 54116 46980
rect 52972 46940 53788 46968
rect 53852 46940 54116 46968
rect 52972 46928 52978 46940
rect 53852 46900 53880 46940
rect 54110 46928 54116 46940
rect 54168 46928 54174 46980
rect 52748 46872 53880 46900
rect 51316 46860 51322 46872
rect 1104 46810 54832 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 54832 46810
rect 1104 46736 54832 46758
rect 30466 46696 30472 46708
rect 30427 46668 30472 46696
rect 30466 46656 30472 46668
rect 30524 46656 30530 46708
rect 34238 46696 34244 46708
rect 33888 46668 34244 46696
rect 29457 46631 29515 46637
rect 29457 46597 29469 46631
rect 29503 46628 29515 46631
rect 30006 46628 30012 46640
rect 29503 46600 30012 46628
rect 29503 46597 29515 46600
rect 29457 46591 29515 46597
rect 30006 46588 30012 46600
rect 30064 46628 30070 46640
rect 32766 46628 32772 46640
rect 30064 46600 32772 46628
rect 30064 46588 30070 46600
rect 2133 46563 2191 46569
rect 2133 46529 2145 46563
rect 2179 46560 2191 46563
rect 2590 46560 2596 46572
rect 2179 46532 2596 46560
rect 2179 46529 2191 46532
rect 2133 46523 2191 46529
rect 2590 46520 2596 46532
rect 2648 46520 2654 46572
rect 32508 46569 32536 46600
rect 32766 46588 32772 46600
rect 32824 46588 32830 46640
rect 32493 46563 32551 46569
rect 32493 46529 32505 46563
rect 32539 46529 32551 46563
rect 32493 46523 32551 46529
rect 32585 46563 32643 46569
rect 32585 46529 32597 46563
rect 32631 46529 32643 46563
rect 32585 46523 32643 46529
rect 32677 46563 32735 46569
rect 32677 46529 32689 46563
rect 32723 46529 32735 46563
rect 32677 46523 32735 46529
rect 32861 46563 32919 46569
rect 32861 46529 32873 46563
rect 32907 46560 32919 46563
rect 33318 46560 33324 46572
rect 32907 46532 33324 46560
rect 32907 46529 32919 46532
rect 32861 46523 32919 46529
rect 2409 46495 2467 46501
rect 2409 46461 2421 46495
rect 2455 46492 2467 46495
rect 2774 46492 2780 46504
rect 2455 46464 2780 46492
rect 2455 46461 2467 46464
rect 2409 46455 2467 46461
rect 2774 46452 2780 46464
rect 2832 46492 2838 46504
rect 2869 46495 2927 46501
rect 2869 46492 2881 46495
rect 2832 46464 2881 46492
rect 2832 46452 2838 46464
rect 2869 46461 2881 46464
rect 2915 46461 2927 46495
rect 32600 46492 32628 46523
rect 2869 46455 2927 46461
rect 32140 46464 32628 46492
rect 32692 46492 32720 46523
rect 33318 46520 33324 46532
rect 33376 46560 33382 46572
rect 33888 46560 33916 46668
rect 34238 46656 34244 46668
rect 34296 46656 34302 46708
rect 34330 46656 34336 46708
rect 34388 46656 34394 46708
rect 34057 46631 34115 46637
rect 34057 46597 34069 46631
rect 34103 46628 34115 46631
rect 34348 46628 34376 46656
rect 34103 46600 34376 46628
rect 34103 46597 34115 46600
rect 34057 46591 34115 46597
rect 47026 46588 47032 46640
rect 47084 46628 47090 46640
rect 47084 46600 53788 46628
rect 47084 46588 47090 46600
rect 33376 46532 33916 46560
rect 33376 46520 33382 46532
rect 33962 46520 33968 46572
rect 34020 46560 34026 46572
rect 34149 46563 34207 46569
rect 34020 46532 34065 46560
rect 34020 46520 34026 46532
rect 34149 46529 34161 46563
rect 34195 46560 34207 46563
rect 34238 46560 34244 46572
rect 34195 46532 34244 46560
rect 34195 46529 34207 46532
rect 34149 46523 34207 46529
rect 34164 46492 34192 46523
rect 34238 46520 34244 46532
rect 34296 46520 34302 46572
rect 53760 46569 53788 46600
rect 34333 46563 34391 46569
rect 34333 46529 34345 46563
rect 34379 46560 34391 46563
rect 50525 46563 50583 46569
rect 34379 46532 35480 46560
rect 34379 46529 34391 46532
rect 34333 46523 34391 46529
rect 32692 46464 34192 46492
rect 2222 46384 2228 46436
rect 2280 46424 2286 46436
rect 31665 46427 31723 46433
rect 31665 46424 31677 46427
rect 2280 46396 31677 46424
rect 2280 46384 2286 46396
rect 31665 46393 31677 46396
rect 31711 46424 31723 46427
rect 32140 46424 32168 46464
rect 32692 46424 32720 46464
rect 31711 46396 32168 46424
rect 32232 46396 32720 46424
rect 31711 46393 31723 46396
rect 31665 46387 31723 46393
rect 31202 46356 31208 46368
rect 31115 46328 31208 46356
rect 31202 46316 31208 46328
rect 31260 46356 31266 46368
rect 32232 46356 32260 46396
rect 33962 46384 33968 46436
rect 34020 46424 34026 46436
rect 34793 46427 34851 46433
rect 34793 46424 34805 46427
rect 34020 46396 34805 46424
rect 34020 46384 34026 46396
rect 34793 46393 34805 46396
rect 34839 46393 34851 46427
rect 34793 46387 34851 46393
rect 31260 46328 32260 46356
rect 32309 46359 32367 46365
rect 31260 46316 31266 46328
rect 32309 46325 32321 46359
rect 32355 46356 32367 46359
rect 33042 46356 33048 46368
rect 32355 46328 33048 46356
rect 32355 46325 32367 46328
rect 32309 46319 32367 46325
rect 33042 46316 33048 46328
rect 33100 46316 33106 46368
rect 33410 46316 33416 46368
rect 33468 46356 33474 46368
rect 35452 46365 35480 46532
rect 50525 46529 50537 46563
rect 50571 46560 50583 46563
rect 53745 46563 53803 46569
rect 50571 46532 53512 46560
rect 50571 46529 50583 46532
rect 50525 46523 50583 46529
rect 53484 46504 53512 46532
rect 53745 46529 53757 46563
rect 53791 46529 53803 46563
rect 53745 46523 53803 46529
rect 51074 46452 51080 46504
rect 51132 46492 51138 46504
rect 52089 46495 52147 46501
rect 52089 46492 52101 46495
rect 51132 46464 52101 46492
rect 51132 46452 51138 46464
rect 52089 46461 52101 46464
rect 52135 46461 52147 46495
rect 52089 46455 52147 46461
rect 52365 46495 52423 46501
rect 52365 46461 52377 46495
rect 52411 46492 52423 46495
rect 53466 46492 53472 46504
rect 52411 46464 53052 46492
rect 53427 46464 53472 46492
rect 52411 46461 52423 46464
rect 52365 46455 52423 46461
rect 53024 46368 53052 46464
rect 53466 46452 53472 46464
rect 53524 46452 53530 46504
rect 33781 46359 33839 46365
rect 33781 46356 33793 46359
rect 33468 46328 33793 46356
rect 33468 46316 33474 46328
rect 33781 46325 33793 46328
rect 33827 46325 33839 46359
rect 33781 46319 33839 46325
rect 35437 46359 35495 46365
rect 35437 46325 35449 46359
rect 35483 46356 35495 46359
rect 48130 46356 48136 46368
rect 35483 46328 48136 46356
rect 35483 46325 35495 46328
rect 35437 46319 35495 46325
rect 48130 46316 48136 46328
rect 48188 46316 48194 46368
rect 51077 46359 51135 46365
rect 51077 46325 51089 46359
rect 51123 46356 51135 46359
rect 51258 46356 51264 46368
rect 51123 46328 51264 46356
rect 51123 46325 51135 46328
rect 51077 46319 51135 46325
rect 51258 46316 51264 46328
rect 51316 46316 51322 46368
rect 53006 46356 53012 46368
rect 52967 46328 53012 46356
rect 53006 46316 53012 46328
rect 53064 46316 53070 46368
rect 1104 46266 54832 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 54832 46266
rect 1104 46192 54832 46214
rect 32953 46155 33011 46161
rect 32953 46121 32965 46155
rect 32999 46152 33011 46155
rect 33134 46152 33140 46164
rect 32999 46124 33140 46152
rect 32999 46121 33011 46124
rect 32953 46115 33011 46121
rect 33134 46112 33140 46124
rect 33192 46112 33198 46164
rect 34977 46155 35035 46161
rect 34977 46121 34989 46155
rect 35023 46152 35035 46155
rect 35618 46152 35624 46164
rect 35023 46124 35624 46152
rect 35023 46121 35035 46124
rect 34977 46115 35035 46121
rect 35618 46112 35624 46124
rect 35676 46112 35682 46164
rect 2406 46044 2412 46096
rect 2464 46084 2470 46096
rect 31386 46084 31392 46096
rect 2464 46056 6914 46084
rect 31299 46056 31392 46084
rect 2464 46044 2470 46056
rect 6886 46016 6914 46056
rect 31386 46044 31392 46056
rect 31444 46084 31450 46096
rect 34057 46087 34115 46093
rect 31444 46056 32352 46084
rect 31444 46044 31450 46056
rect 31849 46019 31907 46025
rect 31849 46016 31861 46019
rect 6886 45988 31861 46016
rect 31849 45985 31861 45988
rect 31895 45985 31907 46019
rect 32324 46016 32352 46056
rect 34057 46053 34069 46087
rect 34103 46084 34115 46087
rect 34238 46084 34244 46096
rect 34103 46056 34244 46084
rect 34103 46053 34115 46056
rect 34057 46047 34115 46053
rect 34238 46044 34244 46056
rect 34296 46084 34302 46096
rect 34296 46056 41414 46084
rect 34296 46044 34302 46056
rect 32324 45988 38654 46016
rect 31849 45979 31907 45985
rect 2133 45951 2191 45957
rect 2133 45917 2145 45951
rect 2179 45948 2191 45951
rect 2314 45948 2320 45960
rect 2179 45920 2320 45948
rect 2179 45917 2191 45920
rect 2133 45911 2191 45917
rect 2314 45908 2320 45920
rect 2372 45908 2378 45960
rect 2409 45951 2467 45957
rect 2409 45917 2421 45951
rect 2455 45948 2467 45951
rect 2774 45948 2780 45960
rect 2455 45920 2780 45948
rect 2455 45917 2467 45920
rect 2409 45911 2467 45917
rect 2774 45908 2780 45920
rect 2832 45948 2838 45960
rect 2869 45951 2927 45957
rect 2869 45948 2881 45951
rect 2832 45920 2881 45948
rect 2832 45908 2838 45920
rect 2869 45917 2881 45920
rect 2915 45917 2927 45951
rect 2869 45911 2927 45917
rect 26786 45840 26792 45892
rect 26844 45880 26850 45892
rect 31386 45880 31392 45892
rect 26844 45852 31392 45880
rect 26844 45840 26850 45852
rect 31386 45840 31392 45852
rect 31444 45840 31450 45892
rect 31864 45880 31892 45979
rect 32398 45948 32404 45960
rect 32359 45920 32404 45948
rect 32398 45908 32404 45920
rect 32456 45908 32462 45960
rect 32600 45957 32628 45988
rect 32585 45951 32643 45957
rect 32585 45917 32597 45951
rect 32631 45917 32643 45951
rect 32766 45948 32772 45960
rect 32727 45920 32772 45948
rect 32585 45911 32643 45917
rect 32766 45908 32772 45920
rect 32824 45908 32830 45960
rect 32677 45883 32735 45889
rect 32677 45880 32689 45883
rect 31864 45852 32689 45880
rect 32677 45849 32689 45852
rect 32723 45849 32735 45883
rect 38626 45880 38654 45988
rect 41386 45948 41414 46056
rect 52638 45976 52644 46028
rect 52696 46016 52702 46028
rect 53745 46019 53803 46025
rect 53745 46016 53757 46019
rect 52696 45988 53757 46016
rect 52696 45976 52702 45988
rect 53745 45985 53757 45988
rect 53791 45985 53803 46019
rect 53745 45979 53803 45985
rect 48222 45948 48228 45960
rect 41386 45920 48228 45948
rect 48222 45908 48228 45920
rect 48280 45908 48286 45960
rect 51721 45951 51779 45957
rect 51721 45917 51733 45951
rect 51767 45948 51779 45951
rect 52178 45948 52184 45960
rect 51767 45920 52184 45948
rect 51767 45917 51779 45920
rect 51721 45911 51779 45917
rect 52178 45908 52184 45920
rect 52236 45908 52242 45960
rect 52457 45951 52515 45957
rect 52457 45917 52469 45951
rect 52503 45948 52515 45951
rect 52546 45948 52552 45960
rect 52503 45920 52552 45948
rect 52503 45917 52515 45920
rect 52457 45911 52515 45917
rect 52546 45908 52552 45920
rect 52604 45908 52610 45960
rect 53374 45908 53380 45960
rect 53432 45948 53438 45960
rect 53469 45951 53527 45957
rect 53469 45948 53481 45951
rect 53432 45920 53481 45948
rect 53432 45908 53438 45920
rect 53469 45917 53481 45920
rect 53515 45917 53527 45951
rect 53469 45911 53527 45917
rect 51169 45883 51227 45889
rect 38626 45852 48314 45880
rect 32677 45843 32735 45849
rect 32398 45772 32404 45824
rect 32456 45812 32462 45824
rect 33502 45812 33508 45824
rect 32456 45784 33508 45812
rect 32456 45772 32462 45784
rect 33502 45772 33508 45784
rect 33560 45772 33566 45824
rect 48286 45812 48314 45852
rect 51169 45849 51181 45883
rect 51215 45880 51227 45883
rect 53392 45880 53420 45908
rect 51215 45852 53420 45880
rect 51215 45849 51227 45852
rect 51169 45843 51227 45849
rect 51258 45812 51264 45824
rect 48286 45784 51264 45812
rect 51258 45772 51264 45784
rect 51316 45772 51322 45824
rect 1104 45722 54832 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 54832 45722
rect 1104 45648 54832 45670
rect 33502 45568 33508 45620
rect 33560 45608 33566 45620
rect 51166 45608 51172 45620
rect 33560 45580 51172 45608
rect 33560 45568 33566 45580
rect 51166 45568 51172 45580
rect 51224 45568 51230 45620
rect 26418 45500 26424 45552
rect 26476 45540 26482 45552
rect 29638 45540 29644 45552
rect 26476 45512 29644 45540
rect 26476 45500 26482 45512
rect 29638 45500 29644 45512
rect 29696 45500 29702 45552
rect 33318 45500 33324 45552
rect 33376 45540 33382 45552
rect 33413 45543 33471 45549
rect 33413 45540 33425 45543
rect 33376 45512 33425 45540
rect 33376 45500 33382 45512
rect 33413 45509 33425 45512
rect 33459 45509 33471 45543
rect 33413 45503 33471 45509
rect 51077 45475 51135 45481
rect 51077 45441 51089 45475
rect 51123 45472 51135 45475
rect 53742 45472 53748 45484
rect 51123 45444 53512 45472
rect 53703 45444 53748 45472
rect 51123 45441 51135 45444
rect 51077 45435 51135 45441
rect 2133 45407 2191 45413
rect 2133 45373 2145 45407
rect 2179 45373 2191 45407
rect 2133 45367 2191 45373
rect 2409 45407 2467 45413
rect 2409 45373 2421 45407
rect 2455 45404 2467 45407
rect 2774 45404 2780 45416
rect 2455 45376 2780 45404
rect 2455 45373 2467 45376
rect 2409 45367 2467 45373
rect 2148 45336 2176 45367
rect 2774 45364 2780 45376
rect 2832 45404 2838 45416
rect 2869 45407 2927 45413
rect 2869 45404 2881 45407
rect 2832 45376 2881 45404
rect 2832 45364 2838 45376
rect 2869 45373 2881 45376
rect 2915 45373 2927 45407
rect 2869 45367 2927 45373
rect 28534 45364 28540 45416
rect 28592 45404 28598 45416
rect 53484 45413 53512 45444
rect 53742 45432 53748 45444
rect 53800 45432 53806 45484
rect 52089 45407 52147 45413
rect 52089 45404 52101 45407
rect 28592 45376 52101 45404
rect 28592 45364 28598 45376
rect 52089 45373 52101 45376
rect 52135 45373 52147 45407
rect 52089 45367 52147 45373
rect 52365 45407 52423 45413
rect 52365 45373 52377 45407
rect 52411 45404 52423 45407
rect 53469 45407 53527 45413
rect 52411 45376 53052 45404
rect 52411 45373 52423 45376
rect 52365 45367 52423 45373
rect 22186 45336 22192 45348
rect 2148 45308 22192 45336
rect 22186 45296 22192 45308
rect 22244 45296 22250 45348
rect 53024 45280 53052 45376
rect 53469 45373 53481 45407
rect 53515 45404 53527 45407
rect 53558 45404 53564 45416
rect 53515 45376 53564 45404
rect 53515 45373 53527 45376
rect 53469 45367 53527 45373
rect 53558 45364 53564 45376
rect 53616 45364 53622 45416
rect 31846 45228 31852 45280
rect 31904 45268 31910 45280
rect 32309 45271 32367 45277
rect 32309 45268 32321 45271
rect 31904 45240 32321 45268
rect 31904 45228 31910 45240
rect 32309 45237 32321 45240
rect 32355 45268 32367 45271
rect 32766 45268 32772 45280
rect 32355 45240 32772 45268
rect 32355 45237 32367 45240
rect 32309 45231 32367 45237
rect 32766 45228 32772 45240
rect 32824 45268 32830 45280
rect 32861 45271 32919 45277
rect 32861 45268 32873 45271
rect 32824 45240 32873 45268
rect 32824 45228 32830 45240
rect 32861 45237 32873 45240
rect 32907 45237 32919 45271
rect 53006 45268 53012 45280
rect 52967 45240 53012 45268
rect 32861 45231 32919 45237
rect 53006 45228 53012 45240
rect 53064 45228 53070 45280
rect 1104 45178 54832 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 54832 45178
rect 1104 45104 54832 45126
rect 27430 45064 27436 45076
rect 27343 45036 27436 45064
rect 27430 45024 27436 45036
rect 27488 45064 27494 45076
rect 28077 45067 28135 45073
rect 28077 45064 28089 45067
rect 27488 45036 28089 45064
rect 27488 45024 27494 45036
rect 28077 45033 28089 45036
rect 28123 45064 28135 45067
rect 31202 45064 31208 45076
rect 28123 45036 31208 45064
rect 28123 45033 28135 45036
rect 28077 45027 28135 45033
rect 31202 45024 31208 45036
rect 31260 45024 31266 45076
rect 28626 44956 28632 45008
rect 28684 44996 28690 45008
rect 52914 44996 52920 45008
rect 28684 44968 52920 44996
rect 28684 44956 28690 44968
rect 52914 44956 52920 44968
rect 52972 44956 52978 45008
rect 52454 44928 52460 44940
rect 52415 44900 52460 44928
rect 52454 44888 52460 44900
rect 52512 44888 52518 44940
rect 2133 44863 2191 44869
rect 2133 44829 2145 44863
rect 2179 44829 2191 44863
rect 2133 44823 2191 44829
rect 2409 44863 2467 44869
rect 2409 44829 2421 44863
rect 2455 44860 2467 44863
rect 2774 44860 2780 44872
rect 2455 44832 2780 44860
rect 2455 44829 2467 44832
rect 2409 44823 2467 44829
rect 2148 44792 2176 44823
rect 2774 44820 2780 44832
rect 2832 44860 2838 44872
rect 2869 44863 2927 44869
rect 2869 44860 2881 44863
rect 2832 44832 2881 44860
rect 2832 44820 2838 44832
rect 2869 44829 2881 44832
rect 2915 44829 2927 44863
rect 2869 44823 2927 44829
rect 28350 44820 28356 44872
rect 28408 44860 28414 44872
rect 47026 44860 47032 44872
rect 28408 44832 47032 44860
rect 28408 44820 28414 44832
rect 47026 44820 47032 44832
rect 47084 44820 47090 44872
rect 51721 44863 51779 44869
rect 51721 44829 51733 44863
rect 51767 44860 51779 44863
rect 52178 44860 52184 44872
rect 51767 44832 52184 44860
rect 51767 44829 51779 44832
rect 51721 44823 51779 44829
rect 52178 44820 52184 44832
rect 52236 44820 52242 44872
rect 53469 44863 53527 44869
rect 53469 44829 53481 44863
rect 53515 44860 53527 44863
rect 53650 44860 53656 44872
rect 53515 44832 53656 44860
rect 53515 44829 53527 44832
rect 53469 44823 53527 44829
rect 22922 44792 22928 44804
rect 2148 44764 22928 44792
rect 22922 44752 22928 44764
rect 22980 44752 22986 44804
rect 51169 44795 51227 44801
rect 51169 44761 51181 44795
rect 51215 44792 51227 44795
rect 53484 44792 53512 44823
rect 53650 44820 53656 44832
rect 53708 44820 53714 44872
rect 53742 44820 53748 44872
rect 53800 44860 53806 44872
rect 53800 44832 53845 44860
rect 53800 44820 53806 44832
rect 51215 44764 53512 44792
rect 51215 44761 51227 44764
rect 51169 44755 51227 44761
rect 26878 44724 26884 44736
rect 26839 44696 26884 44724
rect 26878 44684 26884 44696
rect 26936 44684 26942 44736
rect 1104 44634 54832 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 54832 44634
rect 1104 44560 54832 44582
rect 28626 44520 28632 44532
rect 28587 44492 28632 44520
rect 28626 44480 28632 44492
rect 28684 44480 28690 44532
rect 51077 44523 51135 44529
rect 51077 44489 51089 44523
rect 51123 44520 51135 44523
rect 53466 44520 53472 44532
rect 51123 44492 53472 44520
rect 51123 44489 51135 44492
rect 51077 44483 51135 44489
rect 53466 44480 53472 44492
rect 53524 44480 53530 44532
rect 22278 44412 22284 44464
rect 22336 44452 22342 44464
rect 26237 44455 26295 44461
rect 26237 44452 26249 44455
rect 22336 44424 26249 44452
rect 22336 44412 22342 44424
rect 26237 44421 26249 44424
rect 26283 44421 26295 44455
rect 26237 44415 26295 44421
rect 26329 44455 26387 44461
rect 26329 44421 26341 44455
rect 26375 44452 26387 44455
rect 27062 44452 27068 44464
rect 26375 44424 27068 44452
rect 26375 44421 26387 44424
rect 26329 44415 26387 44421
rect 27062 44412 27068 44424
rect 27120 44452 27126 44464
rect 27430 44452 27436 44464
rect 27120 44424 27436 44452
rect 27120 44412 27126 44424
rect 27430 44412 27436 44424
rect 27488 44412 27494 44464
rect 52638 44452 52644 44464
rect 31726 44424 52644 44452
rect 25501 44387 25559 44393
rect 25501 44353 25513 44387
rect 25547 44384 25559 44387
rect 26145 44387 26203 44393
rect 26145 44384 26157 44387
rect 25547 44356 26157 44384
rect 25547 44353 25559 44356
rect 25501 44347 25559 44353
rect 26145 44353 26157 44356
rect 26191 44384 26203 44387
rect 26418 44384 26424 44396
rect 26191 44356 26424 44384
rect 26191 44353 26203 44356
rect 26145 44347 26203 44353
rect 26418 44344 26424 44356
rect 26476 44344 26482 44396
rect 26513 44387 26571 44393
rect 26513 44353 26525 44387
rect 26559 44384 26571 44387
rect 26878 44384 26884 44396
rect 26559 44356 26884 44384
rect 26559 44353 26571 44356
rect 26513 44347 26571 44353
rect 26878 44344 26884 44356
rect 26936 44384 26942 44396
rect 31726 44384 31754 44424
rect 52638 44412 52644 44424
rect 52696 44412 52702 44464
rect 26936 44356 31754 44384
rect 26936 44344 26942 44356
rect 53098 44344 53104 44396
rect 53156 44384 53162 44396
rect 53745 44387 53803 44393
rect 53745 44384 53757 44387
rect 53156 44356 53757 44384
rect 53156 44344 53162 44356
rect 53745 44353 53757 44356
rect 53791 44353 53803 44387
rect 53745 44347 53803 44353
rect 2133 44319 2191 44325
rect 2133 44285 2145 44319
rect 2179 44316 2191 44319
rect 2222 44316 2228 44328
rect 2179 44288 2228 44316
rect 2179 44285 2191 44288
rect 2133 44279 2191 44285
rect 2222 44276 2228 44288
rect 2280 44276 2286 44328
rect 2409 44319 2467 44325
rect 2409 44285 2421 44319
rect 2455 44316 2467 44319
rect 2774 44316 2780 44328
rect 2455 44288 2780 44316
rect 2455 44285 2467 44288
rect 2409 44279 2467 44285
rect 2774 44276 2780 44288
rect 2832 44316 2838 44328
rect 2869 44319 2927 44325
rect 2869 44316 2881 44319
rect 2832 44288 2881 44316
rect 2832 44276 2838 44288
rect 2869 44285 2881 44288
rect 2915 44285 2927 44319
rect 2869 44279 2927 44285
rect 10410 44276 10416 44328
rect 10468 44316 10474 44328
rect 27157 44319 27215 44325
rect 27157 44316 27169 44319
rect 10468 44288 27169 44316
rect 10468 44276 10474 44288
rect 27157 44285 27169 44288
rect 27203 44316 27215 44319
rect 27798 44316 27804 44328
rect 27203 44288 27804 44316
rect 27203 44285 27215 44288
rect 27157 44279 27215 44285
rect 27798 44276 27804 44288
rect 27856 44276 27862 44328
rect 52086 44316 52092 44328
rect 52047 44288 52092 44316
rect 52086 44276 52092 44288
rect 52144 44276 52150 44328
rect 52365 44319 52423 44325
rect 52365 44285 52377 44319
rect 52411 44316 52423 44319
rect 53466 44316 53472 44328
rect 52411 44288 53052 44316
rect 53427 44288 53472 44316
rect 52411 44285 52423 44288
rect 52365 44279 52423 44285
rect 24762 44208 24768 44260
rect 24820 44248 24826 44260
rect 25961 44251 26019 44257
rect 25961 44248 25973 44251
rect 24820 44220 25973 44248
rect 24820 44208 24826 44220
rect 25961 44217 25973 44220
rect 26007 44217 26019 44251
rect 32306 44248 32312 44260
rect 32267 44220 32312 44248
rect 25961 44211 26019 44217
rect 32306 44208 32312 44220
rect 32364 44208 32370 44260
rect 53024 44192 53052 44288
rect 53466 44276 53472 44288
rect 53524 44276 53530 44328
rect 27982 44180 27988 44192
rect 27943 44152 27988 44180
rect 27982 44140 27988 44152
rect 28040 44140 28046 44192
rect 30469 44183 30527 44189
rect 30469 44149 30481 44183
rect 30515 44180 30527 44183
rect 30834 44180 30840 44192
rect 30515 44152 30840 44180
rect 30515 44149 30527 44152
rect 30469 44143 30527 44149
rect 30834 44140 30840 44152
rect 30892 44140 30898 44192
rect 31018 44180 31024 44192
rect 30979 44152 31024 44180
rect 31018 44140 31024 44152
rect 31076 44140 31082 44192
rect 32766 44140 32772 44192
rect 32824 44180 32830 44192
rect 32861 44183 32919 44189
rect 32861 44180 32873 44183
rect 32824 44152 32873 44180
rect 32824 44140 32830 44152
rect 32861 44149 32873 44152
rect 32907 44149 32919 44183
rect 53006 44180 53012 44192
rect 52967 44152 53012 44180
rect 32861 44143 32919 44149
rect 53006 44140 53012 44152
rect 53064 44140 53070 44192
rect 1104 44090 54832 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 54832 44090
rect 1104 44016 54832 44038
rect 32950 43936 32956 43988
rect 33008 43976 33014 43988
rect 34149 43979 34207 43985
rect 34149 43976 34161 43979
rect 33008 43948 34161 43976
rect 33008 43936 33014 43948
rect 34149 43945 34161 43948
rect 34195 43945 34207 43979
rect 34149 43939 34207 43945
rect 12802 43868 12808 43920
rect 12860 43908 12866 43920
rect 29733 43911 29791 43917
rect 29733 43908 29745 43911
rect 12860 43880 29745 43908
rect 12860 43868 12866 43880
rect 29733 43877 29745 43880
rect 29779 43908 29791 43911
rect 30006 43908 30012 43920
rect 29779 43880 30012 43908
rect 29779 43877 29791 43880
rect 29733 43871 29791 43877
rect 30006 43868 30012 43880
rect 30064 43868 30070 43920
rect 51350 43868 51356 43920
rect 51408 43908 51414 43920
rect 53742 43908 53748 43920
rect 51408 43880 53748 43908
rect 51408 43868 51414 43880
rect 53742 43868 53748 43880
rect 53800 43868 53806 43920
rect 2314 43800 2320 43852
rect 2372 43840 2378 43852
rect 25961 43843 26019 43849
rect 25961 43840 25973 43843
rect 2372 43812 25973 43840
rect 2372 43800 2378 43812
rect 25961 43809 25973 43812
rect 26007 43840 26019 43843
rect 28626 43840 28632 43852
rect 26007 43812 27384 43840
rect 26007 43809 26019 43812
rect 25961 43803 26019 43809
rect 2130 43772 2136 43784
rect 2091 43744 2136 43772
rect 2130 43732 2136 43744
rect 2188 43732 2194 43784
rect 2409 43775 2467 43781
rect 2409 43741 2421 43775
rect 2455 43772 2467 43775
rect 2774 43772 2780 43784
rect 2455 43744 2780 43772
rect 2455 43741 2467 43744
rect 2409 43735 2467 43741
rect 2774 43732 2780 43744
rect 2832 43772 2838 43784
rect 27356 43781 27384 43812
rect 27632 43812 28632 43840
rect 2869 43775 2927 43781
rect 2869 43772 2881 43775
rect 2832 43744 2881 43772
rect 2832 43732 2838 43744
rect 2869 43741 2881 43744
rect 2915 43741 2927 43775
rect 27203 43775 27261 43781
rect 27203 43772 27215 43775
rect 2869 43735 2927 43741
rect 26528 43744 27215 43772
rect 25314 43596 25320 43648
rect 25372 43636 25378 43648
rect 26528 43645 26556 43744
rect 27203 43741 27215 43744
rect 27249 43741 27261 43775
rect 27203 43735 27261 43741
rect 27341 43775 27399 43781
rect 27341 43741 27353 43775
rect 27387 43741 27399 43775
rect 27341 43735 27399 43741
rect 27430 43732 27436 43784
rect 27488 43772 27494 43784
rect 27632 43781 27660 43812
rect 28626 43800 28632 43812
rect 28684 43800 28690 43852
rect 52730 43840 52736 43852
rect 31726 43812 52736 43840
rect 27616 43775 27674 43781
rect 27488 43744 27533 43772
rect 27488 43732 27494 43744
rect 27616 43741 27628 43775
rect 27662 43741 27674 43775
rect 27616 43735 27674 43741
rect 27709 43775 27767 43781
rect 27709 43741 27721 43775
rect 27755 43741 27767 43775
rect 27709 43735 27767 43741
rect 27724 43704 27752 43735
rect 28074 43732 28080 43784
rect 28132 43772 28138 43784
rect 28537 43775 28595 43781
rect 28537 43772 28549 43775
rect 28132 43744 28549 43772
rect 28132 43732 28138 43744
rect 28537 43741 28549 43744
rect 28583 43772 28595 43775
rect 31726 43772 31754 43812
rect 52730 43800 52736 43812
rect 52788 43800 52794 43852
rect 28583 43744 31754 43772
rect 51721 43775 51779 43781
rect 28583 43741 28595 43744
rect 28537 43735 28595 43741
rect 51721 43741 51733 43775
rect 51767 43772 51779 43775
rect 53469 43775 53527 43781
rect 53469 43772 53481 43775
rect 51767 43744 53481 43772
rect 51767 43741 51779 43744
rect 51721 43735 51779 43741
rect 53469 43741 53481 43744
rect 53515 43741 53527 43775
rect 53469 43735 53527 43741
rect 28902 43704 28908 43716
rect 27724 43676 28908 43704
rect 28902 43664 28908 43676
rect 28960 43664 28966 43716
rect 30466 43664 30472 43716
rect 30524 43704 30530 43716
rect 31481 43707 31539 43713
rect 31481 43704 31493 43707
rect 30524 43676 31493 43704
rect 30524 43664 30530 43676
rect 31481 43673 31493 43676
rect 31527 43704 31539 43707
rect 52273 43707 52331 43713
rect 31527 43676 45554 43704
rect 31527 43673 31539 43676
rect 31481 43667 31539 43673
rect 26513 43639 26571 43645
rect 26513 43636 26525 43639
rect 25372 43608 26525 43636
rect 25372 43596 25378 43608
rect 26513 43605 26525 43608
rect 26559 43605 26571 43639
rect 26513 43599 26571 43605
rect 26602 43596 26608 43648
rect 26660 43636 26666 43648
rect 27065 43639 27123 43645
rect 27065 43636 27077 43639
rect 26660 43608 27077 43636
rect 26660 43596 26666 43608
rect 27065 43605 27077 43608
rect 27111 43605 27123 43639
rect 28994 43636 29000 43648
rect 28955 43608 29000 43636
rect 27065 43599 27123 43605
rect 28994 43596 29000 43608
rect 29052 43596 29058 43648
rect 30377 43639 30435 43645
rect 30377 43605 30389 43639
rect 30423 43636 30435 43639
rect 30558 43636 30564 43648
rect 30423 43608 30564 43636
rect 30423 43605 30435 43608
rect 30377 43599 30435 43605
rect 30558 43596 30564 43608
rect 30616 43636 30622 43648
rect 30837 43639 30895 43645
rect 30837 43636 30849 43639
rect 30616 43608 30849 43636
rect 30616 43596 30622 43608
rect 30837 43605 30849 43608
rect 30883 43605 30895 43639
rect 31938 43636 31944 43648
rect 31899 43608 31944 43636
rect 30837 43599 30895 43605
rect 31938 43596 31944 43608
rect 31996 43596 32002 43648
rect 32585 43639 32643 43645
rect 32585 43605 32597 43639
rect 32631 43636 32643 43639
rect 32674 43636 32680 43648
rect 32631 43608 32680 43636
rect 32631 43605 32643 43608
rect 32585 43599 32643 43605
rect 32674 43596 32680 43608
rect 32732 43596 32738 43648
rect 32766 43596 32772 43648
rect 32824 43636 32830 43648
rect 33137 43639 33195 43645
rect 33137 43636 33149 43639
rect 32824 43608 33149 43636
rect 32824 43596 32830 43608
rect 33137 43605 33149 43608
rect 33183 43605 33195 43639
rect 33137 43599 33195 43605
rect 33594 43596 33600 43648
rect 33652 43636 33658 43648
rect 33689 43639 33747 43645
rect 33689 43636 33701 43639
rect 33652 43608 33701 43636
rect 33652 43596 33658 43608
rect 33689 43605 33701 43608
rect 33735 43636 33747 43639
rect 33962 43636 33968 43648
rect 33735 43608 33968 43636
rect 33735 43605 33747 43608
rect 33689 43599 33747 43605
rect 33962 43596 33968 43608
rect 34020 43596 34026 43648
rect 45526 43636 45554 43676
rect 52273 43673 52285 43707
rect 52319 43704 52331 43707
rect 52914 43704 52920 43716
rect 52319 43676 52920 43704
rect 52319 43673 52331 43676
rect 52273 43667 52331 43673
rect 52914 43664 52920 43676
rect 52972 43664 52978 43716
rect 52546 43636 52552 43648
rect 45526 43608 52552 43636
rect 52546 43596 52552 43608
rect 52604 43596 52610 43648
rect 52822 43636 52828 43648
rect 52783 43608 52828 43636
rect 52822 43596 52828 43608
rect 52880 43596 52886 43648
rect 53484 43636 53512 43735
rect 53558 43732 53564 43784
rect 53616 43772 53622 43784
rect 53745 43775 53803 43781
rect 53745 43772 53757 43775
rect 53616 43744 53757 43772
rect 53616 43732 53622 43744
rect 53745 43741 53757 43744
rect 53791 43741 53803 43775
rect 53745 43735 53803 43741
rect 53742 43636 53748 43648
rect 53484 43608 53748 43636
rect 53742 43596 53748 43608
rect 53800 43596 53806 43648
rect 1104 43546 54832 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 54832 43546
rect 1104 43472 54832 43494
rect 32674 43432 32680 43444
rect 22066 43404 32680 43432
rect 1854 43324 1860 43376
rect 1912 43364 1918 43376
rect 22066 43364 22094 43404
rect 32674 43392 32680 43404
rect 32732 43392 32738 43444
rect 34606 43432 34612 43444
rect 34567 43404 34612 43432
rect 34606 43392 34612 43404
rect 34664 43392 34670 43444
rect 52086 43432 52092 43444
rect 41386 43404 52092 43432
rect 25406 43364 25412 43376
rect 1912 43336 22094 43364
rect 25367 43336 25412 43364
rect 1912 43324 1918 43336
rect 25406 43324 25412 43336
rect 25464 43324 25470 43376
rect 26050 43364 26056 43376
rect 26011 43336 26056 43364
rect 26050 43324 26056 43336
rect 26108 43324 26114 43376
rect 26605 43367 26663 43373
rect 26605 43333 26617 43367
rect 26651 43364 26663 43367
rect 26786 43364 26792 43376
rect 26651 43336 26792 43364
rect 26651 43333 26663 43336
rect 26605 43327 26663 43333
rect 26786 43324 26792 43336
rect 26844 43364 26850 43376
rect 27246 43364 27252 43376
rect 26844 43336 27252 43364
rect 26844 43324 26850 43336
rect 27246 43324 27252 43336
rect 27304 43324 27310 43376
rect 28258 43364 28264 43376
rect 28219 43336 28264 43364
rect 28258 43324 28264 43336
rect 28316 43324 28322 43376
rect 29178 43324 29184 43376
rect 29236 43364 29242 43376
rect 41386 43364 41414 43404
rect 52086 43392 52092 43404
rect 52144 43392 52150 43444
rect 29236 43336 41414 43364
rect 29236 43324 29242 43336
rect 2133 43299 2191 43305
rect 2133 43265 2145 43299
rect 2179 43296 2191 43299
rect 2498 43296 2504 43308
rect 2179 43268 2504 43296
rect 2179 43265 2191 43268
rect 2133 43259 2191 43265
rect 2498 43256 2504 43268
rect 2556 43256 2562 43308
rect 2682 43256 2688 43308
rect 2740 43296 2746 43308
rect 28994 43296 29000 43308
rect 2740 43268 29000 43296
rect 2740 43256 2746 43268
rect 28994 43256 29000 43268
rect 29052 43256 29058 43308
rect 32030 43256 32036 43308
rect 32088 43296 32094 43308
rect 32582 43296 32588 43308
rect 32088 43268 32588 43296
rect 32088 43256 32094 43268
rect 32582 43256 32588 43268
rect 32640 43296 32646 43308
rect 32861 43299 32919 43305
rect 32861 43296 32873 43299
rect 32640 43268 32873 43296
rect 32640 43256 32646 43268
rect 32861 43265 32873 43268
rect 32907 43265 32919 43299
rect 53558 43296 53564 43308
rect 32861 43259 32919 43265
rect 45526 43268 53564 43296
rect 2409 43231 2467 43237
rect 2409 43197 2421 43231
rect 2455 43228 2467 43231
rect 2774 43228 2780 43240
rect 2455 43200 2780 43228
rect 2455 43197 2467 43200
rect 2409 43191 2467 43197
rect 2774 43188 2780 43200
rect 2832 43228 2838 43240
rect 2869 43231 2927 43237
rect 2869 43228 2881 43231
rect 2832 43200 2881 43228
rect 2832 43188 2838 43200
rect 2869 43197 2881 43200
rect 2915 43197 2927 43231
rect 29638 43228 29644 43240
rect 29599 43200 29644 43228
rect 2869 43191 2927 43197
rect 29638 43188 29644 43200
rect 29696 43188 29702 43240
rect 32398 43228 32404 43240
rect 32311 43200 32404 43228
rect 32398 43188 32404 43200
rect 32456 43228 32462 43240
rect 45526 43228 45554 43268
rect 53558 43256 53564 43268
rect 53616 43256 53622 43308
rect 32456 43200 45554 43228
rect 52365 43231 52423 43237
rect 32456 43188 32462 43200
rect 52365 43197 52377 43231
rect 52411 43228 52423 43231
rect 53469 43231 53527 43237
rect 53469 43228 53481 43231
rect 52411 43200 53481 43228
rect 52411 43197 52423 43200
rect 52365 43191 52423 43197
rect 53469 43197 53481 43200
rect 53515 43228 53527 43231
rect 53650 43228 53656 43240
rect 53515 43200 53656 43228
rect 53515 43197 53527 43200
rect 53469 43191 53527 43197
rect 53650 43188 53656 43200
rect 53708 43188 53714 43240
rect 53745 43231 53803 43237
rect 53745 43197 53757 43231
rect 53791 43197 53803 43231
rect 53745 43191 53803 43197
rect 1762 43120 1768 43172
rect 1820 43160 1826 43172
rect 32582 43160 32588 43172
rect 1820 43132 32588 43160
rect 1820 43120 1826 43132
rect 32582 43120 32588 43132
rect 32640 43160 32646 43172
rect 33505 43163 33563 43169
rect 33505 43160 33517 43163
rect 32640 43132 33517 43160
rect 32640 43120 32646 43132
rect 33505 43129 33517 43132
rect 33551 43129 33563 43163
rect 33505 43123 33563 43129
rect 52638 43120 52644 43172
rect 52696 43160 52702 43172
rect 53760 43160 53788 43191
rect 52696 43132 53788 43160
rect 52696 43120 52702 43132
rect 27617 43095 27675 43101
rect 27617 43061 27629 43095
rect 27663 43092 27675 43095
rect 27706 43092 27712 43104
rect 27663 43064 27712 43092
rect 27663 43061 27675 43064
rect 27617 43055 27675 43061
rect 27706 43052 27712 43064
rect 27764 43092 27770 43104
rect 28442 43092 28448 43104
rect 27764 43064 28448 43092
rect 27764 43052 27770 43064
rect 28442 43052 28448 43064
rect 28500 43052 28506 43104
rect 29086 43092 29092 43104
rect 29047 43064 29092 43092
rect 29086 43052 29092 43064
rect 29144 43052 29150 43104
rect 30190 43092 30196 43104
rect 30151 43064 30196 43092
rect 30190 43052 30196 43064
rect 30248 43052 30254 43104
rect 30742 43092 30748 43104
rect 30703 43064 30748 43092
rect 30742 43052 30748 43064
rect 30800 43052 30806 43104
rect 31389 43095 31447 43101
rect 31389 43061 31401 43095
rect 31435 43092 31447 43095
rect 31478 43092 31484 43104
rect 31435 43064 31484 43092
rect 31435 43061 31447 43064
rect 31389 43055 31447 43061
rect 31478 43052 31484 43064
rect 31536 43052 31542 43104
rect 34057 43095 34115 43101
rect 34057 43061 34069 43095
rect 34103 43092 34115 43095
rect 34330 43092 34336 43104
rect 34103 43064 34336 43092
rect 34103 43061 34115 43064
rect 34057 43055 34115 43061
rect 34330 43052 34336 43064
rect 34388 43052 34394 43104
rect 35161 43095 35219 43101
rect 35161 43061 35173 43095
rect 35207 43092 35219 43095
rect 35434 43092 35440 43104
rect 35207 43064 35440 43092
rect 35207 43061 35219 43064
rect 35161 43055 35219 43061
rect 35434 43052 35440 43064
rect 35492 43052 35498 43104
rect 53009 43095 53067 43101
rect 53009 43061 53021 43095
rect 53055 43092 53067 43095
rect 53374 43092 53380 43104
rect 53055 43064 53380 43092
rect 53055 43061 53067 43064
rect 53009 43055 53067 43061
rect 53374 43052 53380 43064
rect 53432 43052 53438 43104
rect 1104 43002 54832 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 54832 43002
rect 1104 42928 54832 42950
rect 25593 42891 25651 42897
rect 25593 42857 25605 42891
rect 25639 42888 25651 42891
rect 26050 42888 26056 42900
rect 25639 42860 26056 42888
rect 25639 42857 25651 42860
rect 25593 42851 25651 42857
rect 26050 42848 26056 42860
rect 26108 42848 26114 42900
rect 30742 42848 30748 42900
rect 30800 42888 30806 42900
rect 52546 42888 52552 42900
rect 30800 42860 52552 42888
rect 30800 42848 30806 42860
rect 52546 42848 52552 42860
rect 52604 42848 52610 42900
rect 25774 42780 25780 42832
rect 25832 42820 25838 42832
rect 27157 42823 27215 42829
rect 27157 42820 27169 42823
rect 25832 42792 27169 42820
rect 25832 42780 25838 42792
rect 27157 42789 27169 42792
rect 27203 42789 27215 42823
rect 27157 42783 27215 42789
rect 27801 42823 27859 42829
rect 27801 42789 27813 42823
rect 27847 42820 27859 42823
rect 27890 42820 27896 42832
rect 27847 42792 27896 42820
rect 27847 42789 27859 42792
rect 27801 42783 27859 42789
rect 27890 42780 27896 42792
rect 27948 42820 27954 42832
rect 30558 42820 30564 42832
rect 27948 42792 30564 42820
rect 27948 42780 27954 42792
rect 30558 42780 30564 42792
rect 30616 42780 30622 42832
rect 2590 42712 2596 42764
rect 2648 42752 2654 42764
rect 25866 42752 25872 42764
rect 2648 42724 25872 42752
rect 2648 42712 2654 42724
rect 25866 42712 25872 42724
rect 25924 42712 25930 42764
rect 26145 42755 26203 42761
rect 26145 42721 26157 42755
rect 26191 42752 26203 42755
rect 26418 42752 26424 42764
rect 26191 42724 26424 42752
rect 26191 42721 26203 42724
rect 26145 42715 26203 42721
rect 26418 42712 26424 42724
rect 26476 42712 26482 42764
rect 28350 42752 28356 42764
rect 28311 42724 28356 42752
rect 28350 42712 28356 42724
rect 28408 42712 28414 42764
rect 29638 42712 29644 42764
rect 29696 42752 29702 42764
rect 30834 42752 30840 42764
rect 29696 42724 30840 42752
rect 29696 42712 29702 42724
rect 2133 42687 2191 42693
rect 2133 42653 2145 42687
rect 2179 42653 2191 42687
rect 2133 42647 2191 42653
rect 2409 42687 2467 42693
rect 2409 42653 2421 42687
rect 2455 42684 2467 42687
rect 2774 42684 2780 42696
rect 2455 42656 2780 42684
rect 2455 42653 2467 42656
rect 2409 42647 2467 42653
rect 2148 42616 2176 42647
rect 2774 42644 2780 42656
rect 2832 42684 2838 42696
rect 2869 42687 2927 42693
rect 2869 42684 2881 42687
rect 2832 42656 2881 42684
rect 2832 42644 2838 42656
rect 2869 42653 2881 42656
rect 2915 42653 2927 42687
rect 2869 42647 2927 42653
rect 23842 42644 23848 42696
rect 23900 42684 23906 42696
rect 26234 42684 26240 42696
rect 23900 42656 26240 42684
rect 23900 42644 23906 42656
rect 26234 42644 26240 42656
rect 26292 42644 26298 42696
rect 28442 42644 28448 42696
rect 28500 42684 28506 42696
rect 29932 42693 29960 42724
rect 30834 42712 30840 42724
rect 30892 42712 30898 42764
rect 32306 42712 32312 42764
rect 32364 42752 32370 42764
rect 35526 42752 35532 42764
rect 32364 42724 32628 42752
rect 32364 42712 32370 42724
rect 29181 42687 29239 42693
rect 29181 42684 29193 42687
rect 28500 42656 29193 42684
rect 28500 42644 28506 42656
rect 29181 42653 29193 42656
rect 29227 42684 29239 42687
rect 29917 42687 29975 42693
rect 29227 42656 29868 42684
rect 29227 42653 29239 42656
rect 29181 42647 29239 42653
rect 23382 42616 23388 42628
rect 2148 42588 23388 42616
rect 23382 42576 23388 42588
rect 23440 42576 23446 42628
rect 25041 42619 25099 42625
rect 25041 42585 25053 42619
rect 25087 42616 25099 42619
rect 26326 42616 26332 42628
rect 25087 42588 26332 42616
rect 25087 42585 25099 42588
rect 25041 42579 25099 42585
rect 26326 42576 26332 42588
rect 26384 42576 26390 42628
rect 26697 42619 26755 42625
rect 26697 42585 26709 42619
rect 26743 42616 26755 42619
rect 28258 42616 28264 42628
rect 26743 42588 28264 42616
rect 26743 42585 26755 42588
rect 26697 42579 26755 42585
rect 28258 42576 28264 42588
rect 28316 42616 28322 42628
rect 29454 42616 29460 42628
rect 28316 42588 29460 42616
rect 28316 42576 28322 42588
rect 29454 42576 29460 42588
rect 29512 42576 29518 42628
rect 29840 42616 29868 42656
rect 29917 42653 29929 42687
rect 29963 42653 29975 42687
rect 29917 42647 29975 42653
rect 30006 42644 30012 42696
rect 30064 42684 30070 42696
rect 30282 42684 30288 42696
rect 30064 42656 30109 42684
rect 30243 42656 30288 42684
rect 30064 42644 30070 42656
rect 30282 42644 30288 42656
rect 30340 42644 30346 42696
rect 32490 42684 32496 42696
rect 32451 42656 32496 42684
rect 32490 42644 32496 42656
rect 32548 42644 32554 42696
rect 32600 42693 32628 42724
rect 32973 42724 35532 42752
rect 32586 42687 32644 42693
rect 32586 42653 32598 42687
rect 32632 42653 32644 42687
rect 32858 42684 32864 42696
rect 32819 42656 32864 42684
rect 32586 42647 32644 42653
rect 32858 42644 32864 42656
rect 32916 42644 32922 42696
rect 32973 42693 33001 42724
rect 35526 42712 35532 42724
rect 35584 42712 35590 42764
rect 53742 42752 53748 42764
rect 53703 42724 53748 42752
rect 53742 42712 53748 42724
rect 53800 42712 53806 42764
rect 32958 42687 33016 42693
rect 32958 42653 32970 42687
rect 33004 42653 33016 42687
rect 32958 42647 33016 42653
rect 30101 42619 30159 42625
rect 30101 42616 30113 42619
rect 29840 42588 30113 42616
rect 30101 42585 30113 42588
rect 30147 42616 30159 42619
rect 31297 42619 31355 42625
rect 31297 42616 31309 42619
rect 30147 42588 31309 42616
rect 30147 42585 30159 42588
rect 30101 42579 30159 42585
rect 30300 42560 30328 42588
rect 31297 42585 31309 42588
rect 31343 42616 31355 42619
rect 31849 42619 31907 42625
rect 31849 42616 31861 42619
rect 31343 42588 31861 42616
rect 31343 42585 31355 42588
rect 31297 42579 31355 42585
rect 31849 42585 31861 42588
rect 31895 42585 31907 42619
rect 32766 42616 32772 42628
rect 32727 42588 32772 42616
rect 31849 42579 31907 42585
rect 32766 42576 32772 42588
rect 32824 42576 32830 42628
rect 26786 42508 26792 42560
rect 26844 42548 26850 42560
rect 27890 42548 27896 42560
rect 26844 42520 27896 42548
rect 26844 42508 26850 42520
rect 27890 42508 27896 42520
rect 27948 42508 27954 42560
rect 29546 42508 29552 42560
rect 29604 42548 29610 42560
rect 29733 42551 29791 42557
rect 29733 42548 29745 42551
rect 29604 42520 29745 42548
rect 29604 42508 29610 42520
rect 29733 42517 29745 42520
rect 29779 42517 29791 42551
rect 29733 42511 29791 42517
rect 30282 42508 30288 42560
rect 30340 42508 30346 42560
rect 30834 42548 30840 42560
rect 30747 42520 30840 42548
rect 30834 42508 30840 42520
rect 30892 42548 30898 42560
rect 31570 42548 31576 42560
rect 30892 42520 31576 42548
rect 30892 42508 30898 42520
rect 31570 42508 31576 42520
rect 31628 42548 31634 42560
rect 32973 42548 33001 42647
rect 33134 42644 33140 42696
rect 33192 42684 33198 42696
rect 33965 42687 34023 42693
rect 33965 42684 33977 42687
rect 33192 42656 33977 42684
rect 33192 42644 33198 42656
rect 33965 42653 33977 42656
rect 34011 42653 34023 42687
rect 33965 42647 34023 42653
rect 52362 42644 52368 42696
rect 52420 42684 52426 42696
rect 53009 42687 53067 42693
rect 53009 42684 53021 42687
rect 52420 42656 53021 42684
rect 52420 42644 52426 42656
rect 53009 42653 53021 42656
rect 53055 42653 53067 42687
rect 53466 42684 53472 42696
rect 53427 42656 53472 42684
rect 53009 42647 53067 42653
rect 53466 42644 53472 42656
rect 53524 42644 53530 42696
rect 33594 42616 33600 42628
rect 33555 42588 33600 42616
rect 33594 42576 33600 42588
rect 33652 42576 33658 42628
rect 33781 42619 33839 42625
rect 33781 42585 33793 42619
rect 33827 42616 33839 42619
rect 34054 42616 34060 42628
rect 33827 42588 34060 42616
rect 33827 42585 33839 42588
rect 33781 42579 33839 42585
rect 34054 42576 34060 42588
rect 34112 42576 34118 42628
rect 34238 42576 34244 42628
rect 34296 42616 34302 42628
rect 34790 42616 34796 42628
rect 34296 42588 34796 42616
rect 34296 42576 34302 42588
rect 34790 42576 34796 42588
rect 34848 42576 34854 42628
rect 51813 42619 51871 42625
rect 51813 42585 51825 42619
rect 51859 42616 51871 42619
rect 53484 42616 53512 42644
rect 51859 42588 53512 42616
rect 51859 42585 51871 42588
rect 51813 42579 51871 42585
rect 31628 42520 33001 42548
rect 33137 42551 33195 42557
rect 31628 42508 31634 42520
rect 33137 42517 33149 42551
rect 33183 42548 33195 42551
rect 33502 42548 33508 42560
rect 33183 42520 33508 42548
rect 33183 42517 33195 42520
rect 33137 42511 33195 42517
rect 33502 42508 33508 42520
rect 33560 42508 33566 42560
rect 33962 42508 33968 42560
rect 34020 42548 34026 42560
rect 34885 42551 34943 42557
rect 34885 42548 34897 42551
rect 34020 42520 34897 42548
rect 34020 42508 34026 42520
rect 34885 42517 34897 42520
rect 34931 42517 34943 42551
rect 35526 42548 35532 42560
rect 35487 42520 35532 42548
rect 34885 42511 34943 42517
rect 35526 42508 35532 42520
rect 35584 42508 35590 42560
rect 52362 42548 52368 42560
rect 52323 42520 52368 42548
rect 52362 42508 52368 42520
rect 52420 42508 52426 42560
rect 52454 42508 52460 42560
rect 52512 42548 52518 42560
rect 52825 42551 52883 42557
rect 52825 42548 52837 42551
rect 52512 42520 52837 42548
rect 52512 42508 52518 42520
rect 52825 42517 52837 42520
rect 52871 42517 52883 42551
rect 52825 42511 52883 42517
rect 1104 42458 54832 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 54832 42458
rect 1104 42384 54832 42406
rect 25406 42304 25412 42356
rect 25464 42344 25470 42356
rect 29178 42344 29184 42356
rect 25464 42316 26004 42344
rect 25464 42304 25470 42316
rect 25590 42276 25596 42288
rect 25148 42248 25596 42276
rect 24854 42208 24860 42220
rect 24815 42180 24860 42208
rect 24854 42168 24860 42180
rect 24912 42168 24918 42220
rect 25148 42217 25176 42248
rect 25590 42236 25596 42248
rect 25648 42236 25654 42288
rect 25976 42217 26004 42316
rect 26252 42316 29184 42344
rect 26050 42236 26056 42288
rect 26108 42276 26114 42288
rect 26252 42285 26280 42316
rect 29178 42304 29184 42316
rect 29236 42304 29242 42356
rect 29365 42347 29423 42353
rect 29365 42313 29377 42347
rect 29411 42344 29423 42347
rect 29454 42344 29460 42356
rect 29411 42316 29460 42344
rect 29411 42313 29423 42316
rect 29365 42307 29423 42313
rect 29454 42304 29460 42316
rect 29512 42304 29518 42356
rect 30282 42304 30288 42356
rect 30340 42344 30346 42356
rect 30340 42316 30512 42344
rect 30340 42304 30346 42316
rect 26145 42279 26203 42285
rect 26145 42276 26157 42279
rect 26108 42248 26157 42276
rect 26108 42236 26114 42248
rect 26145 42245 26157 42248
rect 26191 42245 26203 42279
rect 26145 42239 26203 42245
rect 26237 42279 26295 42285
rect 26237 42245 26249 42279
rect 26283 42245 26295 42279
rect 28994 42276 29000 42288
rect 26237 42239 26295 42245
rect 28552 42248 29000 42276
rect 24949 42211 25007 42217
rect 24949 42177 24961 42211
rect 24995 42177 25007 42211
rect 24949 42171 25007 42177
rect 25133 42211 25191 42217
rect 25133 42177 25145 42211
rect 25179 42177 25191 42211
rect 25133 42171 25191 42177
rect 25225 42211 25283 42217
rect 25225 42177 25237 42211
rect 25271 42177 25283 42211
rect 25225 42171 25283 42177
rect 25409 42211 25467 42217
rect 25409 42177 25421 42211
rect 25455 42208 25467 42211
rect 25869 42211 25927 42217
rect 25869 42208 25881 42211
rect 25455 42180 25881 42208
rect 25455 42177 25467 42180
rect 25409 42171 25467 42177
rect 25869 42177 25881 42180
rect 25915 42177 25927 42211
rect 25869 42171 25927 42177
rect 25962 42211 26020 42217
rect 25962 42177 25974 42211
rect 26008 42177 26020 42211
rect 25962 42171 26020 42177
rect 2133 42143 2191 42149
rect 2133 42109 2145 42143
rect 2179 42140 2191 42143
rect 2314 42140 2320 42152
rect 2179 42112 2320 42140
rect 2179 42109 2191 42112
rect 2133 42103 2191 42109
rect 2314 42100 2320 42112
rect 2372 42100 2378 42152
rect 2409 42143 2467 42149
rect 2409 42109 2421 42143
rect 2455 42140 2467 42143
rect 2774 42140 2780 42152
rect 2455 42112 2780 42140
rect 2455 42109 2467 42112
rect 2409 42103 2467 42109
rect 2774 42100 2780 42112
rect 2832 42140 2838 42152
rect 2869 42143 2927 42149
rect 2869 42140 2881 42143
rect 2832 42112 2881 42140
rect 2832 42100 2838 42112
rect 2869 42109 2881 42112
rect 2915 42109 2927 42143
rect 2869 42103 2927 42109
rect 24210 42100 24216 42152
rect 24268 42140 24274 42152
rect 24964 42140 24992 42171
rect 25240 42140 25268 42171
rect 24268 42112 24992 42140
rect 25148 42112 25268 42140
rect 24268 42100 24274 42112
rect 25148 42072 25176 42112
rect 23860 42044 25176 42072
rect 23860 42016 23888 42044
rect 23842 42004 23848 42016
rect 23803 41976 23848 42004
rect 23842 41964 23848 41976
rect 23900 41964 23906 42016
rect 24397 42007 24455 42013
rect 24397 41973 24409 42007
rect 24443 42004 24455 42007
rect 26252 42004 26280 42239
rect 26326 42168 26332 42220
rect 26384 42217 26390 42220
rect 26384 42211 26433 42217
rect 26384 42177 26387 42211
rect 26421 42208 26433 42211
rect 27706 42208 27712 42220
rect 26421 42180 27712 42208
rect 26421 42177 26433 42180
rect 26384 42171 26433 42177
rect 26384 42168 26390 42171
rect 27706 42168 27712 42180
rect 27764 42168 27770 42220
rect 27982 42168 27988 42220
rect 28040 42208 28046 42220
rect 28166 42208 28172 42220
rect 28040 42180 28172 42208
rect 28040 42168 28046 42180
rect 28166 42168 28172 42180
rect 28224 42208 28230 42220
rect 28552 42217 28580 42248
rect 28994 42236 29000 42248
rect 29052 42236 29058 42288
rect 30374 42276 30380 42288
rect 30335 42248 30380 42276
rect 30374 42236 30380 42248
rect 30432 42236 30438 42288
rect 30484 42285 30512 42316
rect 31386 42304 31392 42356
rect 31444 42344 31450 42356
rect 31938 42344 31944 42356
rect 31444 42316 31944 42344
rect 31444 42304 31450 42316
rect 31938 42304 31944 42316
rect 31996 42304 32002 42356
rect 33137 42347 33195 42353
rect 32508 42316 32991 42344
rect 30469 42279 30527 42285
rect 30469 42245 30481 42279
rect 30515 42245 30527 42279
rect 32398 42276 32404 42288
rect 30469 42239 30527 42245
rect 30668 42248 32404 42276
rect 28445 42211 28503 42217
rect 28445 42208 28457 42211
rect 28224 42180 28457 42208
rect 28224 42168 28230 42180
rect 28445 42177 28457 42180
rect 28491 42177 28503 42211
rect 28445 42171 28503 42177
rect 28537 42211 28595 42217
rect 28537 42177 28549 42211
rect 28583 42177 28595 42211
rect 28537 42171 28595 42177
rect 28626 42168 28632 42220
rect 28684 42208 28690 42220
rect 28721 42211 28779 42217
rect 28721 42208 28733 42211
rect 28684 42180 28733 42208
rect 28684 42168 28690 42180
rect 28721 42177 28733 42180
rect 28767 42177 28779 42211
rect 28721 42171 28779 42177
rect 28810 42168 28816 42220
rect 28868 42208 28874 42220
rect 30280 42211 30338 42217
rect 28868 42180 28913 42208
rect 28868 42168 28874 42180
rect 30280 42177 30292 42211
rect 30326 42208 30338 42211
rect 30558 42208 30564 42220
rect 30326 42180 30564 42208
rect 30326 42177 30338 42180
rect 30280 42171 30338 42177
rect 30558 42168 30564 42180
rect 30616 42168 30622 42220
rect 30668 42217 30696 42248
rect 32398 42236 32404 42248
rect 32456 42236 32462 42288
rect 32508 42217 32536 42316
rect 32858 42276 32864 42288
rect 32819 42248 32864 42276
rect 32858 42236 32864 42248
rect 32916 42236 32922 42288
rect 32963 42276 32991 42316
rect 33137 42313 33149 42347
rect 33183 42344 33195 42347
rect 33594 42344 33600 42356
rect 33183 42316 33600 42344
rect 33183 42313 33195 42316
rect 33137 42307 33195 42313
rect 33594 42304 33600 42316
rect 33652 42304 33658 42356
rect 34790 42344 34796 42356
rect 33796 42316 34796 42344
rect 32963 42248 33180 42276
rect 30652 42211 30710 42217
rect 30652 42177 30664 42211
rect 30698 42177 30710 42211
rect 30652 42171 30710 42177
rect 30745 42211 30803 42217
rect 30745 42177 30757 42211
rect 30791 42177 30803 42211
rect 30745 42171 30803 42177
rect 32493 42211 32551 42217
rect 32493 42177 32505 42211
rect 32539 42177 32551 42211
rect 32493 42171 32551 42177
rect 28902 42100 28908 42152
rect 28960 42140 28966 42152
rect 30760 42140 30788 42171
rect 32582 42168 32588 42220
rect 32640 42208 32646 42220
rect 32766 42208 32772 42220
rect 32640 42180 32685 42208
rect 32727 42180 32772 42208
rect 32640 42168 32646 42180
rect 32766 42168 32772 42180
rect 32824 42168 32830 42220
rect 32958 42211 33016 42217
rect 32958 42177 32970 42211
rect 33004 42177 33016 42211
rect 32958 42171 33016 42177
rect 31202 42140 31208 42152
rect 28960 42112 31208 42140
rect 28960 42100 28966 42112
rect 31202 42100 31208 42112
rect 31260 42100 31266 42152
rect 31297 42143 31355 42149
rect 31297 42109 31309 42143
rect 31343 42140 31355 42143
rect 31570 42140 31576 42152
rect 31343 42112 31576 42140
rect 31343 42109 31355 42112
rect 31297 42103 31355 42109
rect 31570 42100 31576 42112
rect 31628 42140 31634 42152
rect 32968 42140 32996 42171
rect 31628 42112 32996 42140
rect 33152 42140 33180 42248
rect 33502 42236 33508 42288
rect 33560 42276 33566 42288
rect 33796 42276 33824 42316
rect 34790 42304 34796 42316
rect 34848 42304 34854 42356
rect 35526 42304 35532 42356
rect 35584 42344 35590 42356
rect 35713 42347 35771 42353
rect 35713 42344 35725 42347
rect 35584 42316 35725 42344
rect 35584 42304 35590 42316
rect 35713 42313 35725 42316
rect 35759 42313 35771 42347
rect 35713 42307 35771 42313
rect 36357 42347 36415 42353
rect 36357 42313 36369 42347
rect 36403 42344 36415 42347
rect 38654 42344 38660 42356
rect 36403 42316 38660 42344
rect 36403 42313 36415 42316
rect 36357 42307 36415 42313
rect 33560 42248 33824 42276
rect 33873 42279 33931 42285
rect 33560 42236 33566 42248
rect 33873 42245 33885 42279
rect 33919 42276 33931 42279
rect 35434 42276 35440 42288
rect 33919 42248 35440 42276
rect 33919 42245 33931 42248
rect 33873 42239 33931 42245
rect 35434 42236 35440 42248
rect 35492 42236 35498 42288
rect 33226 42168 33232 42220
rect 33284 42208 33290 42220
rect 33781 42211 33839 42217
rect 33781 42208 33793 42211
rect 33284 42180 33793 42208
rect 33284 42168 33290 42180
rect 33781 42177 33793 42180
rect 33827 42177 33839 42211
rect 33962 42208 33968 42220
rect 33923 42180 33968 42208
rect 33781 42171 33839 42177
rect 33962 42168 33968 42180
rect 34020 42168 34026 42220
rect 34149 42211 34207 42217
rect 34149 42177 34161 42211
rect 34195 42208 34207 42211
rect 36372 42208 36400 42307
rect 38654 42304 38660 42316
rect 38712 42304 38718 42356
rect 34195 42180 36400 42208
rect 34195 42177 34207 42180
rect 34149 42171 34207 42177
rect 52546 42168 52552 42220
rect 52604 42208 52610 42220
rect 53745 42211 53803 42217
rect 53745 42208 53757 42211
rect 52604 42180 53757 42208
rect 52604 42168 52610 42180
rect 53745 42177 53757 42180
rect 53791 42177 53803 42211
rect 53745 42171 53803 42177
rect 53466 42140 53472 42152
rect 33152 42112 33640 42140
rect 53427 42112 53472 42140
rect 31628 42100 31634 42112
rect 27430 42032 27436 42084
rect 27488 42072 27494 42084
rect 29638 42072 29644 42084
rect 27488 42044 29644 42072
rect 27488 42032 27494 42044
rect 29638 42032 29644 42044
rect 29696 42072 29702 42084
rect 30190 42072 30196 42084
rect 29696 42044 30196 42072
rect 29696 42032 29702 42044
rect 30190 42032 30196 42044
rect 30248 42032 30254 42084
rect 33318 42032 33324 42084
rect 33376 42072 33382 42084
rect 33502 42072 33508 42084
rect 33376 42044 33508 42072
rect 33376 42032 33382 42044
rect 33502 42032 33508 42044
rect 33560 42032 33566 42084
rect 33612 42081 33640 42112
rect 53466 42100 53472 42112
rect 53524 42100 53530 42152
rect 33597 42075 33655 42081
rect 33597 42041 33609 42075
rect 33643 42041 33655 42075
rect 34698 42072 34704 42084
rect 34611 42044 34704 42072
rect 33597 42035 33655 42041
rect 34698 42032 34704 42044
rect 34756 42072 34762 42084
rect 48038 42072 48044 42084
rect 34756 42044 48044 42072
rect 34756 42032 34762 42044
rect 48038 42032 48044 42044
rect 48096 42032 48102 42084
rect 51813 42075 51871 42081
rect 51813 42041 51825 42075
rect 51859 42072 51871 42075
rect 54294 42072 54300 42084
rect 51859 42044 54300 42072
rect 51859 42041 51871 42044
rect 51813 42035 51871 42041
rect 54294 42032 54300 42044
rect 54352 42032 54358 42084
rect 26510 42004 26516 42016
rect 24443 41976 26280 42004
rect 26471 41976 26516 42004
rect 24443 41973 24455 41976
rect 24397 41967 24455 41973
rect 26510 41964 26516 41976
rect 26568 41964 26574 42016
rect 27522 41964 27528 42016
rect 27580 42004 27586 42016
rect 27617 42007 27675 42013
rect 27617 42004 27629 42007
rect 27580 41976 27629 42004
rect 27580 41964 27586 41976
rect 27617 41973 27629 41976
rect 27663 42004 27675 42007
rect 27982 42004 27988 42016
rect 27663 41976 27988 42004
rect 27663 41973 27675 41976
rect 27617 41967 27675 41973
rect 27982 41964 27988 41976
rect 28040 41964 28046 42016
rect 28258 42004 28264 42016
rect 28219 41976 28264 42004
rect 28258 41964 28264 41976
rect 28316 41964 28322 42016
rect 30006 41964 30012 42016
rect 30064 42004 30070 42016
rect 30101 42007 30159 42013
rect 30101 42004 30113 42007
rect 30064 41976 30113 42004
rect 30064 41964 30070 41976
rect 30101 41973 30113 41976
rect 30147 41973 30159 42007
rect 30101 41967 30159 41973
rect 31938 41964 31944 42016
rect 31996 42004 32002 42016
rect 32582 42004 32588 42016
rect 31996 41976 32588 42004
rect 31996 41964 32002 41976
rect 32582 41964 32588 41976
rect 32640 42004 32646 42016
rect 32766 42004 32772 42016
rect 32640 41976 32772 42004
rect 32640 41964 32646 41976
rect 32766 41964 32772 41976
rect 32824 41964 32830 42016
rect 32858 41964 32864 42016
rect 32916 42004 32922 42016
rect 34606 42004 34612 42016
rect 32916 41976 34612 42004
rect 32916 41964 32922 41976
rect 34606 41964 34612 41976
rect 34664 41964 34670 42016
rect 35253 42007 35311 42013
rect 35253 41973 35265 42007
rect 35299 42004 35311 42007
rect 35342 42004 35348 42016
rect 35299 41976 35348 42004
rect 35299 41973 35311 41976
rect 35253 41967 35311 41973
rect 35342 41964 35348 41976
rect 35400 41964 35406 42016
rect 52270 42004 52276 42016
rect 52231 41976 52276 42004
rect 52270 41964 52276 41976
rect 52328 41964 52334 42016
rect 53006 42004 53012 42016
rect 52967 41976 53012 42004
rect 53006 41964 53012 41976
rect 53064 41964 53070 42016
rect 1104 41914 54832 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 54832 41914
rect 1104 41840 54832 41862
rect 24854 41760 24860 41812
rect 24912 41800 24918 41812
rect 24912 41772 27845 41800
rect 24912 41760 24918 41772
rect 25038 41692 25044 41744
rect 25096 41732 25102 41744
rect 25961 41735 26019 41741
rect 25961 41732 25973 41735
rect 25096 41704 25973 41732
rect 25096 41692 25102 41704
rect 25961 41701 25973 41704
rect 26007 41732 26019 41735
rect 26786 41732 26792 41744
rect 26007 41704 26792 41732
rect 26007 41701 26019 41704
rect 25961 41695 26019 41701
rect 26786 41692 26792 41704
rect 26844 41692 26850 41744
rect 27817 41732 27845 41772
rect 27982 41760 27988 41812
rect 28040 41800 28046 41812
rect 28353 41803 28411 41809
rect 28353 41800 28365 41803
rect 28040 41772 28365 41800
rect 28040 41760 28046 41772
rect 28353 41769 28365 41772
rect 28399 41769 28411 41803
rect 28353 41763 28411 41769
rect 28534 41760 28540 41812
rect 28592 41800 28598 41812
rect 28813 41803 28871 41809
rect 28813 41800 28825 41803
rect 28592 41772 28825 41800
rect 28592 41760 28598 41772
rect 28813 41769 28825 41772
rect 28859 41769 28871 41803
rect 30837 41803 30895 41809
rect 30837 41800 30849 41803
rect 28813 41763 28871 41769
rect 28920 41772 30849 41800
rect 28920 41732 28948 41772
rect 30837 41769 30849 41772
rect 30883 41769 30895 41803
rect 32030 41800 32036 41812
rect 30837 41763 30895 41769
rect 31128 41772 32036 41800
rect 27817 41704 28948 41732
rect 29822 41692 29828 41744
rect 29880 41732 29886 41744
rect 29880 41704 30420 41732
rect 29880 41692 29886 41704
rect 2133 41667 2191 41673
rect 2133 41633 2145 41667
rect 2179 41664 2191 41667
rect 24486 41664 24492 41676
rect 2179 41636 24492 41664
rect 2179 41633 2191 41636
rect 2133 41627 2191 41633
rect 24486 41624 24492 41636
rect 24544 41624 24550 41676
rect 25866 41624 25872 41676
rect 25924 41664 25930 41676
rect 26142 41664 26148 41676
rect 25924 41636 26148 41664
rect 25924 41624 25930 41636
rect 26142 41624 26148 41636
rect 26200 41664 26206 41676
rect 26421 41667 26479 41673
rect 26421 41664 26433 41667
rect 26200 41636 26433 41664
rect 26200 41624 26206 41636
rect 26421 41633 26433 41636
rect 26467 41633 26479 41667
rect 26421 41627 26479 41633
rect 28810 41624 28816 41676
rect 28868 41664 28874 41676
rect 29454 41664 29460 41676
rect 28868 41636 29460 41664
rect 28868 41624 28874 41636
rect 29454 41624 29460 41636
rect 29512 41624 29518 41676
rect 30098 41624 30104 41676
rect 30156 41624 30162 41676
rect 2409 41599 2467 41605
rect 2409 41565 2421 41599
rect 2455 41596 2467 41599
rect 2774 41596 2780 41608
rect 2455 41568 2780 41596
rect 2455 41565 2467 41568
rect 2409 41559 2467 41565
rect 2774 41556 2780 41568
rect 2832 41596 2838 41608
rect 2869 41599 2927 41605
rect 2869 41596 2881 41599
rect 2832 41568 2881 41596
rect 2832 41556 2838 41568
rect 2869 41565 2881 41568
rect 2915 41565 2927 41599
rect 2869 41559 2927 41565
rect 26878 41556 26884 41608
rect 26936 41596 26942 41608
rect 27246 41596 27252 41608
rect 26936 41568 27252 41596
rect 26936 41556 26942 41568
rect 27246 41556 27252 41568
rect 27304 41556 27310 41608
rect 27709 41599 27767 41605
rect 27709 41565 27721 41599
rect 27755 41565 27767 41599
rect 27709 41559 27767 41565
rect 23477 41531 23535 41537
rect 23477 41497 23489 41531
rect 23523 41528 23535 41531
rect 24670 41528 24676 41540
rect 23523 41500 24676 41528
rect 23523 41497 23535 41500
rect 23477 41491 23535 41497
rect 24670 41488 24676 41500
rect 24728 41488 24734 41540
rect 25406 41488 25412 41540
rect 25464 41528 25470 41540
rect 27724 41528 27752 41559
rect 27798 41556 27804 41608
rect 27856 41596 27862 41608
rect 28074 41596 28080 41608
rect 27856 41568 27901 41596
rect 28035 41568 28080 41596
rect 27856 41556 27862 41568
rect 28074 41556 28080 41568
rect 28132 41556 28138 41608
rect 28215 41599 28273 41605
rect 28215 41565 28227 41599
rect 28261 41596 28273 41599
rect 28442 41596 28448 41608
rect 28261 41568 28448 41596
rect 28261 41565 28273 41568
rect 28215 41559 28273 41565
rect 28442 41556 28448 41568
rect 28500 41556 28506 41608
rect 29270 41556 29276 41608
rect 29328 41596 29334 41608
rect 29873 41599 29931 41605
rect 29873 41596 29885 41599
rect 29328 41568 29885 41596
rect 29328 41556 29334 41568
rect 29873 41565 29885 41568
rect 29919 41565 29931 41599
rect 29873 41559 29931 41565
rect 30009 41599 30067 41605
rect 30009 41565 30021 41599
rect 30055 41596 30067 41599
rect 30116 41596 30144 41624
rect 30392 41605 30420 41704
rect 30055 41568 30144 41596
rect 30284 41599 30342 41605
rect 30055 41565 30067 41568
rect 30009 41559 30067 41565
rect 30284 41565 30296 41599
rect 30330 41565 30342 41599
rect 30284 41559 30342 41565
rect 30370 41599 30428 41605
rect 30370 41565 30382 41599
rect 30416 41565 30428 41599
rect 30370 41559 30428 41565
rect 27982 41528 27988 41540
rect 25464 41500 27752 41528
rect 27943 41500 27988 41528
rect 25464 41488 25470 41500
rect 27982 41488 27988 41500
rect 28040 41488 28046 41540
rect 24029 41463 24087 41469
rect 24029 41429 24041 41463
rect 24075 41460 24087 41463
rect 24394 41460 24400 41472
rect 24075 41432 24400 41460
rect 24075 41429 24087 41432
rect 24029 41423 24087 41429
rect 24394 41420 24400 41432
rect 24452 41420 24458 41472
rect 24946 41460 24952 41472
rect 24907 41432 24952 41460
rect 24946 41420 24952 41432
rect 25004 41420 25010 41472
rect 27065 41463 27123 41469
rect 27065 41429 27077 41463
rect 27111 41460 27123 41463
rect 27246 41460 27252 41472
rect 27111 41432 27252 41460
rect 27111 41429 27123 41432
rect 27065 41423 27123 41429
rect 27246 41420 27252 41432
rect 27304 41420 27310 41472
rect 29730 41460 29736 41472
rect 29691 41432 29736 41460
rect 29730 41420 29736 41432
rect 29788 41420 29794 41472
rect 29886 41460 29914 41559
rect 30098 41528 30104 41540
rect 30059 41500 30104 41528
rect 30098 41488 30104 41500
rect 30156 41488 30162 41540
rect 30299 41528 30327 41559
rect 30558 41556 30564 41608
rect 30616 41596 30622 41608
rect 31128 41605 31156 41772
rect 32030 41760 32036 41772
rect 32088 41760 32094 41812
rect 32490 41760 32496 41812
rect 32548 41800 32554 41812
rect 33505 41803 33563 41809
rect 33505 41800 33517 41803
rect 32548 41772 33517 41800
rect 32548 41760 32554 41772
rect 33505 41769 33517 41772
rect 33551 41769 33563 41803
rect 33505 41763 33563 41769
rect 35342 41760 35348 41812
rect 35400 41800 35406 41812
rect 54113 41803 54171 41809
rect 54113 41800 54125 41803
rect 35400 41772 54125 41800
rect 35400 41760 35406 41772
rect 54113 41769 54125 41772
rect 54159 41769 54171 41803
rect 54113 41763 54171 41769
rect 33870 41732 33876 41744
rect 33520 41704 33876 41732
rect 31202 41624 31208 41676
rect 31260 41664 31266 41676
rect 33318 41664 33324 41676
rect 31260 41636 31524 41664
rect 31260 41624 31266 41636
rect 30975 41599 31033 41605
rect 30975 41596 30987 41599
rect 30616 41568 30987 41596
rect 30616 41556 30622 41568
rect 30975 41565 30987 41568
rect 31021 41565 31033 41599
rect 30975 41559 31033 41565
rect 31113 41599 31171 41605
rect 31113 41565 31125 41599
rect 31159 41565 31171 41599
rect 31386 41596 31392 41608
rect 31347 41568 31392 41596
rect 31113 41559 31171 41565
rect 31386 41556 31392 41568
rect 31444 41556 31450 41608
rect 31496 41605 31524 41636
rect 32967 41636 33324 41664
rect 32582 41605 32588 41608
rect 31481 41599 31539 41605
rect 31481 41565 31493 41599
rect 31527 41565 31539 41599
rect 32580 41596 32588 41605
rect 32543 41568 32588 41596
rect 31481 41559 31539 41565
rect 32580 41559 32588 41568
rect 32582 41556 32588 41559
rect 32640 41556 32646 41608
rect 32674 41556 32680 41608
rect 32732 41596 32738 41608
rect 32967 41605 32995 41636
rect 33318 41624 33324 41636
rect 33376 41624 33382 41676
rect 32952 41599 33010 41605
rect 32732 41568 32777 41596
rect 32732 41556 32738 41568
rect 32952 41565 32964 41599
rect 32998 41565 33010 41599
rect 32952 41559 33010 41565
rect 33045 41599 33103 41605
rect 33045 41565 33057 41599
rect 33091 41596 33103 41599
rect 33520 41596 33548 41704
rect 33870 41692 33876 41704
rect 33928 41692 33934 41744
rect 34330 41692 34336 41744
rect 34388 41732 34394 41744
rect 52825 41735 52883 41741
rect 52825 41732 52837 41735
rect 34388 41704 52837 41732
rect 34388 41692 34394 41704
rect 52825 41701 52837 41704
rect 52871 41701 52883 41735
rect 52825 41695 52883 41701
rect 53282 41692 53288 41744
rect 53340 41732 53346 41744
rect 53469 41735 53527 41741
rect 53469 41732 53481 41735
rect 53340 41704 53481 41732
rect 53340 41692 53346 41704
rect 53469 41701 53481 41704
rect 53515 41701 53527 41735
rect 53469 41695 53527 41701
rect 33796 41636 36400 41664
rect 33091 41568 33548 41596
rect 33091 41565 33103 41568
rect 33045 41559 33103 41565
rect 33594 41556 33600 41608
rect 33652 41596 33658 41608
rect 33796 41605 33824 41636
rect 33689 41599 33747 41605
rect 33689 41596 33701 41599
rect 33652 41568 33701 41596
rect 33652 41556 33658 41568
rect 33689 41565 33701 41568
rect 33735 41565 33747 41599
rect 33689 41559 33747 41565
rect 33781 41599 33839 41605
rect 33781 41565 33793 41599
rect 33827 41565 33839 41599
rect 33781 41559 33839 41565
rect 34057 41599 34115 41605
rect 34057 41565 34069 41599
rect 34103 41565 34115 41599
rect 34057 41559 34115 41565
rect 30466 41528 30472 41540
rect 30299 41500 30472 41528
rect 30466 41488 30472 41500
rect 30524 41488 30530 41540
rect 31205 41531 31263 41537
rect 31205 41497 31217 41531
rect 31251 41528 31263 41531
rect 32769 41531 32827 41537
rect 32769 41528 32781 41531
rect 31251 41500 32781 41528
rect 31251 41497 31263 41500
rect 31205 41491 31263 41497
rect 32769 41497 32781 41500
rect 32815 41528 32827 41531
rect 33226 41528 33232 41540
rect 32815 41500 33232 41528
rect 32815 41497 32827 41500
rect 32769 41491 32827 41497
rect 31220 41460 31248 41491
rect 33226 41488 33232 41500
rect 33284 41488 33290 41540
rect 33870 41528 33876 41540
rect 33831 41500 33876 41528
rect 33870 41488 33876 41500
rect 33928 41488 33934 41540
rect 34072 41528 34100 41559
rect 34790 41556 34796 41608
rect 34848 41596 34854 41608
rect 34885 41599 34943 41605
rect 34885 41596 34897 41599
rect 34848 41568 34897 41596
rect 34848 41556 34854 41568
rect 34885 41565 34897 41568
rect 34931 41565 34943 41599
rect 36262 41596 36268 41608
rect 34885 41559 34943 41565
rect 34992 41568 36268 41596
rect 34992 41528 35020 41568
rect 36262 41556 36268 41568
rect 36320 41556 36326 41608
rect 36372 41605 36400 41636
rect 36814 41624 36820 41676
rect 36872 41664 36878 41676
rect 38746 41664 38752 41676
rect 36872 41636 38752 41664
rect 36872 41624 36878 41636
rect 38746 41624 38752 41636
rect 38804 41624 38810 41676
rect 52454 41664 52460 41676
rect 45526 41636 52460 41664
rect 36357 41599 36415 41605
rect 36357 41565 36369 41599
rect 36403 41596 36415 41599
rect 45526 41596 45554 41636
rect 52454 41624 52460 41636
rect 52512 41624 52518 41676
rect 36403 41568 45554 41596
rect 51721 41599 51779 41605
rect 36403 41565 36415 41568
rect 36357 41559 36415 41565
rect 51721 41565 51733 41599
rect 51767 41596 51779 41599
rect 52362 41596 52368 41608
rect 51767 41568 52368 41596
rect 51767 41565 51779 41568
rect 51721 41559 51779 41565
rect 52362 41556 52368 41568
rect 52420 41556 52426 41608
rect 53006 41596 53012 41608
rect 52967 41568 53012 41596
rect 53006 41556 53012 41568
rect 53064 41556 53070 41608
rect 53653 41599 53711 41605
rect 53653 41596 53665 41599
rect 53576 41568 53665 41596
rect 34072 41500 35020 41528
rect 35069 41531 35127 41537
rect 35069 41497 35081 41531
rect 35115 41497 35127 41531
rect 35069 41491 35127 41497
rect 29886 41432 31248 41460
rect 32401 41463 32459 41469
rect 32401 41429 32413 41463
rect 32447 41460 32459 41463
rect 33318 41460 33324 41472
rect 32447 41432 33324 41460
rect 32447 41429 32459 41432
rect 32401 41423 32459 41429
rect 33318 41420 33324 41432
rect 33376 41420 33382 41472
rect 34054 41420 34060 41472
rect 34112 41460 34118 41472
rect 35084 41460 35112 41491
rect 35434 41488 35440 41540
rect 35492 41528 35498 41540
rect 35492 41500 52224 41528
rect 35492 41488 35498 41500
rect 34112 41432 35112 41460
rect 35253 41463 35311 41469
rect 34112 41420 34118 41432
rect 35253 41429 35265 41463
rect 35299 41460 35311 41463
rect 35342 41460 35348 41472
rect 35299 41432 35348 41460
rect 35299 41429 35311 41432
rect 35253 41423 35311 41429
rect 35342 41420 35348 41432
rect 35400 41420 35406 41472
rect 35618 41420 35624 41472
rect 35676 41460 35682 41472
rect 35713 41463 35771 41469
rect 35713 41460 35725 41463
rect 35676 41432 35725 41460
rect 35676 41420 35682 41432
rect 35713 41429 35725 41432
rect 35759 41429 35771 41463
rect 35713 41423 35771 41429
rect 36262 41420 36268 41472
rect 36320 41460 36326 41472
rect 36814 41460 36820 41472
rect 36320 41432 36820 41460
rect 36320 41420 36326 41432
rect 36814 41420 36820 41432
rect 36872 41420 36878 41472
rect 52196 41469 52224 41500
rect 52181 41463 52239 41469
rect 52181 41429 52193 41463
rect 52227 41429 52239 41463
rect 52181 41423 52239 41429
rect 52270 41420 52276 41472
rect 52328 41460 52334 41472
rect 53576 41460 53604 41568
rect 53653 41565 53665 41568
rect 53699 41565 53711 41599
rect 54294 41596 54300 41608
rect 54255 41568 54300 41596
rect 53653 41559 53711 41565
rect 54294 41556 54300 41568
rect 54352 41556 54358 41608
rect 53650 41460 53656 41472
rect 52328 41432 53656 41460
rect 52328 41420 52334 41432
rect 53650 41420 53656 41432
rect 53708 41420 53714 41472
rect 1104 41370 54832 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 54832 41370
rect 1104 41296 54832 41318
rect 24486 41256 24492 41268
rect 24447 41228 24492 41256
rect 24486 41216 24492 41228
rect 24544 41216 24550 41268
rect 26326 41256 26332 41268
rect 26287 41228 26332 41256
rect 26326 41216 26332 41228
rect 26384 41216 26390 41268
rect 26510 41216 26516 41268
rect 26568 41256 26574 41268
rect 28261 41259 28319 41265
rect 26568 41228 27568 41256
rect 26568 41216 26574 41228
rect 24394 41148 24400 41200
rect 24452 41188 24458 41200
rect 27540 41197 27568 41228
rect 28261 41225 28273 41259
rect 28307 41256 28319 41259
rect 28626 41256 28632 41268
rect 28307 41228 28632 41256
rect 28307 41225 28319 41228
rect 28261 41219 28319 41225
rect 28626 41216 28632 41228
rect 28684 41216 28690 41268
rect 29362 41216 29368 41268
rect 29420 41216 29426 41268
rect 30558 41216 30564 41268
rect 30616 41256 30622 41268
rect 30929 41259 30987 41265
rect 30929 41256 30941 41259
rect 30616 41228 30941 41256
rect 30616 41216 30622 41228
rect 30929 41225 30941 41228
rect 30975 41225 30987 41259
rect 30929 41219 30987 41225
rect 31573 41259 31631 41265
rect 31573 41225 31585 41259
rect 31619 41256 31631 41259
rect 32214 41256 32220 41268
rect 31619 41228 32220 41256
rect 31619 41225 31631 41228
rect 31573 41219 31631 41225
rect 32214 41216 32220 41228
rect 32272 41216 32278 41268
rect 32674 41216 32680 41268
rect 32732 41256 32738 41268
rect 32732 41228 33180 41256
rect 32732 41216 32738 41228
rect 26237 41191 26295 41197
rect 26237 41188 26249 41191
rect 24452 41160 26249 41188
rect 24452 41148 24458 41160
rect 26237 41157 26249 41160
rect 26283 41157 26295 41191
rect 27433 41191 27491 41197
rect 27433 41188 27445 41191
rect 26237 41151 26295 41157
rect 26344 41160 27445 41188
rect 2133 41123 2191 41129
rect 2133 41089 2145 41123
rect 2179 41120 2191 41123
rect 24026 41120 24032 41132
rect 2179 41092 6914 41120
rect 23939 41092 24032 41120
rect 2179 41089 2191 41092
rect 2133 41083 2191 41089
rect 2409 41055 2467 41061
rect 2409 41021 2421 41055
rect 2455 41052 2467 41055
rect 2774 41052 2780 41064
rect 2455 41024 2780 41052
rect 2455 41021 2467 41024
rect 2409 41015 2467 41021
rect 2774 41012 2780 41024
rect 2832 41052 2838 41064
rect 2869 41055 2927 41061
rect 2869 41052 2881 41055
rect 2832 41024 2881 41052
rect 2832 41012 2838 41024
rect 2869 41021 2881 41024
rect 2915 41021 2927 41055
rect 2869 41015 2927 41021
rect 6886 40984 6914 41092
rect 24026 41080 24032 41092
rect 24084 41120 24090 41132
rect 26344 41120 26372 41160
rect 27433 41157 27445 41160
rect 27479 41157 27491 41191
rect 27433 41151 27491 41157
rect 27525 41191 27583 41197
rect 27525 41157 27537 41191
rect 27571 41157 27583 41191
rect 27525 41151 27583 41157
rect 28537 41191 28595 41197
rect 28537 41157 28549 41191
rect 28583 41188 28595 41191
rect 28718 41188 28724 41200
rect 28583 41160 28724 41188
rect 28583 41157 28595 41160
rect 28537 41151 28595 41157
rect 28718 41148 28724 41160
rect 28776 41148 28782 41200
rect 29380 41188 29408 41216
rect 29641 41191 29699 41197
rect 29641 41188 29653 41191
rect 29380 41160 29653 41188
rect 29641 41157 29653 41160
rect 29687 41157 29699 41191
rect 29641 41151 29699 41157
rect 32766 41148 32772 41200
rect 32824 41188 32830 41200
rect 33152 41197 33180 41228
rect 33226 41216 33232 41268
rect 33284 41256 33290 41268
rect 35250 41256 35256 41268
rect 33284 41228 35256 41256
rect 33284 41216 33290 41228
rect 35250 41216 35256 41228
rect 35308 41216 35314 41268
rect 36538 41216 36544 41268
rect 36596 41256 36602 41268
rect 50154 41256 50160 41268
rect 36596 41228 50160 41256
rect 36596 41216 36602 41228
rect 50154 41216 50160 41228
rect 50212 41216 50218 41268
rect 33045 41191 33103 41197
rect 33045 41188 33057 41191
rect 32824 41160 33057 41188
rect 32824 41148 32830 41160
rect 33045 41157 33057 41160
rect 33091 41157 33103 41191
rect 33045 41151 33103 41157
rect 33137 41191 33195 41197
rect 33137 41157 33149 41191
rect 33183 41157 33195 41191
rect 33137 41151 33195 41157
rect 33686 41148 33692 41200
rect 33744 41188 33750 41200
rect 33873 41191 33931 41197
rect 33873 41188 33885 41191
rect 33744 41160 33885 41188
rect 33744 41148 33750 41160
rect 33873 41157 33885 41160
rect 33919 41157 33931 41191
rect 33873 41151 33931 41157
rect 51166 41148 51172 41200
rect 51224 41188 51230 41200
rect 51224 41160 53788 41188
rect 51224 41148 51230 41160
rect 24084 41092 26372 41120
rect 24084 41080 24090 41092
rect 26418 41080 26424 41132
rect 26476 41120 26482 41132
rect 27062 41120 27068 41132
rect 26476 41092 27068 41120
rect 26476 41080 26482 41092
rect 27062 41080 27068 41092
rect 27120 41120 27126 41132
rect 27341 41123 27399 41129
rect 27341 41120 27353 41123
rect 27120 41092 27353 41120
rect 27120 41080 27126 41092
rect 27341 41089 27353 41092
rect 27387 41089 27399 41123
rect 27706 41120 27712 41132
rect 27667 41092 27712 41120
rect 27341 41083 27399 41089
rect 27706 41080 27712 41092
rect 27764 41080 27770 41132
rect 28445 41123 28503 41129
rect 28445 41089 28457 41123
rect 28491 41089 28503 41123
rect 28626 41120 28632 41132
rect 28587 41092 28632 41120
rect 28445 41083 28503 41089
rect 25133 41055 25191 41061
rect 25133 41021 25145 41055
rect 25179 41052 25191 41055
rect 27724 41052 27752 41080
rect 25179 41024 27752 41052
rect 25179 41021 25191 41024
rect 25133 41015 25191 41021
rect 25774 40984 25780 40996
rect 6886 40956 25780 40984
rect 25774 40944 25780 40956
rect 25832 40944 25838 40996
rect 27430 40944 27436 40996
rect 27488 40984 27494 40996
rect 28460 40984 28488 41083
rect 28626 41080 28632 41092
rect 28684 41080 28690 41132
rect 28813 41123 28871 41129
rect 28813 41089 28825 41123
rect 28859 41120 28871 41123
rect 29086 41120 29092 41132
rect 28859 41092 29092 41120
rect 28859 41089 28871 41092
rect 28813 41083 28871 41089
rect 29086 41080 29092 41092
rect 29144 41080 29150 41132
rect 29178 41080 29184 41132
rect 29236 41120 29242 41132
rect 29273 41123 29331 41129
rect 29273 41120 29285 41123
rect 29236 41092 29285 41120
rect 29236 41080 29242 41092
rect 29273 41089 29285 41092
rect 29319 41089 29331 41123
rect 29273 41083 29331 41089
rect 29421 41123 29479 41129
rect 29421 41089 29433 41123
rect 29467 41120 29479 41123
rect 29549 41123 29607 41129
rect 29467 41089 29500 41120
rect 29421 41083 29500 41089
rect 29549 41089 29561 41123
rect 29595 41089 29607 41123
rect 29549 41083 29607 41089
rect 29779 41123 29837 41129
rect 29779 41089 29791 41123
rect 29825 41120 29837 41123
rect 30190 41120 30196 41132
rect 29825 41092 30196 41120
rect 29825 41089 29837 41092
rect 29779 41083 29837 41089
rect 27488 40956 28488 40984
rect 27488 40944 27494 40956
rect 28626 40944 28632 40996
rect 28684 40984 28690 40996
rect 29270 40984 29276 40996
rect 28684 40956 29276 40984
rect 28684 40944 28690 40956
rect 29270 40944 29276 40956
rect 29328 40944 29334 40996
rect 29472 40984 29500 41083
rect 29564 41052 29592 41083
rect 30190 41080 30196 41092
rect 30248 41080 30254 41132
rect 31846 41080 31852 41132
rect 31904 41080 31910 41132
rect 32948 41123 33006 41129
rect 32948 41089 32960 41123
rect 32994 41089 33006 41123
rect 32948 41083 33006 41089
rect 30098 41052 30104 41064
rect 29564 41024 30104 41052
rect 30098 41012 30104 41024
rect 30156 41012 30162 41064
rect 30742 40984 30748 40996
rect 29472 40956 30748 40984
rect 30742 40944 30748 40956
rect 30800 40944 30806 40996
rect 31864 40984 31892 41080
rect 32973 40984 33001 41083
rect 33226 41080 33232 41132
rect 33284 41120 33290 41132
rect 33320 41123 33378 41129
rect 33320 41120 33332 41123
rect 33284 41092 33332 41120
rect 33284 41080 33290 41092
rect 33320 41089 33332 41092
rect 33366 41089 33378 41123
rect 33320 41083 33378 41089
rect 33413 41123 33471 41129
rect 33413 41089 33425 41123
rect 33459 41089 33471 41123
rect 33413 41083 33471 41089
rect 33428 41052 33456 41083
rect 33962 41080 33968 41132
rect 34020 41120 34026 41132
rect 34057 41123 34115 41129
rect 34057 41120 34069 41123
rect 34020 41092 34069 41120
rect 34020 41080 34026 41092
rect 34057 41089 34069 41092
rect 34103 41089 34115 41123
rect 35250 41120 35256 41132
rect 35211 41092 35256 41120
rect 34057 41083 34115 41089
rect 35250 41080 35256 41092
rect 35308 41080 35314 41132
rect 53098 41120 53104 41132
rect 45526 41092 53104 41120
rect 31864 40956 33001 40984
rect 33336 41024 33456 41052
rect 33336 40984 33364 41024
rect 33870 41012 33876 41064
rect 33928 41052 33934 41064
rect 34701 41055 34759 41061
rect 34701 41052 34713 41055
rect 33928 41024 34713 41052
rect 33928 41012 33934 41024
rect 34701 41021 34713 41024
rect 34747 41021 34759 41055
rect 34701 41015 34759 41021
rect 35805 41055 35863 41061
rect 35805 41021 35817 41055
rect 35851 41021 35863 41055
rect 35805 41015 35863 41021
rect 33410 40984 33416 40996
rect 33336 40956 33416 40984
rect 31956 40928 31984 40956
rect 25685 40919 25743 40925
rect 25685 40885 25697 40919
rect 25731 40916 25743 40919
rect 25866 40916 25872 40928
rect 25731 40888 25872 40916
rect 25731 40885 25743 40888
rect 25685 40879 25743 40885
rect 25866 40876 25872 40888
rect 25924 40876 25930 40928
rect 26510 40876 26516 40928
rect 26568 40916 26574 40928
rect 27157 40919 27215 40925
rect 27157 40916 27169 40919
rect 26568 40888 27169 40916
rect 26568 40876 26574 40888
rect 27157 40885 27169 40888
rect 27203 40885 27215 40919
rect 27157 40879 27215 40885
rect 27246 40876 27252 40928
rect 27304 40916 27310 40928
rect 27706 40916 27712 40928
rect 27304 40888 27712 40916
rect 27304 40876 27310 40888
rect 27706 40876 27712 40888
rect 27764 40916 27770 40928
rect 29454 40916 29460 40928
rect 27764 40888 29460 40916
rect 27764 40876 27770 40888
rect 29454 40876 29460 40888
rect 29512 40876 29518 40928
rect 29914 40916 29920 40928
rect 29875 40888 29920 40916
rect 29914 40876 29920 40888
rect 29972 40876 29978 40928
rect 30190 40876 30196 40928
rect 30248 40916 30254 40928
rect 30377 40919 30435 40925
rect 30377 40916 30389 40919
rect 30248 40888 30389 40916
rect 30248 40876 30254 40888
rect 30377 40885 30389 40888
rect 30423 40916 30435 40919
rect 31754 40916 31760 40928
rect 30423 40888 31760 40916
rect 30423 40885 30435 40888
rect 30377 40879 30435 40885
rect 31754 40876 31760 40888
rect 31812 40876 31818 40928
rect 31938 40876 31944 40928
rect 31996 40876 32002 40928
rect 32766 40916 32772 40928
rect 32727 40888 32772 40916
rect 32766 40876 32772 40888
rect 32824 40876 32830 40928
rect 32973 40916 33001 40956
rect 33410 40944 33416 40956
rect 33468 40944 33474 40996
rect 35820 40984 35848 41015
rect 33520 40956 35848 40984
rect 33520 40916 33548 40956
rect 35894 40944 35900 40996
rect 35952 40984 35958 40996
rect 45526 40984 45554 41092
rect 53098 41080 53104 41092
rect 53156 41080 53162 41132
rect 53760 41129 53788 41160
rect 53745 41123 53803 41129
rect 53745 41089 53757 41123
rect 53791 41089 53803 41123
rect 53745 41083 53803 41089
rect 51813 41055 51871 41061
rect 51813 41021 51825 41055
rect 51859 41052 51871 41055
rect 53466 41052 53472 41064
rect 51859 41024 53472 41052
rect 51859 41021 51871 41024
rect 51813 41015 51871 41021
rect 53466 41012 53472 41024
rect 53524 41012 53530 41064
rect 35952 40956 45554 40984
rect 52365 40987 52423 40993
rect 35952 40944 35958 40956
rect 52365 40953 52377 40987
rect 52411 40984 52423 40987
rect 54294 40984 54300 40996
rect 52411 40956 54300 40984
rect 52411 40953 52423 40956
rect 52365 40947 52423 40953
rect 54294 40944 54300 40956
rect 54352 40944 54358 40996
rect 34238 40916 34244 40928
rect 32973 40888 33548 40916
rect 34199 40888 34244 40916
rect 34238 40876 34244 40888
rect 34296 40876 34302 40928
rect 52914 40916 52920 40928
rect 52875 40888 52920 40916
rect 52914 40876 52920 40888
rect 52972 40876 52978 40928
rect 1104 40826 54832 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 54832 40826
rect 1104 40752 54832 40774
rect 23382 40712 23388 40724
rect 23343 40684 23388 40712
rect 23382 40672 23388 40684
rect 23440 40672 23446 40724
rect 24949 40715 25007 40721
rect 24949 40681 24961 40715
rect 24995 40712 25007 40715
rect 36538 40712 36544 40724
rect 24995 40684 36544 40712
rect 24995 40681 25007 40684
rect 24949 40675 25007 40681
rect 23400 40644 23428 40672
rect 23400 40616 26281 40644
rect 2130 40508 2136 40520
rect 2091 40480 2136 40508
rect 2130 40468 2136 40480
rect 2188 40468 2194 40520
rect 2409 40511 2467 40517
rect 2409 40477 2421 40511
rect 2455 40508 2467 40511
rect 2774 40508 2780 40520
rect 2455 40480 2780 40508
rect 2455 40477 2467 40480
rect 2409 40471 2467 40477
rect 2774 40468 2780 40480
rect 2832 40508 2838 40520
rect 2869 40511 2927 40517
rect 2869 40508 2881 40511
rect 2832 40480 2881 40508
rect 2832 40468 2838 40480
rect 2869 40477 2881 40480
rect 2915 40477 2927 40511
rect 2869 40471 2927 40477
rect 24670 40468 24676 40520
rect 24728 40508 24734 40520
rect 26142 40508 26148 40520
rect 24728 40480 26148 40508
rect 24728 40468 24734 40480
rect 26142 40468 26148 40480
rect 26200 40468 26206 40520
rect 26253 40517 26281 40616
rect 26253 40511 26327 40517
rect 26253 40480 26281 40511
rect 26269 40477 26281 40480
rect 26315 40477 26327 40511
rect 26418 40508 26424 40520
rect 26379 40480 26424 40508
rect 26269 40471 26327 40477
rect 26418 40468 26424 40480
rect 26476 40468 26482 40520
rect 26510 40468 26516 40520
rect 26568 40508 26574 40520
rect 26568 40480 26613 40508
rect 26568 40468 26574 40480
rect 26878 40468 26884 40520
rect 26936 40508 26942 40520
rect 27632 40517 27660 40684
rect 36538 40672 36544 40684
rect 36596 40672 36602 40724
rect 41386 40684 45554 40712
rect 27890 40644 27896 40656
rect 27851 40616 27896 40644
rect 27890 40604 27896 40616
rect 27948 40604 27954 40656
rect 28810 40604 28816 40656
rect 28868 40644 28874 40656
rect 28997 40647 29055 40653
rect 28868 40604 28902 40644
rect 28997 40613 29009 40647
rect 29043 40644 29055 40647
rect 30282 40644 30288 40656
rect 29043 40616 30288 40644
rect 29043 40613 29055 40616
rect 28997 40607 29055 40613
rect 30282 40604 30288 40616
rect 30340 40604 30346 40656
rect 30377 40647 30435 40653
rect 30377 40613 30389 40647
rect 30423 40644 30435 40647
rect 30558 40644 30564 40656
rect 30423 40616 30564 40644
rect 30423 40613 30435 40616
rect 30377 40607 30435 40613
rect 30558 40604 30564 40616
rect 30616 40604 30622 40656
rect 33134 40644 33140 40656
rect 31772 40616 33140 40644
rect 28718 40576 28724 40588
rect 28644 40548 28724 40576
rect 27249 40511 27307 40517
rect 27249 40508 27261 40511
rect 26936 40480 27261 40508
rect 26936 40468 26942 40480
rect 27249 40477 27261 40480
rect 27295 40477 27307 40511
rect 27249 40471 27307 40477
rect 27342 40511 27400 40517
rect 27342 40477 27354 40511
rect 27388 40477 27400 40511
rect 27342 40471 27400 40477
rect 27617 40511 27675 40517
rect 27617 40477 27629 40511
rect 27663 40477 27675 40511
rect 27617 40471 27675 40477
rect 27755 40511 27813 40517
rect 27755 40477 27767 40511
rect 27801 40508 27813 40511
rect 27801 40480 28028 40508
rect 27801 40477 27813 40480
rect 27755 40471 27813 40477
rect 24486 40400 24492 40452
rect 24544 40440 24550 40452
rect 27356 40440 27384 40471
rect 24544 40412 27384 40440
rect 24544 40400 24550 40412
rect 27522 40400 27528 40452
rect 27580 40440 27586 40452
rect 27580 40412 27625 40440
rect 27580 40400 27586 40412
rect 23566 40332 23572 40384
rect 23624 40372 23630 40384
rect 23937 40375 23995 40381
rect 23937 40372 23949 40375
rect 23624 40344 23949 40372
rect 23624 40332 23630 40344
rect 23937 40341 23949 40344
rect 23983 40341 23995 40375
rect 25498 40372 25504 40384
rect 25459 40344 25504 40372
rect 23937 40335 23995 40341
rect 25498 40332 25504 40344
rect 25556 40332 25562 40384
rect 25590 40332 25596 40384
rect 25648 40372 25654 40384
rect 25961 40375 26019 40381
rect 25961 40372 25973 40375
rect 25648 40344 25973 40372
rect 25648 40332 25654 40344
rect 25961 40341 25973 40344
rect 26007 40341 26019 40375
rect 25961 40335 26019 40341
rect 26142 40332 26148 40384
rect 26200 40372 26206 40384
rect 26878 40372 26884 40384
rect 26200 40344 26884 40372
rect 26200 40332 26206 40344
rect 26878 40332 26884 40344
rect 26936 40332 26942 40384
rect 28000 40372 28028 40480
rect 28258 40468 28264 40520
rect 28316 40502 28322 40520
rect 28644 40517 28672 40548
rect 28718 40536 28724 40548
rect 28776 40536 28782 40588
rect 28874 40576 28902 40604
rect 30098 40576 30104 40588
rect 28874 40548 30104 40576
rect 30098 40536 30104 40548
rect 30156 40576 30162 40588
rect 30837 40579 30895 40585
rect 30837 40576 30849 40579
rect 30156 40548 30849 40576
rect 30156 40536 30162 40548
rect 30837 40545 30849 40548
rect 30883 40545 30895 40579
rect 30837 40539 30895 40545
rect 28353 40511 28411 40517
rect 28353 40502 28365 40511
rect 28316 40477 28365 40502
rect 28399 40477 28411 40511
rect 28316 40474 28411 40477
rect 28316 40468 28322 40474
rect 28353 40471 28411 40474
rect 28501 40511 28559 40517
rect 28501 40477 28513 40511
rect 28547 40508 28559 40511
rect 28629 40511 28687 40517
rect 28547 40477 28580 40508
rect 28501 40471 28580 40477
rect 28629 40477 28641 40511
rect 28675 40477 28687 40511
rect 28629 40471 28687 40477
rect 28859 40511 28917 40517
rect 28859 40477 28871 40511
rect 28905 40508 28917 40511
rect 29086 40508 29092 40520
rect 28905 40480 29092 40508
rect 28905 40477 28917 40480
rect 28859 40471 28917 40477
rect 28074 40400 28080 40452
rect 28132 40440 28138 40452
rect 28552 40440 28580 40471
rect 29086 40468 29092 40480
rect 29144 40468 29150 40520
rect 31772 40517 31800 40616
rect 33134 40604 33140 40616
rect 33192 40604 33198 40656
rect 33226 40604 33232 40656
rect 33284 40644 33290 40656
rect 33870 40644 33876 40656
rect 33284 40616 33876 40644
rect 33284 40604 33290 40616
rect 33870 40604 33876 40616
rect 33928 40604 33934 40656
rect 35802 40604 35808 40656
rect 35860 40644 35866 40656
rect 41386 40644 41414 40684
rect 35860 40616 41414 40644
rect 45526 40644 45554 40684
rect 51902 40672 51908 40724
rect 51960 40712 51966 40724
rect 52181 40715 52239 40721
rect 52181 40712 52193 40715
rect 51960 40684 52193 40712
rect 51960 40672 51966 40684
rect 52181 40681 52193 40684
rect 52227 40681 52239 40715
rect 52181 40675 52239 40681
rect 53009 40715 53067 40721
rect 53009 40681 53021 40715
rect 53055 40712 53067 40715
rect 53190 40712 53196 40724
rect 53055 40684 53196 40712
rect 53055 40681 53067 40684
rect 53009 40675 53067 40681
rect 53190 40672 53196 40684
rect 53248 40672 53254 40724
rect 54110 40712 54116 40724
rect 54071 40684 54116 40712
rect 54110 40672 54116 40684
rect 54168 40672 54174 40724
rect 52638 40644 52644 40656
rect 45526 40616 52644 40644
rect 35860 40604 35866 40616
rect 52638 40604 52644 40616
rect 52696 40604 52702 40656
rect 32674 40536 32680 40588
rect 32732 40536 32738 40588
rect 32967 40548 36308 40576
rect 31757 40511 31815 40517
rect 31757 40477 31769 40511
rect 31803 40477 31815 40511
rect 32214 40508 32220 40520
rect 31757 40471 31815 40477
rect 31864 40480 32220 40508
rect 28132 40412 28580 40440
rect 28721 40443 28779 40449
rect 28132 40400 28138 40412
rect 28721 40409 28733 40443
rect 28767 40440 28779 40443
rect 31864 40440 31892 40480
rect 32214 40468 32220 40480
rect 32272 40468 32278 40520
rect 32582 40517 32588 40520
rect 32580 40508 32588 40517
rect 32543 40480 32588 40508
rect 32580 40471 32588 40480
rect 32582 40468 32588 40471
rect 32640 40468 32646 40520
rect 32692 40508 32720 40536
rect 32967 40517 32995 40548
rect 32769 40511 32827 40517
rect 32769 40508 32781 40511
rect 32692 40480 32781 40508
rect 32769 40477 32781 40480
rect 32815 40477 32827 40511
rect 32769 40471 32827 40477
rect 32952 40511 33010 40517
rect 32952 40477 32964 40511
rect 32998 40477 33010 40511
rect 32952 40471 33010 40477
rect 33042 40468 33048 40520
rect 33100 40508 33106 40520
rect 33100 40480 33145 40508
rect 33100 40468 33106 40480
rect 33318 40468 33324 40520
rect 33376 40508 33382 40520
rect 33505 40511 33563 40517
rect 33505 40508 33517 40511
rect 33376 40480 33517 40508
rect 33376 40468 33382 40480
rect 33505 40477 33517 40480
rect 33551 40477 33563 40511
rect 33505 40471 33563 40477
rect 35069 40511 35127 40517
rect 35069 40477 35081 40511
rect 35115 40508 35127 40511
rect 35342 40508 35348 40520
rect 35115 40480 35348 40508
rect 35115 40477 35127 40480
rect 35069 40471 35127 40477
rect 35342 40468 35348 40480
rect 35400 40468 35406 40520
rect 28767 40412 31892 40440
rect 28767 40409 28779 40412
rect 28721 40403 28779 40409
rect 32122 40400 32128 40452
rect 32180 40440 32186 40452
rect 32677 40443 32735 40449
rect 32677 40440 32689 40443
rect 32180 40412 32689 40440
rect 32180 40400 32186 40412
rect 32677 40409 32689 40412
rect 32723 40409 32735 40443
rect 33686 40440 33692 40452
rect 33647 40412 33692 40440
rect 32677 40403 32735 40409
rect 33686 40400 33692 40412
rect 33744 40400 33750 40452
rect 34790 40400 34796 40452
rect 34848 40440 34854 40452
rect 36280 40449 36308 40548
rect 51721 40511 51779 40517
rect 51721 40477 51733 40511
rect 51767 40508 51779 40511
rect 52362 40508 52368 40520
rect 51767 40480 52368 40508
rect 51767 40477 51779 40480
rect 51721 40471 51779 40477
rect 52362 40468 52368 40480
rect 52420 40468 52426 40520
rect 52825 40511 52883 40517
rect 52825 40477 52837 40511
rect 52871 40508 52883 40511
rect 52914 40508 52920 40520
rect 52871 40480 52920 40508
rect 52871 40477 52883 40480
rect 52825 40471 52883 40477
rect 52914 40468 52920 40480
rect 52972 40468 52978 40520
rect 53650 40508 53656 40520
rect 53611 40480 53656 40508
rect 53650 40468 53656 40480
rect 53708 40468 53714 40520
rect 54294 40508 54300 40520
rect 54255 40480 54300 40508
rect 54294 40468 54300 40480
rect 54352 40468 54358 40520
rect 34885 40443 34943 40449
rect 34885 40440 34897 40443
rect 34848 40412 34897 40440
rect 34848 40400 34854 40412
rect 34885 40409 34897 40412
rect 34931 40409 34943 40443
rect 34885 40403 34943 40409
rect 36265 40443 36323 40449
rect 36265 40409 36277 40443
rect 36311 40440 36323 40443
rect 36311 40412 53512 40440
rect 36311 40409 36323 40412
rect 36265 40403 36323 40409
rect 29086 40372 29092 40384
rect 28000 40344 29092 40372
rect 29086 40332 29092 40344
rect 29144 40332 29150 40384
rect 29638 40332 29644 40384
rect 29696 40372 29702 40384
rect 29733 40375 29791 40381
rect 29733 40372 29745 40375
rect 29696 40344 29745 40372
rect 29696 40332 29702 40344
rect 29733 40341 29745 40344
rect 29779 40372 29791 40375
rect 29822 40372 29828 40384
rect 29779 40344 29828 40372
rect 29779 40341 29791 40344
rect 29733 40335 29791 40341
rect 29822 40332 29828 40344
rect 29880 40332 29886 40384
rect 31849 40375 31907 40381
rect 31849 40341 31861 40375
rect 31895 40372 31907 40375
rect 32214 40372 32220 40384
rect 31895 40344 32220 40372
rect 31895 40341 31907 40344
rect 31849 40335 31907 40341
rect 32214 40332 32220 40344
rect 32272 40332 32278 40384
rect 32398 40372 32404 40384
rect 32359 40344 32404 40372
rect 32398 40332 32404 40344
rect 32456 40332 32462 40384
rect 32490 40332 32496 40384
rect 32548 40372 32554 40384
rect 33594 40372 33600 40384
rect 32548 40344 33600 40372
rect 32548 40332 32554 40344
rect 33594 40332 33600 40344
rect 33652 40332 33658 40384
rect 33870 40372 33876 40384
rect 33831 40344 33876 40372
rect 33870 40332 33876 40344
rect 33928 40332 33934 40384
rect 34606 40332 34612 40384
rect 34664 40372 34670 40384
rect 53484 40381 53512 40412
rect 35621 40375 35679 40381
rect 35621 40372 35633 40375
rect 34664 40344 35633 40372
rect 34664 40332 34670 40344
rect 35621 40341 35633 40344
rect 35667 40341 35679 40375
rect 35621 40335 35679 40341
rect 53469 40375 53527 40381
rect 53469 40341 53481 40375
rect 53515 40341 53527 40375
rect 53469 40335 53527 40341
rect 1104 40282 54832 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 54832 40282
rect 1104 40208 54832 40230
rect 24394 40168 24400 40180
rect 24355 40140 24400 40168
rect 24394 40128 24400 40140
rect 24452 40128 24458 40180
rect 25038 40168 25044 40180
rect 24999 40140 25044 40168
rect 25038 40128 25044 40140
rect 25096 40128 25102 40180
rect 25498 40128 25504 40180
rect 25556 40168 25562 40180
rect 26234 40168 26240 40180
rect 25556 40140 26240 40168
rect 25556 40128 25562 40140
rect 26234 40128 26240 40140
rect 26292 40128 26298 40180
rect 26694 40128 26700 40180
rect 26752 40168 26758 40180
rect 26752 40140 27292 40168
rect 26752 40128 26758 40140
rect 25056 40100 25084 40128
rect 24964 40072 25084 40100
rect 2133 40035 2191 40041
rect 2133 40001 2145 40035
rect 2179 40032 2191 40035
rect 23382 40032 23388 40044
rect 2179 40004 23388 40032
rect 2179 40001 2191 40004
rect 2133 39995 2191 40001
rect 23382 39992 23388 40004
rect 23440 39992 23446 40044
rect 23842 40032 23848 40044
rect 23803 40004 23848 40032
rect 23842 39992 23848 40004
rect 23900 39992 23906 40044
rect 2409 39967 2467 39973
rect 2409 39933 2421 39967
rect 2455 39964 2467 39967
rect 2774 39964 2780 39976
rect 2455 39936 2780 39964
rect 2455 39933 2467 39936
rect 2409 39927 2467 39933
rect 2774 39924 2780 39936
rect 2832 39964 2838 39976
rect 2869 39967 2927 39973
rect 2869 39964 2881 39967
rect 2832 39936 2881 39964
rect 2832 39924 2838 39936
rect 2869 39933 2881 39936
rect 2915 39933 2927 39967
rect 2869 39927 2927 39933
rect 19334 39924 19340 39976
rect 19392 39964 19398 39976
rect 23860 39964 23888 39992
rect 19392 39936 23888 39964
rect 24964 39964 24992 40072
rect 25682 40060 25688 40112
rect 25740 40100 25746 40112
rect 27264 40100 27292 40140
rect 28442 40128 28448 40180
rect 28500 40168 28506 40180
rect 28902 40168 28908 40180
rect 28500 40140 28908 40168
rect 28500 40128 28506 40140
rect 28902 40128 28908 40140
rect 28960 40168 28966 40180
rect 28960 40140 29868 40168
rect 28960 40128 28966 40140
rect 27525 40103 27583 40109
rect 27525 40100 27537 40103
rect 25740 40072 27200 40100
rect 27264 40072 27537 40100
rect 25740 40060 25746 40072
rect 25038 39992 25044 40044
rect 25096 40032 25102 40044
rect 25593 40035 25651 40041
rect 25593 40032 25605 40035
rect 25096 40004 25605 40032
rect 25096 39992 25102 40004
rect 25593 40001 25605 40004
rect 25639 40032 25651 40035
rect 26142 40032 26148 40044
rect 25639 40004 26148 40032
rect 25639 40001 25651 40004
rect 25593 39995 25651 40001
rect 26142 39992 26148 40004
rect 26200 39992 26206 40044
rect 26326 39992 26332 40044
rect 26384 40032 26390 40044
rect 26421 40035 26479 40041
rect 26421 40032 26433 40035
rect 26384 40004 26433 40032
rect 26384 39992 26390 40004
rect 26421 40001 26433 40004
rect 26467 40001 26479 40035
rect 26421 39995 26479 40001
rect 26510 39992 26516 40044
rect 26568 40032 26574 40044
rect 27172 40041 27200 40072
rect 27525 40069 27537 40072
rect 27571 40069 27583 40103
rect 27525 40063 27583 40069
rect 27798 40060 27804 40112
rect 27856 40100 27862 40112
rect 29730 40100 29736 40112
rect 27856 40072 28856 40100
rect 27856 40060 27862 40072
rect 27338 40041 27344 40044
rect 26605 40035 26663 40041
rect 26605 40032 26617 40035
rect 26568 40004 26617 40032
rect 26568 39992 26574 40004
rect 26605 40001 26617 40004
rect 26651 40001 26663 40035
rect 26605 39995 26663 40001
rect 27157 40035 27215 40041
rect 27157 40001 27169 40035
rect 27203 40001 27215 40035
rect 27157 39995 27215 40001
rect 27305 40035 27344 40041
rect 27305 40001 27317 40035
rect 27305 39995 27344 40001
rect 25774 39964 25780 39976
rect 24964 39936 25780 39964
rect 19392 39924 19398 39936
rect 25774 39924 25780 39936
rect 25832 39924 25838 39976
rect 26620 39964 26648 39995
rect 27338 39992 27344 39995
rect 27396 39992 27402 40044
rect 27430 39992 27436 40044
rect 27488 40032 27494 40044
rect 27663 40035 27721 40041
rect 27488 40004 27533 40032
rect 27488 39992 27494 40004
rect 27663 40001 27675 40035
rect 27709 40032 27721 40035
rect 28074 40032 28080 40044
rect 27709 40004 28080 40032
rect 27709 40001 27721 40004
rect 27663 39995 27721 40001
rect 28074 39992 28080 40004
rect 28132 39992 28138 40044
rect 28166 39992 28172 40044
rect 28224 40032 28230 40044
rect 28828 40041 28856 40072
rect 29104 40072 29736 40100
rect 29104 40041 29132 40072
rect 29730 40060 29736 40072
rect 29788 40060 29794 40112
rect 29840 40041 29868 40140
rect 30098 40128 30104 40180
rect 30156 40128 30162 40180
rect 32490 40168 32496 40180
rect 30208 40140 32496 40168
rect 30116 40100 30144 40128
rect 30208 40109 30236 40140
rect 32490 40128 32496 40140
rect 32548 40128 32554 40180
rect 35805 40171 35863 40177
rect 35805 40168 35817 40171
rect 32601 40140 35817 40168
rect 30024 40072 30144 40100
rect 30193 40103 30251 40109
rect 30024 40041 30052 40072
rect 30193 40069 30205 40103
rect 30239 40069 30251 40103
rect 31294 40100 31300 40112
rect 31255 40072 31300 40100
rect 30193 40063 30251 40069
rect 31294 40060 31300 40072
rect 31352 40060 31358 40112
rect 32601 40109 32629 40140
rect 35805 40137 35817 40140
rect 35851 40168 35863 40171
rect 35851 40140 38654 40168
rect 35851 40137 35863 40140
rect 35805 40131 35863 40137
rect 32585 40103 32643 40109
rect 32585 40069 32597 40103
rect 32631 40069 32643 40103
rect 33226 40100 33232 40112
rect 32585 40063 32643 40069
rect 32692 40072 33232 40100
rect 28721 40035 28779 40041
rect 28721 40032 28733 40035
rect 28224 40004 28733 40032
rect 28224 39992 28230 40004
rect 28721 40001 28733 40004
rect 28767 40001 28779 40035
rect 28721 39995 28779 40001
rect 28813 40035 28871 40041
rect 28813 40001 28825 40035
rect 28859 40001 28871 40035
rect 28813 39995 28871 40001
rect 28997 40035 29055 40041
rect 28997 40001 29009 40035
rect 29043 40001 29055 40035
rect 28997 39995 29055 40001
rect 29089 40035 29147 40041
rect 29089 40001 29101 40035
rect 29135 40001 29147 40035
rect 29089 39995 29147 40001
rect 29825 40035 29883 40041
rect 29825 40001 29837 40035
rect 29871 40001 29883 40035
rect 29825 39995 29883 40001
rect 29973 40035 30052 40041
rect 29973 40001 29985 40035
rect 30019 40004 30052 40035
rect 30101 40035 30159 40041
rect 30019 40001 30031 40004
rect 29973 39995 30031 40001
rect 30101 40001 30113 40035
rect 30147 40001 30159 40035
rect 30101 39995 30159 40001
rect 30331 40035 30389 40041
rect 30331 40001 30343 40035
rect 30377 40032 30389 40035
rect 30558 40032 30564 40044
rect 30377 40004 30564 40032
rect 30377 40001 30389 40004
rect 30331 39995 30389 40001
rect 28442 39964 28448 39976
rect 26620 39936 28448 39964
rect 28442 39924 28448 39936
rect 28500 39924 28506 39976
rect 22738 39856 22744 39908
rect 22796 39896 22802 39908
rect 23293 39899 23351 39905
rect 23293 39896 23305 39899
rect 22796 39868 23305 39896
rect 22796 39856 22802 39868
rect 23293 39865 23305 39868
rect 23339 39865 23351 39899
rect 28350 39896 28356 39908
rect 23293 39859 23351 39865
rect 25700 39868 28356 39896
rect 17218 39788 17224 39840
rect 17276 39828 17282 39840
rect 22833 39831 22891 39837
rect 22833 39828 22845 39831
rect 17276 39800 22845 39828
rect 17276 39788 17282 39800
rect 22833 39797 22845 39800
rect 22879 39828 22891 39831
rect 25222 39828 25228 39840
rect 22879 39800 25228 39828
rect 22879 39797 22891 39800
rect 22833 39791 22891 39797
rect 25222 39788 25228 39800
rect 25280 39788 25286 39840
rect 25406 39788 25412 39840
rect 25464 39828 25470 39840
rect 25700 39837 25728 39868
rect 28350 39856 28356 39868
rect 28408 39856 28414 39908
rect 28736 39896 28764 39995
rect 29012 39964 29040 39995
rect 29454 39964 29460 39976
rect 29012 39936 29460 39964
rect 29454 39924 29460 39936
rect 29512 39924 29518 39976
rect 30116 39964 30144 39995
rect 30558 39992 30564 40004
rect 30616 39992 30622 40044
rect 31478 40032 31484 40044
rect 31439 40004 31484 40032
rect 31478 39992 31484 40004
rect 31536 39992 31542 40044
rect 32490 40041 32496 40044
rect 32488 40032 32496 40041
rect 32451 40004 32496 40032
rect 32488 39995 32496 40004
rect 32490 39992 32496 39995
rect 32548 39992 32554 40044
rect 32692 40041 32720 40072
rect 33226 40060 33232 40072
rect 33284 40060 33290 40112
rect 33413 40103 33471 40109
rect 33413 40069 33425 40103
rect 33459 40100 33471 40103
rect 33502 40100 33508 40112
rect 33459 40072 33508 40100
rect 33459 40069 33471 40072
rect 33413 40063 33471 40069
rect 33502 40060 33508 40072
rect 33560 40060 33566 40112
rect 33597 40103 33655 40109
rect 33597 40069 33609 40103
rect 33643 40100 33655 40103
rect 33962 40100 33968 40112
rect 33643 40072 33968 40100
rect 33643 40069 33655 40072
rect 33597 40063 33655 40069
rect 33962 40060 33968 40072
rect 34020 40100 34026 40112
rect 34020 40072 34100 40100
rect 34020 40060 34026 40072
rect 32858 40041 32864 40044
rect 32677 40035 32735 40041
rect 32677 40001 32689 40035
rect 32723 40001 32735 40035
rect 32677 39995 32735 40001
rect 32815 40035 32864 40041
rect 32815 40001 32827 40035
rect 32861 40001 32864 40035
rect 32815 39995 32864 40001
rect 30190 39964 30196 39976
rect 30116 39936 30196 39964
rect 28902 39896 28908 39908
rect 28736 39868 28908 39896
rect 28902 39856 28908 39868
rect 28960 39896 28966 39908
rect 30116 39896 30144 39936
rect 30190 39924 30196 39936
rect 30248 39924 30254 39976
rect 31846 39924 31852 39976
rect 31904 39964 31910 39976
rect 32692 39964 32720 39995
rect 32858 39992 32864 39995
rect 32916 39992 32922 40044
rect 32964 40035 33022 40041
rect 32964 40001 32976 40035
rect 33010 40032 33022 40035
rect 34072 40032 34100 40072
rect 34146 40060 34152 40112
rect 34204 40100 34210 40112
rect 34241 40103 34299 40109
rect 34241 40100 34253 40103
rect 34204 40072 34253 40100
rect 34204 40060 34210 40072
rect 34241 40069 34253 40072
rect 34287 40069 34299 40103
rect 34241 40063 34299 40069
rect 34425 40035 34483 40041
rect 34425 40032 34437 40035
rect 33010 40004 33088 40032
rect 34072 40004 34437 40032
rect 33010 40001 33022 40004
rect 32964 39995 33022 40001
rect 31904 39936 32720 39964
rect 31904 39924 31910 39936
rect 28960 39868 30144 39896
rect 28960 39856 28966 39868
rect 30926 39856 30932 39908
rect 30984 39896 30990 39908
rect 33060 39896 33088 40004
rect 34425 40001 34437 40004
rect 34471 40001 34483 40035
rect 34425 39995 34483 40001
rect 34609 40035 34667 40041
rect 34609 40001 34621 40035
rect 34655 40032 34667 40035
rect 35161 40035 35219 40041
rect 35161 40032 35173 40035
rect 34655 40004 35173 40032
rect 34655 40001 34667 40004
rect 34609 39995 34667 40001
rect 35161 40001 35173 40004
rect 35207 40001 35219 40035
rect 38626 40032 38654 40140
rect 46106 40032 46112 40044
rect 38626 40004 46112 40032
rect 35161 39995 35219 40001
rect 46106 39992 46112 40004
rect 46164 39992 46170 40044
rect 53745 40035 53803 40041
rect 53745 40032 53757 40035
rect 46216 40004 53757 40032
rect 35526 39924 35532 39976
rect 35584 39964 35590 39976
rect 46216 39964 46244 40004
rect 53745 40001 53757 40004
rect 53791 40001 53803 40035
rect 53745 39995 53803 40001
rect 35584 39936 46244 39964
rect 51813 39967 51871 39973
rect 35584 39924 35590 39936
rect 51813 39933 51825 39967
rect 51859 39964 51871 39967
rect 53469 39967 53527 39973
rect 53469 39964 53481 39967
rect 51859 39936 53481 39964
rect 51859 39933 51871 39936
rect 51813 39927 51871 39933
rect 53469 39933 53481 39936
rect 53515 39964 53527 39967
rect 53558 39964 53564 39976
rect 53515 39936 53564 39964
rect 53515 39933 53527 39936
rect 53469 39927 53527 39933
rect 53558 39924 53564 39936
rect 53616 39924 53622 39976
rect 30984 39868 33088 39896
rect 35345 39899 35403 39905
rect 30984 39856 30990 39868
rect 35345 39865 35357 39899
rect 35391 39896 35403 39899
rect 36078 39896 36084 39908
rect 35391 39868 36084 39896
rect 35391 39865 35403 39868
rect 35345 39859 35403 39865
rect 36078 39856 36084 39868
rect 36136 39856 36142 39908
rect 52365 39899 52423 39905
rect 52365 39865 52377 39899
rect 52411 39896 52423 39899
rect 53650 39896 53656 39908
rect 52411 39868 53656 39896
rect 52411 39865 52423 39868
rect 52365 39859 52423 39865
rect 53650 39856 53656 39868
rect 53708 39856 53714 39908
rect 25685 39831 25743 39837
rect 25685 39828 25697 39831
rect 25464 39800 25697 39828
rect 25464 39788 25470 39800
rect 25685 39797 25697 39800
rect 25731 39797 25743 39831
rect 25685 39791 25743 39797
rect 26237 39831 26295 39837
rect 26237 39797 26249 39831
rect 26283 39828 26295 39831
rect 27522 39828 27528 39840
rect 26283 39800 27528 39828
rect 26283 39797 26295 39800
rect 26237 39791 26295 39797
rect 27522 39788 27528 39800
rect 27580 39788 27586 39840
rect 27798 39828 27804 39840
rect 27759 39800 27804 39828
rect 27798 39788 27804 39800
rect 27856 39788 27862 39840
rect 28537 39831 28595 39837
rect 28537 39797 28549 39831
rect 28583 39828 28595 39831
rect 28994 39828 29000 39840
rect 28583 39800 29000 39828
rect 28583 39797 28595 39800
rect 28537 39791 28595 39797
rect 28994 39788 29000 39800
rect 29052 39788 29058 39840
rect 30466 39828 30472 39840
rect 30427 39800 30472 39828
rect 30466 39788 30472 39800
rect 30524 39788 30530 39840
rect 31662 39828 31668 39840
rect 31623 39800 31668 39828
rect 31662 39788 31668 39800
rect 31720 39788 31726 39840
rect 32306 39828 32312 39840
rect 32267 39800 32312 39828
rect 32306 39788 32312 39800
rect 32364 39788 32370 39840
rect 32674 39788 32680 39840
rect 32732 39828 32738 39840
rect 33781 39831 33839 39837
rect 33781 39828 33793 39831
rect 32732 39800 33793 39828
rect 32732 39788 32738 39800
rect 33781 39797 33793 39800
rect 33827 39797 33839 39831
rect 33781 39791 33839 39797
rect 53009 39831 53067 39837
rect 53009 39797 53021 39831
rect 53055 39828 53067 39831
rect 53374 39828 53380 39840
rect 53055 39800 53380 39828
rect 53055 39797 53067 39800
rect 53009 39791 53067 39797
rect 53374 39788 53380 39800
rect 53432 39788 53438 39840
rect 1104 39738 54832 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 54832 39738
rect 1104 39664 54832 39686
rect 22186 39584 22192 39636
rect 22244 39624 22250 39636
rect 22281 39627 22339 39633
rect 22281 39624 22293 39627
rect 22244 39596 22293 39624
rect 22244 39584 22250 39596
rect 22281 39593 22293 39596
rect 22327 39624 22339 39627
rect 25682 39624 25688 39636
rect 22327 39596 25549 39624
rect 25643 39596 25688 39624
rect 22327 39593 22339 39596
rect 22281 39587 22339 39593
rect 24578 39556 24584 39568
rect 6886 39528 24584 39556
rect 2133 39491 2191 39497
rect 2133 39457 2145 39491
rect 2179 39488 2191 39491
rect 6886 39488 6914 39528
rect 24578 39516 24584 39528
rect 24636 39516 24642 39568
rect 2179 39460 6914 39488
rect 22925 39491 22983 39497
rect 2179 39457 2191 39460
rect 2133 39451 2191 39457
rect 22925 39457 22937 39491
rect 22971 39488 22983 39491
rect 25314 39488 25320 39500
rect 22971 39460 25320 39488
rect 22971 39457 22983 39460
rect 22925 39451 22983 39457
rect 25314 39448 25320 39460
rect 25372 39448 25378 39500
rect 25521 39488 25549 39596
rect 25682 39584 25688 39596
rect 25740 39584 25746 39636
rect 27614 39584 27620 39636
rect 27672 39624 27678 39636
rect 28166 39624 28172 39636
rect 27672 39596 28172 39624
rect 27672 39584 27678 39596
rect 28166 39584 28172 39596
rect 28224 39584 28230 39636
rect 31386 39584 31392 39636
rect 31444 39624 31450 39636
rect 31444 39596 41414 39624
rect 31444 39584 31450 39596
rect 26234 39516 26240 39568
rect 26292 39556 26298 39568
rect 34422 39556 34428 39568
rect 26292 39528 34428 39556
rect 26292 39516 26298 39528
rect 25521 39460 25636 39488
rect 2409 39423 2467 39429
rect 2409 39389 2421 39423
rect 2455 39420 2467 39423
rect 2774 39420 2780 39432
rect 2455 39392 2780 39420
rect 2455 39389 2467 39392
rect 2409 39383 2467 39389
rect 2774 39380 2780 39392
rect 2832 39420 2838 39432
rect 2869 39423 2927 39429
rect 2869 39420 2881 39423
rect 2832 39392 2881 39420
rect 2832 39380 2838 39392
rect 2869 39389 2881 39392
rect 2915 39389 2927 39423
rect 25038 39420 25044 39432
rect 24999 39392 25044 39420
rect 2869 39383 2927 39389
rect 25038 39380 25044 39392
rect 25096 39380 25102 39432
rect 25134 39423 25192 39429
rect 25134 39389 25146 39423
rect 25180 39389 25192 39423
rect 25134 39383 25192 39389
rect 22922 39312 22928 39364
rect 22980 39352 22986 39364
rect 25148 39352 25176 39383
rect 25222 39380 25228 39432
rect 25280 39420 25286 39432
rect 25409 39423 25467 39429
rect 25409 39420 25421 39423
rect 25280 39392 25421 39420
rect 25280 39380 25286 39392
rect 25409 39389 25421 39392
rect 25455 39389 25467 39423
rect 25409 39383 25467 39389
rect 25506 39423 25564 39429
rect 25506 39389 25518 39423
rect 25552 39389 25564 39423
rect 25506 39383 25564 39389
rect 25314 39352 25320 39364
rect 22980 39324 25176 39352
rect 25275 39324 25320 39352
rect 22980 39312 22986 39324
rect 25314 39312 25320 39324
rect 25372 39312 25378 39364
rect 23474 39284 23480 39296
rect 23435 39256 23480 39284
rect 23474 39244 23480 39256
rect 23532 39244 23538 39296
rect 23934 39284 23940 39296
rect 23895 39256 23940 39284
rect 23934 39244 23940 39256
rect 23992 39244 23998 39296
rect 24302 39244 24308 39296
rect 24360 39284 24366 39296
rect 25222 39284 25228 39296
rect 24360 39256 25228 39284
rect 24360 39244 24366 39256
rect 25222 39244 25228 39256
rect 25280 39284 25286 39296
rect 25516 39284 25544 39383
rect 25608 39352 25636 39460
rect 25958 39448 25964 39500
rect 26016 39488 26022 39500
rect 27246 39488 27252 39500
rect 26016 39460 26556 39488
rect 26016 39448 26022 39460
rect 26142 39420 26148 39432
rect 26103 39392 26148 39420
rect 26142 39380 26148 39392
rect 26200 39380 26206 39432
rect 26528 39429 26556 39460
rect 26896 39460 27252 39488
rect 26238 39423 26296 39429
rect 26238 39389 26250 39423
rect 26284 39389 26296 39423
rect 26238 39383 26296 39389
rect 26513 39423 26571 39429
rect 26513 39389 26525 39423
rect 26559 39389 26571 39423
rect 26513 39383 26571 39389
rect 26610 39423 26668 39429
rect 26610 39389 26622 39423
rect 26656 39420 26668 39423
rect 26896 39420 26924 39460
rect 27246 39448 27252 39460
rect 27304 39448 27310 39500
rect 26656 39392 26924 39420
rect 26656 39389 26668 39392
rect 26610 39383 26668 39389
rect 26253 39352 26281 39383
rect 27062 39380 27068 39432
rect 27120 39420 27126 39432
rect 27338 39420 27344 39432
rect 27120 39392 27344 39420
rect 27120 39380 27126 39392
rect 27338 39380 27344 39392
rect 27396 39420 27402 39432
rect 27525 39423 27583 39429
rect 27525 39420 27537 39423
rect 27396 39392 27537 39420
rect 27396 39380 27402 39392
rect 27525 39389 27537 39392
rect 27571 39389 27583 39423
rect 27706 39420 27712 39432
rect 27667 39392 27712 39420
rect 27525 39383 27583 39389
rect 27706 39380 27712 39392
rect 27764 39380 27770 39432
rect 27908 39429 27936 39528
rect 34422 39516 34428 39528
rect 34480 39516 34486 39568
rect 41386 39556 41414 39596
rect 46106 39584 46112 39636
rect 46164 39624 46170 39636
rect 52825 39627 52883 39633
rect 52825 39624 52837 39627
rect 46164 39596 52837 39624
rect 46164 39584 46170 39596
rect 52825 39593 52837 39596
rect 52871 39593 52883 39627
rect 52825 39587 52883 39593
rect 53742 39556 53748 39568
rect 41386 39528 53748 39556
rect 53742 39516 53748 39528
rect 53800 39516 53806 39568
rect 32674 39488 32680 39500
rect 30668 39460 32680 39488
rect 27893 39423 27951 39429
rect 27893 39389 27905 39423
rect 27939 39389 27951 39423
rect 27893 39383 27951 39389
rect 28258 39380 28264 39432
rect 28316 39420 28322 39432
rect 28353 39423 28411 39429
rect 28353 39420 28365 39423
rect 28316 39392 28365 39420
rect 28316 39380 28322 39392
rect 28353 39389 28365 39392
rect 28399 39389 28411 39423
rect 28353 39383 28411 39389
rect 28537 39423 28595 39429
rect 28537 39389 28549 39423
rect 28583 39420 28595 39423
rect 29086 39420 29092 39432
rect 28583 39392 29092 39420
rect 28583 39389 28595 39392
rect 28537 39383 28595 39389
rect 29086 39380 29092 39392
rect 29144 39420 29150 39432
rect 29270 39420 29276 39432
rect 29144 39392 29276 39420
rect 29144 39380 29150 39392
rect 29270 39380 29276 39392
rect 29328 39420 29334 39432
rect 30558 39420 30564 39432
rect 29328 39392 30564 39420
rect 29328 39380 29334 39392
rect 30558 39380 30564 39392
rect 30616 39380 30622 39432
rect 30668 39429 30696 39460
rect 32674 39448 32680 39460
rect 32732 39448 32738 39500
rect 33594 39448 33600 39500
rect 33652 39488 33658 39500
rect 34149 39491 34207 39497
rect 34149 39488 34161 39491
rect 33652 39460 34161 39488
rect 33652 39448 33658 39460
rect 34149 39457 34161 39460
rect 34195 39488 34207 39491
rect 46290 39488 46296 39500
rect 34195 39460 46296 39488
rect 34195 39457 34207 39460
rect 34149 39451 34207 39457
rect 46290 39448 46296 39460
rect 46348 39448 46354 39500
rect 30653 39423 30711 39429
rect 30653 39389 30665 39423
rect 30699 39389 30711 39423
rect 30653 39383 30711 39389
rect 31573 39423 31631 39429
rect 31573 39389 31585 39423
rect 31619 39420 31631 39423
rect 32306 39420 32312 39432
rect 31619 39392 32312 39420
rect 31619 39389 31631 39392
rect 31573 39383 31631 39389
rect 32306 39380 32312 39392
rect 32364 39380 32370 39432
rect 32398 39380 32404 39432
rect 32456 39420 32462 39432
rect 32493 39423 32551 39429
rect 32493 39420 32505 39423
rect 32456 39392 32505 39420
rect 32456 39380 32462 39392
rect 32493 39389 32505 39392
rect 32539 39389 32551 39423
rect 32493 39383 32551 39389
rect 32858 39380 32864 39432
rect 32916 39420 32922 39432
rect 33689 39423 33747 39429
rect 32916 39392 33645 39420
rect 32916 39380 32922 39392
rect 25608 39324 26281 39352
rect 26421 39355 26479 39361
rect 26421 39321 26433 39355
rect 26467 39321 26479 39355
rect 26421 39315 26479 39321
rect 25280 39256 25544 39284
rect 25280 39244 25286 39256
rect 26050 39244 26056 39296
rect 26108 39284 26114 39296
rect 26436 39284 26464 39315
rect 26970 39312 26976 39364
rect 27028 39352 27034 39364
rect 27617 39355 27675 39361
rect 27617 39352 27629 39355
rect 27028 39324 27629 39352
rect 27028 39312 27034 39324
rect 27617 39321 27629 39324
rect 27663 39321 27675 39355
rect 31389 39355 31447 39361
rect 31389 39352 31401 39355
rect 27617 39315 27675 39321
rect 28644 39324 31401 39352
rect 26786 39284 26792 39296
rect 26108 39256 26464 39284
rect 26747 39256 26792 39284
rect 26108 39244 26114 39256
rect 26786 39244 26792 39256
rect 26844 39244 26850 39296
rect 26878 39244 26884 39296
rect 26936 39284 26942 39296
rect 27341 39287 27399 39293
rect 27341 39284 27353 39287
rect 26936 39256 27353 39284
rect 26936 39244 26942 39256
rect 27341 39253 27353 39256
rect 27387 39253 27399 39287
rect 27341 39247 27399 39253
rect 27522 39244 27528 39296
rect 27580 39284 27586 39296
rect 28644 39284 28672 39324
rect 31389 39321 31401 39324
rect 31435 39352 31447 39355
rect 32677 39355 32735 39361
rect 32677 39352 32689 39355
rect 31435 39324 32689 39352
rect 31435 39321 31447 39324
rect 31389 39315 31447 39321
rect 32677 39321 32689 39324
rect 32723 39352 32735 39355
rect 33505 39355 33563 39361
rect 33505 39352 33517 39355
rect 32723 39324 33517 39352
rect 32723 39321 32735 39324
rect 32677 39315 32735 39321
rect 33505 39321 33517 39324
rect 33551 39321 33563 39355
rect 33505 39315 33563 39321
rect 27580 39256 28672 39284
rect 28721 39287 28779 39293
rect 27580 39244 27586 39256
rect 28721 39253 28733 39287
rect 28767 39284 28779 39287
rect 29454 39284 29460 39296
rect 28767 39256 29460 39284
rect 28767 39253 28779 39256
rect 28721 39247 28779 39253
rect 29454 39244 29460 39256
rect 29512 39244 29518 39296
rect 29730 39284 29736 39296
rect 29691 39256 29736 39284
rect 29730 39244 29736 39256
rect 29788 39244 29794 39296
rect 30561 39287 30619 39293
rect 30561 39253 30573 39287
rect 30607 39284 30619 39287
rect 30742 39284 30748 39296
rect 30607 39256 30748 39284
rect 30607 39253 30619 39256
rect 30561 39247 30619 39253
rect 30742 39244 30748 39256
rect 30800 39244 30806 39296
rect 31202 39284 31208 39296
rect 31163 39256 31208 39284
rect 31202 39244 31208 39256
rect 31260 39244 31266 39296
rect 32858 39284 32864 39296
rect 32819 39256 32864 39284
rect 32858 39244 32864 39256
rect 32916 39244 32922 39296
rect 33318 39284 33324 39296
rect 33279 39256 33324 39284
rect 33318 39244 33324 39256
rect 33376 39244 33382 39296
rect 33617 39284 33645 39392
rect 33689 39389 33701 39423
rect 33735 39420 33747 39423
rect 33778 39420 33784 39432
rect 33735 39392 33784 39420
rect 33735 39389 33747 39392
rect 33689 39383 33747 39389
rect 33778 39380 33784 39392
rect 33836 39380 33842 39432
rect 34238 39380 34244 39432
rect 34296 39420 34302 39432
rect 34977 39423 35035 39429
rect 34977 39420 34989 39423
rect 34296 39392 34989 39420
rect 34296 39380 34302 39392
rect 34977 39389 34989 39392
rect 35023 39389 35035 39423
rect 34977 39383 35035 39389
rect 52365 39423 52423 39429
rect 52365 39389 52377 39423
rect 52411 39420 52423 39423
rect 53006 39420 53012 39432
rect 52411 39392 53012 39420
rect 52411 39389 52423 39392
rect 52365 39383 52423 39389
rect 53006 39380 53012 39392
rect 53064 39380 53070 39432
rect 53466 39420 53472 39432
rect 53427 39392 53472 39420
rect 53466 39380 53472 39392
rect 53524 39380 53530 39432
rect 53650 39380 53656 39432
rect 53708 39420 53714 39432
rect 53745 39423 53803 39429
rect 53745 39420 53757 39423
rect 53708 39392 53757 39420
rect 53708 39380 53714 39392
rect 53745 39389 53757 39392
rect 53791 39389 53803 39423
rect 53745 39383 53803 39389
rect 35161 39355 35219 39361
rect 35161 39321 35173 39355
rect 35207 39352 35219 39355
rect 36538 39352 36544 39364
rect 35207 39324 36544 39352
rect 35207 39321 35219 39324
rect 35161 39315 35219 39321
rect 36538 39312 36544 39324
rect 36596 39312 36602 39364
rect 51813 39355 51871 39361
rect 51813 39321 51825 39355
rect 51859 39352 51871 39355
rect 53484 39352 53512 39380
rect 51859 39324 53512 39352
rect 51859 39321 51871 39324
rect 51813 39315 51871 39321
rect 35621 39287 35679 39293
rect 35621 39284 35633 39287
rect 33617 39256 35633 39284
rect 35621 39253 35633 39256
rect 35667 39284 35679 39287
rect 51074 39284 51080 39296
rect 35667 39256 51080 39284
rect 35667 39253 35679 39256
rect 35621 39247 35679 39253
rect 51074 39244 51080 39256
rect 51132 39244 51138 39296
rect 1104 39194 54832 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 54832 39194
rect 1104 39120 54832 39142
rect 11698 39040 11704 39092
rect 11756 39080 11762 39092
rect 16209 39083 16267 39089
rect 16209 39080 16221 39083
rect 11756 39052 16221 39080
rect 11756 39040 11762 39052
rect 16209 39049 16221 39052
rect 16255 39049 16267 39083
rect 16209 39043 16267 39049
rect 17405 39083 17463 39089
rect 17405 39049 17417 39083
rect 17451 39080 17463 39083
rect 22922 39080 22928 39092
rect 17451 39052 22094 39080
rect 22883 39052 22928 39080
rect 17451 39049 17463 39052
rect 17405 39043 17463 39049
rect 2133 38947 2191 38953
rect 2133 38913 2145 38947
rect 2179 38944 2191 38947
rect 16224 38944 16252 39043
rect 17129 39015 17187 39021
rect 17129 39012 17141 39015
rect 16960 38984 17141 39012
rect 16853 38947 16911 38953
rect 16853 38944 16865 38947
rect 2179 38916 6914 38944
rect 16224 38916 16865 38944
rect 2179 38913 2191 38916
rect 2133 38907 2191 38913
rect 2409 38879 2467 38885
rect 2409 38845 2421 38879
rect 2455 38876 2467 38879
rect 2774 38876 2780 38888
rect 2455 38848 2780 38876
rect 2455 38845 2467 38848
rect 2409 38839 2467 38845
rect 2774 38836 2780 38848
rect 2832 38876 2838 38888
rect 2869 38879 2927 38885
rect 2869 38876 2881 38879
rect 2832 38848 2881 38876
rect 2832 38836 2838 38848
rect 2869 38845 2881 38848
rect 2915 38845 2927 38879
rect 2869 38839 2927 38845
rect 6886 38808 6914 38916
rect 16853 38913 16865 38916
rect 16899 38913 16911 38947
rect 16853 38907 16911 38913
rect 14826 38836 14832 38888
rect 14884 38876 14890 38888
rect 16960 38876 16988 38984
rect 17129 38981 17141 38984
rect 17175 38981 17187 39015
rect 17129 38975 17187 38981
rect 17037 38947 17095 38953
rect 17037 38913 17049 38947
rect 17083 38913 17095 38947
rect 17037 38907 17095 38913
rect 17221 38947 17279 38953
rect 17221 38913 17233 38947
rect 17267 38944 17279 38947
rect 17310 38944 17316 38956
rect 17267 38916 17316 38944
rect 17267 38913 17279 38916
rect 17221 38907 17279 38913
rect 14884 38848 16988 38876
rect 17052 38876 17080 38907
rect 17310 38904 17316 38916
rect 17368 38904 17374 38956
rect 22066 38944 22094 39052
rect 22922 39040 22928 39052
rect 22980 39040 22986 39092
rect 23566 39080 23572 39092
rect 23527 39052 23572 39080
rect 23566 39040 23572 39052
rect 23624 39080 23630 39092
rect 24302 39080 24308 39092
rect 23624 39052 24308 39080
rect 23624 39040 23630 39052
rect 24302 39040 24308 39052
rect 24360 39040 24366 39092
rect 24946 39080 24952 39092
rect 24504 39052 24952 39080
rect 22738 38972 22744 39024
rect 22796 39012 22802 39024
rect 24504 39012 24532 39052
rect 24946 39040 24952 39052
rect 25004 39080 25010 39092
rect 25133 39083 25191 39089
rect 25133 39080 25145 39083
rect 25004 39052 25145 39080
rect 25004 39040 25010 39052
rect 25133 39049 25145 39052
rect 25179 39080 25191 39083
rect 26050 39080 26056 39092
rect 25179 39052 26056 39080
rect 25179 39049 25191 39052
rect 25133 39043 25191 39049
rect 26050 39040 26056 39052
rect 26108 39040 26114 39092
rect 26142 39040 26148 39092
rect 26200 39080 26206 39092
rect 27157 39083 27215 39089
rect 27157 39080 27169 39083
rect 26200 39052 27169 39080
rect 26200 39040 26206 39052
rect 27157 39049 27169 39052
rect 27203 39049 27215 39083
rect 27157 39043 27215 39049
rect 27801 39083 27859 39089
rect 27801 39049 27813 39083
rect 27847 39080 27859 39083
rect 27982 39080 27988 39092
rect 27847 39052 27988 39080
rect 27847 39049 27859 39052
rect 27801 39043 27859 39049
rect 27982 39040 27988 39052
rect 28040 39040 28046 39092
rect 28902 39040 28908 39092
rect 28960 39080 28966 39092
rect 30469 39083 30527 39089
rect 28960 39052 29132 39080
rect 28960 39040 28966 39052
rect 22796 38984 24532 39012
rect 22796 38972 22802 38984
rect 24578 38972 24584 39024
rect 24636 39012 24642 39024
rect 29104 39021 29132 39052
rect 30469 39049 30481 39083
rect 30515 39080 30527 39083
rect 30650 39080 30656 39092
rect 30515 39052 30656 39080
rect 30515 39049 30527 39052
rect 30469 39043 30527 39049
rect 30650 39040 30656 39052
rect 30708 39040 30714 39092
rect 29089 39015 29147 39021
rect 24636 38984 28949 39012
rect 24636 38972 24642 38984
rect 26421 38947 26479 38953
rect 26421 38944 26433 38947
rect 22066 38916 26433 38944
rect 26421 38913 26433 38916
rect 26467 38913 26479 38947
rect 26602 38944 26608 38956
rect 26563 38916 26608 38944
rect 26421 38907 26479 38913
rect 26602 38904 26608 38916
rect 26660 38904 26666 38956
rect 27522 38944 27528 38956
rect 27483 38916 27528 38944
rect 27522 38904 27528 38916
rect 27580 38904 27586 38956
rect 27614 38904 27620 38956
rect 27672 38944 27678 38956
rect 27893 38947 27951 38953
rect 27893 38944 27905 38947
rect 27672 38916 27905 38944
rect 27672 38904 27678 38916
rect 27893 38913 27905 38916
rect 27939 38944 27951 38947
rect 28258 38944 28264 38956
rect 27939 38916 28264 38944
rect 27939 38913 27951 38916
rect 27893 38907 27951 38913
rect 28258 38904 28264 38916
rect 28316 38904 28322 38956
rect 28350 38904 28356 38956
rect 28408 38944 28414 38956
rect 28810 38944 28816 38956
rect 28408 38916 28816 38944
rect 28408 38904 28414 38916
rect 28810 38904 28816 38916
rect 28868 38904 28874 38956
rect 28921 38953 28949 38984
rect 29089 38981 29101 39015
rect 29135 38981 29147 39015
rect 29089 38975 29147 38981
rect 29181 39015 29239 39021
rect 29181 38981 29193 39015
rect 29227 39012 29239 39015
rect 29638 39012 29644 39024
rect 29227 38984 29644 39012
rect 29227 38981 29239 38984
rect 29181 38975 29239 38981
rect 29638 38972 29644 38984
rect 29696 38972 29702 39024
rect 29730 38972 29736 39024
rect 29788 39012 29794 39024
rect 30558 39012 30564 39024
rect 29788 38984 30564 39012
rect 29788 38972 29794 38984
rect 30558 38972 30564 38984
rect 30616 38972 30622 39024
rect 31662 39012 31668 39024
rect 31623 38984 31668 39012
rect 31662 38972 31668 38984
rect 31720 38972 31726 39024
rect 32766 38972 32772 39024
rect 32824 39012 32830 39024
rect 32861 39015 32919 39021
rect 32861 39012 32873 39015
rect 32824 38984 32873 39012
rect 32824 38972 32830 38984
rect 32861 38981 32873 38984
rect 32907 38981 32919 39015
rect 32861 38975 32919 38981
rect 33045 39015 33103 39021
rect 33045 38981 33057 39015
rect 33091 39012 33103 39015
rect 33686 39012 33692 39024
rect 33091 38984 33692 39012
rect 33091 38981 33103 38984
rect 33045 38975 33103 38981
rect 28906 38947 28964 38953
rect 28906 38913 28918 38947
rect 28952 38913 28964 38947
rect 28906 38907 28964 38913
rect 29270 38904 29276 38956
rect 29328 38953 29334 38956
rect 29328 38944 29336 38953
rect 29328 38916 29373 38944
rect 29328 38907 29336 38916
rect 29328 38904 29334 38907
rect 29454 38904 29460 38956
rect 29512 38944 29518 38956
rect 33060 38944 33088 38975
rect 33686 38972 33692 38984
rect 33744 38972 33750 39024
rect 33870 39012 33876 39024
rect 33831 38984 33876 39012
rect 33870 38972 33876 38984
rect 33928 38972 33934 39024
rect 29512 38916 33088 38944
rect 33229 38947 33287 38953
rect 29512 38904 29518 38916
rect 33229 38913 33241 38947
rect 33275 38944 33287 38947
rect 34517 38947 34575 38953
rect 34517 38944 34529 38947
rect 33275 38916 34529 38944
rect 33275 38913 33287 38916
rect 33229 38907 33287 38913
rect 34517 38913 34529 38916
rect 34563 38913 34575 38947
rect 52086 38944 52092 38956
rect 52047 38916 52092 38944
rect 34517 38907 34575 38913
rect 52086 38904 52092 38916
rect 52144 38904 52150 38956
rect 53745 38947 53803 38953
rect 53745 38944 53757 38947
rect 52196 38916 53757 38944
rect 17957 38879 18015 38885
rect 17957 38876 17969 38879
rect 17052 38848 17969 38876
rect 14884 38836 14890 38848
rect 17957 38845 17969 38848
rect 18003 38876 18015 38879
rect 23014 38876 23020 38888
rect 18003 38848 23020 38876
rect 18003 38845 18015 38848
rect 17957 38839 18015 38845
rect 23014 38836 23020 38848
rect 23072 38836 23078 38888
rect 29730 38876 29736 38888
rect 23860 38848 29736 38876
rect 23860 38808 23888 38848
rect 29730 38836 29736 38848
rect 29788 38836 29794 38888
rect 52196 38876 52224 38916
rect 53745 38913 53757 38916
rect 53791 38913 53803 38947
rect 53745 38907 53803 38913
rect 29932 38848 52224 38876
rect 52365 38879 52423 38885
rect 6886 38780 23888 38808
rect 23934 38768 23940 38820
rect 23992 38808 23998 38820
rect 26970 38808 26976 38820
rect 23992 38780 26976 38808
rect 23992 38768 23998 38780
rect 26970 38768 26976 38780
rect 27028 38768 27034 38820
rect 28718 38768 28724 38820
rect 28776 38808 28782 38820
rect 28776 38780 29776 38808
rect 28776 38768 28782 38780
rect 29748 38752 29776 38780
rect 24121 38743 24179 38749
rect 24121 38709 24133 38743
rect 24167 38740 24179 38743
rect 24394 38740 24400 38752
rect 24167 38712 24400 38740
rect 24167 38709 24179 38712
rect 24121 38703 24179 38709
rect 24394 38700 24400 38712
rect 24452 38740 24458 38752
rect 24854 38740 24860 38752
rect 24452 38712 24860 38740
rect 24452 38700 24458 38712
rect 24854 38700 24860 38712
rect 24912 38700 24918 38752
rect 25314 38700 25320 38752
rect 25372 38740 25378 38752
rect 25498 38740 25504 38752
rect 25372 38712 25504 38740
rect 25372 38700 25378 38712
rect 25498 38700 25504 38712
rect 25556 38700 25562 38752
rect 25777 38743 25835 38749
rect 25777 38709 25789 38743
rect 25823 38740 25835 38743
rect 25866 38740 25872 38752
rect 25823 38712 25872 38740
rect 25823 38709 25835 38712
rect 25777 38703 25835 38709
rect 25866 38700 25872 38712
rect 25924 38740 25930 38752
rect 26050 38740 26056 38752
rect 25924 38712 26056 38740
rect 25924 38700 25930 38712
rect 26050 38700 26056 38712
rect 26108 38700 26114 38752
rect 26234 38740 26240 38752
rect 26195 38712 26240 38740
rect 26234 38700 26240 38712
rect 26292 38700 26298 38752
rect 26605 38743 26663 38749
rect 26605 38709 26617 38743
rect 26651 38740 26663 38743
rect 26878 38740 26884 38752
rect 26651 38712 26884 38740
rect 26651 38709 26663 38712
rect 26605 38703 26663 38709
rect 26878 38700 26884 38712
rect 26936 38700 26942 38752
rect 27246 38700 27252 38752
rect 27304 38740 27310 38752
rect 27433 38743 27491 38749
rect 27433 38740 27445 38743
rect 27304 38712 27445 38740
rect 27304 38700 27310 38712
rect 27433 38709 27445 38712
rect 27479 38709 27491 38743
rect 27433 38703 27491 38709
rect 27617 38743 27675 38749
rect 27617 38709 27629 38743
rect 27663 38740 27675 38743
rect 27982 38740 27988 38752
rect 27663 38712 27988 38740
rect 27663 38709 27675 38712
rect 27617 38703 27675 38709
rect 27982 38700 27988 38712
rect 28040 38700 28046 38752
rect 29362 38700 29368 38752
rect 29420 38740 29426 38752
rect 29457 38743 29515 38749
rect 29457 38740 29469 38743
rect 29420 38712 29469 38740
rect 29420 38700 29426 38712
rect 29457 38709 29469 38712
rect 29503 38709 29515 38743
rect 29457 38703 29515 38709
rect 29730 38700 29736 38752
rect 29788 38700 29794 38752
rect 29822 38700 29828 38752
rect 29880 38740 29886 38752
rect 29932 38749 29960 38848
rect 52365 38845 52377 38879
rect 52411 38876 52423 38879
rect 52411 38848 53052 38876
rect 52411 38845 52423 38848
rect 52365 38839 52423 38845
rect 34701 38811 34759 38817
rect 34701 38777 34713 38811
rect 34747 38808 34759 38811
rect 35986 38808 35992 38820
rect 34747 38780 35992 38808
rect 34747 38777 34759 38780
rect 34701 38771 34759 38777
rect 35986 38768 35992 38780
rect 36044 38768 36050 38820
rect 53024 38752 53052 38848
rect 53374 38836 53380 38888
rect 53432 38876 53438 38888
rect 53469 38879 53527 38885
rect 53469 38876 53481 38879
rect 53432 38848 53481 38876
rect 53432 38836 53438 38848
rect 53469 38845 53481 38848
rect 53515 38845 53527 38879
rect 53469 38839 53527 38845
rect 29917 38743 29975 38749
rect 29917 38740 29929 38743
rect 29880 38712 29929 38740
rect 29880 38700 29886 38712
rect 29917 38709 29929 38712
rect 29963 38709 29975 38743
rect 29917 38703 29975 38709
rect 31573 38743 31631 38749
rect 31573 38709 31585 38743
rect 31619 38740 31631 38743
rect 32030 38740 32036 38752
rect 31619 38712 32036 38740
rect 31619 38709 31631 38712
rect 31573 38703 31631 38709
rect 32030 38700 32036 38712
rect 32088 38700 32094 38752
rect 32122 38700 32128 38752
rect 32180 38740 32186 38752
rect 32309 38743 32367 38749
rect 32309 38740 32321 38743
rect 32180 38712 32321 38740
rect 32180 38700 32186 38712
rect 32309 38709 32321 38712
rect 32355 38709 32367 38743
rect 32309 38703 32367 38709
rect 33781 38743 33839 38749
rect 33781 38709 33793 38743
rect 33827 38740 33839 38743
rect 34514 38740 34520 38752
rect 33827 38712 34520 38740
rect 33827 38709 33839 38712
rect 33781 38703 33839 38709
rect 34514 38700 34520 38712
rect 34572 38700 34578 38752
rect 53006 38740 53012 38752
rect 52967 38712 53012 38740
rect 53006 38700 53012 38712
rect 53064 38700 53070 38752
rect 1104 38650 54832 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 54832 38650
rect 1104 38576 54832 38598
rect 24854 38536 24860 38548
rect 24815 38508 24860 38536
rect 24854 38496 24860 38508
rect 24912 38496 24918 38548
rect 26973 38539 27031 38545
rect 26973 38505 26985 38539
rect 27019 38536 27031 38539
rect 27246 38536 27252 38548
rect 27019 38508 27252 38536
rect 27019 38505 27031 38508
rect 26973 38499 27031 38505
rect 27246 38496 27252 38508
rect 27304 38496 27310 38548
rect 27525 38539 27583 38545
rect 27525 38505 27537 38539
rect 27571 38536 27583 38539
rect 29454 38536 29460 38548
rect 27571 38508 29460 38536
rect 27571 38505 27583 38508
rect 27525 38499 27583 38505
rect 29454 38496 29460 38508
rect 29512 38496 29518 38548
rect 29822 38496 29828 38548
rect 29880 38536 29886 38548
rect 31573 38539 31631 38545
rect 31573 38536 31585 38539
rect 29880 38508 31585 38536
rect 29880 38496 29886 38508
rect 31573 38505 31585 38508
rect 31619 38536 31631 38539
rect 31846 38536 31852 38548
rect 31619 38508 31852 38536
rect 31619 38505 31631 38508
rect 31573 38499 31631 38505
rect 31846 38496 31852 38508
rect 31904 38496 31910 38548
rect 26234 38428 26240 38480
rect 26292 38468 26298 38480
rect 26292 38440 28488 38468
rect 26292 38428 26298 38440
rect 21910 38360 21916 38412
rect 21968 38400 21974 38412
rect 25869 38403 25927 38409
rect 25869 38400 25881 38403
rect 21968 38372 25881 38400
rect 21968 38360 21974 38372
rect 25869 38369 25881 38372
rect 25915 38400 25927 38403
rect 27617 38403 27675 38409
rect 25915 38372 27568 38400
rect 25915 38369 25927 38372
rect 25869 38363 25927 38369
rect 23477 38335 23535 38341
rect 23477 38301 23489 38335
rect 23523 38332 23535 38335
rect 26418 38332 26424 38344
rect 23523 38304 26424 38332
rect 23523 38301 23535 38304
rect 23477 38295 23535 38301
rect 26418 38292 26424 38304
rect 26476 38292 26482 38344
rect 26602 38332 26608 38344
rect 26563 38304 26608 38332
rect 26602 38292 26608 38304
rect 26660 38292 26666 38344
rect 26786 38332 26792 38344
rect 26747 38304 26792 38332
rect 26786 38292 26792 38304
rect 26844 38292 26850 38344
rect 1670 38264 1676 38276
rect 1631 38236 1676 38264
rect 1670 38224 1676 38236
rect 1728 38264 1734 38276
rect 2317 38267 2375 38273
rect 2317 38264 2329 38267
rect 1728 38236 2329 38264
rect 1728 38224 1734 38236
rect 2317 38233 2329 38236
rect 2363 38233 2375 38267
rect 2317 38227 2375 38233
rect 5534 38224 5540 38276
rect 5592 38264 5598 38276
rect 22833 38267 22891 38273
rect 22833 38264 22845 38267
rect 5592 38236 22845 38264
rect 5592 38224 5598 38236
rect 22833 38233 22845 38236
rect 22879 38264 22891 38267
rect 26050 38264 26056 38276
rect 22879 38236 26056 38264
rect 22879 38233 22891 38236
rect 22833 38227 22891 38233
rect 26050 38224 26056 38236
rect 26108 38224 26114 38276
rect 26697 38267 26755 38273
rect 26697 38233 26709 38267
rect 26743 38264 26755 38267
rect 26970 38264 26976 38276
rect 26743 38236 26976 38264
rect 26743 38233 26755 38236
rect 26697 38227 26755 38233
rect 26970 38224 26976 38236
rect 27028 38224 27034 38276
rect 27430 38264 27436 38276
rect 27391 38236 27436 38264
rect 27430 38224 27436 38236
rect 27488 38224 27494 38276
rect 27540 38264 27568 38372
rect 27617 38369 27629 38403
rect 27663 38400 27675 38403
rect 28166 38400 28172 38412
rect 27663 38372 28172 38400
rect 27663 38369 27675 38372
rect 27617 38363 27675 38369
rect 28166 38360 28172 38372
rect 28224 38360 28230 38412
rect 27706 38332 27712 38344
rect 27667 38304 27712 38332
rect 27706 38292 27712 38304
rect 27764 38292 27770 38344
rect 28460 38341 28488 38440
rect 28534 38428 28540 38480
rect 28592 38468 28598 38480
rect 28948 38468 28954 38480
rect 28592 38440 28954 38468
rect 28592 38428 28598 38440
rect 28948 38428 28954 38440
rect 29006 38428 29012 38480
rect 29181 38471 29239 38477
rect 29181 38437 29193 38471
rect 29227 38468 29239 38471
rect 29730 38468 29736 38480
rect 29227 38440 29736 38468
rect 29227 38437 29239 38440
rect 29181 38431 29239 38437
rect 29730 38428 29736 38440
rect 29788 38428 29794 38480
rect 28810 38360 28816 38412
rect 28868 38400 28874 38412
rect 30926 38400 30932 38412
rect 28868 38372 29132 38400
rect 28868 38360 28874 38372
rect 28445 38335 28503 38341
rect 28445 38301 28457 38335
rect 28491 38301 28503 38335
rect 28445 38295 28503 38301
rect 28629 38335 28687 38341
rect 28629 38301 28641 38335
rect 28675 38332 28687 38335
rect 28994 38332 29000 38344
rect 28675 38304 29000 38332
rect 28675 38301 28687 38304
rect 28629 38295 28687 38301
rect 28994 38292 29000 38304
rect 29052 38292 29058 38344
rect 29104 38332 29132 38372
rect 29472 38372 30932 38400
rect 29472 38332 29500 38372
rect 30926 38360 30932 38372
rect 30984 38400 30990 38412
rect 31478 38400 31484 38412
rect 30984 38372 31484 38400
rect 30984 38360 30990 38372
rect 31478 38360 31484 38372
rect 31536 38360 31542 38412
rect 31570 38360 31576 38412
rect 31628 38400 31634 38412
rect 32674 38400 32680 38412
rect 31628 38372 32680 38400
rect 31628 38360 31634 38372
rect 32674 38360 32680 38372
rect 32732 38360 32738 38412
rect 34422 38360 34428 38412
rect 34480 38400 34486 38412
rect 52457 38403 52515 38409
rect 52457 38400 52469 38403
rect 34480 38372 52469 38400
rect 34480 38360 34486 38372
rect 52457 38369 52469 38372
rect 52503 38369 52515 38403
rect 53742 38400 53748 38412
rect 53703 38372 53748 38400
rect 52457 38363 52515 38369
rect 53742 38360 53748 38372
rect 53800 38360 53806 38412
rect 29104 38304 29500 38332
rect 29825 38335 29883 38341
rect 29825 38301 29837 38335
rect 29871 38332 29883 38335
rect 29914 38332 29920 38344
rect 29871 38304 29920 38332
rect 29871 38301 29883 38304
rect 29825 38295 29883 38301
rect 29914 38292 29920 38304
rect 29972 38292 29978 38344
rect 30837 38335 30895 38341
rect 30837 38301 30849 38335
rect 30883 38332 30895 38335
rect 31202 38332 31208 38344
rect 30883 38304 31208 38332
rect 30883 38301 30895 38304
rect 30837 38295 30895 38301
rect 31202 38292 31208 38304
rect 31260 38292 31266 38344
rect 31395 38335 31453 38341
rect 31395 38301 31407 38335
rect 31441 38332 31453 38335
rect 32769 38335 32827 38341
rect 31441 38304 31524 38332
rect 31441 38301 31453 38304
rect 31395 38295 31453 38301
rect 31496 38276 31524 38304
rect 32769 38301 32781 38335
rect 32815 38332 32827 38335
rect 32858 38332 32864 38344
rect 32815 38304 32864 38332
rect 32815 38301 32827 38304
rect 32769 38295 32827 38301
rect 32858 38292 32864 38304
rect 32916 38292 32922 38344
rect 33318 38292 33324 38344
rect 33376 38332 33382 38344
rect 33505 38335 33563 38341
rect 33505 38332 33517 38335
rect 33376 38304 33517 38332
rect 33376 38292 33382 38304
rect 33505 38301 33517 38304
rect 33551 38301 33563 38335
rect 33505 38295 33563 38301
rect 51721 38335 51779 38341
rect 51721 38301 51733 38335
rect 51767 38332 51779 38335
rect 52178 38332 52184 38344
rect 51767 38304 52184 38332
rect 51767 38301 51779 38304
rect 51721 38295 51779 38301
rect 52178 38292 52184 38304
rect 52236 38292 52242 38344
rect 53469 38335 53527 38341
rect 53469 38301 53481 38335
rect 53515 38332 53527 38335
rect 53515 38304 53788 38332
rect 53515 38301 53527 38304
rect 53469 38295 53527 38301
rect 28810 38264 28816 38276
rect 27540 38236 28816 38264
rect 28810 38224 28816 38236
rect 28868 38224 28874 38276
rect 30009 38267 30067 38273
rect 30009 38233 30021 38267
rect 30055 38264 30067 38267
rect 30098 38264 30104 38276
rect 30055 38236 30104 38264
rect 30055 38233 30067 38236
rect 30009 38227 30067 38233
rect 30098 38224 30104 38236
rect 30156 38224 30162 38276
rect 31478 38224 31484 38276
rect 31536 38264 31542 38276
rect 34057 38267 34115 38273
rect 34057 38264 34069 38267
rect 31536 38236 34069 38264
rect 31536 38224 31542 38236
rect 34057 38233 34069 38236
rect 34103 38233 34115 38267
rect 34057 38227 34115 38233
rect 51169 38267 51227 38273
rect 51169 38233 51181 38267
rect 51215 38264 51227 38267
rect 53484 38264 53512 38295
rect 53760 38276 53788 38304
rect 51215 38236 53512 38264
rect 51215 38233 51227 38236
rect 51169 38227 51227 38233
rect 53742 38224 53748 38276
rect 53800 38224 53806 38276
rect 1765 38199 1823 38205
rect 1765 38165 1777 38199
rect 1811 38196 1823 38199
rect 4338 38196 4344 38208
rect 1811 38168 4344 38196
rect 1811 38165 1823 38168
rect 1765 38159 1823 38165
rect 4338 38156 4344 38168
rect 4396 38156 4402 38208
rect 17310 38156 17316 38208
rect 17368 38196 17374 38208
rect 17497 38199 17555 38205
rect 17497 38196 17509 38199
rect 17368 38168 17509 38196
rect 17368 38156 17374 38168
rect 17497 38165 17509 38168
rect 17543 38165 17555 38199
rect 17497 38159 17555 38165
rect 21450 38156 21456 38208
rect 21508 38196 21514 38208
rect 24026 38196 24032 38208
rect 21508 38168 24032 38196
rect 21508 38156 21514 38168
rect 24026 38156 24032 38168
rect 24084 38156 24090 38208
rect 25222 38156 25228 38208
rect 25280 38196 25286 38208
rect 25409 38199 25467 38205
rect 25409 38196 25421 38199
rect 25280 38168 25421 38196
rect 25280 38156 25286 38168
rect 25409 38165 25421 38168
rect 25455 38196 25467 38199
rect 25866 38196 25872 38208
rect 25455 38168 25872 38196
rect 25455 38165 25467 38168
rect 25409 38159 25467 38165
rect 25866 38156 25872 38168
rect 25924 38196 25930 38208
rect 26786 38196 26792 38208
rect 25924 38168 26792 38196
rect 25924 38156 25930 38168
rect 26786 38156 26792 38168
rect 26844 38156 26850 38208
rect 27893 38199 27951 38205
rect 27893 38165 27905 38199
rect 27939 38196 27951 38199
rect 28350 38196 28356 38208
rect 27939 38168 28356 38196
rect 27939 38165 27951 38168
rect 27893 38159 27951 38165
rect 28350 38156 28356 38168
rect 28408 38156 28414 38208
rect 28534 38156 28540 38208
rect 28592 38196 28598 38208
rect 28718 38196 28724 38208
rect 28592 38168 28724 38196
rect 28592 38156 28598 38168
rect 28718 38156 28724 38168
rect 28776 38156 28782 38208
rect 28994 38156 29000 38208
rect 29052 38196 29058 38208
rect 29914 38196 29920 38208
rect 29052 38168 29920 38196
rect 29052 38156 29058 38168
rect 29914 38156 29920 38168
rect 29972 38156 29978 38208
rect 30190 38196 30196 38208
rect 30151 38168 30196 38196
rect 30190 38156 30196 38168
rect 30248 38156 30254 38208
rect 30745 38199 30803 38205
rect 30745 38165 30757 38199
rect 30791 38196 30803 38199
rect 31662 38196 31668 38208
rect 30791 38168 31668 38196
rect 30791 38165 30803 38168
rect 30745 38159 30803 38165
rect 31662 38156 31668 38168
rect 31720 38156 31726 38208
rect 32677 38199 32735 38205
rect 32677 38165 32689 38199
rect 32723 38196 32735 38199
rect 32858 38196 32864 38208
rect 32723 38168 32864 38196
rect 32723 38165 32735 38168
rect 32677 38159 32735 38165
rect 32858 38156 32864 38168
rect 32916 38156 32922 38208
rect 33410 38196 33416 38208
rect 33371 38168 33416 38196
rect 33410 38156 33416 38168
rect 33468 38156 33474 38208
rect 1104 38106 54832 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 54832 38106
rect 1104 38032 54832 38054
rect 24121 37995 24179 38001
rect 24121 37961 24133 37995
rect 24167 37992 24179 37995
rect 25682 37992 25688 38004
rect 24167 37964 25688 37992
rect 24167 37961 24179 37964
rect 24121 37955 24179 37961
rect 25682 37952 25688 37964
rect 25740 37992 25746 38004
rect 25740 37964 26439 37992
rect 25740 37952 25746 37964
rect 2130 37884 2136 37936
rect 2188 37924 2194 37936
rect 2188 37896 6914 37924
rect 2188 37884 2194 37896
rect 1578 37856 1584 37868
rect 1539 37828 1584 37856
rect 1578 37816 1584 37828
rect 1636 37856 1642 37868
rect 2777 37859 2835 37865
rect 2777 37856 2789 37859
rect 1636 37828 2789 37856
rect 1636 37816 1642 37828
rect 2777 37825 2789 37828
rect 2823 37825 2835 37859
rect 6886 37856 6914 37896
rect 23106 37884 23112 37936
rect 23164 37924 23170 37936
rect 26411 37924 26439 37964
rect 26602 37952 26608 38004
rect 26660 37992 26666 38004
rect 27893 37995 27951 38001
rect 26660 37964 26705 37992
rect 27448 37964 27845 37992
rect 26660 37952 26666 37964
rect 27448 37924 27476 37964
rect 27525 37927 27583 37933
rect 27525 37924 27537 37927
rect 23164 37896 24164 37924
rect 26411 37896 27537 37924
rect 23164 37884 23170 37896
rect 22002 37856 22008 37868
rect 6886 37828 22008 37856
rect 2777 37819 2835 37825
rect 22002 37816 22008 37828
rect 22060 37816 22066 37868
rect 24136 37856 24164 37896
rect 27525 37893 27537 37896
rect 27571 37893 27583 37927
rect 27817 37924 27845 37964
rect 27893 37961 27905 37995
rect 27939 37992 27951 37995
rect 28166 37992 28172 38004
rect 27939 37964 28172 37992
rect 27939 37961 27951 37964
rect 27893 37955 27951 37961
rect 28166 37952 28172 37964
rect 28224 37952 28230 38004
rect 28997 37995 29055 38001
rect 28997 37961 29009 37995
rect 29043 37961 29055 37995
rect 29822 37992 29828 38004
rect 28997 37955 29055 37961
rect 29472 37964 29828 37992
rect 28902 37924 28908 37936
rect 27817 37896 28908 37924
rect 27525 37887 27583 37893
rect 28902 37884 28908 37896
rect 28960 37884 28966 37936
rect 24136 37828 24716 37856
rect 4338 37748 4344 37800
rect 4396 37788 4402 37800
rect 24302 37788 24308 37800
rect 4396 37760 24308 37788
rect 4396 37748 4402 37760
rect 24302 37748 24308 37760
rect 24360 37748 24366 37800
rect 24688 37788 24716 37828
rect 24762 37816 24768 37868
rect 24820 37856 24826 37868
rect 25406 37856 25412 37868
rect 24820 37828 24865 37856
rect 25367 37828 25412 37856
rect 24820 37816 24826 37828
rect 25406 37816 25412 37828
rect 25464 37816 25470 37868
rect 25590 37856 25596 37868
rect 25551 37828 25596 37856
rect 25590 37816 25596 37828
rect 25648 37816 25654 37868
rect 26050 37856 26056 37868
rect 26011 37828 26056 37856
rect 26050 37816 26056 37828
rect 26108 37816 26114 37868
rect 26237 37859 26295 37865
rect 26237 37825 26249 37859
rect 26283 37825 26295 37859
rect 26237 37819 26295 37825
rect 26329 37859 26387 37865
rect 26329 37825 26341 37859
rect 26375 37825 26387 37859
rect 26329 37819 26387 37825
rect 26421 37859 26479 37865
rect 26421 37825 26433 37859
rect 26467 37825 26479 37859
rect 27338 37856 27344 37868
rect 27299 37828 27344 37856
rect 26421 37819 26479 37825
rect 25958 37788 25964 37800
rect 24688 37760 25964 37788
rect 25958 37748 25964 37760
rect 26016 37788 26022 37800
rect 26252 37788 26280 37819
rect 26016 37760 26280 37788
rect 26016 37748 26022 37760
rect 1765 37723 1823 37729
rect 1765 37689 1777 37723
rect 1811 37720 1823 37723
rect 14826 37720 14832 37732
rect 1811 37692 14832 37720
rect 1811 37689 1823 37692
rect 1765 37683 1823 37689
rect 14826 37680 14832 37692
rect 14884 37680 14890 37732
rect 23106 37720 23112 37732
rect 23067 37692 23112 37720
rect 23106 37680 23112 37692
rect 23164 37680 23170 37732
rect 23661 37723 23719 37729
rect 23661 37689 23673 37723
rect 23707 37720 23719 37723
rect 26234 37720 26240 37732
rect 23707 37692 26240 37720
rect 23707 37689 23719 37692
rect 23661 37683 23719 37689
rect 26234 37680 26240 37692
rect 26292 37720 26298 37732
rect 26344 37720 26372 37819
rect 26436 37788 26464 37819
rect 27338 37816 27344 37828
rect 27396 37816 27402 37868
rect 27617 37859 27675 37865
rect 27617 37846 27629 37859
rect 27540 37825 27629 37846
rect 27663 37825 27675 37859
rect 27540 37819 27675 37825
rect 27755 37859 27813 37865
rect 27755 37825 27767 37859
rect 27801 37856 27813 37859
rect 28074 37856 28080 37868
rect 27801 37828 28080 37856
rect 27801 37825 27813 37828
rect 27755 37819 27813 37825
rect 27540 37818 27660 37819
rect 26694 37788 26700 37800
rect 26436 37760 26700 37788
rect 26694 37748 26700 37760
rect 26752 37748 26758 37800
rect 27154 37748 27160 37800
rect 27212 37788 27218 37800
rect 27540 37788 27568 37818
rect 28074 37816 28080 37828
rect 28132 37816 28138 37868
rect 28718 37816 28724 37868
rect 28776 37856 28782 37868
rect 29012 37856 29040 37955
rect 29472 37936 29500 37964
rect 29822 37952 29828 37964
rect 29880 37952 29886 38004
rect 30098 37992 30104 38004
rect 30059 37964 30104 37992
rect 30098 37952 30104 37964
rect 30156 37952 30162 38004
rect 32582 37992 32588 38004
rect 30392 37964 32588 37992
rect 29270 37924 29276 37936
rect 29231 37896 29276 37924
rect 29270 37884 29276 37896
rect 29328 37884 29334 37936
rect 29365 37927 29423 37933
rect 29365 37893 29377 37927
rect 29411 37924 29423 37927
rect 29454 37924 29460 37936
rect 29411 37896 29460 37924
rect 29411 37893 29423 37896
rect 29365 37887 29423 37893
rect 29454 37884 29460 37896
rect 29512 37884 29518 37936
rect 29730 37924 29736 37936
rect 29564 37896 29736 37924
rect 28776 37828 29040 37856
rect 28776 37816 28782 37828
rect 29086 37816 29092 37868
rect 29144 37865 29150 37868
rect 29564 37865 29592 37896
rect 29730 37884 29736 37896
rect 29788 37884 29794 37936
rect 30392 37933 30420 37964
rect 32582 37952 32588 37964
rect 32640 37952 32646 38004
rect 32674 37952 32680 38004
rect 32732 37992 32738 38004
rect 34330 37992 34336 38004
rect 32732 37964 32777 37992
rect 34291 37964 34336 37992
rect 32732 37952 32738 37964
rect 34330 37952 34336 37964
rect 34388 37952 34394 38004
rect 51350 37992 51356 38004
rect 45526 37964 51356 37992
rect 30377 37927 30435 37933
rect 30377 37893 30389 37927
rect 30423 37893 30435 37927
rect 30377 37887 30435 37893
rect 30469 37927 30527 37933
rect 30469 37893 30481 37927
rect 30515 37924 30527 37927
rect 30834 37924 30840 37936
rect 30515 37896 30840 37924
rect 30515 37893 30527 37896
rect 30469 37887 30527 37893
rect 30834 37884 30840 37896
rect 30892 37884 30898 37936
rect 31018 37884 31024 37936
rect 31076 37924 31082 37936
rect 33781 37927 33839 37933
rect 33781 37924 33793 37927
rect 31076 37896 33793 37924
rect 31076 37884 31082 37896
rect 33781 37893 33793 37896
rect 33827 37924 33839 37927
rect 33827 37896 37274 37924
rect 33827 37893 33839 37896
rect 33781 37887 33839 37893
rect 29144 37859 29193 37865
rect 29144 37825 29147 37859
rect 29181 37825 29193 37859
rect 29144 37819 29193 37825
rect 29548 37859 29606 37865
rect 29548 37825 29560 37859
rect 29594 37825 29606 37859
rect 29548 37819 29606 37825
rect 29144 37816 29150 37819
rect 29638 37816 29644 37868
rect 29696 37856 29702 37868
rect 29696 37828 29741 37856
rect 29696 37816 29702 37828
rect 29822 37816 29828 37868
rect 29880 37856 29886 37868
rect 30239 37859 30297 37865
rect 30239 37856 30251 37859
rect 29880 37828 30251 37856
rect 29880 37816 29886 37828
rect 30239 37825 30251 37828
rect 30285 37825 30297 37859
rect 30239 37819 30297 37825
rect 30558 37816 30564 37868
rect 30616 37865 30622 37868
rect 30616 37859 30655 37865
rect 30643 37825 30655 37859
rect 30616 37819 30655 37825
rect 30745 37859 30803 37865
rect 30745 37825 30757 37859
rect 30791 37856 30803 37859
rect 30926 37856 30932 37868
rect 30791 37828 30932 37856
rect 30791 37825 30803 37828
rect 30745 37819 30803 37825
rect 30616 37816 30622 37819
rect 30926 37816 30932 37828
rect 30984 37816 30990 37868
rect 31202 37856 31208 37868
rect 31163 37828 31208 37856
rect 31202 37816 31208 37828
rect 31260 37816 31266 37868
rect 32401 37859 32459 37865
rect 32401 37825 32413 37859
rect 32447 37856 32459 37859
rect 33042 37856 33048 37868
rect 32447 37828 33048 37856
rect 32447 37825 32459 37828
rect 32401 37819 32459 37825
rect 33042 37816 33048 37828
rect 33100 37816 33106 37868
rect 33226 37856 33232 37868
rect 33187 37828 33232 37856
rect 33226 37816 33232 37828
rect 33284 37816 33290 37868
rect 37246 37856 37274 37896
rect 45526 37856 45554 37964
rect 51350 37952 51356 37964
rect 51408 37952 51414 38004
rect 51077 37927 51135 37933
rect 51077 37893 51089 37927
rect 51123 37924 51135 37927
rect 53650 37924 53656 37936
rect 51123 37896 53656 37924
rect 51123 37893 51135 37896
rect 51077 37887 51135 37893
rect 53650 37884 53656 37896
rect 53708 37884 53714 37936
rect 53745 37859 53803 37865
rect 53745 37856 53757 37859
rect 37246 37828 45554 37856
rect 49528 37828 53757 37856
rect 49528 37788 49556 37828
rect 53745 37825 53757 37828
rect 53791 37825 53803 37859
rect 53745 37819 53803 37825
rect 27212 37760 27568 37788
rect 27724 37760 29040 37788
rect 27212 37748 27218 37760
rect 27724 37720 27752 37760
rect 29012 37720 29040 37760
rect 29564 37760 49556 37788
rect 52089 37791 52147 37797
rect 29564 37720 29592 37760
rect 52089 37757 52101 37791
rect 52135 37757 52147 37791
rect 52089 37751 52147 37757
rect 52365 37791 52423 37797
rect 52365 37757 52377 37791
rect 52411 37788 52423 37791
rect 53469 37791 53527 37797
rect 52411 37760 53052 37788
rect 52411 37757 52423 37760
rect 52365 37751 52423 37757
rect 52104 37720 52132 37751
rect 26292 37692 26372 37720
rect 26411 37692 27752 37720
rect 28184 37692 28949 37720
rect 29012 37692 29592 37720
rect 29748 37692 52132 37720
rect 26292 37680 26298 37692
rect 2317 37655 2375 37661
rect 2317 37621 2329 37655
rect 2363 37652 2375 37655
rect 2774 37652 2780 37664
rect 2363 37624 2780 37652
rect 2363 37621 2375 37624
rect 2317 37615 2375 37621
rect 2774 37612 2780 37624
rect 2832 37612 2838 37664
rect 22557 37655 22615 37661
rect 22557 37621 22569 37655
rect 22603 37652 22615 37655
rect 23566 37652 23572 37664
rect 22603 37624 23572 37652
rect 22603 37621 22615 37624
rect 22557 37615 22615 37621
rect 23566 37612 23572 37624
rect 23624 37612 23630 37664
rect 25222 37652 25228 37664
rect 25183 37624 25228 37652
rect 25222 37612 25228 37624
rect 25280 37612 25286 37664
rect 25590 37652 25596 37664
rect 25551 37624 25596 37652
rect 25590 37612 25596 37624
rect 25648 37612 25654 37664
rect 26142 37612 26148 37664
rect 26200 37652 26206 37664
rect 26411 37652 26439 37692
rect 26200 37624 26439 37652
rect 26200 37612 26206 37624
rect 26694 37612 26700 37664
rect 26752 37652 26758 37664
rect 28184 37652 28212 37692
rect 26752 37624 28212 37652
rect 26752 37612 26758 37624
rect 28258 37612 28264 37664
rect 28316 37652 28322 37664
rect 28353 37655 28411 37661
rect 28353 37652 28365 37655
rect 28316 37624 28365 37652
rect 28316 37612 28322 37624
rect 28353 37621 28365 37624
rect 28399 37621 28411 37655
rect 28921 37652 28949 37692
rect 29748 37652 29776 37692
rect 53024 37664 53052 37760
rect 53469 37757 53481 37791
rect 53515 37788 53527 37791
rect 53650 37788 53656 37800
rect 53515 37760 53656 37788
rect 53515 37757 53527 37760
rect 53469 37751 53527 37757
rect 53650 37748 53656 37760
rect 53708 37748 53714 37800
rect 28921 37624 29776 37652
rect 28353 37615 28411 37621
rect 29822 37612 29828 37664
rect 29880 37652 29886 37664
rect 32122 37652 32128 37664
rect 29880 37624 32128 37652
rect 29880 37612 29886 37624
rect 32122 37612 32128 37624
rect 32180 37612 32186 37664
rect 33042 37612 33048 37664
rect 33100 37652 33106 37664
rect 34606 37652 34612 37664
rect 33100 37624 34612 37652
rect 33100 37612 33106 37624
rect 34606 37612 34612 37624
rect 34664 37652 34670 37664
rect 34885 37655 34943 37661
rect 34885 37652 34897 37655
rect 34664 37624 34897 37652
rect 34664 37612 34670 37624
rect 34885 37621 34897 37624
rect 34931 37621 34943 37655
rect 53006 37652 53012 37664
rect 52967 37624 53012 37652
rect 34885 37615 34943 37621
rect 53006 37612 53012 37624
rect 53064 37612 53070 37664
rect 1104 37562 54832 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 54832 37562
rect 1104 37488 54832 37510
rect 2314 37408 2320 37460
rect 2372 37448 2378 37460
rect 24026 37448 24032 37460
rect 2372 37420 6914 37448
rect 23987 37420 24032 37448
rect 2372 37408 2378 37420
rect 6886 37380 6914 37420
rect 24026 37408 24032 37420
rect 24084 37408 24090 37460
rect 24670 37448 24676 37460
rect 24631 37420 24676 37448
rect 24670 37408 24676 37420
rect 24728 37408 24734 37460
rect 24762 37408 24768 37460
rect 24820 37448 24826 37460
rect 27338 37448 27344 37460
rect 24820 37420 27344 37448
rect 24820 37408 24826 37420
rect 27338 37408 27344 37420
rect 27396 37408 27402 37460
rect 27430 37408 27436 37460
rect 27488 37448 27494 37460
rect 27617 37451 27675 37457
rect 27617 37448 27629 37451
rect 27488 37420 27629 37448
rect 27488 37408 27494 37420
rect 27617 37417 27629 37420
rect 27663 37417 27675 37451
rect 27617 37411 27675 37417
rect 28166 37408 28172 37460
rect 28224 37448 28230 37460
rect 28721 37451 28779 37457
rect 28721 37448 28733 37451
rect 28224 37420 28733 37448
rect 28224 37408 28230 37420
rect 28721 37417 28733 37420
rect 28767 37417 28779 37451
rect 28721 37411 28779 37417
rect 30098 37408 30104 37460
rect 30156 37448 30162 37460
rect 30374 37448 30380 37460
rect 30156 37420 30380 37448
rect 30156 37408 30162 37420
rect 30374 37408 30380 37420
rect 30432 37448 30438 37460
rect 31573 37451 31631 37457
rect 31573 37448 31585 37451
rect 30432 37420 31585 37448
rect 30432 37408 30438 37420
rect 31573 37417 31585 37420
rect 31619 37417 31631 37451
rect 32122 37448 32128 37460
rect 32083 37420 32128 37448
rect 31573 37411 31631 37417
rect 32122 37408 32128 37420
rect 32180 37448 32186 37460
rect 32306 37448 32312 37460
rect 32180 37420 32312 37448
rect 32180 37408 32186 37420
rect 32306 37408 32312 37420
rect 32364 37408 32370 37460
rect 53558 37448 53564 37460
rect 41386 37420 53564 37448
rect 25225 37383 25283 37389
rect 25225 37380 25237 37383
rect 6886 37352 25237 37380
rect 25225 37349 25237 37352
rect 25271 37349 25283 37383
rect 25225 37343 25283 37349
rect 2409 37315 2467 37321
rect 2409 37281 2421 37315
rect 2455 37312 2467 37315
rect 2774 37312 2780 37324
rect 2455 37284 2780 37312
rect 2455 37281 2467 37284
rect 2409 37275 2467 37281
rect 2774 37272 2780 37284
rect 2832 37272 2838 37324
rect 22370 37312 22376 37324
rect 22331 37284 22376 37312
rect 22370 37272 22376 37284
rect 22428 37272 22434 37324
rect 25240 37312 25268 37343
rect 26418 37340 26424 37392
rect 26476 37380 26482 37392
rect 41386 37380 41414 37420
rect 53558 37408 53564 37420
rect 53616 37408 53622 37460
rect 26476 37352 31708 37380
rect 26476 37340 26482 37352
rect 27430 37312 27436 37324
rect 25240 37284 27436 37312
rect 27430 37272 27436 37284
rect 27488 37272 27494 37324
rect 28442 37312 28448 37324
rect 28000 37284 28448 37312
rect 2133 37247 2191 37253
rect 2133 37213 2145 37247
rect 2179 37213 2191 37247
rect 23934 37244 23940 37256
rect 2133 37207 2191 37213
rect 6886 37216 23940 37244
rect 2148 37176 2176 37207
rect 6886 37176 6914 37216
rect 23934 37204 23940 37216
rect 23992 37204 23998 37256
rect 25222 37204 25228 37256
rect 25280 37244 25286 37256
rect 25869 37247 25927 37253
rect 25869 37244 25881 37247
rect 25280 37216 25881 37244
rect 25280 37204 25286 37216
rect 25869 37213 25881 37216
rect 25915 37213 25927 37247
rect 26651 37247 26709 37253
rect 26651 37244 26663 37247
rect 25869 37207 25927 37213
rect 25976 37216 26663 37244
rect 25976 37176 26004 37216
rect 26651 37213 26663 37216
rect 26697 37213 26709 37247
rect 26878 37244 26884 37256
rect 26839 37216 26884 37244
rect 26651 37207 26709 37213
rect 26878 37204 26884 37216
rect 26936 37204 26942 37256
rect 27062 37244 27068 37256
rect 27023 37216 27068 37244
rect 27062 37204 27068 37216
rect 27120 37204 27126 37256
rect 27154 37204 27160 37256
rect 27212 37244 27218 37256
rect 27212 37216 27257 37244
rect 27212 37204 27218 37216
rect 27338 37204 27344 37256
rect 27396 37244 27402 37256
rect 27614 37244 27620 37256
rect 27396 37216 27620 37244
rect 27396 37204 27402 37216
rect 27614 37204 27620 37216
rect 27672 37244 27678 37256
rect 28000 37253 28028 37284
rect 28442 37272 28448 37284
rect 28500 37272 28506 37324
rect 28810 37312 28816 37324
rect 28771 37284 28816 37312
rect 28810 37272 28816 37284
rect 28868 37272 28874 37324
rect 28902 37272 28908 37324
rect 28960 37312 28966 37324
rect 29822 37312 29828 37324
rect 28960 37284 29828 37312
rect 28960 37272 28966 37284
rect 29822 37272 29828 37284
rect 29880 37272 29886 37324
rect 30190 37272 30196 37324
rect 30248 37312 30254 37324
rect 31113 37315 31171 37321
rect 30248 37284 30604 37312
rect 30248 37272 30254 37284
rect 27755 37247 27813 37253
rect 27755 37244 27767 37247
rect 27672 37216 27767 37244
rect 27672 37204 27678 37216
rect 27755 37213 27767 37216
rect 27801 37213 27813 37247
rect 27755 37207 27813 37213
rect 27985 37247 28043 37253
rect 27985 37213 27997 37247
rect 28031 37213 28043 37247
rect 28166 37244 28172 37256
rect 28127 37216 28172 37244
rect 27985 37207 28043 37213
rect 28166 37204 28172 37216
rect 28224 37204 28230 37256
rect 28261 37247 28319 37253
rect 28261 37213 28273 37247
rect 28307 37244 28319 37247
rect 28718 37244 28724 37256
rect 28307 37216 28396 37244
rect 28679 37216 28724 37244
rect 28307 37213 28319 37216
rect 28261 37207 28319 37213
rect 2148 37148 6914 37176
rect 23032 37148 26004 37176
rect 23032 37120 23060 37148
rect 26050 37136 26056 37188
rect 26108 37176 26114 37188
rect 26786 37176 26792 37188
rect 26108 37148 26153 37176
rect 26747 37148 26792 37176
rect 26108 37136 26114 37148
rect 26786 37136 26792 37148
rect 26844 37136 26850 37188
rect 27890 37136 27896 37188
rect 27948 37176 27954 37188
rect 27948 37148 27993 37176
rect 27948 37136 27954 37148
rect 22925 37111 22983 37117
rect 22925 37077 22937 37111
rect 22971 37108 22983 37111
rect 23014 37108 23020 37120
rect 22971 37080 23020 37108
rect 22971 37077 22983 37080
rect 22925 37071 22983 37077
rect 23014 37068 23020 37080
rect 23072 37068 23078 37120
rect 23477 37111 23535 37117
rect 23477 37077 23489 37111
rect 23523 37108 23535 37111
rect 25498 37108 25504 37120
rect 23523 37080 25504 37108
rect 23523 37077 23535 37080
rect 23477 37071 23535 37077
rect 25498 37068 25504 37080
rect 25556 37068 25562 37120
rect 25590 37068 25596 37120
rect 25648 37108 25654 37120
rect 26513 37111 26571 37117
rect 26513 37108 26525 37111
rect 25648 37080 26525 37108
rect 25648 37068 25654 37080
rect 26513 37077 26525 37080
rect 26559 37077 26571 37111
rect 26513 37071 26571 37077
rect 26694 37068 26700 37120
rect 26752 37108 26758 37120
rect 28368 37108 28396 37216
rect 28718 37204 28724 37216
rect 28776 37204 28782 37256
rect 29840 37244 29868 37272
rect 29912 37247 29970 37253
rect 29912 37244 29924 37247
rect 29840 37216 29924 37244
rect 29912 37213 29924 37216
rect 29958 37213 29970 37247
rect 29912 37207 29970 37213
rect 30284 37247 30342 37253
rect 30284 37213 30296 37247
rect 30330 37213 30342 37247
rect 30284 37207 30342 37213
rect 30009 37179 30067 37185
rect 30009 37145 30021 37179
rect 30055 37145 30067 37179
rect 30009 37139 30067 37145
rect 29086 37108 29092 37120
rect 26752 37080 28396 37108
rect 29047 37080 29092 37108
rect 26752 37068 26758 37080
rect 29086 37068 29092 37080
rect 29144 37068 29150 37120
rect 29733 37111 29791 37117
rect 29733 37077 29745 37111
rect 29779 37108 29791 37111
rect 29822 37108 29828 37120
rect 29779 37080 29828 37108
rect 29779 37077 29791 37080
rect 29733 37071 29791 37077
rect 29822 37068 29828 37080
rect 29880 37068 29886 37120
rect 30024 37108 30052 37139
rect 30098 37136 30104 37188
rect 30156 37176 30162 37188
rect 30299 37176 30327 37207
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30576 37244 30604 37284
rect 31113 37281 31125 37315
rect 31159 37312 31171 37315
rect 31570 37312 31576 37324
rect 31159 37284 31576 37312
rect 31159 37281 31171 37284
rect 31113 37275 31171 37281
rect 31570 37272 31576 37284
rect 31628 37272 31634 37324
rect 31680 37312 31708 37352
rect 31772 37352 41414 37380
rect 31772 37312 31800 37352
rect 33778 37312 33784 37324
rect 31680 37284 31800 37312
rect 33739 37284 33784 37312
rect 33778 37272 33784 37284
rect 33836 37272 33842 37324
rect 51721 37315 51779 37321
rect 51721 37281 51733 37315
rect 51767 37312 51779 37315
rect 53466 37312 53472 37324
rect 51767 37284 53472 37312
rect 51767 37281 51779 37284
rect 51721 37275 51779 37281
rect 53466 37272 53472 37284
rect 53524 37272 53530 37324
rect 30929 37247 30987 37253
rect 30929 37244 30941 37247
rect 30432 37216 30477 37244
rect 30576 37216 30941 37244
rect 30432 37204 30438 37216
rect 30929 37213 30941 37216
rect 30975 37213 30987 37247
rect 30929 37207 30987 37213
rect 44174 37204 44180 37256
rect 44232 37244 44238 37256
rect 52733 37247 52791 37253
rect 52733 37244 52745 37247
rect 44232 37216 52745 37244
rect 44232 37204 44238 37216
rect 52733 37213 52745 37216
rect 52779 37213 52791 37247
rect 53006 37244 53012 37256
rect 52967 37216 53012 37244
rect 52733 37207 52791 37213
rect 53006 37204 53012 37216
rect 53064 37204 53070 37256
rect 53558 37204 53564 37256
rect 53616 37244 53622 37256
rect 53745 37247 53803 37253
rect 53745 37244 53757 37247
rect 53616 37216 53757 37244
rect 53616 37204 53622 37216
rect 53745 37213 53757 37216
rect 53791 37213 53803 37247
rect 53745 37207 53803 37213
rect 30834 37176 30840 37188
rect 30156 37148 30201 37176
rect 30299 37148 30840 37176
rect 30156 37136 30162 37148
rect 30834 37136 30840 37148
rect 30892 37136 30898 37188
rect 32953 37179 33011 37185
rect 32953 37145 32965 37179
rect 32999 37176 33011 37179
rect 33226 37176 33232 37188
rect 32999 37148 33232 37176
rect 32999 37145 33011 37148
rect 32953 37139 33011 37145
rect 33226 37136 33232 37148
rect 33284 37136 33290 37188
rect 30282 37108 30288 37120
rect 30024 37080 30288 37108
rect 30282 37068 30288 37080
rect 30340 37068 30346 37120
rect 33042 37108 33048 37120
rect 33003 37080 33048 37108
rect 33042 37068 33048 37080
rect 33100 37068 33106 37120
rect 1104 37018 54832 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 54832 37018
rect 1104 36944 54832 36966
rect 23658 36864 23664 36916
rect 23716 36904 23722 36916
rect 26421 36907 26479 36913
rect 23716 36876 26280 36904
rect 23716 36864 23722 36876
rect 22097 36839 22155 36845
rect 22097 36836 22109 36839
rect 19306 36808 22109 36836
rect 2133 36771 2191 36777
rect 2133 36737 2145 36771
rect 2179 36768 2191 36771
rect 17218 36768 17224 36780
rect 2179 36740 17224 36768
rect 2179 36737 2191 36740
rect 2133 36731 2191 36737
rect 17218 36728 17224 36740
rect 17276 36728 17282 36780
rect 2409 36703 2467 36709
rect 2409 36669 2421 36703
rect 2455 36700 2467 36703
rect 2774 36700 2780 36712
rect 2455 36672 2780 36700
rect 2455 36669 2467 36672
rect 2409 36663 2467 36669
rect 2774 36660 2780 36672
rect 2832 36700 2838 36712
rect 2869 36703 2927 36709
rect 2869 36700 2881 36703
rect 2832 36672 2881 36700
rect 2832 36660 2838 36672
rect 2869 36669 2881 36672
rect 2915 36669 2927 36703
rect 2869 36663 2927 36669
rect 13446 36524 13452 36576
rect 13504 36564 13510 36576
rect 19306 36564 19334 36808
rect 22097 36805 22109 36808
rect 22143 36836 22155 36839
rect 26145 36839 26203 36845
rect 26145 36836 26157 36839
rect 22143 36808 26157 36836
rect 22143 36805 22155 36808
rect 22097 36799 22155 36805
rect 26145 36805 26157 36808
rect 26191 36805 26203 36839
rect 26252 36836 26280 36876
rect 26421 36873 26433 36907
rect 26467 36904 26479 36907
rect 26694 36904 26700 36916
rect 26467 36876 26700 36904
rect 26467 36873 26479 36876
rect 26421 36867 26479 36873
rect 26694 36864 26700 36876
rect 26752 36864 26758 36916
rect 27709 36907 27767 36913
rect 27709 36873 27721 36907
rect 27755 36904 27767 36907
rect 28718 36904 28724 36916
rect 27755 36876 28212 36904
rect 28679 36876 28724 36904
rect 27755 36873 27767 36876
rect 27709 36867 27767 36873
rect 27433 36839 27491 36845
rect 27433 36836 27445 36839
rect 26252 36808 27445 36836
rect 26145 36799 26203 36805
rect 27433 36805 27445 36808
rect 27479 36805 27491 36839
rect 27433 36799 27491 36805
rect 28184 36799 28212 36876
rect 28718 36864 28724 36876
rect 28776 36864 28782 36916
rect 31846 36864 31852 36916
rect 31904 36904 31910 36916
rect 32309 36907 32367 36913
rect 32309 36904 32321 36907
rect 31904 36876 32321 36904
rect 31904 36864 31910 36876
rect 32309 36873 32321 36876
rect 32355 36873 32367 36907
rect 32309 36867 32367 36873
rect 32953 36907 33011 36913
rect 32953 36873 32965 36907
rect 32999 36904 33011 36907
rect 35894 36904 35900 36916
rect 32999 36876 35900 36904
rect 32999 36873 33011 36876
rect 32953 36867 33011 36873
rect 28159 36793 28217 36799
rect 28350 36796 28356 36848
rect 28408 36836 28414 36848
rect 29365 36839 29423 36845
rect 29365 36836 29377 36839
rect 28408 36808 29377 36836
rect 28408 36796 28414 36808
rect 29365 36805 29377 36808
rect 29411 36805 29423 36839
rect 29365 36799 29423 36805
rect 30834 36796 30840 36848
rect 30892 36836 30898 36848
rect 32968 36836 32996 36867
rect 35894 36864 35900 36876
rect 35952 36864 35958 36916
rect 53006 36904 53012 36916
rect 52967 36876 53012 36904
rect 53006 36864 53012 36876
rect 53064 36864 53070 36916
rect 30892 36808 32996 36836
rect 30892 36796 30898 36808
rect 25406 36728 25412 36780
rect 25464 36768 25470 36780
rect 25866 36768 25872 36780
rect 25464 36740 25509 36768
rect 25827 36740 25872 36768
rect 25464 36728 25470 36740
rect 25866 36728 25872 36740
rect 25924 36728 25930 36780
rect 26050 36768 26056 36780
rect 26011 36740 26056 36768
rect 26050 36728 26056 36740
rect 26108 36728 26114 36780
rect 26234 36728 26240 36780
rect 26292 36768 26298 36780
rect 27157 36771 27215 36777
rect 26292 36740 26337 36768
rect 26292 36728 26298 36740
rect 27157 36737 27169 36771
rect 27203 36737 27215 36771
rect 27338 36768 27344 36780
rect 27299 36740 27344 36768
rect 27157 36731 27215 36737
rect 24305 36703 24363 36709
rect 24305 36669 24317 36703
rect 24351 36700 24363 36703
rect 27172 36700 27200 36731
rect 27338 36728 27344 36740
rect 27396 36728 27402 36780
rect 27525 36771 27583 36777
rect 27525 36737 27537 36771
rect 27571 36768 27583 36771
rect 27614 36768 27620 36780
rect 27571 36740 27620 36768
rect 27571 36737 27583 36740
rect 27525 36731 27583 36737
rect 27614 36728 27620 36740
rect 27672 36728 27678 36780
rect 28159 36759 28171 36793
rect 28205 36759 28217 36793
rect 28159 36753 28217 36759
rect 28258 36728 28264 36780
rect 28316 36768 28322 36780
rect 28445 36771 28503 36777
rect 28316 36740 28361 36768
rect 28316 36728 28322 36740
rect 28445 36737 28457 36771
rect 28491 36737 28503 36771
rect 28445 36731 28503 36737
rect 27890 36700 27896 36712
rect 24351 36672 27896 36700
rect 24351 36669 24363 36672
rect 24305 36663 24363 36669
rect 27890 36660 27896 36672
rect 27948 36660 27954 36712
rect 22554 36632 22560 36644
rect 22515 36604 22560 36632
rect 22554 36592 22560 36604
rect 22612 36592 22618 36644
rect 24857 36635 24915 36641
rect 24857 36601 24869 36635
rect 24903 36632 24915 36635
rect 26142 36632 26148 36644
rect 24903 36604 26148 36632
rect 24903 36601 24915 36604
rect 24857 36595 24915 36601
rect 26142 36592 26148 36604
rect 26200 36592 26206 36644
rect 27430 36592 27436 36644
rect 27488 36632 27494 36644
rect 28460 36632 28488 36731
rect 28534 36728 28540 36780
rect 28592 36768 28598 36780
rect 28592 36740 28685 36768
rect 28592 36728 28598 36740
rect 29730 36728 29736 36780
rect 29788 36768 29794 36780
rect 30285 36771 30343 36777
rect 30285 36768 30297 36771
rect 29788 36740 30297 36768
rect 29788 36728 29794 36740
rect 30285 36737 30297 36740
rect 30331 36768 30343 36771
rect 31757 36771 31815 36777
rect 31757 36768 31769 36771
rect 30331 36740 31769 36768
rect 30331 36737 30343 36740
rect 30285 36731 30343 36737
rect 31757 36737 31769 36740
rect 31803 36768 31815 36771
rect 31938 36768 31944 36780
rect 31803 36740 31944 36768
rect 31803 36737 31815 36740
rect 31757 36731 31815 36737
rect 31938 36728 31944 36740
rect 31996 36728 32002 36780
rect 53558 36768 53564 36780
rect 45526 36740 53564 36768
rect 27488 36604 28488 36632
rect 28552 36632 28580 36728
rect 28718 36660 28724 36712
rect 28776 36700 28782 36712
rect 45526 36700 45554 36740
rect 53558 36728 53564 36740
rect 53616 36728 53622 36780
rect 28776 36672 45554 36700
rect 52365 36703 52423 36709
rect 28776 36660 28782 36672
rect 52365 36669 52377 36703
rect 52411 36700 52423 36703
rect 53469 36703 53527 36709
rect 53469 36700 53481 36703
rect 52411 36672 53481 36700
rect 52411 36669 52423 36672
rect 52365 36663 52423 36669
rect 53469 36669 53481 36672
rect 53515 36700 53527 36703
rect 53742 36700 53748 36712
rect 53515 36672 53604 36700
rect 53703 36672 53748 36700
rect 53515 36669 53527 36672
rect 53469 36663 53527 36669
rect 53576 36644 53604 36672
rect 53742 36660 53748 36672
rect 53800 36660 53806 36712
rect 28902 36632 28908 36644
rect 28552 36604 28908 36632
rect 27488 36592 27494 36604
rect 28902 36592 28908 36604
rect 28960 36632 28966 36644
rect 30469 36635 30527 36641
rect 30469 36632 30481 36635
rect 28960 36604 30481 36632
rect 28960 36592 28966 36604
rect 30469 36601 30481 36604
rect 30515 36601 30527 36635
rect 31202 36632 31208 36644
rect 31115 36604 31208 36632
rect 30469 36595 30527 36601
rect 31202 36592 31208 36604
rect 31260 36632 31266 36644
rect 49602 36632 49608 36644
rect 31260 36604 49608 36632
rect 31260 36592 31266 36604
rect 49602 36592 49608 36604
rect 49660 36592 49666 36644
rect 53558 36592 53564 36644
rect 53616 36592 53622 36644
rect 13504 36536 19334 36564
rect 13504 36524 13510 36536
rect 22646 36524 22652 36576
rect 22704 36564 22710 36576
rect 23109 36567 23167 36573
rect 23109 36564 23121 36567
rect 22704 36536 23121 36564
rect 22704 36524 22710 36536
rect 23109 36533 23121 36536
rect 23155 36564 23167 36567
rect 23658 36564 23664 36576
rect 23155 36536 23664 36564
rect 23155 36533 23167 36536
rect 23109 36527 23167 36533
rect 23658 36524 23664 36536
rect 23716 36524 23722 36576
rect 23753 36567 23811 36573
rect 23753 36533 23765 36567
rect 23799 36564 23811 36567
rect 24670 36564 24676 36576
rect 23799 36536 24676 36564
rect 23799 36533 23811 36536
rect 23753 36527 23811 36533
rect 24670 36524 24676 36536
rect 24728 36564 24734 36576
rect 26694 36564 26700 36576
rect 24728 36536 26700 36564
rect 24728 36524 24734 36536
rect 26694 36524 26700 36536
rect 26752 36524 26758 36576
rect 29270 36564 29276 36576
rect 29231 36536 29276 36564
rect 29270 36524 29276 36536
rect 29328 36524 29334 36576
rect 33226 36524 33232 36576
rect 33284 36564 33290 36576
rect 33413 36567 33471 36573
rect 33413 36564 33425 36567
rect 33284 36536 33425 36564
rect 33284 36524 33290 36536
rect 33413 36533 33425 36536
rect 33459 36533 33471 36567
rect 33413 36527 33471 36533
rect 1104 36474 54832 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 54832 36474
rect 1104 36400 54832 36422
rect 23474 36320 23480 36372
rect 23532 36360 23538 36372
rect 25130 36360 25136 36372
rect 23532 36332 25136 36360
rect 23532 36320 23538 36332
rect 25130 36320 25136 36332
rect 25188 36320 25194 36372
rect 25222 36320 25228 36372
rect 25280 36360 25286 36372
rect 26329 36363 26387 36369
rect 26329 36360 26341 36363
rect 25280 36332 26341 36360
rect 25280 36320 25286 36332
rect 26329 36329 26341 36332
rect 26375 36329 26387 36363
rect 26329 36323 26387 36329
rect 26418 36320 26424 36372
rect 26476 36360 26482 36372
rect 27614 36360 27620 36372
rect 26476 36332 27620 36360
rect 26476 36320 26482 36332
rect 27614 36320 27620 36332
rect 27672 36320 27678 36372
rect 28902 36320 28908 36372
rect 28960 36360 28966 36372
rect 31938 36360 31944 36372
rect 28960 36332 29776 36360
rect 31899 36332 31944 36360
rect 28960 36320 28966 36332
rect 13446 36292 13452 36304
rect 6886 36264 13452 36292
rect 2133 36227 2191 36233
rect 2133 36193 2145 36227
rect 2179 36224 2191 36227
rect 6886 36224 6914 36264
rect 13446 36252 13452 36264
rect 13504 36252 13510 36304
rect 17310 36252 17316 36304
rect 17368 36292 17374 36304
rect 22278 36292 22284 36304
rect 17368 36264 22284 36292
rect 17368 36252 17374 36264
rect 22278 36252 22284 36264
rect 22336 36252 22342 36304
rect 29748 36301 29776 36332
rect 31938 36320 31944 36332
rect 31996 36360 32002 36372
rect 33042 36360 33048 36372
rect 31996 36332 33048 36360
rect 31996 36320 32002 36332
rect 33042 36320 33048 36332
rect 33100 36320 33106 36372
rect 53742 36360 53748 36372
rect 38626 36332 53748 36360
rect 24765 36295 24823 36301
rect 24765 36261 24777 36295
rect 24811 36292 24823 36295
rect 29733 36295 29791 36301
rect 24811 36264 29684 36292
rect 24811 36261 24823 36264
rect 24765 36255 24823 36261
rect 21821 36227 21879 36233
rect 21821 36224 21833 36227
rect 2179 36196 6914 36224
rect 19306 36196 21833 36224
rect 2179 36193 2191 36196
rect 2133 36187 2191 36193
rect 2409 36159 2467 36165
rect 2409 36125 2421 36159
rect 2455 36156 2467 36159
rect 2774 36156 2780 36168
rect 2455 36128 2780 36156
rect 2455 36125 2467 36128
rect 2409 36119 2467 36125
rect 2774 36116 2780 36128
rect 2832 36156 2838 36168
rect 2869 36159 2927 36165
rect 2869 36156 2881 36159
rect 2832 36128 2881 36156
rect 2832 36116 2838 36128
rect 2869 36125 2881 36128
rect 2915 36125 2927 36159
rect 2869 36119 2927 36125
rect 2038 36048 2044 36100
rect 2096 36088 2102 36100
rect 19306 36088 19334 36196
rect 21821 36193 21833 36196
rect 21867 36224 21879 36227
rect 26694 36224 26700 36236
rect 21867 36196 25361 36224
rect 26655 36196 26700 36224
rect 21867 36193 21879 36196
rect 21821 36187 21879 36193
rect 25222 36156 25228 36168
rect 25183 36128 25228 36156
rect 25222 36116 25228 36128
rect 25280 36116 25286 36168
rect 25333 36165 25361 36196
rect 26694 36184 26700 36196
rect 26752 36184 26758 36236
rect 25318 36159 25376 36165
rect 25318 36125 25330 36159
rect 25364 36125 25376 36159
rect 25318 36119 25376 36125
rect 25590 36116 25596 36168
rect 25648 36156 25654 36168
rect 25731 36159 25789 36165
rect 25648 36128 25693 36156
rect 25648 36116 25654 36128
rect 25731 36125 25743 36159
rect 25777 36156 25789 36159
rect 25958 36156 25964 36168
rect 25777 36128 25964 36156
rect 25777 36125 25789 36128
rect 25731 36119 25789 36125
rect 25958 36116 25964 36128
rect 26016 36156 26022 36168
rect 26418 36156 26424 36168
rect 26016 36128 26424 36156
rect 26016 36116 26022 36128
rect 26418 36116 26424 36128
rect 26476 36116 26482 36168
rect 27172 36165 27200 36264
rect 27890 36184 27896 36236
rect 27948 36224 27954 36236
rect 27948 36196 28488 36224
rect 27948 36184 27954 36196
rect 26513 36159 26571 36165
rect 26513 36125 26525 36159
rect 26559 36125 26571 36159
rect 26513 36119 26571 36125
rect 27157 36159 27215 36165
rect 27157 36125 27169 36159
rect 27203 36125 27215 36159
rect 27157 36119 27215 36125
rect 21266 36088 21272 36100
rect 2096 36060 19334 36088
rect 21227 36060 21272 36088
rect 2096 36048 2102 36060
rect 21266 36048 21272 36060
rect 21324 36048 21330 36100
rect 25406 36048 25412 36100
rect 25464 36088 25470 36100
rect 25501 36091 25559 36097
rect 25501 36088 25513 36091
rect 25464 36060 25513 36088
rect 25464 36048 25470 36060
rect 25501 36057 25513 36060
rect 25547 36057 25559 36091
rect 26528 36088 26556 36119
rect 27338 36116 27344 36168
rect 27396 36156 27402 36168
rect 27396 36128 27441 36156
rect 27396 36116 27402 36128
rect 27522 36116 27528 36168
rect 27580 36156 27586 36168
rect 27580 36128 27625 36156
rect 27580 36116 27586 36128
rect 28074 36116 28080 36168
rect 28132 36156 28138 36168
rect 28460 36165 28488 36196
rect 28810 36184 28816 36236
rect 28868 36224 28874 36236
rect 28994 36224 29000 36236
rect 28868 36196 29000 36224
rect 28868 36184 28874 36196
rect 28994 36184 29000 36196
rect 29052 36184 29058 36236
rect 29656 36224 29684 36264
rect 29733 36261 29745 36295
rect 29779 36261 29791 36295
rect 29733 36255 29791 36261
rect 31481 36295 31539 36301
rect 31481 36261 31493 36295
rect 31527 36292 31539 36295
rect 31754 36292 31760 36304
rect 31527 36264 31760 36292
rect 31527 36261 31539 36264
rect 31481 36255 31539 36261
rect 31754 36252 31760 36264
rect 31812 36292 31818 36304
rect 32306 36292 32312 36304
rect 31812 36264 32312 36292
rect 31812 36252 31818 36264
rect 32306 36252 32312 36264
rect 32364 36252 32370 36304
rect 38626 36224 38654 36332
rect 53742 36320 53748 36332
rect 53800 36320 53806 36372
rect 51813 36295 51871 36301
rect 51813 36261 51825 36295
rect 51859 36292 51871 36295
rect 51859 36264 53880 36292
rect 51859 36261 51871 36264
rect 51813 36255 51871 36261
rect 29656 36196 38654 36224
rect 49602 36184 49608 36236
rect 49660 36224 49666 36236
rect 53745 36227 53803 36233
rect 53745 36224 53757 36227
rect 49660 36196 53757 36224
rect 49660 36184 49666 36196
rect 53745 36193 53757 36196
rect 53791 36193 53803 36227
rect 53745 36187 53803 36193
rect 28353 36159 28411 36165
rect 28353 36156 28365 36159
rect 28132 36128 28365 36156
rect 28132 36116 28138 36128
rect 28353 36125 28365 36128
rect 28399 36125 28411 36159
rect 28353 36119 28411 36125
rect 28445 36159 28503 36165
rect 28445 36125 28457 36159
rect 28491 36125 28503 36159
rect 28445 36119 28503 36125
rect 28537 36159 28595 36165
rect 28537 36125 28549 36159
rect 28583 36156 28595 36159
rect 28626 36156 28632 36168
rect 28583 36128 28632 36156
rect 28583 36125 28595 36128
rect 28537 36119 28595 36125
rect 26878 36088 26884 36100
rect 26528 36060 26884 36088
rect 25501 36051 25559 36057
rect 26878 36048 26884 36060
rect 26936 36048 26942 36100
rect 27430 36088 27436 36100
rect 27391 36060 27436 36088
rect 27430 36048 27436 36060
rect 27488 36048 27494 36100
rect 28368 36088 28396 36119
rect 28626 36116 28632 36128
rect 28684 36116 28690 36168
rect 28721 36159 28779 36165
rect 28721 36125 28733 36159
rect 28767 36156 28779 36159
rect 29454 36156 29460 36168
rect 28767 36128 29460 36156
rect 28767 36125 28779 36128
rect 28721 36119 28779 36125
rect 29454 36116 29460 36128
rect 29512 36116 29518 36168
rect 52362 36156 52368 36168
rect 52275 36128 52368 36156
rect 52362 36116 52368 36128
rect 52420 36156 52426 36168
rect 53009 36159 53067 36165
rect 53009 36156 53021 36159
rect 52420 36128 53021 36156
rect 52420 36116 52426 36128
rect 53009 36125 53021 36128
rect 53055 36125 53067 36159
rect 53466 36156 53472 36168
rect 53379 36128 53472 36156
rect 53009 36119 53067 36125
rect 53466 36116 53472 36128
rect 53524 36156 53530 36168
rect 53852 36156 53880 36264
rect 53524 36128 53880 36156
rect 53524 36116 53530 36128
rect 28994 36088 29000 36100
rect 28368 36060 29000 36088
rect 28994 36048 29000 36060
rect 29052 36048 29058 36100
rect 32306 36048 32312 36100
rect 32364 36088 32370 36100
rect 32364 36060 52868 36088
rect 32364 36048 32370 36060
rect 15102 35980 15108 36032
rect 15160 36020 15166 36032
rect 21284 36020 21312 36048
rect 22922 36020 22928 36032
rect 15160 35992 21312 36020
rect 22883 35992 22928 36020
rect 15160 35980 15166 35992
rect 22922 35980 22928 35992
rect 22980 35980 22986 36032
rect 23566 35980 23572 36032
rect 23624 36020 23630 36032
rect 24029 36023 24087 36029
rect 24029 36020 24041 36023
rect 23624 35992 24041 36020
rect 23624 35980 23630 35992
rect 24029 35989 24041 35992
rect 24075 36020 24087 36023
rect 25590 36020 25596 36032
rect 24075 35992 25596 36020
rect 24075 35989 24087 35992
rect 24029 35983 24087 35989
rect 25590 35980 25596 35992
rect 25648 35980 25654 36032
rect 25869 36023 25927 36029
rect 25869 35989 25881 36023
rect 25915 36020 25927 36023
rect 25958 36020 25964 36032
rect 25915 35992 25964 36020
rect 25915 35989 25927 35992
rect 25869 35983 25927 35989
rect 25958 35980 25964 35992
rect 26016 35980 26022 36032
rect 27709 36023 27767 36029
rect 27709 35989 27721 36023
rect 27755 36020 27767 36023
rect 27890 36020 27896 36032
rect 27755 35992 27896 36020
rect 27755 35989 27767 35992
rect 27709 35983 27767 35989
rect 27890 35980 27896 35992
rect 27948 35980 27954 36032
rect 28166 36020 28172 36032
rect 28127 35992 28172 36020
rect 28166 35980 28172 35992
rect 28224 35980 28230 36032
rect 28718 35980 28724 36032
rect 28776 36020 28782 36032
rect 29638 36020 29644 36032
rect 28776 35992 29644 36020
rect 28776 35980 28782 35992
rect 29638 35980 29644 35992
rect 29696 35980 29702 36032
rect 29730 35980 29736 36032
rect 29788 36020 29794 36032
rect 30285 36023 30343 36029
rect 30285 36020 30297 36023
rect 29788 35992 30297 36020
rect 29788 35980 29794 35992
rect 30285 35989 30297 35992
rect 30331 35989 30343 36023
rect 30285 35983 30343 35989
rect 30929 36023 30987 36029
rect 30929 35989 30941 36023
rect 30975 36020 30987 36023
rect 31202 36020 31208 36032
rect 30975 35992 31208 36020
rect 30975 35989 30987 35992
rect 30929 35983 30987 35989
rect 31202 35980 31208 35992
rect 31260 35980 31266 36032
rect 32582 36020 32588 36032
rect 32543 35992 32588 36020
rect 32582 35980 32588 35992
rect 32640 35980 32646 36032
rect 52840 36029 52868 36060
rect 52825 36023 52883 36029
rect 52825 35989 52837 36023
rect 52871 35989 52883 36023
rect 52825 35983 52883 35989
rect 1104 35930 54832 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 54832 35930
rect 1104 35856 54832 35878
rect 20806 35776 20812 35828
rect 20864 35816 20870 35828
rect 20864 35788 22094 35816
rect 20864 35776 20870 35788
rect 22066 35748 22094 35788
rect 22278 35776 22284 35828
rect 22336 35816 22342 35828
rect 23017 35819 23075 35825
rect 23017 35816 23029 35819
rect 22336 35788 23029 35816
rect 22336 35776 22342 35788
rect 23017 35785 23029 35788
rect 23063 35816 23075 35819
rect 23290 35816 23296 35828
rect 23063 35788 23296 35816
rect 23063 35785 23075 35788
rect 23017 35779 23075 35785
rect 23290 35776 23296 35788
rect 23348 35776 23354 35828
rect 23658 35776 23664 35828
rect 23716 35816 23722 35828
rect 24026 35816 24032 35828
rect 23716 35788 23888 35816
rect 23716 35776 23722 35788
rect 23474 35748 23480 35760
rect 22066 35720 23480 35748
rect 23474 35708 23480 35720
rect 23532 35708 23538 35760
rect 23860 35757 23888 35788
rect 23952 35788 24032 35816
rect 23952 35757 23980 35788
rect 24026 35776 24032 35788
rect 24084 35776 24090 35828
rect 24210 35816 24216 35828
rect 24171 35788 24216 35816
rect 24210 35776 24216 35788
rect 24268 35776 24274 35828
rect 25314 35776 25320 35828
rect 25372 35816 25378 35828
rect 26605 35819 26663 35825
rect 25372 35788 26556 35816
rect 25372 35776 25378 35788
rect 23845 35751 23903 35757
rect 23845 35717 23857 35751
rect 23891 35717 23903 35751
rect 23845 35711 23903 35717
rect 23937 35751 23995 35757
rect 23937 35717 23949 35751
rect 23983 35717 23995 35751
rect 23937 35711 23995 35717
rect 24394 35708 24400 35760
rect 24452 35748 24458 35760
rect 25038 35748 25044 35760
rect 24452 35720 24809 35748
rect 24999 35720 25044 35748
rect 24452 35708 24458 35720
rect 2133 35683 2191 35689
rect 2133 35649 2145 35683
rect 2179 35680 2191 35683
rect 15102 35680 15108 35692
rect 2179 35652 15108 35680
rect 2179 35649 2191 35652
rect 2133 35643 2191 35649
rect 15102 35640 15108 35652
rect 15160 35640 15166 35692
rect 23566 35680 23572 35692
rect 23527 35652 23572 35680
rect 23566 35640 23572 35652
rect 23624 35640 23630 35692
rect 23662 35683 23720 35689
rect 23662 35649 23674 35683
rect 23708 35649 23720 35683
rect 23662 35643 23720 35649
rect 2409 35615 2467 35621
rect 2409 35581 2421 35615
rect 2455 35612 2467 35615
rect 2774 35612 2780 35624
rect 2455 35584 2780 35612
rect 2455 35581 2467 35584
rect 2409 35575 2467 35581
rect 2774 35572 2780 35584
rect 2832 35612 2838 35624
rect 2869 35615 2927 35621
rect 2869 35612 2881 35615
rect 2832 35584 2881 35612
rect 2832 35572 2838 35584
rect 2869 35581 2881 35584
rect 2915 35581 2927 35615
rect 23676 35612 23704 35643
rect 23750 35640 23756 35692
rect 23808 35680 23814 35692
rect 24034 35683 24092 35689
rect 24034 35680 24046 35683
rect 23808 35652 24046 35680
rect 23808 35640 23814 35652
rect 24034 35649 24046 35652
rect 24080 35649 24092 35683
rect 24034 35643 24092 35649
rect 2869 35575 2927 35581
rect 20272 35584 23704 35612
rect 24049 35612 24077 35643
rect 24578 35640 24584 35692
rect 24636 35680 24642 35692
rect 24781 35689 24809 35720
rect 25038 35708 25044 35720
rect 25096 35708 25102 35760
rect 26329 35751 26387 35757
rect 26329 35748 26341 35751
rect 25240 35720 26341 35748
rect 24673 35683 24731 35689
rect 24673 35680 24685 35683
rect 24636 35652 24685 35680
rect 24636 35640 24642 35652
rect 24673 35649 24685 35652
rect 24719 35649 24731 35683
rect 24673 35643 24731 35649
rect 24766 35683 24824 35689
rect 24766 35649 24778 35683
rect 24812 35649 24824 35683
rect 24766 35643 24824 35649
rect 24854 35640 24860 35692
rect 24912 35680 24918 35692
rect 24949 35683 25007 35689
rect 24949 35680 24961 35683
rect 24912 35652 24961 35680
rect 24912 35640 24918 35652
rect 24949 35649 24961 35652
rect 24995 35649 25007 35683
rect 24949 35643 25007 35649
rect 25138 35683 25196 35689
rect 25138 35649 25150 35683
rect 25184 35649 25196 35683
rect 25138 35643 25196 35649
rect 25153 35612 25181 35643
rect 24049 35584 25181 35612
rect 2498 35436 2504 35488
rect 2556 35476 2562 35488
rect 20272 35485 20300 35584
rect 22554 35544 22560 35556
rect 22467 35516 22560 35544
rect 22554 35504 22560 35516
rect 22612 35544 22618 35556
rect 25240 35544 25268 35720
rect 26329 35717 26341 35720
rect 26375 35717 26387 35751
rect 26329 35711 26387 35717
rect 26053 35683 26111 35689
rect 26053 35649 26065 35683
rect 26099 35680 26111 35683
rect 26142 35680 26148 35692
rect 26099 35652 26148 35680
rect 26099 35649 26111 35652
rect 26053 35643 26111 35649
rect 26142 35640 26148 35652
rect 26200 35640 26206 35692
rect 26237 35683 26295 35689
rect 26237 35649 26249 35683
rect 26283 35649 26295 35683
rect 26418 35680 26424 35692
rect 26379 35652 26424 35680
rect 26237 35643 26295 35649
rect 25590 35572 25596 35624
rect 25648 35612 25654 35624
rect 26252 35612 26280 35643
rect 26418 35640 26424 35652
rect 26476 35640 26482 35692
rect 26528 35680 26556 35788
rect 26605 35785 26617 35819
rect 26651 35816 26663 35819
rect 27154 35816 27160 35828
rect 26651 35788 27160 35816
rect 26651 35785 26663 35788
rect 26605 35779 26663 35785
rect 27154 35776 27160 35788
rect 27212 35776 27218 35828
rect 27632 35788 31616 35816
rect 27522 35748 27528 35760
rect 27483 35720 27528 35748
rect 27522 35708 27528 35720
rect 27580 35708 27586 35760
rect 27295 35683 27353 35689
rect 27295 35680 27307 35683
rect 26528 35652 27307 35680
rect 27295 35649 27307 35652
rect 27341 35649 27353 35683
rect 27430 35680 27436 35692
rect 27391 35652 27436 35680
rect 27295 35643 27353 35649
rect 27430 35640 27436 35652
rect 27488 35640 27494 35692
rect 27632 35680 27660 35788
rect 28718 35708 28724 35760
rect 28776 35748 28782 35760
rect 28776 35720 28821 35748
rect 28776 35708 28782 35720
rect 29086 35708 29092 35760
rect 29144 35748 29150 35760
rect 29365 35751 29423 35757
rect 29365 35748 29377 35751
rect 29144 35720 29377 35748
rect 29144 35708 29150 35720
rect 29365 35717 29377 35720
rect 29411 35717 29423 35751
rect 29365 35711 29423 35717
rect 29564 35720 31524 35748
rect 27708 35683 27766 35689
rect 27708 35680 27720 35683
rect 27632 35652 27720 35680
rect 27708 35649 27720 35652
rect 27754 35649 27766 35683
rect 27708 35643 27766 35649
rect 27801 35683 27859 35689
rect 27801 35649 27813 35683
rect 27847 35649 27859 35683
rect 28350 35680 28356 35692
rect 28311 35652 28356 35680
rect 27801 35643 27859 35649
rect 27816 35612 27844 35643
rect 28350 35640 28356 35652
rect 28408 35640 28414 35692
rect 28534 35640 28540 35692
rect 28592 35680 28598 35692
rect 29564 35680 29592 35720
rect 28592 35652 29592 35680
rect 28592 35640 28598 35652
rect 29638 35640 29644 35692
rect 29696 35680 29702 35692
rect 29917 35683 29975 35689
rect 29917 35680 29929 35683
rect 29696 35652 29929 35680
rect 29696 35640 29702 35652
rect 29917 35649 29929 35652
rect 29963 35649 29975 35683
rect 29917 35643 29975 35649
rect 30006 35640 30012 35692
rect 30064 35680 30070 35692
rect 30193 35683 30251 35689
rect 30064 35652 30109 35680
rect 30064 35640 30070 35652
rect 30193 35649 30205 35683
rect 30239 35649 30251 35683
rect 30193 35643 30251 35649
rect 25648 35584 26280 35612
rect 26436 35584 27844 35612
rect 25648 35572 25654 35584
rect 26160 35556 26188 35584
rect 22612 35516 25268 35544
rect 22612 35504 22618 35516
rect 26142 35504 26148 35556
rect 26200 35504 26206 35556
rect 20257 35479 20315 35485
rect 20257 35476 20269 35479
rect 2556 35448 20269 35476
rect 2556 35436 2562 35448
rect 20257 35445 20269 35448
rect 20303 35445 20315 35479
rect 20806 35476 20812 35488
rect 20767 35448 20812 35476
rect 20257 35439 20315 35445
rect 20806 35436 20812 35448
rect 20864 35436 20870 35488
rect 21453 35479 21511 35485
rect 21453 35445 21465 35479
rect 21499 35476 21511 35479
rect 23014 35476 23020 35488
rect 21499 35448 23020 35476
rect 21499 35445 21511 35448
rect 21453 35439 21511 35445
rect 23014 35436 23020 35448
rect 23072 35436 23078 35488
rect 23290 35436 23296 35488
rect 23348 35476 23354 35488
rect 24210 35476 24216 35488
rect 23348 35448 24216 35476
rect 23348 35436 23354 35448
rect 24210 35436 24216 35448
rect 24268 35436 24274 35488
rect 25317 35479 25375 35485
rect 25317 35445 25329 35479
rect 25363 35476 25375 35479
rect 25866 35476 25872 35488
rect 25363 35448 25872 35476
rect 25363 35445 25375 35448
rect 25317 35439 25375 35445
rect 25866 35436 25872 35448
rect 25924 35436 25930 35488
rect 25958 35436 25964 35488
rect 26016 35476 26022 35488
rect 26436 35476 26464 35584
rect 28626 35572 28632 35624
rect 28684 35612 28690 35624
rect 29454 35612 29460 35624
rect 28684 35584 29460 35612
rect 28684 35572 28690 35584
rect 29454 35572 29460 35584
rect 29512 35612 29518 35624
rect 30208 35612 30236 35643
rect 30282 35640 30288 35692
rect 30340 35680 30346 35692
rect 30340 35652 30385 35680
rect 30340 35640 30346 35652
rect 30469 35615 30527 35621
rect 29512 35584 30144 35612
rect 30208 35584 30420 35612
rect 29512 35572 29518 35584
rect 26510 35504 26516 35556
rect 26568 35544 26574 35556
rect 30116 35544 30144 35584
rect 30282 35544 30288 35556
rect 26568 35516 29409 35544
rect 30116 35516 30288 35544
rect 26568 35504 26574 35516
rect 27154 35476 27160 35488
rect 26016 35448 26464 35476
rect 27115 35448 27160 35476
rect 26016 35436 26022 35448
rect 27154 35436 27160 35448
rect 27212 35436 27218 35488
rect 28626 35436 28632 35488
rect 28684 35476 28690 35488
rect 28902 35476 28908 35488
rect 28684 35448 28908 35476
rect 28684 35436 28690 35448
rect 28902 35436 28908 35448
rect 28960 35436 28966 35488
rect 29086 35436 29092 35488
rect 29144 35476 29150 35488
rect 29273 35479 29331 35485
rect 29273 35476 29285 35479
rect 29144 35448 29285 35476
rect 29144 35436 29150 35448
rect 29273 35445 29285 35448
rect 29319 35445 29331 35479
rect 29381 35476 29409 35516
rect 30282 35504 30288 35516
rect 30340 35504 30346 35556
rect 30392 35544 30420 35584
rect 30469 35581 30481 35615
rect 30515 35612 30527 35615
rect 31386 35612 31392 35624
rect 30515 35584 31392 35612
rect 30515 35581 30527 35584
rect 30469 35575 30527 35581
rect 31386 35572 31392 35584
rect 31444 35572 31450 35624
rect 31496 35612 31524 35720
rect 31588 35680 31616 35788
rect 33686 35776 33692 35828
rect 33744 35816 33750 35828
rect 54018 35816 54024 35828
rect 33744 35788 54024 35816
rect 33744 35776 33750 35788
rect 54018 35776 54024 35788
rect 54076 35776 54082 35828
rect 32401 35683 32459 35689
rect 32401 35680 32413 35683
rect 31588 35652 32413 35680
rect 32401 35649 32413 35652
rect 32447 35680 32459 35683
rect 44174 35680 44180 35692
rect 32447 35652 44180 35680
rect 32447 35649 32459 35652
rect 32401 35643 32459 35649
rect 44174 35640 44180 35652
rect 44232 35640 44238 35692
rect 33686 35612 33692 35624
rect 31496 35584 33692 35612
rect 33686 35572 33692 35584
rect 33744 35572 33750 35624
rect 52365 35615 52423 35621
rect 52365 35581 52377 35615
rect 52411 35612 52423 35615
rect 53466 35612 53472 35624
rect 52411 35584 53472 35612
rect 52411 35581 52423 35584
rect 52365 35575 52423 35581
rect 53466 35572 53472 35584
rect 53524 35572 53530 35624
rect 53745 35615 53803 35621
rect 53745 35581 53757 35615
rect 53791 35581 53803 35615
rect 53745 35575 53803 35581
rect 32953 35547 33011 35553
rect 30392 35516 31754 35544
rect 29638 35476 29644 35488
rect 29381 35448 29644 35476
rect 29273 35439 29331 35445
rect 29638 35436 29644 35448
rect 29696 35436 29702 35488
rect 30300 35476 30328 35504
rect 30834 35476 30840 35488
rect 30300 35448 30840 35476
rect 30834 35436 30840 35448
rect 30892 35436 30898 35488
rect 31018 35476 31024 35488
rect 30979 35448 31024 35476
rect 31018 35436 31024 35448
rect 31076 35436 31082 35488
rect 31478 35436 31484 35488
rect 31536 35476 31542 35488
rect 31573 35479 31631 35485
rect 31573 35476 31585 35479
rect 31536 35448 31585 35476
rect 31536 35436 31542 35448
rect 31573 35445 31585 35448
rect 31619 35445 31631 35479
rect 31726 35476 31754 35516
rect 32953 35513 32965 35547
rect 32999 35544 33011 35547
rect 53760 35544 53788 35575
rect 32999 35516 53788 35544
rect 32999 35513 33011 35516
rect 32953 35507 33011 35513
rect 32968 35476 32996 35507
rect 31726 35448 32996 35476
rect 53009 35479 53067 35485
rect 31573 35439 31631 35445
rect 53009 35445 53021 35479
rect 53055 35476 53067 35479
rect 53558 35476 53564 35488
rect 53055 35448 53564 35476
rect 53055 35445 53067 35448
rect 53009 35439 53067 35445
rect 53558 35436 53564 35448
rect 53616 35436 53622 35488
rect 1104 35386 54832 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 54832 35386
rect 1104 35312 54832 35334
rect 15102 35232 15108 35284
rect 15160 35272 15166 35284
rect 16577 35275 16635 35281
rect 16577 35272 16589 35275
rect 15160 35244 16589 35272
rect 15160 35232 15166 35244
rect 16577 35241 16589 35244
rect 16623 35241 16635 35275
rect 16577 35235 16635 35241
rect 16666 35232 16672 35284
rect 16724 35272 16730 35284
rect 27614 35272 27620 35284
rect 16724 35244 27620 35272
rect 16724 35232 16730 35244
rect 27614 35232 27620 35244
rect 27672 35232 27678 35284
rect 27985 35275 28043 35281
rect 27985 35241 27997 35275
rect 28031 35272 28043 35275
rect 28442 35272 28448 35284
rect 28031 35244 28448 35272
rect 28031 35241 28043 35244
rect 27985 35235 28043 35241
rect 28442 35232 28448 35244
rect 28500 35232 28506 35284
rect 29178 35272 29184 35284
rect 28552 35244 28949 35272
rect 29139 35244 29184 35272
rect 15010 35164 15016 35216
rect 15068 35164 15074 35216
rect 15473 35207 15531 35213
rect 15473 35173 15485 35207
rect 15519 35204 15531 35207
rect 26510 35204 26516 35216
rect 15519 35176 26516 35204
rect 15519 35173 15531 35176
rect 15473 35167 15531 35173
rect 26510 35164 26516 35176
rect 26568 35164 26574 35216
rect 27062 35204 27068 35216
rect 27023 35176 27068 35204
rect 27062 35164 27068 35176
rect 27120 35164 27126 35216
rect 14550 35096 14556 35148
rect 14608 35136 14614 35148
rect 15028 35136 15056 35164
rect 15933 35139 15991 35145
rect 15933 35136 15945 35139
rect 14608 35108 14964 35136
rect 15028 35108 15945 35136
rect 14608 35096 14614 35108
rect 1578 35068 1584 35080
rect 1539 35040 1584 35068
rect 1578 35028 1584 35040
rect 1636 35068 1642 35080
rect 14936 35077 14964 35108
rect 15212 35077 15240 35108
rect 15933 35105 15945 35108
rect 15979 35105 15991 35139
rect 21174 35136 21180 35148
rect 21135 35108 21180 35136
rect 15933 35099 15991 35105
rect 21174 35096 21180 35108
rect 21232 35096 21238 35148
rect 22281 35139 22339 35145
rect 22281 35105 22293 35139
rect 22327 35136 22339 35139
rect 25590 35136 25596 35148
rect 22327 35108 23336 35136
rect 22327 35105 22339 35108
rect 22281 35099 22339 35105
rect 23308 35080 23336 35108
rect 23768 35108 25596 35136
rect 2777 35071 2835 35077
rect 2777 35068 2789 35071
rect 1636 35040 2789 35068
rect 1636 35028 1642 35040
rect 2777 35037 2789 35040
rect 2823 35037 2835 35071
rect 2777 35031 2835 35037
rect 14829 35071 14887 35077
rect 14829 35037 14841 35071
rect 14875 35037 14887 35071
rect 14829 35031 14887 35037
rect 14922 35071 14980 35077
rect 14922 35037 14934 35071
rect 14968 35037 14980 35071
rect 14922 35031 14980 35037
rect 15197 35071 15255 35077
rect 15197 35037 15209 35071
rect 15243 35037 15255 35071
rect 15197 35031 15255 35037
rect 15335 35071 15393 35077
rect 15335 35037 15347 35071
rect 15381 35068 15393 35071
rect 15654 35068 15660 35080
rect 15381 35040 15660 35068
rect 15381 35037 15393 35040
rect 15335 35031 15393 35037
rect 1762 34932 1768 34944
rect 1723 34904 1768 34932
rect 1762 34892 1768 34904
rect 1820 34892 1826 34944
rect 2317 34935 2375 34941
rect 2317 34901 2329 34935
rect 2363 34932 2375 34935
rect 2774 34932 2780 34944
rect 2363 34904 2780 34932
rect 2363 34901 2375 34904
rect 2317 34895 2375 34901
rect 2774 34892 2780 34904
rect 2832 34892 2838 34944
rect 14369 34935 14427 34941
rect 14369 34901 14381 34935
rect 14415 34932 14427 34935
rect 14550 34932 14556 34944
rect 14415 34904 14556 34932
rect 14415 34901 14427 34904
rect 14369 34895 14427 34901
rect 14550 34892 14556 34904
rect 14608 34892 14614 34944
rect 14844 34932 14872 35031
rect 15654 35028 15660 35040
rect 15712 35068 15718 35080
rect 19334 35068 19340 35080
rect 15712 35040 19340 35068
rect 15712 35028 15718 35040
rect 19334 35028 19340 35040
rect 19392 35028 19398 35080
rect 21726 35068 21732 35080
rect 21687 35040 21732 35068
rect 21726 35028 21732 35040
rect 21784 35028 21790 35080
rect 22833 35071 22891 35077
rect 22833 35037 22845 35071
rect 22879 35068 22891 35071
rect 23106 35068 23112 35080
rect 22879 35040 23112 35068
rect 22879 35037 22891 35040
rect 22833 35031 22891 35037
rect 23106 35028 23112 35040
rect 23164 35028 23170 35080
rect 23290 35028 23296 35080
rect 23348 35028 23354 35080
rect 23474 35077 23480 35080
rect 23453 35071 23480 35077
rect 23453 35037 23465 35071
rect 23532 35068 23538 35080
rect 23768 35068 23796 35108
rect 25590 35096 25596 35108
rect 25648 35096 25654 35148
rect 27154 35136 27160 35148
rect 26068 35108 27160 35136
rect 23532 35040 23796 35068
rect 23453 35031 23480 35037
rect 23474 35028 23480 35031
rect 23532 35028 23538 35040
rect 23842 35028 23848 35080
rect 23900 35068 23906 35080
rect 25133 35071 25191 35077
rect 23900 35040 23945 35068
rect 23900 35028 23906 35040
rect 25133 35037 25145 35071
rect 25179 35068 25191 35071
rect 25685 35071 25743 35077
rect 25685 35068 25697 35071
rect 25179 35040 25697 35068
rect 25179 35037 25191 35040
rect 25133 35031 25191 35037
rect 25685 35037 25697 35040
rect 25731 35037 25743 35071
rect 25866 35068 25872 35080
rect 25827 35040 25872 35068
rect 25685 35031 25743 35037
rect 25866 35028 25872 35040
rect 25924 35028 25930 35080
rect 26068 35077 26096 35108
rect 27154 35096 27160 35108
rect 27212 35096 27218 35148
rect 26053 35071 26111 35077
rect 26053 35037 26065 35071
rect 26099 35037 26111 35071
rect 26510 35068 26516 35080
rect 26471 35040 26516 35068
rect 26053 35031 26111 35037
rect 26510 35028 26516 35040
rect 26568 35028 26574 35080
rect 26694 35068 26700 35080
rect 26655 35040 26700 35068
rect 26694 35028 26700 35040
rect 26752 35028 26758 35080
rect 26786 35028 26792 35080
rect 26844 35068 26850 35080
rect 26933 35071 26991 35077
rect 26844 35040 26889 35068
rect 26844 35028 26850 35040
rect 26933 35037 26945 35071
rect 26979 35068 26991 35071
rect 28552 35068 28580 35244
rect 28921 35136 28949 35244
rect 29178 35232 29184 35244
rect 29236 35232 29242 35284
rect 31018 35272 31024 35284
rect 30300 35244 31024 35272
rect 29086 35164 29092 35216
rect 29144 35204 29150 35216
rect 29638 35204 29644 35216
rect 29144 35176 29644 35204
rect 29144 35164 29150 35176
rect 29638 35164 29644 35176
rect 29696 35164 29702 35216
rect 30300 35136 30328 35244
rect 31018 35232 31024 35244
rect 31076 35272 31082 35284
rect 31076 35244 45554 35272
rect 31076 35232 31082 35244
rect 30374 35164 30380 35216
rect 30432 35204 30438 35216
rect 32217 35207 32275 35213
rect 32217 35204 32229 35207
rect 30432 35176 32229 35204
rect 30432 35164 30438 35176
rect 32217 35173 32229 35176
rect 32263 35173 32275 35207
rect 32217 35167 32275 35173
rect 32861 35207 32919 35213
rect 32861 35173 32873 35207
rect 32907 35204 32919 35207
rect 35802 35204 35808 35216
rect 32907 35176 35808 35204
rect 32907 35173 32919 35176
rect 32861 35167 32919 35173
rect 32876 35136 32904 35167
rect 35802 35164 35808 35176
rect 35860 35164 35866 35216
rect 28921 35108 30328 35136
rect 30504 35108 32904 35136
rect 45526 35136 45554 35244
rect 53745 35139 53803 35145
rect 53745 35136 53757 35139
rect 45526 35108 53757 35136
rect 28629 35071 28687 35077
rect 28629 35068 28641 35071
rect 26979 35040 27200 35068
rect 28552 35040 28641 35068
rect 26979 35037 26991 35040
rect 26933 35031 26991 35037
rect 15010 34960 15016 35012
rect 15068 35000 15074 35012
rect 15105 35003 15163 35009
rect 15105 35000 15117 35003
rect 15068 34972 15117 35000
rect 15068 34960 15074 34972
rect 15105 34969 15117 34972
rect 15151 34969 15163 35003
rect 23308 35000 23336 35028
rect 27172 35012 27200 35040
rect 28629 35037 28641 35040
rect 28675 35037 28687 35071
rect 28629 35031 28687 35037
rect 29043 35071 29101 35077
rect 29043 35037 29055 35071
rect 29089 35068 29101 35071
rect 29089 35040 29592 35068
rect 29089 35037 29101 35040
rect 29043 35031 29101 35037
rect 23569 35003 23627 35009
rect 23569 35000 23581 35003
rect 15105 34963 15163 34969
rect 15396 34972 23152 35000
rect 23308 34972 23581 35000
rect 15396 34932 15424 34972
rect 14844 34904 15424 34932
rect 23124 34932 23152 34972
rect 23569 34969 23581 34972
rect 23615 34969 23627 35003
rect 23569 34963 23627 34969
rect 23658 34960 23664 35012
rect 23716 35000 23722 35012
rect 23716 34972 23761 35000
rect 23716 34960 23722 34972
rect 25958 34960 25964 35012
rect 26016 35000 26022 35012
rect 26326 35000 26332 35012
rect 26016 34972 26332 35000
rect 26016 34960 26022 34972
rect 26326 34960 26332 34972
rect 26384 35000 26390 35012
rect 27062 35000 27068 35012
rect 26384 34972 27068 35000
rect 26384 34960 26390 34972
rect 27062 34960 27068 34972
rect 27120 34960 27126 35012
rect 27154 34960 27160 35012
rect 27212 34960 27218 35012
rect 28077 35003 28135 35009
rect 28077 34969 28089 35003
rect 28123 35000 28135 35003
rect 28258 35000 28264 35012
rect 28123 34972 28264 35000
rect 28123 34969 28135 34972
rect 28077 34963 28135 34969
rect 28258 34960 28264 34972
rect 28316 34960 28322 35012
rect 28718 34960 28724 35012
rect 28776 35000 28782 35012
rect 28813 35003 28871 35009
rect 28813 35000 28825 35003
rect 28776 34972 28825 35000
rect 28776 34960 28782 34972
rect 28813 34969 28825 34972
rect 28859 34969 28871 35003
rect 28813 34963 28871 34969
rect 28905 35003 28963 35009
rect 28905 34969 28917 35003
rect 28951 34969 28963 35003
rect 29564 35000 29592 35040
rect 29638 35028 29644 35080
rect 29696 35068 29702 35080
rect 30101 35071 30159 35077
rect 30101 35068 30113 35071
rect 29696 35040 30113 35068
rect 29696 35028 29702 35040
rect 30101 35037 30113 35040
rect 30147 35037 30159 35071
rect 30101 35031 30159 35037
rect 30249 35071 30307 35077
rect 30249 35037 30261 35071
rect 30295 35068 30307 35071
rect 30504 35068 30532 35108
rect 53745 35105 53757 35108
rect 53791 35105 53803 35139
rect 53745 35099 53803 35105
rect 30650 35077 30656 35080
rect 30295 35040 30532 35068
rect 30607 35071 30656 35077
rect 30295 35037 30307 35040
rect 30249 35031 30307 35037
rect 30607 35037 30619 35071
rect 30653 35037 30656 35071
rect 30607 35031 30656 35037
rect 30650 35028 30656 35031
rect 30708 35028 30714 35080
rect 30926 35068 30932 35080
rect 30760 35040 30932 35068
rect 29730 35000 29736 35012
rect 29564 34972 29736 35000
rect 28905 34963 28963 34969
rect 23293 34935 23351 34941
rect 23293 34932 23305 34935
rect 23124 34904 23305 34932
rect 23293 34901 23305 34904
rect 23339 34901 23351 34935
rect 25038 34932 25044 34944
rect 24999 34904 25044 34932
rect 23293 34895 23351 34901
rect 25038 34892 25044 34904
rect 25096 34892 25102 34944
rect 28920 34932 28948 34963
rect 29730 34960 29736 34972
rect 29788 34960 29794 35012
rect 30374 35000 30380 35012
rect 30116 34972 30380 35000
rect 30116 34944 30144 34972
rect 30374 34960 30380 34972
rect 30432 34960 30438 35012
rect 30469 35003 30527 35009
rect 30469 34969 30481 35003
rect 30515 34969 30527 35003
rect 30469 34963 30527 34969
rect 28994 34932 29000 34944
rect 28920 34904 29000 34932
rect 28994 34892 29000 34904
rect 29052 34892 29058 34944
rect 30098 34892 30104 34944
rect 30156 34892 30162 34944
rect 30484 34932 30512 34963
rect 30558 34932 30564 34944
rect 30484 34904 30564 34932
rect 30558 34892 30564 34904
rect 30616 34892 30622 34944
rect 30760 34941 30788 35040
rect 30926 35028 30932 35040
rect 30984 35028 30990 35080
rect 31110 35028 31116 35080
rect 31168 35068 31174 35080
rect 31481 35071 31539 35077
rect 31481 35068 31493 35071
rect 31168 35040 31493 35068
rect 31168 35028 31174 35040
rect 31481 35037 31493 35040
rect 31527 35037 31539 35071
rect 31481 35031 31539 35037
rect 53009 35071 53067 35077
rect 53009 35037 53021 35071
rect 53055 35068 53067 35071
rect 53282 35068 53288 35080
rect 53055 35040 53288 35068
rect 53055 35037 53067 35040
rect 53009 35031 53067 35037
rect 53282 35028 53288 35040
rect 53340 35028 53346 35080
rect 53469 35071 53527 35077
rect 53469 35037 53481 35071
rect 53515 35068 53527 35071
rect 53558 35068 53564 35080
rect 53515 35040 53564 35068
rect 53515 35037 53527 35040
rect 53469 35031 53527 35037
rect 53558 35028 53564 35040
rect 53616 35028 53622 35080
rect 30745 34935 30803 34941
rect 30745 34901 30757 34935
rect 30791 34901 30803 34935
rect 30745 34895 30803 34901
rect 30834 34892 30840 34944
rect 30892 34932 30898 34944
rect 31665 34935 31723 34941
rect 31665 34932 31677 34935
rect 30892 34904 31677 34932
rect 30892 34892 30898 34904
rect 31665 34901 31677 34904
rect 31711 34901 31723 34935
rect 31665 34895 31723 34901
rect 33413 34935 33471 34941
rect 33413 34901 33425 34935
rect 33459 34932 33471 34935
rect 33502 34932 33508 34944
rect 33459 34904 33508 34932
rect 33459 34901 33471 34904
rect 33413 34895 33471 34901
rect 33502 34892 33508 34904
rect 33560 34892 33566 34944
rect 1104 34842 54832 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 54832 34842
rect 1104 34768 54832 34790
rect 1762 34688 1768 34740
rect 1820 34728 1826 34740
rect 23474 34728 23480 34740
rect 1820 34700 23480 34728
rect 1820 34688 1826 34700
rect 23474 34688 23480 34700
rect 23532 34688 23538 34740
rect 23566 34688 23572 34740
rect 23624 34728 23630 34740
rect 24581 34731 24639 34737
rect 24581 34728 24593 34731
rect 23624 34700 24593 34728
rect 23624 34688 23630 34700
rect 24581 34697 24593 34700
rect 24627 34697 24639 34731
rect 24581 34691 24639 34697
rect 25593 34731 25651 34737
rect 25593 34697 25605 34731
rect 25639 34728 25651 34731
rect 25682 34728 25688 34740
rect 25639 34700 25688 34728
rect 25639 34697 25651 34700
rect 25593 34691 25651 34697
rect 25682 34688 25688 34700
rect 25740 34688 25746 34740
rect 25774 34688 25780 34740
rect 25832 34728 25838 34740
rect 27341 34731 27399 34737
rect 27341 34728 27353 34731
rect 25832 34700 27353 34728
rect 25832 34688 25838 34700
rect 27341 34697 27353 34700
rect 27387 34697 27399 34731
rect 28534 34728 28540 34740
rect 27341 34691 27399 34697
rect 28276 34700 28540 34728
rect 22554 34660 22560 34672
rect 6886 34632 22560 34660
rect 2133 34595 2191 34601
rect 2133 34561 2145 34595
rect 2179 34592 2191 34595
rect 6886 34592 6914 34632
rect 22554 34620 22560 34632
rect 22612 34620 22618 34672
rect 23934 34660 23940 34672
rect 23032 34632 23940 34660
rect 2179 34564 6914 34592
rect 14001 34595 14059 34601
rect 2179 34561 2191 34564
rect 2133 34555 2191 34561
rect 14001 34561 14013 34595
rect 14047 34561 14059 34595
rect 14001 34555 14059 34561
rect 14185 34595 14243 34601
rect 14185 34561 14197 34595
rect 14231 34561 14243 34595
rect 14185 34555 14243 34561
rect 2409 34527 2467 34533
rect 2409 34493 2421 34527
rect 2455 34524 2467 34527
rect 2774 34524 2780 34536
rect 2455 34496 2780 34524
rect 2455 34493 2467 34496
rect 2409 34487 2467 34493
rect 2774 34484 2780 34496
rect 2832 34484 2838 34536
rect 13446 34524 13452 34536
rect 13407 34496 13452 34524
rect 13446 34484 13452 34496
rect 13504 34524 13510 34536
rect 14016 34524 14044 34555
rect 13504 34496 14044 34524
rect 14200 34524 14228 34555
rect 14274 34552 14280 34604
rect 14332 34592 14338 34604
rect 14415 34595 14473 34601
rect 14332 34564 14377 34592
rect 14332 34552 14338 34564
rect 14415 34561 14427 34595
rect 14461 34592 14473 34595
rect 14734 34592 14740 34604
rect 14461 34564 14740 34592
rect 14461 34561 14473 34564
rect 14415 34555 14473 34561
rect 14734 34552 14740 34564
rect 14792 34592 14798 34604
rect 15654 34592 15660 34604
rect 14792 34564 15660 34592
rect 14792 34552 14798 34564
rect 15654 34552 15660 34564
rect 15712 34552 15718 34604
rect 15010 34524 15016 34536
rect 14200 34496 15016 34524
rect 13504 34484 13510 34496
rect 15010 34484 15016 34496
rect 15068 34484 15074 34536
rect 16666 34524 16672 34536
rect 15120 34496 16672 34524
rect 14553 34459 14611 34465
rect 14553 34425 14565 34459
rect 14599 34456 14611 34459
rect 15120 34456 15148 34496
rect 16666 34484 16672 34496
rect 16724 34484 16730 34536
rect 17862 34484 17868 34536
rect 17920 34524 17926 34536
rect 21361 34527 21419 34533
rect 21361 34524 21373 34527
rect 17920 34496 21373 34524
rect 17920 34484 17926 34496
rect 21361 34493 21373 34496
rect 21407 34524 21419 34527
rect 23032 34524 23060 34632
rect 23934 34620 23940 34632
rect 23992 34620 23998 34672
rect 24210 34660 24216 34672
rect 24171 34632 24216 34660
rect 24210 34620 24216 34632
rect 24268 34620 24274 34672
rect 25314 34660 25320 34672
rect 25275 34632 25320 34660
rect 25314 34620 25320 34632
rect 25372 34620 25378 34672
rect 25700 34660 25728 34688
rect 25958 34660 25964 34672
rect 25700 34632 25964 34660
rect 25958 34620 25964 34632
rect 26016 34620 26022 34672
rect 26234 34660 26240 34672
rect 26195 34632 26240 34660
rect 26234 34620 26240 34632
rect 26292 34620 26298 34672
rect 27614 34660 27620 34672
rect 26344 34632 27620 34660
rect 23474 34552 23480 34604
rect 23532 34592 23538 34604
rect 24029 34595 24087 34601
rect 24029 34592 24041 34595
rect 23532 34564 24041 34592
rect 23532 34552 23538 34564
rect 24029 34561 24041 34564
rect 24075 34561 24087 34595
rect 24029 34555 24087 34561
rect 24302 34552 24308 34604
rect 24360 34592 24366 34604
rect 24443 34595 24501 34601
rect 24360 34564 24405 34592
rect 24360 34552 24366 34564
rect 24443 34561 24455 34595
rect 24489 34592 24501 34595
rect 25332 34592 25360 34620
rect 25498 34592 25504 34604
rect 24489 34564 25504 34592
rect 24489 34561 24501 34564
rect 24443 34555 24501 34561
rect 25498 34552 25504 34564
rect 25556 34552 25562 34604
rect 26344 34592 26372 34632
rect 27614 34620 27620 34632
rect 27672 34660 27678 34672
rect 28276 34660 28304 34700
rect 28534 34688 28540 34700
rect 28592 34688 28598 34740
rect 29730 34688 29736 34740
rect 29788 34728 29794 34740
rect 29914 34728 29920 34740
rect 29788 34700 29920 34728
rect 29788 34688 29794 34700
rect 29914 34688 29920 34700
rect 29972 34688 29978 34740
rect 31478 34728 31484 34740
rect 30612 34700 31484 34728
rect 30612 34660 30640 34700
rect 31478 34688 31484 34700
rect 31536 34688 31542 34740
rect 32401 34731 32459 34737
rect 32401 34697 32413 34731
rect 32447 34728 32459 34731
rect 32447 34700 53788 34728
rect 32447 34697 32459 34700
rect 32401 34691 32459 34697
rect 32306 34660 32312 34672
rect 27672 34632 28304 34660
rect 28368 34632 30640 34660
rect 30668 34632 32312 34660
rect 27672 34620 27678 34632
rect 26068 34564 26372 34592
rect 21407 34496 23060 34524
rect 23569 34527 23627 34533
rect 21407 34493 21419 34496
rect 21361 34487 21419 34493
rect 23569 34493 23581 34527
rect 23615 34524 23627 34527
rect 24320 34524 24348 34552
rect 23615 34496 24348 34524
rect 23615 34493 23627 34496
rect 23569 34487 23627 34493
rect 24578 34484 24584 34536
rect 24636 34524 24642 34536
rect 26068 34524 26096 34564
rect 27062 34552 27068 34604
rect 27120 34592 27126 34604
rect 27249 34595 27307 34601
rect 27249 34592 27261 34595
rect 27120 34564 27261 34592
rect 27120 34552 27126 34564
rect 27249 34561 27261 34564
rect 27295 34561 27307 34595
rect 27249 34555 27307 34561
rect 28074 34552 28080 34604
rect 28132 34592 28138 34604
rect 28368 34601 28396 34632
rect 28261 34595 28319 34601
rect 28261 34592 28273 34595
rect 28132 34564 28273 34592
rect 28132 34552 28138 34564
rect 28261 34561 28273 34564
rect 28307 34561 28319 34595
rect 28261 34555 28319 34561
rect 28353 34595 28411 34601
rect 28353 34561 28365 34595
rect 28399 34561 28411 34595
rect 28534 34592 28540 34604
rect 28495 34564 28540 34592
rect 28353 34555 28411 34561
rect 28534 34552 28540 34564
rect 28592 34552 28598 34604
rect 28626 34552 28632 34604
rect 28684 34592 28690 34604
rect 29270 34592 29276 34604
rect 28684 34564 28777 34592
rect 29231 34564 29276 34592
rect 28684 34552 28690 34564
rect 29270 34552 29276 34564
rect 29328 34552 29334 34604
rect 29366 34595 29424 34601
rect 29366 34561 29378 34595
rect 29412 34561 29424 34595
rect 29366 34555 29424 34561
rect 24636 34496 26096 34524
rect 24636 34484 24642 34496
rect 23014 34456 23020 34468
rect 14599 34428 15148 34456
rect 22975 34428 23020 34456
rect 14599 34425 14611 34428
rect 14553 34419 14611 34425
rect 23014 34416 23020 34428
rect 23072 34416 23078 34468
rect 28644 34456 28672 34552
rect 29381 34524 29409 34555
rect 29454 34552 29460 34604
rect 29512 34592 29518 34604
rect 29549 34595 29607 34601
rect 29549 34592 29561 34595
rect 29512 34564 29561 34592
rect 29512 34552 29518 34564
rect 29549 34561 29561 34564
rect 29595 34561 29607 34595
rect 29549 34555 29607 34561
rect 29638 34552 29644 34604
rect 29696 34592 29702 34604
rect 29779 34595 29837 34601
rect 29696 34564 29741 34592
rect 29696 34552 29702 34564
rect 29779 34561 29791 34595
rect 29825 34592 29837 34595
rect 29914 34592 29920 34604
rect 29825 34564 29920 34592
rect 29825 34561 29837 34564
rect 29779 34555 29837 34561
rect 29914 34552 29920 34564
rect 29972 34552 29978 34604
rect 30374 34592 30380 34604
rect 30335 34564 30380 34592
rect 30374 34552 30380 34564
rect 30432 34552 30438 34604
rect 30466 34552 30472 34604
rect 30524 34592 30530 34604
rect 30668 34601 30696 34632
rect 32306 34620 32312 34632
rect 32364 34620 32370 34672
rect 30653 34595 30711 34601
rect 30524 34564 30569 34592
rect 30524 34552 30530 34564
rect 30653 34561 30665 34595
rect 30699 34561 30711 34595
rect 30653 34555 30711 34561
rect 30745 34595 30803 34601
rect 30745 34561 30757 34595
rect 30791 34592 30803 34595
rect 32416 34592 32444 34691
rect 51721 34663 51779 34669
rect 51721 34629 51733 34663
rect 51767 34660 51779 34663
rect 51767 34632 53512 34660
rect 51767 34629 51779 34632
rect 51721 34623 51779 34629
rect 53484 34604 53512 34632
rect 43898 34592 43904 34604
rect 30791 34564 30880 34592
rect 30791 34561 30803 34564
rect 30745 34555 30803 34561
rect 30852 34524 30880 34564
rect 31036 34564 32444 34592
rect 41386 34564 43904 34592
rect 30926 34524 30932 34536
rect 29381 34496 30512 34524
rect 30852 34496 30932 34524
rect 23676 34428 28672 34456
rect 29917 34459 29975 34465
rect 23676 34400 23704 34428
rect 29917 34425 29929 34459
rect 29963 34456 29975 34459
rect 30374 34456 30380 34468
rect 29963 34428 30380 34456
rect 29963 34425 29975 34428
rect 29917 34419 29975 34425
rect 30374 34416 30380 34428
rect 30432 34416 30438 34468
rect 30484 34456 30512 34496
rect 30926 34484 30932 34496
rect 30984 34484 30990 34536
rect 31036 34456 31064 34564
rect 31478 34484 31484 34536
rect 31536 34524 31542 34536
rect 31573 34527 31631 34533
rect 31573 34524 31585 34527
rect 31536 34496 31585 34524
rect 31536 34484 31542 34496
rect 31573 34493 31585 34496
rect 31619 34524 31631 34527
rect 41386 34524 41414 34564
rect 43898 34552 43904 34564
rect 43956 34552 43962 34604
rect 52181 34595 52239 34601
rect 52181 34561 52193 34595
rect 52227 34592 52239 34595
rect 53466 34592 53472 34604
rect 52227 34564 53052 34592
rect 53427 34564 53472 34592
rect 52227 34561 52239 34564
rect 52181 34555 52239 34561
rect 53024 34536 53052 34564
rect 53466 34552 53472 34564
rect 53524 34552 53530 34604
rect 53760 34601 53788 34700
rect 53745 34595 53803 34601
rect 53745 34561 53757 34595
rect 53791 34561 53803 34595
rect 53745 34555 53803 34561
rect 53006 34524 53012 34536
rect 31619 34496 41414 34524
rect 52967 34496 53012 34524
rect 31619 34493 31631 34496
rect 31573 34487 31631 34493
rect 53006 34484 53012 34496
rect 53064 34484 53070 34536
rect 30484 34428 31064 34456
rect 31110 34416 31116 34468
rect 31168 34456 31174 34468
rect 32861 34459 32919 34465
rect 32861 34456 32873 34459
rect 31168 34428 32873 34456
rect 31168 34416 31174 34428
rect 32861 34425 32873 34428
rect 32907 34425 32919 34459
rect 32861 34419 32919 34425
rect 52365 34459 52423 34465
rect 52365 34425 52377 34459
rect 52411 34456 52423 34459
rect 53650 34456 53656 34468
rect 52411 34428 53656 34456
rect 52411 34425 52423 34428
rect 52365 34419 52423 34425
rect 53650 34416 53656 34428
rect 53708 34416 53714 34468
rect 22465 34391 22523 34397
rect 22465 34357 22477 34391
rect 22511 34388 22523 34391
rect 22830 34388 22836 34400
rect 22511 34360 22836 34388
rect 22511 34357 22523 34360
rect 22465 34351 22523 34357
rect 22830 34348 22836 34360
rect 22888 34388 22894 34400
rect 23658 34388 23664 34400
rect 22888 34360 23664 34388
rect 22888 34348 22894 34360
rect 23658 34348 23664 34360
rect 23716 34348 23722 34400
rect 24210 34348 24216 34400
rect 24268 34388 24274 34400
rect 26329 34391 26387 34397
rect 26329 34388 26341 34391
rect 24268 34360 26341 34388
rect 24268 34348 24274 34360
rect 26329 34357 26341 34360
rect 26375 34388 26387 34391
rect 26418 34388 26424 34400
rect 26375 34360 26424 34388
rect 26375 34357 26387 34360
rect 26329 34351 26387 34357
rect 26418 34348 26424 34360
rect 26476 34348 26482 34400
rect 28813 34391 28871 34397
rect 28813 34357 28825 34391
rect 28859 34388 28871 34391
rect 29086 34388 29092 34400
rect 28859 34360 29092 34388
rect 28859 34357 28871 34360
rect 28813 34351 28871 34357
rect 29086 34348 29092 34360
rect 29144 34348 29150 34400
rect 30926 34348 30932 34400
rect 30984 34388 30990 34400
rect 30984 34360 31029 34388
rect 30984 34348 30990 34360
rect 1104 34298 54832 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 54832 34298
rect 1104 34224 54832 34246
rect 14734 34184 14740 34196
rect 14695 34156 14740 34184
rect 14734 34144 14740 34156
rect 14792 34144 14798 34196
rect 22002 34144 22008 34196
rect 22060 34184 22066 34196
rect 22281 34187 22339 34193
rect 22281 34184 22293 34187
rect 22060 34156 22293 34184
rect 22060 34144 22066 34156
rect 22281 34153 22293 34156
rect 22327 34153 22339 34187
rect 22830 34184 22836 34196
rect 22791 34156 22836 34184
rect 22281 34147 22339 34153
rect 22296 34116 22324 34147
rect 22830 34144 22836 34156
rect 22888 34144 22894 34196
rect 23474 34184 23480 34196
rect 23435 34156 23480 34184
rect 23474 34144 23480 34156
rect 23532 34144 23538 34196
rect 24029 34187 24087 34193
rect 24029 34153 24041 34187
rect 24075 34184 24087 34187
rect 24210 34184 24216 34196
rect 24075 34156 24216 34184
rect 24075 34153 24087 34156
rect 24029 34147 24087 34153
rect 24210 34144 24216 34156
rect 24268 34144 24274 34196
rect 24670 34144 24676 34196
rect 24728 34184 24734 34196
rect 24765 34187 24823 34193
rect 24765 34184 24777 34187
rect 24728 34156 24777 34184
rect 24728 34144 24734 34156
rect 24765 34153 24777 34156
rect 24811 34153 24823 34187
rect 24765 34147 24823 34153
rect 25777 34187 25835 34193
rect 25777 34153 25789 34187
rect 25823 34184 25835 34187
rect 26694 34184 26700 34196
rect 25823 34156 26700 34184
rect 25823 34153 25835 34156
rect 25777 34147 25835 34153
rect 26694 34144 26700 34156
rect 26752 34144 26758 34196
rect 28258 34144 28264 34196
rect 28316 34184 28322 34196
rect 31202 34184 31208 34196
rect 28316 34156 31208 34184
rect 28316 34144 28322 34156
rect 31202 34144 31208 34156
rect 31260 34144 31266 34196
rect 31294 34144 31300 34196
rect 31352 34184 31358 34196
rect 31389 34187 31447 34193
rect 31389 34184 31401 34187
rect 31352 34156 31401 34184
rect 31352 34144 31358 34156
rect 31389 34153 31401 34156
rect 31435 34153 31447 34187
rect 31389 34147 31447 34153
rect 32033 34187 32091 34193
rect 32033 34153 32045 34187
rect 32079 34184 32091 34187
rect 32306 34184 32312 34196
rect 32079 34156 32312 34184
rect 32079 34153 32091 34156
rect 32033 34147 32091 34153
rect 32306 34144 32312 34156
rect 32364 34144 32370 34196
rect 23842 34116 23848 34128
rect 22296 34088 23848 34116
rect 23842 34076 23848 34088
rect 23900 34076 23906 34128
rect 26050 34076 26056 34128
rect 26108 34116 26114 34128
rect 26237 34119 26295 34125
rect 26237 34116 26249 34119
rect 26108 34088 26249 34116
rect 26108 34076 26114 34088
rect 26237 34085 26249 34088
rect 26283 34116 26295 34119
rect 28074 34116 28080 34128
rect 26283 34088 28080 34116
rect 26283 34085 26295 34088
rect 26237 34079 26295 34085
rect 28074 34076 28080 34088
rect 28132 34116 28138 34128
rect 28350 34116 28356 34128
rect 28132 34088 28356 34116
rect 28132 34076 28138 34088
rect 28350 34076 28356 34088
rect 28408 34076 28414 34128
rect 29546 34076 29552 34128
rect 29604 34116 29610 34128
rect 30282 34116 30288 34128
rect 29604 34088 30288 34116
rect 29604 34076 29610 34088
rect 30282 34076 30288 34088
rect 30340 34076 30346 34128
rect 30837 34119 30895 34125
rect 30837 34085 30849 34119
rect 30883 34116 30895 34119
rect 31754 34116 31760 34128
rect 30883 34088 31760 34116
rect 30883 34085 30895 34088
rect 30837 34079 30895 34085
rect 2133 34051 2191 34057
rect 2133 34017 2145 34051
rect 2179 34048 2191 34051
rect 22646 34048 22652 34060
rect 2179 34020 22652 34048
rect 2179 34017 2191 34020
rect 2133 34011 2191 34017
rect 22646 34008 22652 34020
rect 22704 34008 22710 34060
rect 26326 34008 26332 34060
rect 26384 34048 26390 34060
rect 26605 34051 26663 34057
rect 26605 34048 26617 34051
rect 26384 34020 26617 34048
rect 26384 34008 26390 34020
rect 26605 34017 26617 34020
rect 26651 34017 26663 34051
rect 26605 34011 26663 34017
rect 26970 34008 26976 34060
rect 27028 34048 27034 34060
rect 28169 34051 28227 34057
rect 28169 34048 28181 34051
rect 27028 34020 28181 34048
rect 27028 34008 27034 34020
rect 28169 34017 28181 34020
rect 28215 34048 28227 34051
rect 28905 34051 28963 34057
rect 28905 34048 28917 34051
rect 28215 34020 28917 34048
rect 28215 34017 28227 34020
rect 28169 34011 28227 34017
rect 28905 34017 28917 34020
rect 28951 34048 28963 34051
rect 29454 34048 29460 34060
rect 28951 34020 29460 34048
rect 28951 34017 28963 34020
rect 28905 34011 28963 34017
rect 29454 34008 29460 34020
rect 29512 34008 29518 34060
rect 30650 34048 30656 34060
rect 30024 34020 30656 34048
rect 2409 33983 2467 33989
rect 2409 33949 2421 33983
rect 2455 33980 2467 33983
rect 2774 33980 2780 33992
rect 2455 33952 2780 33980
rect 2455 33949 2467 33952
rect 2409 33943 2467 33949
rect 2774 33940 2780 33952
rect 2832 33980 2838 33992
rect 2869 33983 2927 33989
rect 2869 33980 2881 33983
rect 2832 33952 2881 33980
rect 2832 33940 2838 33952
rect 2869 33949 2881 33952
rect 2915 33949 2927 33983
rect 25314 33980 25320 33992
rect 25275 33952 25320 33980
rect 2869 33943 2927 33949
rect 25314 33940 25320 33952
rect 25372 33940 25378 33992
rect 25593 33983 25651 33989
rect 25593 33949 25605 33983
rect 25639 33980 25651 33983
rect 26344 33980 26372 34008
rect 25639 33952 26372 33980
rect 25639 33949 25651 33952
rect 25593 33943 25651 33949
rect 26510 33940 26516 33992
rect 26568 33980 26574 33992
rect 26881 33983 26939 33989
rect 26881 33980 26893 33983
rect 26568 33952 26893 33980
rect 26568 33940 26574 33952
rect 26881 33949 26893 33952
rect 26927 33980 26939 33983
rect 27062 33980 27068 33992
rect 26927 33952 27068 33980
rect 26927 33949 26939 33952
rect 26881 33943 26939 33949
rect 27062 33940 27068 33952
rect 27120 33940 27126 33992
rect 27338 33980 27344 33992
rect 27299 33952 27344 33980
rect 27338 33940 27344 33952
rect 27396 33940 27402 33992
rect 27525 33983 27583 33989
rect 27525 33949 27537 33983
rect 27571 33949 27583 33983
rect 27982 33980 27988 33992
rect 27943 33952 27988 33980
rect 27525 33943 27583 33949
rect 26396 33915 26454 33921
rect 26396 33881 26408 33915
rect 26442 33912 26454 33915
rect 26694 33912 26700 33924
rect 26442 33884 26700 33912
rect 26442 33881 26454 33884
rect 26396 33875 26454 33881
rect 26694 33872 26700 33884
rect 26752 33872 26758 33924
rect 27246 33872 27252 33924
rect 27304 33912 27310 33924
rect 27540 33912 27568 33943
rect 27982 33940 27988 33952
rect 28040 33940 28046 33992
rect 30024 33989 30052 34020
rect 30650 34008 30656 34020
rect 30708 34048 30714 34060
rect 30852 34048 30880 34079
rect 31754 34076 31760 34088
rect 31812 34076 31818 34128
rect 53374 34116 53380 34128
rect 53335 34088 53380 34116
rect 53374 34076 53380 34088
rect 53432 34076 53438 34128
rect 30708 34020 30880 34048
rect 30708 34008 30714 34020
rect 30009 33983 30067 33989
rect 30009 33949 30021 33983
rect 30055 33949 30067 33983
rect 30009 33943 30067 33949
rect 30101 33983 30159 33989
rect 30101 33949 30113 33983
rect 30147 33949 30159 33983
rect 30282 33980 30288 33992
rect 30243 33952 30288 33980
rect 30101 33943 30159 33949
rect 27304 33884 27568 33912
rect 30116 33912 30144 33943
rect 30282 33940 30288 33952
rect 30340 33940 30346 33992
rect 30374 33940 30380 33992
rect 30432 33980 30438 33992
rect 30432 33952 30477 33980
rect 30432 33940 30438 33952
rect 31202 33940 31208 33992
rect 31260 33980 31266 33992
rect 31260 33952 41414 33980
rect 31260 33940 31266 33952
rect 31754 33912 31760 33924
rect 30116 33884 31760 33912
rect 27304 33872 27310 33884
rect 31754 33872 31760 33884
rect 31812 33872 31818 33924
rect 41386 33912 41414 33952
rect 53098 33940 53104 33992
rect 53156 33980 53162 33992
rect 53509 33983 53567 33989
rect 53509 33980 53521 33983
rect 53156 33952 53521 33980
rect 53156 33940 53162 33952
rect 53509 33949 53521 33952
rect 53555 33949 53567 33983
rect 53509 33943 53567 33949
rect 53650 33940 53656 33992
rect 53708 33980 53714 33992
rect 53926 33980 53932 33992
rect 53708 33952 53753 33980
rect 53887 33952 53932 33980
rect 53708 33940 53714 33952
rect 53926 33940 53932 33952
rect 53984 33940 53990 33992
rect 52733 33915 52791 33921
rect 52733 33912 52745 33915
rect 41386 33884 52745 33912
rect 52733 33881 52745 33884
rect 52779 33881 52791 33915
rect 52733 33875 52791 33881
rect 53745 33915 53803 33921
rect 53745 33881 53757 33915
rect 53791 33881 53803 33915
rect 53745 33875 53803 33881
rect 24946 33804 24952 33856
rect 25004 33844 25010 33856
rect 25409 33847 25467 33853
rect 25409 33844 25421 33847
rect 25004 33816 25421 33844
rect 25004 33804 25010 33816
rect 25409 33813 25421 33816
rect 25455 33844 25467 33847
rect 25866 33844 25872 33856
rect 25455 33816 25872 33844
rect 25455 33813 25467 33816
rect 25409 33807 25467 33813
rect 25866 33804 25872 33816
rect 25924 33804 25930 33856
rect 26513 33847 26571 33853
rect 26513 33813 26525 33847
rect 26559 33844 26571 33847
rect 26878 33844 26884 33856
rect 26559 33816 26884 33844
rect 26559 33813 26571 33816
rect 26513 33807 26571 33813
rect 26878 33804 26884 33816
rect 26936 33804 26942 33856
rect 27433 33847 27491 33853
rect 27433 33813 27445 33847
rect 27479 33844 27491 33847
rect 28442 33844 28448 33856
rect 27479 33816 28448 33844
rect 27479 33813 27491 33816
rect 27433 33807 27491 33813
rect 28442 33804 28448 33816
rect 28500 33804 28506 33856
rect 29825 33847 29883 33853
rect 29825 33813 29837 33847
rect 29871 33844 29883 33847
rect 30558 33844 30564 33856
rect 29871 33816 30564 33844
rect 29871 33813 29883 33816
rect 29825 33807 29883 33813
rect 30558 33804 30564 33816
rect 30616 33804 30622 33856
rect 52748 33844 52776 33875
rect 53760 33844 53788 33875
rect 52748 33816 53788 33844
rect 1104 33754 54832 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 54832 33754
rect 1104 33680 54832 33702
rect 23106 33600 23112 33652
rect 23164 33640 23170 33652
rect 24026 33640 24032 33652
rect 23164 33612 24032 33640
rect 23164 33600 23170 33612
rect 23860 33581 23888 33612
rect 24026 33600 24032 33612
rect 24084 33600 24090 33652
rect 24210 33640 24216 33652
rect 24171 33612 24216 33640
rect 24210 33600 24216 33612
rect 24268 33600 24274 33652
rect 24762 33600 24768 33652
rect 24820 33640 24826 33652
rect 26970 33640 26976 33652
rect 24820 33612 26976 33640
rect 24820 33600 24826 33612
rect 26970 33600 26976 33612
rect 27028 33600 27034 33652
rect 27062 33600 27068 33652
rect 27120 33640 27126 33652
rect 27433 33643 27491 33649
rect 27433 33640 27445 33643
rect 27120 33612 27445 33640
rect 27120 33600 27126 33612
rect 27433 33609 27445 33612
rect 27479 33609 27491 33643
rect 27433 33603 27491 33609
rect 27801 33643 27859 33649
rect 27801 33609 27813 33643
rect 27847 33640 27859 33643
rect 28258 33640 28264 33652
rect 27847 33612 28264 33640
rect 27847 33609 27859 33612
rect 27801 33603 27859 33609
rect 28258 33600 28264 33612
rect 28316 33600 28322 33652
rect 51258 33600 51264 33652
rect 51316 33640 51322 33652
rect 53098 33640 53104 33652
rect 51316 33612 53104 33640
rect 51316 33600 51322 33612
rect 53098 33600 53104 33612
rect 53156 33600 53162 33652
rect 23845 33575 23903 33581
rect 23845 33541 23857 33575
rect 23891 33541 23903 33575
rect 26510 33572 26516 33584
rect 23845 33535 23903 33541
rect 24688 33544 26516 33572
rect 6730 33464 6736 33516
rect 6788 33504 6794 33516
rect 23474 33504 23480 33516
rect 6788 33476 23480 33504
rect 6788 33464 6794 33476
rect 23474 33464 23480 33476
rect 23532 33504 23538 33516
rect 24688 33513 24716 33544
rect 26510 33532 26516 33544
rect 26568 33532 26574 33584
rect 26694 33532 26700 33584
rect 26752 33572 26758 33584
rect 27341 33575 27399 33581
rect 27341 33572 27353 33575
rect 26752 33544 27353 33572
rect 26752 33532 26758 33544
rect 27341 33541 27353 33544
rect 27387 33541 27399 33575
rect 27341 33535 27399 33541
rect 23661 33507 23719 33513
rect 23661 33504 23673 33507
rect 23532 33476 23673 33504
rect 23532 33464 23538 33476
rect 23661 33473 23673 33476
rect 23707 33473 23719 33507
rect 23661 33467 23719 33473
rect 23937 33507 23995 33513
rect 23937 33473 23949 33507
rect 23983 33473 23995 33507
rect 23937 33467 23995 33473
rect 24029 33507 24087 33513
rect 24029 33473 24041 33507
rect 24075 33473 24087 33507
rect 24029 33467 24087 33473
rect 24673 33507 24731 33513
rect 24673 33473 24685 33507
rect 24719 33473 24731 33507
rect 24946 33504 24952 33516
rect 24907 33476 24952 33504
rect 24673 33467 24731 33473
rect 2133 33439 2191 33445
rect 2133 33405 2145 33439
rect 2179 33405 2191 33439
rect 2133 33399 2191 33405
rect 2409 33439 2467 33445
rect 2409 33405 2421 33439
rect 2455 33436 2467 33439
rect 2774 33436 2780 33448
rect 2455 33408 2780 33436
rect 2455 33405 2467 33408
rect 2409 33399 2467 33405
rect 2148 33368 2176 33399
rect 2774 33396 2780 33408
rect 2832 33436 2838 33448
rect 2869 33439 2927 33445
rect 2869 33436 2881 33439
rect 2832 33408 2881 33436
rect 2832 33396 2838 33408
rect 2869 33405 2881 33408
rect 2915 33405 2927 33439
rect 23952 33436 23980 33467
rect 2869 33399 2927 33405
rect 23124 33408 23980 33436
rect 13538 33368 13544 33380
rect 2148 33340 13544 33368
rect 13538 33328 13544 33340
rect 13596 33328 13602 33380
rect 15102 33260 15108 33312
rect 15160 33300 15166 33312
rect 23124 33309 23152 33408
rect 24044 33368 24072 33467
rect 24946 33464 24952 33476
rect 25004 33464 25010 33516
rect 25406 33464 25412 33516
rect 25464 33504 25470 33516
rect 25593 33507 25651 33513
rect 25593 33504 25605 33507
rect 25464 33476 25605 33504
rect 25464 33464 25470 33476
rect 25593 33473 25605 33476
rect 25639 33473 25651 33507
rect 25593 33467 25651 33473
rect 25777 33507 25835 33513
rect 25777 33473 25789 33507
rect 25823 33504 25835 33507
rect 26234 33504 26240 33516
rect 25823 33476 26240 33504
rect 25823 33473 25835 33476
rect 25777 33467 25835 33473
rect 26234 33464 26240 33476
rect 26292 33464 26298 33516
rect 26329 33507 26387 33513
rect 26329 33473 26341 33507
rect 26375 33473 26387 33507
rect 26329 33467 26387 33473
rect 25130 33396 25136 33448
rect 25188 33436 25194 33448
rect 25501 33439 25559 33445
rect 25501 33436 25513 33439
rect 25188 33408 25513 33436
rect 25188 33396 25194 33408
rect 25501 33405 25513 33408
rect 25547 33405 25559 33439
rect 25501 33399 25559 33405
rect 25866 33396 25872 33448
rect 25924 33436 25930 33448
rect 26344 33436 26372 33467
rect 26418 33464 26424 33516
rect 26476 33504 26482 33516
rect 27249 33507 27307 33513
rect 27249 33504 27261 33507
rect 26476 33476 27261 33504
rect 26476 33464 26482 33476
rect 27249 33473 27261 33476
rect 27295 33473 27307 33507
rect 29086 33504 29092 33516
rect 29047 33476 29092 33504
rect 27249 33467 27307 33473
rect 29086 33464 29092 33476
rect 29144 33464 29150 33516
rect 29730 33504 29736 33516
rect 29691 33476 29736 33504
rect 29730 33464 29736 33476
rect 29788 33464 29794 33516
rect 27338 33436 27344 33448
rect 25924 33408 27344 33436
rect 25924 33396 25930 33408
rect 27338 33396 27344 33408
rect 27396 33396 27402 33448
rect 27985 33439 28043 33445
rect 27985 33405 27997 33439
rect 28031 33405 28043 33439
rect 27985 33399 28043 33405
rect 29365 33439 29423 33445
rect 29365 33405 29377 33439
rect 29411 33405 29423 33439
rect 29365 33399 29423 33405
rect 24578 33368 24584 33380
rect 24044 33340 24584 33368
rect 24578 33328 24584 33340
rect 24636 33368 24642 33380
rect 24673 33371 24731 33377
rect 24673 33368 24685 33371
rect 24636 33340 24685 33368
rect 24636 33328 24642 33340
rect 24673 33337 24685 33340
rect 24719 33337 24731 33371
rect 24673 33331 24731 33337
rect 24765 33371 24823 33377
rect 24765 33337 24777 33371
rect 24811 33368 24823 33371
rect 25314 33368 25320 33380
rect 24811 33340 25320 33368
rect 24811 33337 24823 33340
rect 24765 33331 24823 33337
rect 25314 33328 25320 33340
rect 25372 33328 25378 33380
rect 26878 33328 26884 33380
rect 26936 33368 26942 33380
rect 28000 33368 28028 33399
rect 26936 33340 28028 33368
rect 26936 33328 26942 33340
rect 28994 33328 29000 33380
rect 29052 33368 29058 33380
rect 29380 33368 29408 33399
rect 29454 33396 29460 33448
rect 29512 33436 29518 33448
rect 29641 33439 29699 33445
rect 29641 33436 29653 33439
rect 29512 33408 29653 33436
rect 29512 33396 29518 33408
rect 29641 33405 29653 33408
rect 29687 33405 29699 33439
rect 30561 33439 30619 33445
rect 30561 33436 30573 33439
rect 29641 33399 29699 33405
rect 29748 33408 30573 33436
rect 29748 33368 29776 33408
rect 30561 33405 30573 33408
rect 30607 33436 30619 33439
rect 30607 33408 31754 33436
rect 30607 33405 30619 33408
rect 30561 33399 30619 33405
rect 29052 33340 29776 33368
rect 30101 33371 30159 33377
rect 29052 33328 29058 33340
rect 30101 33337 30113 33371
rect 30147 33368 30159 33371
rect 30650 33368 30656 33380
rect 30147 33340 30656 33368
rect 30147 33337 30159 33340
rect 30101 33331 30159 33337
rect 30650 33328 30656 33340
rect 30708 33328 30714 33380
rect 31726 33368 31754 33408
rect 53374 33368 53380 33380
rect 31726 33340 53380 33368
rect 53374 33328 53380 33340
rect 53432 33328 53438 33380
rect 23109 33303 23167 33309
rect 23109 33300 23121 33303
rect 15160 33272 23121 33300
rect 15160 33260 15166 33272
rect 23109 33269 23121 33272
rect 23155 33269 23167 33303
rect 23109 33263 23167 33269
rect 31205 33303 31263 33309
rect 31205 33269 31217 33303
rect 31251 33300 31263 33303
rect 31754 33300 31760 33312
rect 31251 33272 31760 33300
rect 31251 33269 31263 33272
rect 31205 33263 31263 33269
rect 31754 33260 31760 33272
rect 31812 33260 31818 33312
rect 54294 33300 54300 33312
rect 54255 33272 54300 33300
rect 54294 33260 54300 33272
rect 54352 33260 54358 33312
rect 1104 33210 54832 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 54832 33210
rect 1104 33136 54832 33158
rect 23385 33099 23443 33105
rect 23385 33065 23397 33099
rect 23431 33096 23443 33099
rect 23474 33096 23480 33108
rect 23431 33068 23480 33096
rect 23431 33065 23443 33068
rect 23385 33059 23443 33065
rect 23474 33056 23480 33068
rect 23532 33056 23538 33108
rect 25593 33099 25651 33105
rect 25593 33065 25605 33099
rect 25639 33096 25651 33099
rect 25774 33096 25780 33108
rect 25639 33068 25780 33096
rect 25639 33065 25651 33068
rect 25593 33059 25651 33065
rect 25774 33056 25780 33068
rect 25832 33056 25838 33108
rect 26053 33099 26111 33105
rect 26053 33065 26065 33099
rect 26099 33096 26111 33099
rect 26142 33096 26148 33108
rect 26099 33068 26148 33096
rect 26099 33065 26111 33068
rect 26053 33059 26111 33065
rect 26142 33056 26148 33068
rect 26200 33056 26206 33108
rect 27893 33099 27951 33105
rect 27893 33065 27905 33099
rect 27939 33096 27951 33099
rect 27982 33096 27988 33108
rect 27939 33068 27988 33096
rect 27939 33065 27951 33068
rect 27893 33059 27951 33065
rect 27982 33056 27988 33068
rect 28040 33056 28046 33108
rect 28994 33096 29000 33108
rect 28955 33068 29000 33096
rect 28994 33056 29000 33068
rect 29052 33056 29058 33108
rect 26694 32988 26700 33040
rect 26752 33028 26758 33040
rect 26789 33031 26847 33037
rect 26789 33028 26801 33031
rect 26752 33000 26801 33028
rect 26752 32988 26758 33000
rect 26789 32997 26801 33000
rect 26835 32997 26847 33031
rect 26789 32991 26847 32997
rect 25314 32960 25320 32972
rect 25227 32932 25320 32960
rect 25314 32920 25320 32932
rect 25372 32960 25378 32972
rect 26418 32960 26424 32972
rect 25372 32932 26424 32960
rect 25372 32920 25378 32932
rect 26418 32920 26424 32932
rect 26476 32920 26482 32972
rect 27433 32963 27491 32969
rect 27433 32929 27445 32963
rect 27479 32960 27491 32963
rect 27614 32960 27620 32972
rect 27479 32932 27620 32960
rect 27479 32929 27491 32932
rect 27433 32923 27491 32929
rect 27614 32920 27620 32932
rect 27672 32960 27678 32972
rect 29012 32960 29040 33056
rect 27672 32932 28212 32960
rect 27672 32920 27678 32932
rect 1578 32892 1584 32904
rect 1539 32864 1584 32892
rect 1578 32852 1584 32864
rect 1636 32892 1642 32904
rect 2777 32895 2835 32901
rect 2777 32892 2789 32895
rect 1636 32864 2789 32892
rect 1636 32852 1642 32864
rect 2777 32861 2789 32864
rect 2823 32861 2835 32895
rect 2777 32855 2835 32861
rect 25225 32895 25283 32901
rect 25225 32861 25237 32895
rect 25271 32861 25283 32895
rect 25225 32855 25283 32861
rect 25409 32895 25467 32901
rect 25409 32861 25421 32895
rect 25455 32892 25467 32895
rect 26234 32892 26240 32904
rect 25455 32864 26240 32892
rect 25455 32861 25467 32864
rect 25409 32855 25467 32861
rect 15102 32824 15108 32836
rect 1780 32796 15108 32824
rect 1780 32765 1808 32796
rect 15102 32784 15108 32796
rect 15160 32784 15166 32836
rect 25240 32824 25268 32855
rect 26234 32852 26240 32864
rect 26292 32852 26298 32904
rect 26878 32892 26884 32904
rect 26712 32864 26884 32892
rect 26712 32824 26740 32864
rect 26878 32852 26884 32864
rect 26936 32892 26942 32904
rect 27338 32892 27344 32904
rect 26936 32864 27344 32892
rect 26936 32852 26942 32864
rect 27338 32852 27344 32864
rect 27396 32852 27402 32904
rect 28074 32892 28080 32904
rect 28035 32864 28080 32892
rect 28074 32852 28080 32864
rect 28132 32852 28138 32904
rect 28184 32901 28212 32932
rect 28368 32932 29040 32960
rect 28368 32901 28396 32932
rect 28169 32895 28227 32901
rect 28169 32861 28181 32895
rect 28215 32861 28227 32895
rect 28169 32855 28227 32861
rect 28353 32895 28411 32901
rect 28353 32861 28365 32895
rect 28399 32861 28411 32895
rect 28353 32855 28411 32861
rect 28442 32852 28448 32904
rect 28500 32892 28506 32904
rect 54294 32892 54300 32904
rect 28500 32864 28545 32892
rect 54255 32864 54300 32892
rect 28500 32852 28506 32864
rect 54294 32852 54300 32864
rect 54352 32852 54358 32904
rect 25240 32796 26740 32824
rect 26789 32827 26847 32833
rect 1765 32759 1823 32765
rect 1765 32725 1777 32759
rect 1811 32725 1823 32759
rect 1765 32719 1823 32725
rect 2317 32759 2375 32765
rect 2317 32725 2329 32759
rect 2363 32756 2375 32759
rect 2774 32756 2780 32768
rect 2363 32728 2780 32756
rect 2363 32725 2375 32728
rect 2317 32719 2375 32725
rect 2774 32716 2780 32728
rect 2832 32716 2838 32768
rect 24026 32716 24032 32768
rect 24084 32756 24090 32768
rect 26252 32765 26280 32796
rect 26789 32793 26801 32827
rect 26835 32824 26847 32827
rect 27062 32824 27068 32836
rect 26835 32796 27068 32824
rect 26835 32793 26847 32796
rect 26789 32787 26847 32793
rect 27062 32784 27068 32796
rect 27120 32784 27126 32836
rect 24581 32759 24639 32765
rect 24581 32756 24593 32759
rect 24084 32728 24593 32756
rect 24084 32716 24090 32728
rect 24581 32725 24593 32728
rect 24627 32725 24639 32759
rect 24581 32719 24639 32725
rect 26237 32759 26295 32765
rect 26237 32725 26249 32759
rect 26283 32725 26295 32759
rect 26237 32719 26295 32725
rect 26326 32716 26332 32768
rect 26384 32756 26390 32768
rect 29825 32759 29883 32765
rect 26384 32728 26429 32756
rect 26384 32716 26390 32728
rect 29825 32725 29837 32759
rect 29871 32756 29883 32759
rect 29914 32756 29920 32768
rect 29871 32728 29920 32756
rect 29871 32725 29883 32728
rect 29825 32719 29883 32725
rect 29914 32716 29920 32728
rect 29972 32716 29978 32768
rect 1104 32666 54832 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 54832 32666
rect 1104 32592 54832 32614
rect 24026 32512 24032 32564
rect 24084 32552 24090 32564
rect 24854 32552 24860 32564
rect 24084 32524 24860 32552
rect 24084 32512 24090 32524
rect 24854 32512 24860 32524
rect 24912 32552 24918 32564
rect 25593 32555 25651 32561
rect 25593 32552 25605 32555
rect 24912 32524 25605 32552
rect 24912 32512 24918 32524
rect 25593 32521 25605 32524
rect 25639 32521 25651 32555
rect 25593 32515 25651 32521
rect 27249 32555 27307 32561
rect 27249 32521 27261 32555
rect 27295 32552 27307 32555
rect 29730 32552 29736 32564
rect 27295 32524 29736 32552
rect 27295 32521 27307 32524
rect 27249 32515 27307 32521
rect 29730 32512 29736 32524
rect 29788 32512 29794 32564
rect 24578 32484 24584 32496
rect 24539 32456 24584 32484
rect 24578 32444 24584 32456
rect 24636 32444 24642 32496
rect 26510 32444 26516 32496
rect 26568 32484 26574 32496
rect 26878 32484 26884 32496
rect 26568 32456 26884 32484
rect 26568 32444 26574 32456
rect 26878 32444 26884 32456
rect 26936 32484 26942 32496
rect 26936 32456 27384 32484
rect 26936 32444 26942 32456
rect 25777 32419 25835 32425
rect 25777 32385 25789 32419
rect 25823 32416 25835 32419
rect 25866 32416 25872 32428
rect 25823 32388 25872 32416
rect 25823 32385 25835 32388
rect 25777 32379 25835 32385
rect 25866 32376 25872 32388
rect 25924 32376 25930 32428
rect 26234 32376 26240 32428
rect 26292 32416 26298 32428
rect 26329 32419 26387 32425
rect 26329 32416 26341 32419
rect 26292 32388 26341 32416
rect 26292 32376 26298 32388
rect 26329 32385 26341 32388
rect 26375 32416 26387 32419
rect 26970 32416 26976 32428
rect 26375 32388 26976 32416
rect 26375 32385 26387 32388
rect 26329 32379 26387 32385
rect 26970 32376 26976 32388
rect 27028 32376 27034 32428
rect 27356 32425 27384 32456
rect 27614 32444 27620 32496
rect 27672 32484 27678 32496
rect 28353 32487 28411 32493
rect 28353 32484 28365 32487
rect 27672 32456 28365 32484
rect 27672 32444 27678 32456
rect 28353 32453 28365 32456
rect 28399 32453 28411 32487
rect 28353 32447 28411 32453
rect 27157 32419 27215 32425
rect 27157 32385 27169 32419
rect 27203 32385 27215 32419
rect 27157 32379 27215 32385
rect 27341 32419 27399 32425
rect 27341 32385 27353 32419
rect 27387 32385 27399 32419
rect 27341 32379 27399 32385
rect 2133 32351 2191 32357
rect 2133 32317 2145 32351
rect 2179 32317 2191 32351
rect 2133 32311 2191 32317
rect 2409 32351 2467 32357
rect 2409 32317 2421 32351
rect 2455 32348 2467 32351
rect 2774 32348 2780 32360
rect 2455 32320 2780 32348
rect 2455 32317 2467 32320
rect 2409 32311 2467 32317
rect 2148 32280 2176 32311
rect 2774 32308 2780 32320
rect 2832 32308 2838 32360
rect 26418 32348 26424 32360
rect 26379 32320 26424 32348
rect 26418 32308 26424 32320
rect 26476 32348 26482 32360
rect 27172 32348 27200 32379
rect 32582 32376 32588 32428
rect 32640 32416 32646 32428
rect 47854 32416 47860 32428
rect 32640 32388 47860 32416
rect 32640 32376 32646 32388
rect 47854 32376 47860 32388
rect 47912 32376 47918 32428
rect 26476 32320 27200 32348
rect 26476 32308 26482 32320
rect 24946 32280 24952 32292
rect 2148 32252 24952 32280
rect 24946 32240 24952 32252
rect 25004 32240 25010 32292
rect 27430 32240 27436 32292
rect 27488 32280 27494 32292
rect 27801 32283 27859 32289
rect 27801 32280 27813 32283
rect 27488 32252 27813 32280
rect 27488 32240 27494 32252
rect 27801 32249 27813 32252
rect 27847 32280 27859 32283
rect 27847 32252 28994 32280
rect 27847 32249 27859 32252
rect 27801 32243 27859 32249
rect 23014 32172 23020 32224
rect 23072 32212 23078 32224
rect 24854 32212 24860 32224
rect 23072 32184 24860 32212
rect 23072 32172 23078 32184
rect 24854 32172 24860 32184
rect 24912 32172 24918 32224
rect 26970 32172 26976 32224
rect 27028 32212 27034 32224
rect 27246 32212 27252 32224
rect 27028 32184 27252 32212
rect 27028 32172 27034 32184
rect 27246 32172 27252 32184
rect 27304 32172 27310 32224
rect 28966 32212 28994 32252
rect 51166 32212 51172 32224
rect 28966 32184 51172 32212
rect 51166 32172 51172 32184
rect 51224 32172 51230 32224
rect 1104 32122 54832 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 54832 32122
rect 1104 32048 54832 32070
rect 24946 32008 24952 32020
rect 24907 31980 24952 32008
rect 24946 31968 24952 31980
rect 25004 31968 25010 32020
rect 25958 31968 25964 32020
rect 26016 32008 26022 32020
rect 26053 32011 26111 32017
rect 26053 32008 26065 32011
rect 26016 31980 26065 32008
rect 26016 31968 26022 31980
rect 26053 31977 26065 31980
rect 26099 31977 26111 32011
rect 27430 32008 27436 32020
rect 26053 31971 26111 31977
rect 26712 31980 27436 32008
rect 2130 31804 2136 31816
rect 2091 31776 2136 31804
rect 2130 31764 2136 31776
rect 2188 31764 2194 31816
rect 2409 31807 2467 31813
rect 2409 31773 2421 31807
rect 2455 31804 2467 31807
rect 2774 31804 2780 31816
rect 2455 31776 2780 31804
rect 2455 31773 2467 31776
rect 2409 31767 2467 31773
rect 2774 31764 2780 31776
rect 2832 31804 2838 31816
rect 2869 31807 2927 31813
rect 2869 31804 2881 31807
rect 2832 31776 2881 31804
rect 2832 31764 2838 31776
rect 2869 31773 2881 31776
rect 2915 31773 2927 31807
rect 26602 31804 26608 31816
rect 26563 31776 26608 31804
rect 2869 31767 2927 31773
rect 26602 31764 26608 31776
rect 26660 31764 26666 31816
rect 26712 31813 26740 31980
rect 27430 31968 27436 31980
rect 27488 31968 27494 32020
rect 27249 31943 27307 31949
rect 27249 31909 27261 31943
rect 27295 31909 27307 31943
rect 27249 31903 27307 31909
rect 26698 31807 26756 31813
rect 26698 31773 26710 31807
rect 26744 31773 26756 31807
rect 26970 31804 26976 31816
rect 26931 31776 26976 31804
rect 26698 31767 26756 31773
rect 26970 31764 26976 31776
rect 27028 31764 27034 31816
rect 27070 31807 27128 31813
rect 27070 31773 27082 31807
rect 27116 31773 27128 31807
rect 27264 31804 27292 31903
rect 27893 31807 27951 31813
rect 27893 31804 27905 31807
rect 27264 31776 27905 31804
rect 27070 31767 27128 31773
rect 27893 31773 27905 31776
rect 27939 31773 27951 31807
rect 54294 31804 54300 31816
rect 54255 31776 54300 31804
rect 27893 31767 27951 31773
rect 25682 31696 25688 31748
rect 25740 31736 25746 31748
rect 25958 31736 25964 31748
rect 25740 31708 25964 31736
rect 25740 31696 25746 31708
rect 25958 31696 25964 31708
rect 26016 31736 26022 31748
rect 26881 31739 26939 31745
rect 26881 31736 26893 31739
rect 26016 31708 26893 31736
rect 26016 31696 26022 31708
rect 26881 31705 26893 31708
rect 26927 31705 26939 31739
rect 26881 31699 26939 31705
rect 24854 31628 24860 31680
rect 24912 31668 24918 31680
rect 25593 31671 25651 31677
rect 25593 31668 25605 31671
rect 24912 31640 25605 31668
rect 24912 31628 24918 31640
rect 25593 31637 25605 31640
rect 25639 31668 25651 31671
rect 26142 31668 26148 31680
rect 25639 31640 26148 31668
rect 25639 31637 25651 31640
rect 25593 31631 25651 31637
rect 26142 31628 26148 31640
rect 26200 31668 26206 31680
rect 27079 31668 27107 31767
rect 54294 31764 54300 31776
rect 54352 31764 54358 31816
rect 27709 31739 27767 31745
rect 27709 31705 27721 31739
rect 27755 31736 27767 31739
rect 27798 31736 27804 31748
rect 27755 31708 27804 31736
rect 27755 31705 27767 31708
rect 27709 31699 27767 31705
rect 27798 31696 27804 31708
rect 27856 31696 27862 31748
rect 26200 31640 27107 31668
rect 28077 31671 28135 31677
rect 26200 31628 26206 31640
rect 28077 31637 28089 31671
rect 28123 31668 28135 31671
rect 28350 31668 28356 31680
rect 28123 31640 28356 31668
rect 28123 31637 28135 31640
rect 28077 31631 28135 31637
rect 28350 31628 28356 31640
rect 28408 31628 28414 31680
rect 1104 31578 54832 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 54832 31578
rect 1104 31504 54832 31526
rect 26418 31464 26424 31476
rect 26379 31436 26424 31464
rect 26418 31424 26424 31436
rect 26476 31424 26482 31476
rect 25866 31356 25872 31408
rect 25924 31396 25930 31408
rect 26326 31396 26332 31408
rect 25924 31368 26332 31396
rect 25924 31356 25930 31368
rect 26326 31356 26332 31368
rect 26384 31356 26390 31408
rect 26513 31399 26571 31405
rect 26513 31365 26525 31399
rect 26559 31396 26571 31399
rect 26602 31396 26608 31408
rect 26559 31368 26608 31396
rect 26559 31365 26571 31368
rect 26513 31359 26571 31365
rect 26602 31356 26608 31368
rect 26660 31396 26666 31408
rect 27062 31396 27068 31408
rect 26660 31368 27068 31396
rect 26660 31356 26666 31368
rect 27062 31356 27068 31368
rect 27120 31356 27126 31408
rect 2133 31331 2191 31337
rect 2133 31297 2145 31331
rect 2179 31328 2191 31331
rect 20806 31328 20812 31340
rect 2179 31300 20812 31328
rect 2179 31297 2191 31300
rect 2133 31291 2191 31297
rect 20806 31288 20812 31300
rect 20864 31288 20870 31340
rect 25498 31288 25504 31340
rect 25556 31328 25562 31340
rect 28350 31328 28356 31340
rect 25556 31300 26004 31328
rect 28311 31300 28356 31328
rect 25556 31288 25562 31300
rect 2409 31263 2467 31269
rect 2409 31229 2421 31263
rect 2455 31260 2467 31263
rect 2774 31260 2780 31272
rect 2455 31232 2780 31260
rect 2455 31229 2467 31232
rect 2409 31223 2467 31229
rect 2774 31220 2780 31232
rect 2832 31260 2838 31272
rect 2869 31263 2927 31269
rect 2869 31260 2881 31263
rect 2832 31232 2881 31260
rect 2832 31220 2838 31232
rect 2869 31229 2881 31232
rect 2915 31229 2927 31263
rect 25774 31260 25780 31272
rect 25735 31232 25780 31260
rect 2869 31223 2927 31229
rect 25774 31220 25780 31232
rect 25832 31220 25838 31272
rect 25976 31269 26004 31300
rect 28350 31288 28356 31300
rect 28408 31288 28414 31340
rect 25961 31263 26019 31269
rect 25961 31229 25973 31263
rect 26007 31260 26019 31263
rect 26050 31260 26056 31272
rect 26007 31232 26056 31260
rect 26007 31229 26019 31232
rect 25961 31223 26019 31229
rect 26050 31220 26056 31232
rect 26108 31220 26114 31272
rect 27982 31220 27988 31272
rect 28040 31260 28046 31272
rect 28077 31263 28135 31269
rect 28077 31260 28089 31263
rect 28040 31232 28089 31260
rect 28040 31220 28046 31232
rect 28077 31229 28089 31232
rect 28123 31229 28135 31263
rect 28077 31223 28135 31229
rect 33778 31152 33784 31204
rect 33836 31192 33842 31204
rect 49326 31192 49332 31204
rect 33836 31164 49332 31192
rect 33836 31152 33842 31164
rect 49326 31152 49332 31164
rect 49384 31152 49390 31204
rect 30374 31084 30380 31136
rect 30432 31124 30438 31136
rect 52822 31124 52828 31136
rect 30432 31096 52828 31124
rect 30432 31084 30438 31096
rect 52822 31084 52828 31096
rect 52880 31084 52886 31136
rect 54294 31124 54300 31136
rect 54255 31096 54300 31124
rect 54294 31084 54300 31096
rect 54352 31084 54358 31136
rect 1104 31034 54832 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 54832 31034
rect 1104 30960 54832 30982
rect 27249 30923 27307 30929
rect 27249 30889 27261 30923
rect 27295 30920 27307 30923
rect 27706 30920 27712 30932
rect 27295 30892 27712 30920
rect 27295 30889 27307 30892
rect 27249 30883 27307 30889
rect 27706 30880 27712 30892
rect 27764 30880 27770 30932
rect 30742 30880 30748 30932
rect 30800 30920 30806 30932
rect 32398 30920 32404 30932
rect 30800 30892 32404 30920
rect 30800 30880 30806 30892
rect 32398 30880 32404 30892
rect 32456 30880 32462 30932
rect 26142 30812 26148 30864
rect 26200 30852 26206 30864
rect 26200 30824 27016 30852
rect 26200 30812 26206 30824
rect 2133 30787 2191 30793
rect 2133 30753 2145 30787
rect 2179 30784 2191 30787
rect 17862 30784 17868 30796
rect 2179 30756 17868 30784
rect 2179 30753 2191 30756
rect 2133 30747 2191 30753
rect 17862 30744 17868 30756
rect 17920 30744 17926 30796
rect 26050 30744 26056 30796
rect 26108 30784 26114 30796
rect 26108 30756 26924 30784
rect 26108 30744 26114 30756
rect 2409 30719 2467 30725
rect 2409 30685 2421 30719
rect 2455 30716 2467 30719
rect 2774 30716 2780 30728
rect 2455 30688 2780 30716
rect 2455 30685 2467 30688
rect 2409 30679 2467 30685
rect 2774 30676 2780 30688
rect 2832 30716 2838 30728
rect 26896 30725 26924 30756
rect 2869 30719 2927 30725
rect 2869 30716 2881 30719
rect 2832 30688 2881 30716
rect 2832 30676 2838 30688
rect 2869 30685 2881 30688
rect 2915 30685 2927 30719
rect 2869 30679 2927 30685
rect 26697 30719 26755 30725
rect 26697 30685 26709 30719
rect 26743 30685 26755 30719
rect 26697 30679 26755 30685
rect 26881 30719 26939 30725
rect 26881 30685 26893 30719
rect 26927 30685 26939 30719
rect 26988 30716 27016 30824
rect 27065 30719 27123 30725
rect 27065 30716 27077 30719
rect 26988 30688 27077 30716
rect 26881 30679 26939 30685
rect 27065 30685 27077 30688
rect 27111 30685 27123 30719
rect 27065 30679 27123 30685
rect 26142 30580 26148 30592
rect 26103 30552 26148 30580
rect 26142 30540 26148 30552
rect 26200 30540 26206 30592
rect 26712 30580 26740 30679
rect 26970 30608 26976 30660
rect 27028 30648 27034 30660
rect 27028 30620 27073 30648
rect 27028 30608 27034 30620
rect 27801 30583 27859 30589
rect 27801 30580 27813 30583
rect 26712 30552 27813 30580
rect 27801 30549 27813 30552
rect 27847 30580 27859 30583
rect 44818 30580 44824 30592
rect 27847 30552 44824 30580
rect 27847 30549 27859 30552
rect 27801 30543 27859 30549
rect 44818 30540 44824 30552
rect 44876 30540 44882 30592
rect 1104 30490 54832 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 54832 30490
rect 1104 30416 54832 30438
rect 2130 30336 2136 30388
rect 2188 30376 2194 30388
rect 26329 30379 26387 30385
rect 26329 30376 26341 30379
rect 2188 30348 26341 30376
rect 2188 30336 2194 30348
rect 26329 30345 26341 30348
rect 26375 30376 26387 30379
rect 26970 30376 26976 30388
rect 26375 30348 26976 30376
rect 26375 30345 26387 30348
rect 26329 30339 26387 30345
rect 26970 30336 26976 30348
rect 27028 30336 27034 30388
rect 2133 30243 2191 30249
rect 2133 30209 2145 30243
rect 2179 30240 2191 30243
rect 22370 30240 22376 30252
rect 2179 30212 22376 30240
rect 2179 30209 2191 30212
rect 2133 30203 2191 30209
rect 22370 30200 22376 30212
rect 22428 30200 22434 30252
rect 54021 30243 54079 30249
rect 54021 30240 54033 30243
rect 53484 30212 54033 30240
rect 2222 30132 2228 30184
rect 2280 30172 2286 30184
rect 2409 30175 2467 30181
rect 2409 30172 2421 30175
rect 2280 30144 2421 30172
rect 2280 30132 2286 30144
rect 2409 30141 2421 30144
rect 2455 30141 2467 30175
rect 2409 30135 2467 30141
rect 37642 29996 37648 30048
rect 37700 30036 37706 30048
rect 53484 30045 53512 30212
rect 54021 30209 54033 30212
rect 54067 30209 54079 30243
rect 54021 30203 54079 30209
rect 53469 30039 53527 30045
rect 53469 30036 53481 30039
rect 37700 30008 53481 30036
rect 37700 29996 37706 30008
rect 53469 30005 53481 30008
rect 53515 30005 53527 30039
rect 54202 30036 54208 30048
rect 54163 30008 54208 30036
rect 53469 29999 53527 30005
rect 54202 29996 54208 30008
rect 54260 29996 54266 30048
rect 1104 29946 54832 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 54832 29946
rect 1104 29872 54832 29894
rect 2222 29832 2228 29844
rect 2183 29804 2228 29832
rect 2222 29792 2228 29804
rect 2280 29792 2286 29844
rect 26881 29835 26939 29841
rect 26881 29801 26893 29835
rect 26927 29832 26939 29835
rect 27338 29832 27344 29844
rect 26927 29804 27344 29832
rect 26927 29801 26939 29804
rect 26881 29795 26939 29801
rect 27338 29792 27344 29804
rect 27396 29832 27402 29844
rect 27798 29832 27804 29844
rect 27396 29804 27804 29832
rect 27396 29792 27402 29804
rect 27798 29792 27804 29804
rect 27856 29792 27862 29844
rect 23290 29656 23296 29708
rect 23348 29696 23354 29708
rect 47578 29696 47584 29708
rect 23348 29668 47584 29696
rect 23348 29656 23354 29668
rect 47578 29656 47584 29668
rect 47636 29656 47642 29708
rect 1578 29628 1584 29640
rect 1539 29600 1584 29628
rect 1578 29588 1584 29600
rect 1636 29628 1642 29640
rect 2777 29631 2835 29637
rect 2777 29628 2789 29631
rect 1636 29600 2789 29628
rect 1636 29588 1642 29600
rect 2777 29597 2789 29600
rect 2823 29597 2835 29631
rect 2777 29591 2835 29597
rect 4522 29588 4528 29640
rect 4580 29628 4586 29640
rect 4580 29600 16574 29628
rect 4580 29588 4586 29600
rect 13814 29560 13820 29572
rect 1780 29532 13820 29560
rect 1780 29501 1808 29532
rect 13814 29520 13820 29532
rect 13872 29520 13878 29572
rect 16546 29560 16574 29600
rect 24302 29588 24308 29640
rect 24360 29628 24366 29640
rect 50798 29628 50804 29640
rect 24360 29600 50804 29628
rect 24360 29588 24366 29600
rect 50798 29588 50804 29600
rect 50856 29588 50862 29640
rect 53561 29631 53619 29637
rect 53561 29597 53573 29631
rect 53607 29628 53619 29631
rect 54202 29628 54208 29640
rect 53607 29600 54208 29628
rect 53607 29597 53619 29600
rect 53561 29591 53619 29597
rect 54202 29588 54208 29600
rect 54260 29588 54266 29640
rect 25958 29560 25964 29572
rect 16546 29532 25964 29560
rect 25958 29520 25964 29532
rect 26016 29520 26022 29572
rect 27798 29520 27804 29572
rect 27856 29560 27862 29572
rect 27893 29563 27951 29569
rect 27893 29560 27905 29563
rect 27856 29532 27905 29560
rect 27856 29520 27862 29532
rect 27893 29529 27905 29532
rect 27939 29560 27951 29563
rect 28350 29560 28356 29572
rect 27939 29532 28356 29560
rect 27939 29529 27951 29532
rect 27893 29523 27951 29529
rect 28350 29520 28356 29532
rect 28408 29560 28414 29572
rect 30098 29560 30104 29572
rect 28408 29532 30104 29560
rect 28408 29520 28414 29532
rect 30098 29520 30104 29532
rect 30156 29520 30162 29572
rect 1765 29495 1823 29501
rect 1765 29461 1777 29495
rect 1811 29461 1823 29495
rect 1765 29455 1823 29461
rect 22738 29452 22744 29504
rect 22796 29492 22802 29504
rect 30466 29492 30472 29504
rect 22796 29464 30472 29492
rect 22796 29452 22802 29464
rect 30466 29452 30472 29464
rect 30524 29452 30530 29504
rect 53558 29452 53564 29504
rect 53616 29492 53622 29504
rect 54113 29495 54171 29501
rect 54113 29492 54125 29495
rect 53616 29464 54125 29492
rect 53616 29452 53622 29464
rect 54113 29461 54125 29464
rect 54159 29461 54171 29495
rect 54113 29455 54171 29461
rect 1104 29402 54832 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 54832 29402
rect 1104 29328 54832 29350
rect 25958 29288 25964 29300
rect 25919 29260 25964 29288
rect 25958 29248 25964 29260
rect 26016 29248 26022 29300
rect 28261 29291 28319 29297
rect 28261 29257 28273 29291
rect 28307 29288 28319 29291
rect 30374 29288 30380 29300
rect 28307 29260 30380 29288
rect 28307 29257 28319 29260
rect 28261 29251 28319 29257
rect 11054 29180 11060 29232
rect 11112 29220 11118 29232
rect 14093 29223 14151 29229
rect 14093 29220 14105 29223
rect 11112 29192 14105 29220
rect 11112 29180 11118 29192
rect 14093 29189 14105 29192
rect 14139 29189 14151 29223
rect 25976 29220 26004 29248
rect 27433 29223 27491 29229
rect 27433 29220 27445 29223
rect 25976 29192 27445 29220
rect 14093 29183 14151 29189
rect 27433 29189 27445 29192
rect 27479 29189 27491 29223
rect 27433 29183 27491 29189
rect 2133 29155 2191 29161
rect 2133 29121 2145 29155
rect 2179 29152 2191 29155
rect 4522 29152 4528 29164
rect 2179 29124 4528 29152
rect 2179 29121 2191 29124
rect 2133 29115 2191 29121
rect 4522 29112 4528 29124
rect 4580 29112 4586 29164
rect 13814 29152 13820 29164
rect 13775 29124 13820 29152
rect 13814 29112 13820 29124
rect 13872 29112 13878 29164
rect 14001 29155 14059 29161
rect 14001 29121 14013 29155
rect 14047 29121 14059 29155
rect 14182 29152 14188 29164
rect 14143 29124 14188 29152
rect 14001 29115 14059 29121
rect 2409 29087 2467 29093
rect 2409 29053 2421 29087
rect 2455 29084 2467 29087
rect 2774 29084 2780 29096
rect 2455 29056 2780 29084
rect 2455 29053 2467 29056
rect 2409 29047 2467 29053
rect 2774 29044 2780 29056
rect 2832 29084 2838 29096
rect 2869 29087 2927 29093
rect 2869 29084 2881 29087
rect 2832 29056 2881 29084
rect 2832 29044 2838 29056
rect 2869 29053 2881 29056
rect 2915 29053 2927 29087
rect 2869 29047 2927 29053
rect 13354 29044 13360 29096
rect 13412 29084 13418 29096
rect 14016 29084 14044 29115
rect 14182 29112 14188 29124
rect 14240 29112 14246 29164
rect 24394 29152 24400 29164
rect 14844 29124 24400 29152
rect 14844 29093 14872 29124
rect 24394 29112 24400 29124
rect 24452 29152 24458 29164
rect 26142 29152 26148 29164
rect 24452 29124 26148 29152
rect 24452 29112 24458 29124
rect 26142 29112 26148 29124
rect 26200 29152 26206 29164
rect 26513 29155 26571 29161
rect 26513 29152 26525 29155
rect 26200 29124 26525 29152
rect 26200 29112 26206 29124
rect 26513 29121 26525 29124
rect 26559 29121 26571 29155
rect 26513 29115 26571 29121
rect 27157 29155 27215 29161
rect 27157 29121 27169 29155
rect 27203 29121 27215 29155
rect 27338 29152 27344 29164
rect 27299 29124 27344 29152
rect 27157 29115 27215 29121
rect 14829 29087 14887 29093
rect 14829 29084 14841 29087
rect 13412 29056 14841 29084
rect 13412 29044 13418 29056
rect 14829 29053 14841 29056
rect 14875 29053 14887 29087
rect 21910 29084 21916 29096
rect 14829 29047 14887 29053
rect 16546 29056 21916 29084
rect 14369 29019 14427 29025
rect 14369 28985 14381 29019
rect 14415 29016 14427 29019
rect 16546 29016 16574 29056
rect 21910 29044 21916 29056
rect 21968 29044 21974 29096
rect 14415 28988 16574 29016
rect 26528 29016 26556 29115
rect 27172 29084 27200 29115
rect 27338 29112 27344 29124
rect 27396 29112 27402 29164
rect 27522 29152 27528 29164
rect 27483 29124 27528 29152
rect 27522 29112 27528 29124
rect 27580 29112 27586 29164
rect 28276 29084 28304 29251
rect 30374 29248 30380 29260
rect 30432 29248 30438 29300
rect 30466 29248 30472 29300
rect 30524 29288 30530 29300
rect 53558 29288 53564 29300
rect 30524 29260 53564 29288
rect 30524 29248 30530 29260
rect 53558 29248 53564 29260
rect 53616 29248 53622 29300
rect 54202 29288 54208 29300
rect 54163 29260 54208 29288
rect 54202 29248 54208 29260
rect 54260 29248 54266 29300
rect 54021 29155 54079 29161
rect 54021 29152 54033 29155
rect 27172 29056 28304 29084
rect 53484 29124 54033 29152
rect 27338 29016 27344 29028
rect 26528 28988 27344 29016
rect 14415 28985 14427 28988
rect 14369 28979 14427 28985
rect 27338 28976 27344 28988
rect 27396 29016 27402 29028
rect 27522 29016 27528 29028
rect 27396 28988 27528 29016
rect 27396 28976 27402 28988
rect 27522 28976 27528 28988
rect 27580 28976 27586 29028
rect 35894 28976 35900 29028
rect 35952 29016 35958 29028
rect 53484 29025 53512 29124
rect 54021 29121 54033 29124
rect 54067 29121 54079 29155
rect 54021 29115 54079 29121
rect 53469 29019 53527 29025
rect 53469 29016 53481 29019
rect 35952 28988 53481 29016
rect 35952 28976 35958 28988
rect 53469 28985 53481 28988
rect 53515 28985 53527 29019
rect 53469 28979 53527 28985
rect 27709 28951 27767 28957
rect 27709 28917 27721 28951
rect 27755 28948 27767 28951
rect 28074 28948 28080 28960
rect 27755 28920 28080 28948
rect 27755 28917 27767 28920
rect 27709 28911 27767 28917
rect 28074 28908 28080 28920
rect 28132 28908 28138 28960
rect 53009 28951 53067 28957
rect 53009 28917 53021 28951
rect 53055 28948 53067 28951
rect 54202 28948 54208 28960
rect 53055 28920 54208 28948
rect 53055 28917 53067 28920
rect 53009 28911 53067 28917
rect 54202 28908 54208 28920
rect 54260 28908 54266 28960
rect 1104 28858 54832 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 54832 28858
rect 1104 28784 54832 28806
rect 25406 28704 25412 28756
rect 25464 28744 25470 28756
rect 27065 28747 27123 28753
rect 27065 28744 27077 28747
rect 25464 28716 27077 28744
rect 25464 28704 25470 28716
rect 27065 28713 27077 28716
rect 27111 28713 27123 28747
rect 28905 28747 28963 28753
rect 28905 28744 28917 28747
rect 27065 28707 27123 28713
rect 28276 28716 28917 28744
rect 26694 28568 26700 28620
rect 26752 28608 26758 28620
rect 28276 28608 28304 28716
rect 28905 28713 28917 28716
rect 28951 28744 28963 28747
rect 29914 28744 29920 28756
rect 28951 28716 29920 28744
rect 28951 28713 28963 28716
rect 28905 28707 28963 28713
rect 29914 28704 29920 28716
rect 29972 28704 29978 28756
rect 28353 28679 28411 28685
rect 28353 28645 28365 28679
rect 28399 28676 28411 28679
rect 29546 28676 29552 28688
rect 28399 28648 29552 28676
rect 28399 28645 28411 28648
rect 28353 28639 28411 28645
rect 29546 28636 29552 28648
rect 29604 28636 29610 28688
rect 26752 28580 27108 28608
rect 26752 28568 26758 28580
rect 2133 28543 2191 28549
rect 2133 28509 2145 28543
rect 2179 28509 2191 28543
rect 2133 28503 2191 28509
rect 2409 28543 2467 28549
rect 2409 28509 2421 28543
rect 2455 28540 2467 28543
rect 2774 28540 2780 28552
rect 2455 28512 2780 28540
rect 2455 28509 2467 28512
rect 2409 28503 2467 28509
rect 2148 28472 2176 28503
rect 2774 28500 2780 28512
rect 2832 28540 2838 28552
rect 2869 28543 2927 28549
rect 2869 28540 2881 28543
rect 2832 28512 2881 28540
rect 2832 28500 2838 28512
rect 2869 28509 2881 28512
rect 2915 28509 2927 28543
rect 2869 28503 2927 28509
rect 24578 28500 24584 28552
rect 24636 28540 24642 28552
rect 27080 28549 27108 28580
rect 28184 28580 28304 28608
rect 28184 28549 28212 28580
rect 25593 28543 25651 28549
rect 25593 28540 25605 28543
rect 24636 28512 25605 28540
rect 24636 28500 24642 28512
rect 25593 28509 25605 28512
rect 25639 28540 25651 28543
rect 27065 28543 27123 28549
rect 25639 28512 27016 28540
rect 25639 28509 25651 28512
rect 25593 28503 25651 28509
rect 24670 28472 24676 28484
rect 2148 28444 24676 28472
rect 24670 28432 24676 28444
rect 24728 28432 24734 28484
rect 26510 28472 26516 28484
rect 26471 28444 26516 28472
rect 26510 28432 26516 28444
rect 26568 28432 26574 28484
rect 26988 28472 27016 28512
rect 27065 28509 27077 28543
rect 27111 28509 27123 28543
rect 28169 28543 28227 28549
rect 28169 28540 28181 28543
rect 27065 28503 27123 28509
rect 27632 28512 28181 28540
rect 27522 28472 27528 28484
rect 26988 28444 27528 28472
rect 27522 28432 27528 28444
rect 27580 28432 27586 28484
rect 27632 28416 27660 28512
rect 28169 28509 28181 28512
rect 28215 28509 28227 28543
rect 28350 28540 28356 28552
rect 28311 28512 28356 28540
rect 28169 28503 28227 28509
rect 28350 28500 28356 28512
rect 28408 28500 28414 28552
rect 29733 28543 29791 28549
rect 29733 28509 29745 28543
rect 29779 28540 29791 28543
rect 29822 28540 29828 28552
rect 29779 28512 29828 28540
rect 29779 28509 29791 28512
rect 29733 28503 29791 28509
rect 29822 28500 29828 28512
rect 29880 28500 29886 28552
rect 54202 28540 54208 28552
rect 54163 28512 54208 28540
rect 54202 28500 54208 28512
rect 54260 28500 54266 28552
rect 27798 28432 27804 28484
rect 27856 28472 27862 28484
rect 29917 28475 29975 28481
rect 29917 28472 29929 28475
rect 27856 28444 29929 28472
rect 27856 28432 27862 28444
rect 29917 28441 29929 28444
rect 29963 28441 29975 28475
rect 29917 28435 29975 28441
rect 33502 28432 33508 28484
rect 33560 28472 33566 28484
rect 48590 28472 48596 28484
rect 33560 28444 48596 28472
rect 33560 28432 33566 28444
rect 48590 28432 48596 28444
rect 48648 28432 48654 28484
rect 52825 28475 52883 28481
rect 52825 28441 52837 28475
rect 52871 28472 52883 28475
rect 53466 28472 53472 28484
rect 52871 28444 53472 28472
rect 52871 28441 52883 28444
rect 52825 28435 52883 28441
rect 53466 28432 53472 28444
rect 53524 28432 53530 28484
rect 14182 28364 14188 28416
rect 14240 28404 14246 28416
rect 14553 28407 14611 28413
rect 14553 28404 14565 28407
rect 14240 28376 14565 28404
rect 14240 28364 14246 28376
rect 14553 28373 14565 28376
rect 14599 28404 14611 28407
rect 15102 28404 15108 28416
rect 14599 28376 15108 28404
rect 14599 28373 14611 28376
rect 14553 28367 14611 28373
rect 15102 28364 15108 28376
rect 15160 28364 15166 28416
rect 25133 28407 25191 28413
rect 25133 28373 25145 28407
rect 25179 28404 25191 28407
rect 25222 28404 25228 28416
rect 25179 28376 25228 28404
rect 25179 28373 25191 28376
rect 25133 28367 25191 28373
rect 25222 28364 25228 28376
rect 25280 28404 25286 28416
rect 26421 28407 26479 28413
rect 26421 28404 26433 28407
rect 25280 28376 26433 28404
rect 25280 28364 25286 28376
rect 26421 28373 26433 28376
rect 26467 28404 26479 28407
rect 27062 28404 27068 28416
rect 26467 28376 27068 28404
rect 26467 28373 26479 28376
rect 26421 28367 26479 28373
rect 27062 28364 27068 28376
rect 27120 28404 27126 28416
rect 27614 28404 27620 28416
rect 27120 28376 27620 28404
rect 27120 28364 27126 28376
rect 27614 28364 27620 28376
rect 27672 28364 27678 28416
rect 30098 28404 30104 28416
rect 30059 28376 30104 28404
rect 30098 28364 30104 28376
rect 30156 28364 30162 28416
rect 53190 28364 53196 28416
rect 53248 28404 53254 28416
rect 53377 28407 53435 28413
rect 53377 28404 53389 28407
rect 53248 28376 53389 28404
rect 53248 28364 53254 28376
rect 53377 28373 53389 28376
rect 53423 28373 53435 28407
rect 53377 28367 53435 28373
rect 53558 28364 53564 28416
rect 53616 28404 53622 28416
rect 54113 28407 54171 28413
rect 54113 28404 54125 28407
rect 53616 28376 54125 28404
rect 53616 28364 53622 28376
rect 54113 28373 54125 28376
rect 54159 28373 54171 28407
rect 54113 28367 54171 28373
rect 1104 28314 54832 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 54832 28314
rect 1104 28240 54832 28262
rect 24670 28200 24676 28212
rect 24631 28172 24676 28200
rect 24670 28160 24676 28172
rect 24728 28200 24734 28212
rect 24728 28172 26464 28200
rect 24728 28160 24734 28172
rect 25222 28132 25228 28144
rect 25183 28104 25228 28132
rect 25222 28092 25228 28104
rect 25280 28092 25286 28144
rect 25866 28132 25872 28144
rect 25827 28104 25872 28132
rect 25866 28092 25872 28104
rect 25924 28092 25930 28144
rect 26436 28132 26464 28172
rect 26510 28160 26516 28212
rect 26568 28200 26574 28212
rect 26605 28203 26663 28209
rect 26605 28200 26617 28203
rect 26568 28172 26617 28200
rect 26568 28160 26574 28172
rect 26605 28169 26617 28172
rect 26651 28169 26663 28203
rect 27798 28200 27804 28212
rect 27759 28172 27804 28200
rect 26605 28163 26663 28169
rect 27798 28160 27804 28172
rect 27856 28160 27862 28212
rect 33042 28160 33048 28212
rect 33100 28200 33106 28212
rect 53558 28200 53564 28212
rect 33100 28172 53564 28200
rect 33100 28160 33106 28172
rect 53558 28160 53564 28172
rect 53616 28160 53622 28212
rect 54202 28200 54208 28212
rect 54163 28172 54208 28200
rect 54202 28160 54208 28172
rect 54260 28160 54266 28212
rect 27522 28132 27528 28144
rect 26436 28104 27292 28132
rect 27483 28104 27528 28132
rect 2133 28067 2191 28073
rect 2133 28033 2145 28067
rect 2179 28064 2191 28067
rect 2682 28064 2688 28076
rect 2179 28036 2688 28064
rect 2179 28033 2191 28036
rect 2133 28027 2191 28033
rect 2682 28024 2688 28036
rect 2740 28024 2746 28076
rect 26418 28064 26424 28076
rect 26379 28036 26424 28064
rect 26418 28024 26424 28036
rect 26476 28024 26482 28076
rect 27264 28073 27292 28104
rect 27522 28092 27528 28104
rect 27580 28092 27586 28144
rect 27157 28067 27215 28073
rect 27157 28033 27169 28067
rect 27203 28033 27215 28067
rect 27157 28027 27215 28033
rect 27250 28067 27308 28073
rect 27250 28033 27262 28067
rect 27296 28033 27308 28067
rect 27250 28027 27308 28033
rect 2222 27956 2228 28008
rect 2280 27996 2286 28008
rect 2409 27999 2467 28005
rect 2409 27996 2421 27999
rect 2280 27968 2421 27996
rect 2280 27956 2286 27968
rect 2409 27965 2421 27968
rect 2455 27965 2467 27999
rect 2409 27959 2467 27965
rect 15102 27956 15108 28008
rect 15160 27996 15166 28008
rect 25222 27996 25228 28008
rect 15160 27968 25228 27996
rect 15160 27956 15166 27968
rect 25222 27956 25228 27968
rect 25280 27956 25286 28008
rect 25774 27956 25780 28008
rect 25832 27996 25838 28008
rect 26329 27999 26387 28005
rect 26329 27996 26341 27999
rect 25832 27968 26341 27996
rect 25832 27956 25838 27968
rect 26329 27965 26341 27968
rect 26375 27965 26387 27999
rect 27172 27996 27200 28027
rect 27338 28024 27344 28076
rect 27396 28064 27402 28076
rect 27433 28067 27491 28073
rect 27433 28064 27445 28067
rect 27396 28036 27445 28064
rect 27396 28024 27402 28036
rect 27433 28033 27445 28036
rect 27479 28033 27491 28067
rect 27433 28027 27491 28033
rect 27614 28024 27620 28076
rect 27672 28073 27678 28076
rect 27672 28064 27680 28073
rect 28258 28064 28264 28076
rect 27672 28036 27717 28064
rect 28219 28036 28264 28064
rect 27672 28027 27680 28036
rect 27672 28024 27678 28027
rect 28258 28024 28264 28036
rect 28316 28024 28322 28076
rect 53285 28067 53343 28073
rect 53285 28064 53297 28067
rect 52288 28036 53297 28064
rect 28166 27996 28172 28008
rect 27172 27968 28172 27996
rect 26329 27959 26387 27965
rect 28166 27956 28172 27968
rect 28224 27956 28230 28008
rect 28350 27996 28356 28008
rect 28311 27968 28356 27996
rect 28350 27956 28356 27968
rect 28408 27956 28414 28008
rect 25869 27931 25927 27937
rect 25869 27897 25881 27931
rect 25915 27928 25927 27931
rect 26602 27928 26608 27940
rect 25915 27900 26608 27928
rect 25915 27897 25927 27900
rect 25869 27891 25927 27897
rect 26602 27888 26608 27900
rect 26660 27888 26666 27940
rect 27338 27888 27344 27940
rect 27396 27928 27402 27940
rect 29089 27931 29147 27937
rect 29089 27928 29101 27931
rect 27396 27900 29101 27928
rect 27396 27888 27402 27900
rect 29089 27897 29101 27900
rect 29135 27897 29147 27931
rect 29089 27891 29147 27897
rect 28074 27820 28080 27872
rect 28132 27860 28138 27872
rect 28261 27863 28319 27869
rect 28261 27860 28273 27863
rect 28132 27832 28273 27860
rect 28132 27820 28138 27832
rect 28261 27829 28273 27832
rect 28307 27829 28319 27863
rect 28626 27860 28632 27872
rect 28587 27832 28632 27860
rect 28261 27823 28319 27829
rect 28626 27820 28632 27832
rect 28684 27820 28690 27872
rect 37458 27820 37464 27872
rect 37516 27860 37522 27872
rect 52288 27869 52316 28036
rect 53285 28033 53297 28036
rect 53331 28033 53343 28067
rect 53285 28027 53343 28033
rect 54021 28067 54079 28073
rect 54021 28033 54033 28067
rect 54067 28033 54079 28067
rect 54021 28027 54079 28033
rect 52822 27956 52828 28008
rect 52880 27996 52886 28008
rect 54036 27996 54064 28027
rect 52880 27968 54064 27996
rect 52880 27956 52886 27968
rect 52273 27863 52331 27869
rect 52273 27860 52285 27863
rect 37516 27832 52285 27860
rect 37516 27820 37522 27832
rect 52273 27829 52285 27832
rect 52319 27829 52331 27863
rect 53466 27860 53472 27872
rect 53427 27832 53472 27860
rect 52273 27823 52331 27829
rect 53466 27820 53472 27832
rect 53524 27820 53530 27872
rect 1104 27770 54832 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 54832 27770
rect 1104 27696 54832 27718
rect 2222 27656 2228 27668
rect 2183 27628 2228 27656
rect 2222 27616 2228 27628
rect 2280 27616 2286 27668
rect 25041 27659 25099 27665
rect 25041 27656 25053 27659
rect 24780 27628 25053 27656
rect 24394 27548 24400 27600
rect 24452 27588 24458 27600
rect 24780 27588 24808 27628
rect 25041 27625 25053 27628
rect 25087 27625 25099 27659
rect 25041 27619 25099 27625
rect 26418 27588 26424 27600
rect 24452 27560 24808 27588
rect 26379 27560 26424 27588
rect 24452 27548 24458 27560
rect 26418 27548 26424 27560
rect 26476 27548 26482 27600
rect 27157 27591 27215 27597
rect 27157 27557 27169 27591
rect 27203 27588 27215 27591
rect 28350 27588 28356 27600
rect 27203 27560 28356 27588
rect 27203 27557 27215 27560
rect 27157 27551 27215 27557
rect 28350 27548 28356 27560
rect 28408 27548 28414 27600
rect 23934 27480 23940 27532
rect 23992 27520 23998 27532
rect 24029 27523 24087 27529
rect 24029 27520 24041 27523
rect 23992 27492 24041 27520
rect 23992 27480 23998 27492
rect 24029 27489 24041 27492
rect 24075 27520 24087 27523
rect 28261 27523 28319 27529
rect 24075 27492 27476 27520
rect 24075 27489 24087 27492
rect 24029 27483 24087 27489
rect 1578 27452 1584 27464
rect 1539 27424 1584 27452
rect 1578 27412 1584 27424
rect 1636 27452 1642 27464
rect 2777 27455 2835 27461
rect 2777 27452 2789 27455
rect 1636 27424 2789 27452
rect 1636 27412 1642 27424
rect 2777 27421 2789 27424
rect 2823 27421 2835 27455
rect 2777 27415 2835 27421
rect 25041 27455 25099 27461
rect 25041 27421 25053 27455
rect 25087 27421 25099 27455
rect 25222 27452 25228 27464
rect 25183 27424 25228 27452
rect 25041 27415 25099 27421
rect 11054 27384 11060 27396
rect 1780 27356 11060 27384
rect 1780 27325 1808 27356
rect 11054 27344 11060 27356
rect 11112 27344 11118 27396
rect 25056 27384 25084 27415
rect 25222 27412 25228 27424
rect 25280 27412 25286 27464
rect 25866 27452 25872 27464
rect 25827 27424 25872 27452
rect 25866 27412 25872 27424
rect 25924 27412 25930 27464
rect 26237 27455 26295 27461
rect 26237 27421 26249 27455
rect 26283 27452 26295 27455
rect 26510 27452 26516 27464
rect 26283 27424 26516 27452
rect 26283 27421 26295 27424
rect 26237 27415 26295 27421
rect 26510 27412 26516 27424
rect 26568 27412 26574 27464
rect 27062 27412 27068 27464
rect 27120 27452 27126 27464
rect 27448 27461 27476 27492
rect 28261 27489 28273 27523
rect 28307 27520 28319 27523
rect 28626 27520 28632 27532
rect 28307 27492 28632 27520
rect 28307 27489 28319 27492
rect 28261 27483 28319 27489
rect 28626 27480 28632 27492
rect 28684 27480 28690 27532
rect 27295 27455 27353 27461
rect 27295 27452 27307 27455
rect 27120 27424 27307 27452
rect 27120 27412 27126 27424
rect 27295 27421 27307 27424
rect 27341 27421 27353 27455
rect 27295 27415 27353 27421
rect 27433 27455 27491 27461
rect 27433 27421 27445 27455
rect 27479 27421 27491 27455
rect 27706 27452 27712 27464
rect 27667 27424 27712 27452
rect 27433 27415 27491 27421
rect 27706 27412 27712 27424
rect 27764 27412 27770 27464
rect 27801 27455 27859 27461
rect 27801 27421 27813 27455
rect 27847 27452 27859 27455
rect 27890 27452 27896 27464
rect 27847 27424 27896 27452
rect 27847 27421 27859 27424
rect 27801 27415 27859 27421
rect 27890 27412 27896 27424
rect 27948 27412 27954 27464
rect 28537 27455 28595 27461
rect 28537 27421 28549 27455
rect 28583 27452 28595 27455
rect 29822 27452 29828 27464
rect 28583 27424 29828 27452
rect 28583 27421 28595 27424
rect 28537 27415 28595 27421
rect 29822 27412 29828 27424
rect 29880 27412 29886 27464
rect 29917 27455 29975 27461
rect 29917 27421 29929 27455
rect 29963 27452 29975 27455
rect 30098 27452 30104 27464
rect 29963 27424 30104 27452
rect 29963 27421 29975 27424
rect 29917 27415 29975 27421
rect 30098 27412 30104 27424
rect 30156 27412 30162 27464
rect 52457 27455 52515 27461
rect 52457 27421 52469 27455
rect 52503 27452 52515 27455
rect 53466 27452 53472 27464
rect 52503 27424 53472 27452
rect 52503 27421 52515 27424
rect 52457 27415 52515 27421
rect 53466 27412 53472 27424
rect 53524 27412 53530 27464
rect 53650 27412 53656 27464
rect 53708 27452 53714 27464
rect 53745 27455 53803 27461
rect 53745 27452 53757 27455
rect 53708 27424 53757 27452
rect 53708 27412 53714 27424
rect 53745 27421 53757 27424
rect 53791 27421 53803 27455
rect 53745 27415 53803 27421
rect 26050 27384 26056 27396
rect 25056 27356 26056 27384
rect 26050 27344 26056 27356
rect 26108 27344 26114 27396
rect 26142 27344 26148 27396
rect 26200 27384 26206 27396
rect 27525 27387 27583 27393
rect 26200 27356 26245 27384
rect 26200 27344 26206 27356
rect 27525 27353 27537 27387
rect 27571 27353 27583 27387
rect 27525 27347 27583 27353
rect 1765 27319 1823 27325
rect 1765 27285 1777 27319
rect 1811 27285 1823 27319
rect 25406 27316 25412 27328
rect 25367 27288 25412 27316
rect 1765 27279 1823 27285
rect 25406 27276 25412 27288
rect 25464 27276 25470 27328
rect 27062 27276 27068 27328
rect 27120 27316 27126 27328
rect 27540 27316 27568 27347
rect 27120 27288 27568 27316
rect 29825 27319 29883 27325
rect 27120 27276 27126 27288
rect 29825 27285 29837 27319
rect 29871 27316 29883 27319
rect 33778 27316 33784 27328
rect 29871 27288 33784 27316
rect 29871 27285 29883 27288
rect 29825 27279 29883 27285
rect 33778 27276 33784 27288
rect 33836 27276 33842 27328
rect 52822 27276 52828 27328
rect 52880 27316 52886 27328
rect 52917 27319 52975 27325
rect 52917 27316 52929 27319
rect 52880 27288 52929 27316
rect 52880 27276 52886 27288
rect 52917 27285 52929 27288
rect 52963 27285 52975 27319
rect 52917 27279 52975 27285
rect 1104 27226 54832 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 54832 27226
rect 1104 27152 54832 27174
rect 24394 27112 24400 27124
rect 24355 27084 24400 27112
rect 24394 27072 24400 27084
rect 24452 27072 24458 27124
rect 25222 27072 25228 27124
rect 25280 27112 25286 27124
rect 25501 27115 25559 27121
rect 25501 27112 25513 27115
rect 25280 27084 25513 27112
rect 25280 27072 25286 27084
rect 25501 27081 25513 27084
rect 25547 27081 25559 27115
rect 25501 27075 25559 27081
rect 25866 27072 25872 27124
rect 25924 27112 25930 27124
rect 28813 27115 28871 27121
rect 28813 27112 28825 27115
rect 25924 27084 28825 27112
rect 25924 27072 25930 27084
rect 28813 27081 28825 27084
rect 28859 27081 28871 27115
rect 34514 27112 34520 27124
rect 34475 27084 34520 27112
rect 28813 27075 28871 27081
rect 25406 27004 25412 27056
rect 25464 27044 25470 27056
rect 25464 27016 28120 27044
rect 25464 27004 25470 27016
rect 25958 26936 25964 26988
rect 26016 26976 26022 26988
rect 26053 26979 26111 26985
rect 26053 26976 26065 26979
rect 26016 26948 26065 26976
rect 26016 26936 26022 26948
rect 26053 26945 26065 26948
rect 26099 26945 26111 26979
rect 27062 26976 27068 26988
rect 26053 26939 26111 26945
rect 26344 26948 27068 26976
rect 2133 26911 2191 26917
rect 2133 26877 2145 26911
rect 2179 26877 2191 26911
rect 2133 26871 2191 26877
rect 2409 26911 2467 26917
rect 2409 26877 2421 26911
rect 2455 26908 2467 26911
rect 2774 26908 2780 26920
rect 2455 26880 2780 26908
rect 2455 26877 2467 26880
rect 2409 26871 2467 26877
rect 2148 26840 2176 26871
rect 2774 26868 2780 26880
rect 2832 26908 2838 26920
rect 2869 26911 2927 26917
rect 2869 26908 2881 26911
rect 2832 26880 2881 26908
rect 2832 26868 2838 26880
rect 2869 26877 2881 26880
rect 2915 26877 2927 26911
rect 2869 26871 2927 26877
rect 25041 26911 25099 26917
rect 25041 26877 25053 26911
rect 25087 26908 25099 26911
rect 25682 26908 25688 26920
rect 25087 26880 25688 26908
rect 25087 26877 25099 26880
rect 25041 26871 25099 26877
rect 25682 26868 25688 26880
rect 25740 26908 25746 26920
rect 26344 26908 26372 26948
rect 27062 26936 27068 26948
rect 27120 26936 27126 26988
rect 27430 26936 27436 26988
rect 27488 26976 27494 26988
rect 28092 26985 28120 27016
rect 27525 26979 27583 26985
rect 27525 26976 27537 26979
rect 27488 26948 27537 26976
rect 27488 26936 27494 26948
rect 27525 26945 27537 26948
rect 27571 26945 27583 26979
rect 27525 26939 27583 26945
rect 28077 26979 28135 26985
rect 28077 26945 28089 26979
rect 28123 26945 28135 26979
rect 28077 26939 28135 26945
rect 26510 26908 26516 26920
rect 25740 26880 26372 26908
rect 26423 26880 26516 26908
rect 25740 26868 25746 26880
rect 26510 26868 26516 26880
rect 26568 26908 26574 26920
rect 26878 26908 26884 26920
rect 26568 26880 26884 26908
rect 26568 26868 26574 26880
rect 26878 26868 26884 26880
rect 26936 26868 26942 26920
rect 23934 26840 23940 26852
rect 2148 26812 23940 26840
rect 23934 26800 23940 26812
rect 23992 26800 23998 26852
rect 25774 26800 25780 26852
rect 25832 26840 25838 26852
rect 27249 26843 27307 26849
rect 27249 26840 27261 26843
rect 25832 26812 27261 26840
rect 25832 26800 25838 26812
rect 27249 26809 27261 26812
rect 27295 26809 27307 26843
rect 28828 26840 28856 27075
rect 34514 27072 34520 27084
rect 34572 27072 34578 27124
rect 35897 27115 35955 27121
rect 35897 27081 35909 27115
rect 35943 27112 35955 27115
rect 36078 27112 36084 27124
rect 35943 27084 36084 27112
rect 35943 27081 35955 27084
rect 35897 27075 35955 27081
rect 36078 27072 36084 27084
rect 36136 27072 36142 27124
rect 51813 27047 51871 27053
rect 51813 27013 51825 27047
rect 51859 27044 51871 27047
rect 54202 27044 54208 27056
rect 51859 27016 54208 27044
rect 51859 27013 51871 27016
rect 51813 27007 51871 27013
rect 54202 27004 54208 27016
rect 54260 27004 54266 27056
rect 52365 26979 52423 26985
rect 52365 26945 52377 26979
rect 52411 26976 52423 26979
rect 53469 26979 53527 26985
rect 53469 26976 53481 26979
rect 52411 26948 53481 26976
rect 52411 26945 52423 26948
rect 52365 26939 52423 26945
rect 53469 26945 53481 26948
rect 53515 26976 53527 26979
rect 53558 26976 53564 26988
rect 53515 26948 53564 26976
rect 53515 26945 53527 26948
rect 53469 26939 53527 26945
rect 53558 26936 53564 26948
rect 53616 26936 53622 26988
rect 31754 26868 31760 26920
rect 31812 26908 31818 26920
rect 48498 26908 48504 26920
rect 31812 26880 48504 26908
rect 31812 26868 31818 26880
rect 48498 26868 48504 26880
rect 48556 26868 48562 26920
rect 39574 26840 39580 26852
rect 28828 26812 39580 26840
rect 27249 26803 27307 26809
rect 39574 26800 39580 26812
rect 39632 26800 39638 26852
rect 52546 26800 52552 26852
rect 52604 26840 52610 26852
rect 54021 26843 54079 26849
rect 54021 26840 54033 26843
rect 52604 26812 54033 26840
rect 52604 26800 52610 26812
rect 54021 26809 54033 26812
rect 54067 26809 54079 26843
rect 54021 26803 54079 26809
rect 26329 26775 26387 26781
rect 26329 26741 26341 26775
rect 26375 26772 26387 26775
rect 26418 26772 26424 26784
rect 26375 26744 26424 26772
rect 26375 26741 26387 26744
rect 26329 26735 26387 26741
rect 26418 26732 26424 26744
rect 26476 26772 26482 26784
rect 26602 26772 26608 26784
rect 26476 26744 26608 26772
rect 26476 26732 26482 26744
rect 26602 26732 26608 26744
rect 26660 26732 26666 26784
rect 28258 26772 28264 26784
rect 28219 26744 28264 26772
rect 28258 26732 28264 26744
rect 28316 26732 28322 26784
rect 34330 26732 34336 26784
rect 34388 26772 34394 26784
rect 35069 26775 35127 26781
rect 35069 26772 35081 26775
rect 34388 26744 35081 26772
rect 34388 26732 34394 26744
rect 35069 26741 35081 26744
rect 35115 26772 35127 26775
rect 35710 26772 35716 26784
rect 35115 26744 35716 26772
rect 35115 26741 35127 26744
rect 35069 26735 35127 26741
rect 35710 26732 35716 26744
rect 35768 26732 35774 26784
rect 52362 26732 52368 26784
rect 52420 26772 52426 26784
rect 53377 26775 53435 26781
rect 53377 26772 53389 26775
rect 52420 26744 53389 26772
rect 52420 26732 52426 26744
rect 53377 26741 53389 26744
rect 53423 26741 53435 26775
rect 53377 26735 53435 26741
rect 1104 26682 54832 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 54832 26682
rect 1104 26608 54832 26630
rect 23658 26528 23664 26580
rect 23716 26568 23722 26580
rect 26053 26571 26111 26577
rect 26053 26568 26065 26571
rect 23716 26540 26065 26568
rect 23716 26528 23722 26540
rect 26053 26537 26065 26540
rect 26099 26568 26111 26571
rect 27154 26568 27160 26580
rect 26099 26540 27160 26568
rect 26099 26537 26111 26540
rect 26053 26531 26111 26537
rect 27154 26528 27160 26540
rect 27212 26528 27218 26580
rect 34330 26568 34336 26580
rect 34291 26540 34336 26568
rect 34330 26528 34336 26540
rect 34388 26528 34394 26580
rect 35986 26568 35992 26580
rect 35947 26540 35992 26568
rect 35986 26528 35992 26540
rect 36044 26528 36050 26580
rect 36170 26528 36176 26580
rect 36228 26568 36234 26580
rect 36538 26568 36544 26580
rect 36228 26540 36544 26568
rect 36228 26528 36234 26540
rect 36538 26528 36544 26540
rect 36596 26528 36602 26580
rect 37185 26571 37243 26577
rect 37185 26537 37197 26571
rect 37231 26568 37243 26571
rect 37458 26568 37464 26580
rect 37231 26540 37464 26568
rect 37231 26537 37243 26540
rect 37185 26531 37243 26537
rect 37458 26528 37464 26540
rect 37516 26528 37522 26580
rect 42610 26528 42616 26580
rect 42668 26568 42674 26580
rect 52362 26568 52368 26580
rect 42668 26540 52368 26568
rect 42668 26528 42674 26540
rect 52362 26528 52368 26540
rect 52420 26528 52426 26580
rect 54202 26568 54208 26580
rect 54163 26540 54208 26568
rect 54202 26528 54208 26540
rect 54260 26528 54266 26580
rect 2682 26460 2688 26512
rect 2740 26500 2746 26512
rect 2740 26472 16574 26500
rect 2740 26460 2746 26472
rect 2133 26435 2191 26441
rect 2133 26401 2145 26435
rect 2179 26432 2191 26435
rect 16546 26432 16574 26472
rect 26694 26460 26700 26512
rect 26752 26500 26758 26512
rect 26789 26503 26847 26509
rect 26789 26500 26801 26503
rect 26752 26472 26801 26500
rect 26752 26460 26758 26472
rect 26789 26469 26801 26472
rect 26835 26469 26847 26503
rect 26789 26463 26847 26469
rect 28258 26460 28264 26512
rect 28316 26500 28322 26512
rect 35529 26503 35587 26509
rect 28316 26472 35388 26500
rect 28316 26460 28322 26472
rect 25501 26435 25559 26441
rect 25501 26432 25513 26435
rect 2179 26404 6914 26432
rect 16546 26404 25513 26432
rect 2179 26401 2191 26404
rect 2133 26395 2191 26401
rect 2222 26324 2228 26376
rect 2280 26364 2286 26376
rect 2409 26367 2467 26373
rect 2409 26364 2421 26367
rect 2280 26336 2421 26364
rect 2280 26324 2286 26336
rect 2409 26333 2421 26336
rect 2455 26333 2467 26367
rect 6886 26364 6914 26404
rect 25501 26401 25513 26404
rect 25547 26432 25559 26435
rect 26142 26432 26148 26444
rect 25547 26404 26148 26432
rect 25547 26401 25559 26404
rect 25501 26395 25559 26401
rect 26142 26392 26148 26404
rect 26200 26392 26206 26444
rect 26237 26435 26295 26441
rect 26237 26401 26249 26435
rect 26283 26432 26295 26435
rect 26602 26432 26608 26444
rect 26283 26404 26608 26432
rect 26283 26401 26295 26404
rect 26237 26395 26295 26401
rect 26602 26392 26608 26404
rect 26660 26432 26666 26444
rect 27430 26432 27436 26444
rect 26660 26404 27436 26432
rect 26660 26392 26666 26404
rect 27430 26392 27436 26404
rect 27488 26392 27494 26444
rect 24578 26364 24584 26376
rect 6886 26336 24584 26364
rect 2409 26327 2467 26333
rect 24578 26324 24584 26336
rect 24636 26324 24642 26376
rect 26329 26367 26387 26373
rect 26329 26333 26341 26367
rect 26375 26364 26387 26367
rect 26418 26364 26424 26376
rect 26375 26336 26424 26364
rect 26375 26333 26387 26336
rect 26329 26327 26387 26333
rect 26418 26324 26424 26336
rect 26476 26324 26482 26376
rect 27706 26324 27712 26376
rect 27764 26364 27770 26376
rect 28169 26367 28227 26373
rect 28169 26364 28181 26367
rect 27764 26336 28181 26364
rect 27764 26324 27770 26336
rect 28169 26333 28181 26336
rect 28215 26364 28227 26367
rect 35360 26364 35388 26472
rect 35529 26469 35541 26503
rect 35575 26500 35587 26503
rect 35894 26500 35900 26512
rect 35575 26472 35900 26500
rect 35575 26469 35587 26472
rect 35529 26463 35587 26469
rect 35894 26460 35900 26472
rect 35952 26460 35958 26512
rect 43346 26460 43352 26512
rect 43404 26500 43410 26512
rect 52546 26500 52552 26512
rect 43404 26472 52552 26500
rect 43404 26460 43410 26472
rect 52546 26460 52552 26472
rect 52604 26460 52610 26512
rect 53377 26503 53435 26509
rect 53377 26469 53389 26503
rect 53423 26469 53435 26503
rect 53377 26463 53435 26469
rect 44082 26392 44088 26444
rect 44140 26432 44146 26444
rect 53392 26432 53420 26463
rect 44140 26404 53420 26432
rect 44140 26392 44146 26404
rect 42426 26364 42432 26376
rect 28215 26336 33456 26364
rect 35360 26336 42432 26364
rect 28215 26333 28227 26336
rect 28169 26327 28227 26333
rect 25958 26256 25964 26308
rect 26016 26296 26022 26308
rect 26234 26296 26240 26308
rect 26016 26268 26240 26296
rect 26016 26256 26022 26268
rect 26234 26256 26240 26268
rect 26292 26296 26298 26308
rect 26789 26299 26847 26305
rect 26789 26296 26801 26299
rect 26292 26268 26801 26296
rect 26292 26256 26298 26268
rect 26789 26265 26801 26268
rect 26835 26296 26847 26299
rect 27341 26299 27399 26305
rect 27341 26296 27353 26299
rect 26835 26268 27353 26296
rect 26835 26265 26847 26268
rect 26789 26259 26847 26265
rect 27341 26265 27353 26268
rect 27387 26265 27399 26299
rect 27522 26296 27528 26308
rect 27483 26268 27528 26296
rect 27341 26259 27399 26265
rect 27522 26256 27528 26268
rect 27580 26256 27586 26308
rect 33428 26296 33456 26336
rect 42426 26324 42432 26336
rect 42484 26324 42490 26376
rect 52825 26367 52883 26373
rect 52825 26333 52837 26367
rect 52871 26364 52883 26367
rect 53558 26364 53564 26376
rect 52871 26336 53564 26364
rect 52871 26333 52883 26336
rect 52825 26327 52883 26333
rect 53558 26324 53564 26336
rect 53616 26324 53622 26376
rect 54021 26367 54079 26373
rect 54021 26333 54033 26367
rect 54067 26333 54079 26367
rect 54021 26327 54079 26333
rect 44910 26296 44916 26308
rect 33428 26268 44916 26296
rect 44910 26256 44916 26268
rect 44968 26256 44974 26308
rect 52914 26256 52920 26308
rect 52972 26296 52978 26308
rect 54036 26296 54064 26327
rect 52972 26268 54064 26296
rect 52972 26256 52978 26268
rect 31938 26188 31944 26240
rect 31996 26228 32002 26240
rect 33321 26231 33379 26237
rect 33321 26228 33333 26231
rect 31996 26200 33333 26228
rect 31996 26188 32002 26200
rect 33321 26197 33333 26200
rect 33367 26197 33379 26231
rect 33321 26191 33379 26197
rect 34422 26188 34428 26240
rect 34480 26228 34486 26240
rect 34885 26231 34943 26237
rect 34885 26228 34897 26231
rect 34480 26200 34897 26228
rect 34480 26188 34486 26200
rect 34885 26197 34897 26200
rect 34931 26197 34943 26231
rect 34885 26191 34943 26197
rect 1104 26138 54832 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 54832 26138
rect 1104 26064 54832 26086
rect 2222 26024 2228 26036
rect 2183 25996 2228 26024
rect 2222 25984 2228 25996
rect 2280 25984 2286 26036
rect 26326 25984 26332 26036
rect 26384 26024 26390 26036
rect 26421 26027 26479 26033
rect 26421 26024 26433 26027
rect 26384 25996 26433 26024
rect 26384 25984 26390 25996
rect 26421 25993 26433 25996
rect 26467 25993 26479 26027
rect 27246 26024 27252 26036
rect 27207 25996 27252 26024
rect 26421 25987 26479 25993
rect 27246 25984 27252 25996
rect 27304 25984 27310 26036
rect 32585 26027 32643 26033
rect 32585 25993 32597 26027
rect 32631 26024 32643 26027
rect 32858 26024 32864 26036
rect 32631 25996 32864 26024
rect 32631 25993 32643 25996
rect 32585 25987 32643 25993
rect 32858 25984 32864 25996
rect 32916 26024 32922 26036
rect 33410 26024 33416 26036
rect 32916 25996 33416 26024
rect 32916 25984 32922 25996
rect 33410 25984 33416 25996
rect 33468 25984 33474 26036
rect 33594 26024 33600 26036
rect 33555 25996 33600 26024
rect 33594 25984 33600 25996
rect 33652 25984 33658 26036
rect 35710 25984 35716 26036
rect 35768 26024 35774 26036
rect 35805 26027 35863 26033
rect 35805 26024 35817 26027
rect 35768 25996 35817 26024
rect 35768 25984 35774 25996
rect 35805 25993 35817 25996
rect 35851 26024 35863 26027
rect 37461 26027 37519 26033
rect 37461 26024 37473 26027
rect 35851 25996 37473 26024
rect 35851 25993 35863 25996
rect 35805 25987 35863 25993
rect 37461 25993 37473 25996
rect 37507 26024 37519 26027
rect 38194 26024 38200 26036
rect 37507 25996 38200 26024
rect 37507 25993 37519 25996
rect 37461 25987 37519 25993
rect 38194 25984 38200 25996
rect 38252 25984 38258 26036
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 25406 25888 25412 25900
rect 25367 25860 25412 25888
rect 25406 25848 25412 25860
rect 25464 25848 25470 25900
rect 26237 25891 26295 25897
rect 26237 25857 26249 25891
rect 26283 25888 26295 25891
rect 26694 25888 26700 25900
rect 26283 25860 26700 25888
rect 26283 25857 26295 25860
rect 26237 25851 26295 25857
rect 26694 25848 26700 25860
rect 26752 25848 26758 25900
rect 27525 25891 27583 25897
rect 27525 25857 27537 25891
rect 27571 25888 27583 25891
rect 28994 25888 29000 25900
rect 27571 25860 29000 25888
rect 27571 25857 27583 25860
rect 27525 25851 27583 25857
rect 28994 25848 29000 25860
rect 29052 25848 29058 25900
rect 34514 25888 34520 25900
rect 34475 25860 34520 25888
rect 34514 25848 34520 25860
rect 34572 25848 34578 25900
rect 35345 25891 35403 25897
rect 35345 25857 35357 25891
rect 35391 25888 35403 25891
rect 35434 25888 35440 25900
rect 35391 25860 35440 25888
rect 35391 25857 35403 25860
rect 35345 25851 35403 25857
rect 35434 25848 35440 25860
rect 35492 25848 35498 25900
rect 21634 25780 21640 25832
rect 21692 25820 21698 25832
rect 33042 25820 33048 25832
rect 21692 25792 33048 25820
rect 21692 25780 21698 25792
rect 33042 25780 33048 25792
rect 33100 25780 33106 25832
rect 33137 25823 33195 25829
rect 33137 25789 33149 25823
rect 33183 25820 33195 25823
rect 34333 25823 34391 25829
rect 34333 25820 34345 25823
rect 33183 25792 34345 25820
rect 33183 25789 33195 25792
rect 33137 25783 33195 25789
rect 34333 25789 34345 25792
rect 34379 25820 34391 25823
rect 34422 25820 34428 25832
rect 34379 25792 34428 25820
rect 34379 25789 34391 25792
rect 34333 25783 34391 25789
rect 1765 25755 1823 25761
rect 1765 25721 1777 25755
rect 1811 25752 1823 25755
rect 14550 25752 14556 25764
rect 1811 25724 14556 25752
rect 1811 25721 1823 25724
rect 1765 25715 1823 25721
rect 14550 25712 14556 25724
rect 14608 25712 14614 25764
rect 14918 25712 14924 25764
rect 14976 25752 14982 25764
rect 28258 25752 28264 25764
rect 14976 25724 28264 25752
rect 14976 25712 14982 25724
rect 28258 25712 28264 25724
rect 28316 25712 28322 25764
rect 32858 25712 32864 25764
rect 32916 25752 32922 25764
rect 33152 25752 33180 25783
rect 34422 25780 34428 25792
rect 34480 25780 34486 25832
rect 52365 25823 52423 25829
rect 52365 25789 52377 25823
rect 52411 25820 52423 25823
rect 53466 25820 53472 25832
rect 52411 25792 53472 25820
rect 52411 25789 52423 25792
rect 52365 25783 52423 25789
rect 53466 25780 53472 25792
rect 53524 25780 53530 25832
rect 53742 25820 53748 25832
rect 53703 25792 53748 25820
rect 53742 25780 53748 25792
rect 53800 25780 53806 25832
rect 32916 25724 33180 25752
rect 32916 25712 32922 25724
rect 35526 25712 35532 25764
rect 35584 25752 35590 25764
rect 36449 25755 36507 25761
rect 36449 25752 36461 25755
rect 35584 25724 36461 25752
rect 35584 25712 35590 25724
rect 36449 25721 36461 25724
rect 36495 25752 36507 25755
rect 52822 25752 52828 25764
rect 36495 25724 52828 25752
rect 36495 25721 36507 25724
rect 36449 25715 36507 25721
rect 52822 25712 52828 25724
rect 52880 25712 52886 25764
rect 25222 25684 25228 25696
rect 25183 25656 25228 25684
rect 25222 25644 25228 25656
rect 25280 25644 25286 25696
rect 34698 25684 34704 25696
rect 34659 25656 34704 25684
rect 34698 25644 34704 25656
rect 34756 25644 34762 25696
rect 35161 25687 35219 25693
rect 35161 25653 35173 25687
rect 35207 25684 35219 25687
rect 35342 25684 35348 25696
rect 35207 25656 35348 25684
rect 35207 25653 35219 25656
rect 35161 25647 35219 25653
rect 35342 25644 35348 25656
rect 35400 25644 35406 25696
rect 38841 25687 38899 25693
rect 38841 25653 38853 25687
rect 38887 25684 38899 25687
rect 39022 25684 39028 25696
rect 38887 25656 39028 25684
rect 38887 25653 38899 25656
rect 38841 25647 38899 25653
rect 39022 25644 39028 25656
rect 39080 25644 39086 25696
rect 52914 25684 52920 25696
rect 52875 25656 52920 25684
rect 52914 25644 52920 25656
rect 52972 25644 52978 25696
rect 1104 25594 54832 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 54832 25594
rect 1104 25520 54832 25542
rect 1578 25440 1584 25492
rect 1636 25480 1642 25492
rect 2225 25483 2283 25489
rect 2225 25480 2237 25483
rect 1636 25452 2237 25480
rect 1636 25440 1642 25452
rect 2225 25449 2237 25452
rect 2271 25449 2283 25483
rect 2225 25443 2283 25449
rect 25685 25483 25743 25489
rect 25685 25449 25697 25483
rect 25731 25480 25743 25483
rect 26234 25480 26240 25492
rect 25731 25452 26240 25480
rect 25731 25449 25743 25452
rect 25685 25443 25743 25449
rect 26234 25440 26240 25452
rect 26292 25440 26298 25492
rect 28994 25480 29000 25492
rect 28955 25452 29000 25480
rect 28994 25440 29000 25452
rect 29052 25440 29058 25492
rect 31938 25480 31944 25492
rect 31899 25452 31944 25480
rect 31938 25440 31944 25452
rect 31996 25440 32002 25492
rect 32398 25480 32404 25492
rect 32359 25452 32404 25480
rect 32398 25440 32404 25452
rect 32456 25440 32462 25492
rect 35253 25483 35311 25489
rect 35253 25449 35265 25483
rect 35299 25480 35311 25483
rect 35434 25480 35440 25492
rect 35299 25452 35440 25480
rect 35299 25449 35311 25452
rect 35253 25443 35311 25449
rect 35434 25440 35440 25452
rect 35492 25440 35498 25492
rect 37642 25480 37648 25492
rect 37603 25452 37648 25480
rect 37642 25440 37648 25452
rect 37700 25440 37706 25492
rect 39022 25440 39028 25492
rect 39080 25480 39086 25492
rect 52733 25483 52791 25489
rect 52733 25480 52745 25483
rect 39080 25452 52745 25480
rect 39080 25440 39086 25452
rect 52733 25449 52745 25452
rect 52779 25449 52791 25483
rect 54202 25480 54208 25492
rect 54163 25452 54208 25480
rect 52733 25443 52791 25449
rect 35802 25412 35808 25424
rect 34072 25384 35808 25412
rect 25685 25347 25743 25353
rect 25685 25313 25697 25347
rect 25731 25344 25743 25347
rect 25774 25344 25780 25356
rect 25731 25316 25780 25344
rect 25731 25313 25743 25316
rect 25685 25307 25743 25313
rect 25774 25304 25780 25316
rect 25832 25304 25838 25356
rect 26053 25347 26111 25353
rect 26053 25313 26065 25347
rect 26099 25344 26111 25347
rect 26418 25344 26424 25356
rect 26099 25316 26424 25344
rect 26099 25313 26111 25316
rect 26053 25307 26111 25313
rect 26418 25304 26424 25316
rect 26476 25304 26482 25356
rect 28994 25304 29000 25356
rect 29052 25344 29058 25356
rect 30006 25344 30012 25356
rect 29052 25316 30012 25344
rect 29052 25304 29058 25316
rect 30006 25304 30012 25316
rect 30064 25304 30070 25356
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25276 1642 25288
rect 2777 25279 2835 25285
rect 2777 25276 2789 25279
rect 1636 25248 2789 25276
rect 1636 25236 1642 25248
rect 2777 25245 2789 25248
rect 2823 25245 2835 25279
rect 24854 25276 24860 25288
rect 24815 25248 24860 25276
rect 2777 25239 2835 25245
rect 24854 25236 24860 25248
rect 24912 25236 24918 25288
rect 26602 25276 26608 25288
rect 26563 25248 26608 25276
rect 26602 25236 26608 25248
rect 26660 25236 26666 25288
rect 26694 25236 26700 25288
rect 26752 25276 26758 25288
rect 26973 25279 27031 25285
rect 26973 25276 26985 25279
rect 26752 25248 26985 25276
rect 26752 25236 26758 25248
rect 26973 25245 26985 25248
rect 27019 25245 27031 25279
rect 27522 25276 27528 25288
rect 27483 25248 27528 25276
rect 26973 25239 27031 25245
rect 27522 25236 27528 25248
rect 27580 25236 27586 25288
rect 28166 25276 28172 25288
rect 28127 25248 28172 25276
rect 28166 25236 28172 25248
rect 28224 25276 28230 25288
rect 28813 25279 28871 25285
rect 28813 25276 28825 25279
rect 28224 25248 28825 25276
rect 28224 25236 28230 25248
rect 28813 25245 28825 25248
rect 28859 25245 28871 25279
rect 33134 25276 33140 25288
rect 33095 25248 33140 25276
rect 28813 25239 28871 25245
rect 33134 25236 33140 25248
rect 33192 25236 33198 25288
rect 33594 25236 33600 25288
rect 33652 25276 33658 25288
rect 34072 25285 34100 25384
rect 35802 25372 35808 25384
rect 35860 25372 35866 25424
rect 39209 25415 39267 25421
rect 39209 25381 39221 25415
rect 39255 25412 39267 25415
rect 40126 25412 40132 25424
rect 39255 25384 40132 25412
rect 39255 25381 39267 25384
rect 39209 25375 39267 25381
rect 40126 25372 40132 25384
rect 40184 25372 40190 25424
rect 34698 25304 34704 25356
rect 34756 25344 34762 25356
rect 52748 25344 52776 25443
rect 54202 25440 54208 25452
rect 54260 25440 54266 25492
rect 34756 25316 35940 25344
rect 52748 25316 54064 25344
rect 34756 25304 34762 25316
rect 33781 25279 33839 25285
rect 33781 25276 33793 25279
rect 33652 25248 33793 25276
rect 33652 25236 33658 25248
rect 33781 25245 33793 25248
rect 33827 25245 33839 25279
rect 33781 25239 33839 25245
rect 34057 25279 34115 25285
rect 34057 25245 34069 25279
rect 34103 25245 34115 25279
rect 34057 25239 34115 25245
rect 34149 25279 34207 25285
rect 34149 25245 34161 25279
rect 34195 25276 34207 25279
rect 34330 25276 34336 25288
rect 34195 25248 34336 25276
rect 34195 25245 34207 25248
rect 34149 25239 34207 25245
rect 13446 25208 13452 25220
rect 1780 25180 13452 25208
rect 1780 25149 1808 25180
rect 13446 25168 13452 25180
rect 13504 25168 13510 25220
rect 27540 25208 27568 25236
rect 28534 25208 28540 25220
rect 27540 25180 28540 25208
rect 28534 25168 28540 25180
rect 28592 25208 28598 25220
rect 28629 25211 28687 25217
rect 28629 25208 28641 25211
rect 28592 25180 28641 25208
rect 28592 25168 28598 25180
rect 28629 25177 28641 25180
rect 28675 25177 28687 25211
rect 28629 25171 28687 25177
rect 31389 25211 31447 25217
rect 31389 25177 31401 25211
rect 31435 25208 31447 25211
rect 32582 25208 32588 25220
rect 31435 25180 32588 25208
rect 31435 25177 31447 25180
rect 31389 25171 31447 25177
rect 32582 25168 32588 25180
rect 32640 25168 32646 25220
rect 33962 25208 33968 25220
rect 33923 25180 33968 25208
rect 33962 25168 33968 25180
rect 34020 25168 34026 25220
rect 1765 25143 1823 25149
rect 1765 25109 1777 25143
rect 1811 25109 1823 25143
rect 25038 25140 25044 25152
rect 24999 25112 25044 25140
rect 1765 25103 1823 25109
rect 25038 25100 25044 25112
rect 25096 25100 25102 25152
rect 25866 25140 25872 25152
rect 25827 25112 25872 25140
rect 25866 25100 25872 25112
rect 25924 25100 25930 25152
rect 26605 25143 26663 25149
rect 26605 25109 26617 25143
rect 26651 25140 26663 25143
rect 26786 25140 26792 25152
rect 26651 25112 26792 25140
rect 26651 25109 26663 25112
rect 26605 25103 26663 25109
rect 26786 25100 26792 25112
rect 26844 25100 26850 25152
rect 33318 25140 33324 25152
rect 33279 25112 33324 25140
rect 33318 25100 33324 25112
rect 33376 25100 33382 25152
rect 33870 25100 33876 25152
rect 33928 25140 33934 25152
rect 34164 25140 34192 25239
rect 34330 25236 34336 25248
rect 34388 25236 34394 25288
rect 34422 25236 34428 25288
rect 34480 25276 34486 25288
rect 34974 25276 34980 25288
rect 34480 25248 34980 25276
rect 34480 25236 34486 25248
rect 34974 25236 34980 25248
rect 35032 25236 35038 25288
rect 35912 25285 35940 25316
rect 35069 25279 35127 25285
rect 35069 25245 35081 25279
rect 35115 25245 35127 25279
rect 35069 25239 35127 25245
rect 35897 25279 35955 25285
rect 35897 25245 35909 25279
rect 35943 25245 35955 25279
rect 35897 25239 35955 25245
rect 36357 25279 36415 25285
rect 36357 25245 36369 25279
rect 36403 25245 36415 25279
rect 38378 25276 38384 25288
rect 38339 25248 38384 25276
rect 36357 25239 36415 25245
rect 35084 25208 35112 25239
rect 36372 25208 36400 25239
rect 38378 25236 38384 25248
rect 38436 25236 38442 25288
rect 39025 25279 39083 25285
rect 39025 25245 39037 25279
rect 39071 25276 39083 25279
rect 39758 25276 39764 25288
rect 39071 25248 39764 25276
rect 39071 25245 39083 25248
rect 39025 25239 39083 25245
rect 39758 25236 39764 25248
rect 39816 25236 39822 25288
rect 41414 25236 41420 25288
rect 41472 25276 41478 25288
rect 54036 25285 54064 25316
rect 53285 25279 53343 25285
rect 53285 25276 53297 25279
rect 41472 25248 53297 25276
rect 41472 25236 41478 25248
rect 53285 25245 53297 25248
rect 53331 25245 53343 25279
rect 53285 25239 53343 25245
rect 54021 25279 54079 25285
rect 54021 25245 54033 25279
rect 54067 25245 54079 25279
rect 54021 25239 54079 25245
rect 34348 25180 35112 25208
rect 35820 25180 36400 25208
rect 34348 25149 34376 25180
rect 35820 25152 35848 25180
rect 38194 25168 38200 25220
rect 38252 25208 38258 25220
rect 40037 25211 40095 25217
rect 40037 25208 40049 25211
rect 38252 25180 40049 25208
rect 38252 25168 38258 25180
rect 40037 25177 40049 25180
rect 40083 25177 40095 25211
rect 40037 25171 40095 25177
rect 33928 25112 34192 25140
rect 34333 25143 34391 25149
rect 33928 25100 33934 25112
rect 34333 25109 34345 25143
rect 34379 25109 34391 25143
rect 35710 25140 35716 25152
rect 35671 25112 35716 25140
rect 34333 25103 34391 25109
rect 35710 25100 35716 25112
rect 35768 25100 35774 25152
rect 35802 25100 35808 25152
rect 35860 25100 35866 25152
rect 36541 25143 36599 25149
rect 36541 25109 36553 25143
rect 36587 25140 36599 25143
rect 36814 25140 36820 25152
rect 36587 25112 36820 25140
rect 36587 25109 36599 25112
rect 36541 25103 36599 25109
rect 36814 25100 36820 25112
rect 36872 25100 36878 25152
rect 37093 25143 37151 25149
rect 37093 25109 37105 25143
rect 37139 25140 37151 25143
rect 37826 25140 37832 25152
rect 37139 25112 37832 25140
rect 37139 25109 37151 25112
rect 37093 25103 37151 25109
rect 37826 25100 37832 25112
rect 37884 25100 37890 25152
rect 38565 25143 38623 25149
rect 38565 25109 38577 25143
rect 38611 25140 38623 25143
rect 38654 25140 38660 25152
rect 38611 25112 38660 25140
rect 38611 25109 38623 25112
rect 38565 25103 38623 25109
rect 38654 25100 38660 25112
rect 38712 25100 38718 25152
rect 53466 25140 53472 25152
rect 53427 25112 53472 25140
rect 53466 25100 53472 25112
rect 53524 25100 53530 25152
rect 1104 25050 54832 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 54832 25050
rect 1104 24976 54832 24998
rect 26421 24939 26479 24945
rect 26421 24905 26433 24939
rect 26467 24936 26479 24939
rect 26602 24936 26608 24948
rect 26467 24908 26608 24936
rect 26467 24905 26479 24908
rect 26421 24899 26479 24905
rect 26602 24896 26608 24908
rect 26660 24896 26666 24948
rect 28534 24936 28540 24948
rect 28495 24908 28540 24936
rect 28534 24896 28540 24908
rect 28592 24896 28598 24948
rect 31481 24939 31539 24945
rect 31481 24905 31493 24939
rect 31527 24936 31539 24939
rect 31938 24936 31944 24948
rect 31527 24908 31944 24936
rect 31527 24905 31539 24908
rect 31481 24899 31539 24905
rect 31938 24896 31944 24908
rect 31996 24896 32002 24948
rect 33134 24936 33140 24948
rect 33095 24908 33140 24936
rect 33134 24896 33140 24908
rect 33192 24896 33198 24948
rect 34977 24939 35035 24945
rect 34977 24905 34989 24939
rect 35023 24936 35035 24939
rect 35526 24936 35532 24948
rect 35023 24908 35532 24936
rect 35023 24905 35035 24908
rect 34977 24899 35035 24905
rect 25038 24828 25044 24880
rect 25096 24868 25102 24880
rect 25286 24871 25344 24877
rect 25286 24868 25298 24871
rect 25096 24840 25298 24868
rect 25096 24828 25102 24840
rect 25286 24837 25298 24840
rect 25332 24837 25344 24871
rect 25286 24831 25344 24837
rect 33318 24828 33324 24880
rect 33376 24868 33382 24880
rect 33842 24871 33900 24877
rect 33842 24868 33854 24871
rect 33376 24840 33854 24868
rect 33376 24828 33382 24840
rect 33842 24837 33854 24840
rect 33888 24837 33900 24871
rect 33842 24831 33900 24837
rect 1670 24800 1676 24812
rect 1631 24772 1676 24800
rect 1670 24760 1676 24772
rect 1728 24800 1734 24812
rect 2317 24803 2375 24809
rect 2317 24800 2329 24803
rect 1728 24772 2329 24800
rect 1728 24760 1734 24772
rect 2317 24769 2329 24772
rect 2363 24769 2375 24803
rect 2317 24763 2375 24769
rect 24397 24803 24455 24809
rect 24397 24769 24409 24803
rect 24443 24769 24455 24803
rect 27413 24803 27471 24809
rect 27413 24800 27425 24803
rect 24397 24763 24455 24769
rect 24596 24772 27425 24800
rect 1765 24599 1823 24605
rect 1765 24565 1777 24599
rect 1811 24596 1823 24599
rect 4062 24596 4068 24608
rect 1811 24568 4068 24596
rect 1811 24565 1823 24568
rect 1765 24559 1823 24565
rect 4062 24556 4068 24568
rect 4120 24556 4126 24608
rect 23937 24599 23995 24605
rect 23937 24565 23949 24599
rect 23983 24596 23995 24599
rect 24302 24596 24308 24608
rect 23983 24568 24308 24596
rect 23983 24565 23995 24568
rect 23937 24559 23995 24565
rect 24302 24556 24308 24568
rect 24360 24556 24366 24608
rect 24412 24596 24440 24763
rect 24596 24673 24624 24772
rect 27413 24769 27425 24772
rect 27459 24769 27471 24803
rect 27413 24763 27471 24769
rect 28166 24760 28172 24812
rect 28224 24800 28230 24812
rect 29181 24803 29239 24809
rect 29181 24800 29193 24803
rect 28224 24772 29193 24800
rect 28224 24760 28230 24772
rect 29181 24769 29193 24772
rect 29227 24769 29239 24803
rect 29181 24763 29239 24769
rect 30745 24803 30803 24809
rect 30745 24769 30757 24803
rect 30791 24800 30803 24803
rect 30926 24800 30932 24812
rect 30791 24772 30932 24800
rect 30791 24769 30803 24772
rect 30745 24763 30803 24769
rect 30926 24760 30932 24772
rect 30984 24760 30990 24812
rect 32858 24800 32864 24812
rect 32819 24772 32864 24800
rect 32858 24760 32864 24772
rect 32916 24760 32922 24812
rect 32953 24803 33011 24809
rect 32953 24769 32965 24803
rect 32999 24800 33011 24803
rect 33686 24800 33692 24812
rect 32999 24772 33692 24800
rect 32999 24769 33011 24772
rect 32953 24763 33011 24769
rect 33686 24760 33692 24772
rect 33744 24760 33750 24812
rect 34146 24760 34152 24812
rect 34204 24800 34210 24812
rect 34992 24800 35020 24899
rect 35526 24896 35532 24908
rect 35584 24896 35590 24948
rect 35710 24877 35716 24880
rect 35704 24868 35716 24877
rect 35671 24840 35716 24868
rect 35704 24831 35716 24840
rect 35710 24828 35716 24831
rect 35768 24828 35774 24880
rect 36262 24828 36268 24880
rect 36320 24868 36326 24880
rect 36320 24840 38792 24868
rect 36320 24828 36326 24840
rect 37734 24800 37740 24812
rect 34204 24772 35020 24800
rect 37695 24772 37740 24800
rect 34204 24760 34210 24772
rect 37734 24760 37740 24772
rect 37792 24760 37798 24812
rect 38654 24809 38660 24812
rect 38648 24800 38660 24809
rect 38615 24772 38660 24800
rect 38648 24763 38660 24772
rect 38654 24760 38660 24763
rect 38712 24760 38718 24812
rect 38764 24800 38792 24840
rect 40402 24800 40408 24812
rect 38764 24772 39436 24800
rect 40363 24772 40408 24800
rect 25038 24732 25044 24744
rect 24999 24704 25044 24732
rect 25038 24692 25044 24704
rect 25096 24692 25102 24744
rect 26878 24692 26884 24744
rect 26936 24732 26942 24744
rect 27157 24735 27215 24741
rect 27157 24732 27169 24735
rect 26936 24704 27169 24732
rect 26936 24692 26942 24704
rect 27157 24701 27169 24704
rect 27203 24701 27215 24735
rect 33594 24732 33600 24744
rect 33555 24704 33600 24732
rect 27157 24695 27215 24701
rect 33594 24692 33600 24704
rect 33652 24692 33658 24744
rect 35437 24735 35495 24741
rect 35437 24732 35449 24735
rect 34900 24704 35449 24732
rect 24581 24667 24639 24673
rect 24581 24633 24593 24667
rect 24627 24633 24639 24667
rect 24581 24627 24639 24633
rect 25774 24596 25780 24608
rect 24412 24568 25780 24596
rect 25774 24556 25780 24568
rect 25832 24556 25838 24608
rect 26418 24556 26424 24608
rect 26476 24596 26482 24608
rect 29089 24599 29147 24605
rect 29089 24596 29101 24599
rect 26476 24568 29101 24596
rect 26476 24556 26482 24568
rect 29089 24565 29101 24568
rect 29135 24565 29147 24599
rect 29089 24559 29147 24565
rect 30929 24599 30987 24605
rect 30929 24565 30941 24599
rect 30975 24596 30987 24599
rect 31294 24596 31300 24608
rect 30975 24568 31300 24596
rect 30975 24565 30987 24568
rect 30929 24559 30987 24565
rect 31294 24556 31300 24568
rect 31352 24556 31358 24608
rect 33594 24556 33600 24608
rect 33652 24596 33658 24608
rect 34900 24596 34928 24704
rect 35437 24701 35449 24704
rect 35483 24701 35495 24735
rect 35437 24695 35495 24701
rect 38286 24692 38292 24744
rect 38344 24732 38350 24744
rect 38381 24735 38439 24741
rect 38381 24732 38393 24735
rect 38344 24704 38393 24732
rect 38344 24692 38350 24704
rect 38381 24701 38393 24704
rect 38427 24701 38439 24735
rect 39408 24732 39436 24772
rect 40402 24760 40408 24772
rect 40460 24760 40466 24812
rect 42058 24760 42064 24812
rect 42116 24800 42122 24812
rect 53285 24803 53343 24809
rect 53285 24800 53297 24803
rect 42116 24772 53297 24800
rect 42116 24760 42122 24772
rect 53285 24769 53297 24772
rect 53331 24769 53343 24803
rect 53285 24763 53343 24769
rect 53558 24760 53564 24812
rect 53616 24800 53622 24812
rect 54205 24803 54263 24809
rect 54205 24800 54217 24803
rect 53616 24772 54217 24800
rect 53616 24760 53622 24772
rect 54205 24769 54217 24772
rect 54251 24769 54263 24803
rect 54205 24763 54263 24769
rect 42886 24732 42892 24744
rect 39408 24704 42892 24732
rect 38381 24695 38439 24701
rect 42886 24692 42892 24704
rect 42944 24732 42950 24744
rect 44082 24732 44088 24744
rect 42944 24704 44088 24732
rect 42944 24692 42950 24704
rect 44082 24692 44088 24704
rect 44140 24692 44146 24744
rect 36817 24667 36875 24673
rect 36817 24633 36829 24667
rect 36863 24664 36875 24667
rect 37274 24664 37280 24676
rect 36863 24636 37280 24664
rect 36863 24633 36875 24636
rect 36817 24627 36875 24633
rect 37274 24624 37280 24636
rect 37332 24664 37338 24676
rect 37642 24664 37648 24676
rect 37332 24636 37648 24664
rect 37332 24624 37338 24636
rect 37642 24624 37648 24636
rect 37700 24624 37706 24676
rect 37752 24636 38056 24664
rect 33652 24568 34928 24596
rect 33652 24556 33658 24568
rect 34974 24556 34980 24608
rect 35032 24596 35038 24608
rect 35618 24596 35624 24608
rect 35032 24568 35624 24596
rect 35032 24556 35038 24568
rect 35618 24556 35624 24568
rect 35676 24556 35682 24608
rect 35710 24556 35716 24608
rect 35768 24596 35774 24608
rect 37752 24596 37780 24636
rect 37918 24596 37924 24608
rect 35768 24568 37780 24596
rect 37879 24568 37924 24596
rect 35768 24556 35774 24568
rect 37918 24556 37924 24568
rect 37976 24556 37982 24608
rect 38028 24596 38056 24636
rect 49878 24624 49884 24676
rect 49936 24664 49942 24676
rect 54021 24667 54079 24673
rect 54021 24664 54033 24667
rect 49936 24636 54033 24664
rect 49936 24624 49942 24636
rect 54021 24633 54033 24636
rect 54067 24633 54079 24667
rect 54021 24627 54079 24633
rect 38562 24596 38568 24608
rect 38028 24568 38568 24596
rect 38562 24556 38568 24568
rect 38620 24556 38626 24608
rect 39022 24556 39028 24608
rect 39080 24596 39086 24608
rect 39761 24599 39819 24605
rect 39761 24596 39773 24599
rect 39080 24568 39773 24596
rect 39080 24556 39086 24568
rect 39761 24565 39773 24568
rect 39807 24565 39819 24599
rect 40586 24596 40592 24608
rect 40547 24568 40592 24596
rect 39761 24559 39819 24565
rect 40586 24556 40592 24568
rect 40644 24556 40650 24608
rect 53466 24596 53472 24608
rect 53427 24568 53472 24596
rect 53466 24556 53472 24568
rect 53524 24556 53530 24608
rect 1104 24506 54832 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 54832 24506
rect 1104 24432 54832 24454
rect 14642 24392 14648 24404
rect 14603 24364 14648 24392
rect 14642 24352 14648 24364
rect 14700 24352 14706 24404
rect 15102 24352 15108 24404
rect 15160 24392 15166 24404
rect 15197 24395 15255 24401
rect 15197 24392 15209 24395
rect 15160 24364 15209 24392
rect 15160 24352 15166 24364
rect 15197 24361 15209 24364
rect 15243 24361 15255 24395
rect 15197 24355 15255 24361
rect 24029 24395 24087 24401
rect 24029 24361 24041 24395
rect 24075 24392 24087 24395
rect 24578 24392 24584 24404
rect 24075 24364 24584 24392
rect 24075 24361 24087 24364
rect 24029 24355 24087 24361
rect 24578 24352 24584 24364
rect 24636 24352 24642 24404
rect 25682 24392 25688 24404
rect 24872 24364 25688 24392
rect 23109 24259 23167 24265
rect 23109 24225 23121 24259
rect 23155 24256 23167 24259
rect 23382 24256 23388 24268
rect 23155 24228 23388 24256
rect 23155 24225 23167 24228
rect 23109 24219 23167 24225
rect 23382 24216 23388 24228
rect 23440 24256 23446 24268
rect 23845 24259 23903 24265
rect 23845 24256 23857 24259
rect 23440 24228 23857 24256
rect 23440 24216 23446 24228
rect 23845 24225 23857 24228
rect 23891 24225 23903 24259
rect 23845 24219 23903 24225
rect 14737 24191 14795 24197
rect 14737 24157 14749 24191
rect 14783 24188 14795 24191
rect 15102 24188 15108 24200
rect 14783 24160 15108 24188
rect 14783 24157 14795 24160
rect 14737 24151 14795 24157
rect 15102 24148 15108 24160
rect 15160 24148 15166 24200
rect 23753 24191 23811 24197
rect 23753 24157 23765 24191
rect 23799 24188 23811 24191
rect 24872 24188 24900 24364
rect 25682 24352 25688 24364
rect 25740 24352 25746 24404
rect 26329 24395 26387 24401
rect 26329 24361 26341 24395
rect 26375 24392 26387 24395
rect 26694 24392 26700 24404
rect 26375 24364 26700 24392
rect 26375 24361 26387 24364
rect 26329 24355 26387 24361
rect 26694 24352 26700 24364
rect 26752 24352 26758 24404
rect 28166 24352 28172 24404
rect 28224 24392 28230 24404
rect 28261 24395 28319 24401
rect 28261 24392 28273 24395
rect 28224 24364 28273 24392
rect 28224 24352 28230 24364
rect 28261 24361 28273 24364
rect 28307 24361 28319 24395
rect 30926 24392 30932 24404
rect 30887 24364 30932 24392
rect 28261 24355 28319 24361
rect 30926 24352 30932 24364
rect 30984 24352 30990 24404
rect 33686 24392 33692 24404
rect 33647 24364 33692 24392
rect 33686 24352 33692 24364
rect 33744 24352 33750 24404
rect 33870 24352 33876 24404
rect 33928 24392 33934 24404
rect 34238 24392 34244 24404
rect 33928 24364 34244 24392
rect 33928 24352 33934 24364
rect 34238 24352 34244 24364
rect 34296 24352 34302 24404
rect 35894 24352 35900 24404
rect 35952 24392 35958 24404
rect 36265 24395 36323 24401
rect 36265 24392 36277 24395
rect 35952 24364 36277 24392
rect 35952 24352 35958 24364
rect 36265 24361 36277 24364
rect 36311 24361 36323 24395
rect 36265 24355 36323 24361
rect 37458 24352 37464 24404
rect 37516 24392 37522 24404
rect 37516 24364 37688 24392
rect 37516 24352 37522 24364
rect 31202 24324 31208 24336
rect 27908 24296 31208 24324
rect 23799 24160 24900 24188
rect 24949 24191 25007 24197
rect 23799 24157 23811 24160
rect 23753 24151 23811 24157
rect 24949 24157 24961 24191
rect 24995 24188 25007 24191
rect 25038 24188 25044 24200
rect 24995 24160 25044 24188
rect 24995 24157 25007 24160
rect 24949 24151 25007 24157
rect 25038 24148 25044 24160
rect 25096 24188 25102 24200
rect 26878 24188 26884 24200
rect 25096 24160 26884 24188
rect 25096 24148 25102 24160
rect 26878 24148 26884 24160
rect 26936 24148 26942 24200
rect 27908 24188 27936 24296
rect 31202 24284 31208 24296
rect 31260 24284 31266 24336
rect 34698 24324 34704 24336
rect 33060 24296 34704 24324
rect 29638 24216 29644 24268
rect 29696 24256 29702 24268
rect 30561 24259 30619 24265
rect 30561 24256 30573 24259
rect 29696 24228 30573 24256
rect 29696 24216 29702 24228
rect 30561 24225 30573 24228
rect 30607 24256 30619 24259
rect 31389 24259 31447 24265
rect 31389 24256 31401 24259
rect 30607 24228 31401 24256
rect 30607 24225 30619 24228
rect 30561 24219 30619 24225
rect 31389 24225 31401 24228
rect 31435 24256 31447 24259
rect 31938 24256 31944 24268
rect 31435 24228 31944 24256
rect 31435 24225 31447 24228
rect 31389 24219 31447 24225
rect 31938 24216 31944 24228
rect 31996 24256 32002 24268
rect 32861 24259 32919 24265
rect 32861 24256 32873 24259
rect 31996 24228 32873 24256
rect 31996 24216 32002 24228
rect 32861 24225 32873 24228
rect 32907 24225 32919 24259
rect 32861 24219 32919 24225
rect 26988 24160 27936 24188
rect 30745 24191 30803 24197
rect 1670 24120 1676 24132
rect 1631 24092 1676 24120
rect 1670 24080 1676 24092
rect 1728 24120 1734 24132
rect 25222 24129 25228 24132
rect 2317 24123 2375 24129
rect 2317 24120 2329 24123
rect 1728 24092 2329 24120
rect 1728 24080 1734 24092
rect 2317 24089 2329 24092
rect 2363 24089 2375 24123
rect 2317 24083 2375 24089
rect 24029 24123 24087 24129
rect 24029 24089 24041 24123
rect 24075 24089 24087 24123
rect 25216 24120 25228 24129
rect 25183 24092 25228 24120
rect 24029 24083 24087 24089
rect 25216 24083 25228 24092
rect 1762 24052 1768 24064
rect 1723 24024 1768 24052
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 14277 24055 14335 24061
rect 14277 24021 14289 24055
rect 14323 24052 14335 24055
rect 14458 24052 14464 24064
rect 14323 24024 14464 24052
rect 14323 24021 14335 24024
rect 14277 24015 14335 24021
rect 14458 24012 14464 24024
rect 14516 24012 14522 24064
rect 23566 24052 23572 24064
rect 23527 24024 23572 24052
rect 23566 24012 23572 24024
rect 23624 24012 23630 24064
rect 24044 24052 24072 24083
rect 25222 24080 25228 24083
rect 25280 24080 25286 24132
rect 25314 24080 25320 24132
rect 25372 24120 25378 24132
rect 26988 24120 27016 24160
rect 30745 24157 30757 24191
rect 30791 24157 30803 24191
rect 31570 24188 31576 24200
rect 31531 24160 31576 24188
rect 30745 24151 30803 24157
rect 27154 24129 27160 24132
rect 25372 24092 27016 24120
rect 25372 24080 25378 24092
rect 27148 24083 27160 24129
rect 27212 24120 27218 24132
rect 30760 24120 30788 24151
rect 31570 24148 31576 24160
rect 31628 24148 31634 24200
rect 33060 24197 33088 24296
rect 34698 24284 34704 24296
rect 34756 24284 34762 24336
rect 37660 24324 37688 24364
rect 37734 24352 37740 24404
rect 37792 24392 37798 24404
rect 38565 24395 38623 24401
rect 38565 24392 38577 24395
rect 37792 24364 38577 24392
rect 37792 24352 37798 24364
rect 38565 24361 38577 24364
rect 38611 24361 38623 24395
rect 38565 24355 38623 24361
rect 38746 24352 38752 24404
rect 38804 24392 38810 24404
rect 40310 24392 40316 24404
rect 38804 24364 40316 24392
rect 38804 24352 38810 24364
rect 40310 24352 40316 24364
rect 40368 24352 40374 24404
rect 41414 24352 41420 24404
rect 41472 24392 41478 24404
rect 53558 24392 53564 24404
rect 41472 24364 41517 24392
rect 53519 24364 53564 24392
rect 41472 24352 41478 24364
rect 53558 24352 53564 24364
rect 53616 24352 53622 24404
rect 38105 24327 38163 24333
rect 38105 24324 38117 24327
rect 37660 24296 38117 24324
rect 38105 24293 38117 24296
rect 38151 24293 38163 24327
rect 39393 24327 39451 24333
rect 39393 24324 39405 24327
rect 38105 24287 38163 24293
rect 38212 24296 39405 24324
rect 33594 24216 33600 24268
rect 33652 24256 33658 24268
rect 34885 24259 34943 24265
rect 34885 24256 34897 24259
rect 33652 24228 34897 24256
rect 33652 24216 33658 24228
rect 34885 24225 34897 24228
rect 34931 24225 34943 24259
rect 34885 24219 34943 24225
rect 31757 24191 31815 24197
rect 31757 24157 31769 24191
rect 31803 24188 31815 24191
rect 32401 24191 32459 24197
rect 32401 24188 32413 24191
rect 31803 24160 32413 24188
rect 31803 24157 31815 24160
rect 31757 24151 31815 24157
rect 32401 24157 32413 24160
rect 32447 24157 32459 24191
rect 32401 24151 32459 24157
rect 33045 24191 33103 24197
rect 33045 24157 33057 24191
rect 33091 24157 33103 24191
rect 33870 24188 33876 24200
rect 33831 24160 33876 24188
rect 33045 24151 33103 24157
rect 33870 24148 33876 24160
rect 33928 24148 33934 24200
rect 33965 24191 34023 24197
rect 33965 24157 33977 24191
rect 34011 24188 34023 24191
rect 34146 24188 34152 24200
rect 34011 24160 34152 24188
rect 34011 24157 34023 24160
rect 33965 24151 34023 24157
rect 34146 24148 34152 24160
rect 34204 24148 34210 24200
rect 34241 24191 34299 24197
rect 34241 24157 34253 24191
rect 34287 24188 34299 24191
rect 34606 24188 34612 24200
rect 34287 24160 34612 24188
rect 34287 24157 34299 24160
rect 34241 24151 34299 24157
rect 32306 24120 32312 24132
rect 27212 24092 27248 24120
rect 30760 24092 32312 24120
rect 27154 24080 27160 24083
rect 27212 24080 27218 24092
rect 32306 24080 32312 24092
rect 32364 24080 32370 24132
rect 34054 24080 34060 24132
rect 34112 24120 34118 24132
rect 34112 24092 34157 24120
rect 34112 24080 34118 24092
rect 26510 24052 26516 24064
rect 24044 24024 26516 24052
rect 26510 24012 26516 24024
rect 26568 24012 26574 24064
rect 30101 24055 30159 24061
rect 30101 24021 30113 24055
rect 30147 24052 30159 24055
rect 31386 24052 31392 24064
rect 30147 24024 31392 24052
rect 30147 24021 30159 24024
rect 30101 24015 30159 24021
rect 31386 24012 31392 24024
rect 31444 24012 31450 24064
rect 32214 24052 32220 24064
rect 32175 24024 32220 24052
rect 32214 24012 32220 24024
rect 32272 24012 32278 24064
rect 33226 24052 33232 24064
rect 33187 24024 33232 24052
rect 33226 24012 33232 24024
rect 33284 24012 33290 24064
rect 33870 24012 33876 24064
rect 33928 24052 33934 24064
rect 34256 24052 34284 24151
rect 34606 24148 34612 24160
rect 34664 24148 34670 24200
rect 34900 24188 34928 24219
rect 37826 24216 37832 24268
rect 37884 24256 37890 24268
rect 38212 24256 38240 24296
rect 39393 24293 39405 24296
rect 39439 24293 39451 24327
rect 39393 24287 39451 24293
rect 37884 24228 38240 24256
rect 37884 24216 37890 24228
rect 38286 24216 38292 24268
rect 38344 24256 38350 24268
rect 40034 24256 40040 24268
rect 38344 24228 40040 24256
rect 38344 24216 38350 24228
rect 40034 24216 40040 24228
rect 40092 24216 40098 24268
rect 36354 24188 36360 24200
rect 34900 24160 36360 24188
rect 36354 24148 36360 24160
rect 36412 24188 36418 24200
rect 36725 24191 36783 24197
rect 36725 24188 36737 24191
rect 36412 24160 36737 24188
rect 36412 24148 36418 24160
rect 36725 24157 36737 24160
rect 36771 24157 36783 24191
rect 36725 24151 36783 24157
rect 36814 24148 36820 24200
rect 36872 24188 36878 24200
rect 36981 24191 37039 24197
rect 36981 24188 36993 24191
rect 36872 24160 36993 24188
rect 36872 24148 36878 24160
rect 36981 24157 36993 24160
rect 37027 24157 37039 24191
rect 38746 24188 38752 24200
rect 38707 24160 38752 24188
rect 36981 24151 37039 24157
rect 38746 24148 38752 24160
rect 38804 24148 38810 24200
rect 38933 24191 38991 24197
rect 38933 24157 38945 24191
rect 38979 24157 38991 24191
rect 38933 24151 38991 24157
rect 35152 24123 35210 24129
rect 35152 24089 35164 24123
rect 35198 24120 35210 24123
rect 35342 24120 35348 24132
rect 35198 24092 35348 24120
rect 35198 24089 35210 24092
rect 35152 24083 35210 24089
rect 35342 24080 35348 24092
rect 35400 24080 35406 24132
rect 38948 24120 38976 24151
rect 40126 24148 40132 24200
rect 40184 24188 40190 24200
rect 40293 24191 40351 24197
rect 40293 24188 40305 24191
rect 40184 24160 40305 24188
rect 40184 24148 40190 24160
rect 40293 24157 40305 24160
rect 40339 24157 40351 24191
rect 40293 24151 40351 24157
rect 53009 24191 53067 24197
rect 53009 24157 53021 24191
rect 53055 24188 53067 24191
rect 54202 24188 54208 24200
rect 53055 24160 54208 24188
rect 53055 24157 53067 24160
rect 53009 24151 53067 24157
rect 54202 24148 54208 24160
rect 54260 24148 54266 24200
rect 38948 24092 40172 24120
rect 40144 24064 40172 24092
rect 44082 24080 44088 24132
rect 44140 24120 44146 24132
rect 52914 24120 52920 24132
rect 44140 24092 52920 24120
rect 44140 24080 44146 24092
rect 52914 24080 52920 24092
rect 52972 24080 52978 24132
rect 33928 24024 34284 24052
rect 33928 24012 33934 24024
rect 34330 24012 34336 24064
rect 34388 24052 34394 24064
rect 34790 24052 34796 24064
rect 34388 24024 34796 24052
rect 34388 24012 34394 24024
rect 34790 24012 34796 24024
rect 34848 24052 34854 24064
rect 39298 24052 39304 24064
rect 34848 24024 39304 24052
rect 34848 24012 34854 24024
rect 39298 24012 39304 24024
rect 39356 24012 39362 24064
rect 40126 24012 40132 24064
rect 40184 24012 40190 24064
rect 54110 24052 54116 24064
rect 54071 24024 54116 24052
rect 54110 24012 54116 24024
rect 54168 24012 54174 24064
rect 1104 23962 54832 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 54832 23962
rect 1104 23888 54832 23910
rect 4062 23808 4068 23860
rect 4120 23848 4126 23860
rect 24949 23851 25007 23857
rect 4120 23820 24440 23848
rect 4120 23808 4126 23820
rect 1762 23740 1768 23792
rect 1820 23780 1826 23792
rect 1820 23752 24164 23780
rect 1820 23740 1826 23752
rect 1857 23715 1915 23721
rect 1857 23681 1869 23715
rect 1903 23712 1915 23715
rect 22741 23715 22799 23721
rect 1903 23684 2452 23712
rect 1903 23681 1915 23684
rect 1857 23675 1915 23681
rect 2424 23585 2452 23684
rect 22741 23681 22753 23715
rect 22787 23712 22799 23715
rect 23658 23712 23664 23724
rect 22787 23684 23244 23712
rect 23619 23684 23664 23712
rect 22787 23681 22799 23684
rect 22741 23675 22799 23681
rect 23216 23653 23244 23684
rect 23658 23672 23664 23684
rect 23716 23672 23722 23724
rect 23201 23647 23259 23653
rect 23201 23613 23213 23647
rect 23247 23613 23259 23647
rect 23201 23607 23259 23613
rect 2409 23579 2467 23585
rect 2409 23545 2421 23579
rect 2455 23576 2467 23579
rect 22557 23579 22615 23585
rect 22557 23576 22569 23579
rect 2455 23548 22569 23576
rect 2455 23545 2467 23548
rect 2409 23539 2467 23545
rect 22557 23545 22569 23548
rect 22603 23545 22615 23579
rect 22557 23539 22615 23545
rect 1670 23508 1676 23520
rect 1631 23480 1676 23508
rect 1670 23468 1676 23480
rect 1728 23468 1734 23520
rect 14642 23468 14648 23520
rect 14700 23508 14706 23520
rect 14829 23511 14887 23517
rect 14829 23508 14841 23511
rect 14700 23480 14841 23508
rect 14700 23468 14706 23480
rect 14829 23477 14841 23480
rect 14875 23477 14887 23511
rect 14829 23471 14887 23477
rect 22097 23511 22155 23517
rect 22097 23477 22109 23511
rect 22143 23508 22155 23511
rect 23382 23508 23388 23520
rect 22143 23480 23388 23508
rect 22143 23477 22155 23480
rect 22097 23471 22155 23477
rect 23382 23468 23388 23480
rect 23440 23468 23446 23520
rect 24136 23508 24164 23752
rect 24412 23712 24440 23820
rect 24949 23817 24961 23851
rect 24995 23848 25007 23851
rect 25406 23848 25412 23860
rect 24995 23820 25412 23848
rect 24995 23817 25007 23820
rect 24949 23811 25007 23817
rect 25406 23808 25412 23820
rect 25464 23808 25470 23860
rect 26418 23808 26424 23860
rect 26476 23848 26482 23860
rect 27525 23851 27583 23857
rect 27525 23848 27537 23851
rect 26476 23820 27537 23848
rect 26476 23808 26482 23820
rect 27525 23817 27537 23820
rect 27571 23817 27583 23851
rect 27525 23811 27583 23817
rect 31202 23808 31208 23860
rect 31260 23848 31266 23860
rect 31754 23848 31760 23860
rect 31260 23820 31760 23848
rect 31260 23808 31266 23820
rect 31754 23808 31760 23820
rect 31812 23808 31818 23860
rect 31938 23808 31944 23860
rect 31996 23848 32002 23860
rect 32398 23848 32404 23860
rect 31996 23820 32404 23848
rect 31996 23808 32002 23820
rect 32398 23808 32404 23820
rect 32456 23848 32462 23860
rect 32585 23851 32643 23857
rect 32585 23848 32597 23851
rect 32456 23820 32597 23848
rect 32456 23808 32462 23820
rect 32585 23817 32597 23820
rect 32631 23817 32643 23851
rect 32585 23811 32643 23817
rect 34425 23851 34483 23857
rect 34425 23817 34437 23851
rect 34471 23848 34483 23851
rect 34514 23848 34520 23860
rect 34471 23820 34520 23848
rect 34471 23817 34483 23820
rect 34425 23811 34483 23817
rect 34514 23808 34520 23820
rect 34572 23808 34578 23860
rect 35713 23851 35771 23857
rect 35713 23817 35725 23851
rect 35759 23848 35771 23851
rect 35802 23848 35808 23860
rect 35759 23820 35808 23848
rect 35759 23817 35771 23820
rect 35713 23811 35771 23817
rect 35802 23808 35808 23820
rect 35860 23808 35866 23860
rect 37458 23848 37464 23860
rect 36464 23820 37464 23848
rect 24578 23780 24584 23792
rect 24491 23752 24584 23780
rect 24578 23740 24584 23752
rect 24636 23780 24642 23792
rect 26326 23780 26332 23792
rect 24636 23752 26332 23780
rect 24636 23740 24642 23752
rect 26326 23740 26332 23752
rect 26384 23740 26390 23792
rect 36464 23789 36492 23820
rect 37458 23808 37464 23820
rect 37516 23808 37522 23860
rect 37829 23851 37887 23857
rect 37829 23817 37841 23851
rect 37875 23848 37887 23851
rect 38378 23848 38384 23860
rect 37875 23820 38384 23848
rect 37875 23817 37887 23820
rect 37829 23811 37887 23817
rect 38378 23808 38384 23820
rect 38436 23808 38442 23860
rect 39298 23808 39304 23860
rect 39356 23848 39362 23860
rect 40221 23851 40279 23857
rect 40221 23848 40233 23851
rect 39356 23820 40233 23848
rect 39356 23808 39362 23820
rect 40221 23817 40233 23820
rect 40267 23817 40279 23851
rect 40221 23811 40279 23817
rect 40310 23808 40316 23860
rect 40368 23848 40374 23860
rect 54018 23848 54024 23860
rect 40368 23820 54024 23848
rect 40368 23808 40374 23820
rect 54018 23808 54024 23820
rect 54076 23808 54082 23860
rect 36449 23783 36507 23789
rect 29472 23752 31524 23780
rect 25314 23712 25320 23724
rect 24412 23684 25320 23712
rect 25314 23672 25320 23684
rect 25372 23672 25378 23724
rect 25685 23715 25743 23721
rect 25685 23681 25697 23715
rect 25731 23712 25743 23715
rect 25866 23712 25872 23724
rect 25731 23684 25872 23712
rect 25731 23681 25743 23684
rect 25685 23675 25743 23681
rect 25866 23672 25872 23684
rect 25924 23672 25930 23724
rect 26145 23715 26203 23721
rect 26145 23681 26157 23715
rect 26191 23712 26203 23715
rect 27246 23712 27252 23724
rect 26191 23684 27252 23712
rect 26191 23681 26203 23684
rect 26145 23675 26203 23681
rect 27246 23672 27252 23684
rect 27304 23672 27310 23724
rect 24302 23644 24308 23656
rect 24263 23616 24308 23644
rect 24302 23604 24308 23616
rect 24360 23604 24366 23656
rect 24489 23647 24547 23653
rect 24489 23613 24501 23647
rect 24535 23644 24547 23647
rect 25406 23644 25412 23656
rect 24535 23616 25412 23644
rect 24535 23613 24547 23616
rect 24489 23607 24547 23613
rect 25406 23604 25412 23616
rect 25464 23604 25470 23656
rect 25498 23604 25504 23656
rect 25556 23644 25562 23656
rect 26329 23647 26387 23653
rect 26329 23644 26341 23647
rect 25556 23616 26341 23644
rect 25556 23604 25562 23616
rect 26329 23613 26341 23616
rect 26375 23613 26387 23647
rect 26329 23607 26387 23613
rect 26970 23604 26976 23656
rect 27028 23644 27034 23656
rect 27617 23647 27675 23653
rect 27617 23644 27629 23647
rect 27028 23616 27629 23644
rect 27028 23604 27034 23616
rect 27617 23613 27629 23616
rect 27663 23613 27675 23647
rect 27617 23607 27675 23613
rect 27706 23604 27712 23656
rect 27764 23644 27770 23656
rect 28353 23647 28411 23653
rect 28353 23644 28365 23647
rect 27764 23616 28365 23644
rect 27764 23604 27770 23616
rect 28353 23613 28365 23616
rect 28399 23613 28411 23647
rect 28353 23607 28411 23613
rect 24394 23536 24400 23588
rect 24452 23576 24458 23588
rect 25593 23579 25651 23585
rect 25593 23576 25605 23579
rect 24452 23548 25605 23576
rect 24452 23536 24458 23548
rect 25593 23545 25605 23548
rect 25639 23545 25651 23579
rect 25593 23539 25651 23545
rect 25700 23548 27384 23576
rect 25700 23508 25728 23548
rect 24136 23480 25728 23508
rect 27157 23511 27215 23517
rect 27157 23477 27169 23511
rect 27203 23508 27215 23511
rect 27246 23508 27252 23520
rect 27203 23480 27252 23508
rect 27203 23477 27215 23480
rect 27157 23471 27215 23477
rect 27246 23468 27252 23480
rect 27304 23468 27310 23520
rect 27356 23508 27384 23548
rect 27430 23536 27436 23588
rect 27488 23576 27494 23588
rect 29472 23585 29500 23752
rect 30006 23712 30012 23724
rect 29967 23684 30012 23712
rect 30006 23672 30012 23684
rect 30064 23672 30070 23724
rect 31113 23715 31171 23721
rect 31113 23681 31125 23715
rect 31159 23712 31171 23715
rect 31202 23712 31208 23724
rect 31159 23684 31208 23712
rect 31159 23681 31171 23684
rect 31113 23675 31171 23681
rect 31202 23672 31208 23684
rect 31260 23672 31266 23724
rect 31496 23644 31524 23752
rect 35452 23752 36400 23780
rect 31754 23672 31760 23724
rect 31812 23712 31818 23724
rect 32677 23715 32735 23721
rect 32677 23712 32689 23715
rect 31812 23684 32689 23712
rect 31812 23672 31818 23684
rect 32677 23681 32689 23684
rect 32723 23681 32735 23715
rect 32677 23675 32735 23681
rect 33873 23715 33931 23721
rect 33873 23681 33885 23715
rect 33919 23681 33931 23715
rect 34054 23712 34060 23724
rect 34015 23684 34060 23712
rect 33873 23675 33931 23681
rect 32122 23644 32128 23656
rect 31496 23616 32128 23644
rect 32122 23604 32128 23616
rect 32180 23604 32186 23656
rect 32398 23644 32404 23656
rect 32359 23616 32404 23644
rect 32398 23604 32404 23616
rect 32456 23604 32462 23656
rect 33888 23644 33916 23675
rect 34054 23672 34060 23684
rect 34112 23672 34118 23724
rect 34149 23715 34207 23721
rect 34149 23681 34161 23715
rect 34195 23681 34207 23715
rect 34149 23675 34207 23681
rect 34164 23644 34192 23675
rect 34238 23672 34244 23724
rect 34296 23712 34302 23724
rect 35452 23712 35480 23752
rect 34296 23684 35480 23712
rect 34296 23672 34302 23684
rect 35526 23672 35532 23724
rect 35584 23712 35590 23724
rect 36372 23721 36400 23752
rect 36449 23749 36461 23783
rect 36495 23749 36507 23783
rect 36449 23743 36507 23749
rect 36541 23783 36599 23789
rect 36541 23749 36553 23783
rect 36587 23780 36599 23783
rect 37734 23780 37740 23792
rect 36587 23752 37740 23780
rect 36587 23749 36599 23752
rect 36541 23743 36599 23749
rect 37734 23740 37740 23752
rect 37792 23740 37798 23792
rect 37918 23740 37924 23792
rect 37976 23780 37982 23792
rect 38534 23783 38592 23789
rect 38534 23780 38546 23783
rect 37976 23752 38546 23780
rect 37976 23740 37982 23752
rect 38534 23749 38546 23752
rect 38580 23749 38592 23783
rect 40126 23780 40132 23792
rect 38534 23743 38592 23749
rect 39408 23752 40132 23780
rect 36357 23715 36415 23721
rect 35584 23684 35629 23712
rect 35584 23672 35590 23684
rect 36357 23681 36369 23715
rect 36403 23681 36415 23715
rect 36722 23712 36728 23724
rect 36683 23684 36728 23712
rect 36357 23675 36415 23681
rect 36722 23672 36728 23684
rect 36780 23672 36786 23724
rect 37642 23712 37648 23724
rect 37603 23684 37648 23712
rect 37642 23672 37648 23684
rect 37700 23672 37706 23724
rect 38286 23712 38292 23724
rect 38247 23684 38292 23712
rect 38286 23672 38292 23684
rect 38344 23672 38350 23724
rect 39408 23712 39436 23752
rect 40126 23740 40132 23752
rect 40184 23740 40190 23792
rect 40586 23740 40592 23792
rect 40644 23780 40650 23792
rect 40926 23783 40984 23789
rect 40926 23780 40938 23783
rect 40644 23752 40938 23780
rect 40644 23740 40650 23752
rect 40926 23749 40938 23752
rect 40972 23749 40984 23783
rect 40926 23743 40984 23749
rect 43990 23740 43996 23792
rect 44048 23780 44054 23792
rect 54110 23780 54116 23792
rect 44048 23752 54116 23780
rect 44048 23740 44054 23752
rect 54110 23740 54116 23752
rect 54168 23740 54174 23792
rect 54202 23740 54208 23792
rect 54260 23780 54266 23792
rect 54260 23752 54305 23780
rect 54260 23740 54266 23752
rect 38396 23684 39436 23712
rect 35345 23647 35403 23653
rect 33888 23616 34008 23644
rect 34164 23616 34560 23644
rect 29457 23579 29515 23585
rect 29457 23576 29469 23579
rect 27488 23548 29469 23576
rect 27488 23536 27494 23548
rect 29457 23545 29469 23548
rect 29503 23545 29515 23579
rect 33980 23576 34008 23616
rect 34330 23576 34336 23588
rect 33980 23548 34336 23576
rect 29457 23539 29515 23545
rect 34330 23536 34336 23548
rect 34388 23536 34394 23588
rect 28902 23508 28908 23520
rect 27356 23480 28908 23508
rect 28902 23468 28908 23480
rect 28960 23468 28966 23520
rect 28997 23511 29055 23517
rect 28997 23477 29009 23511
rect 29043 23508 29055 23511
rect 29178 23508 29184 23520
rect 29043 23480 29184 23508
rect 29043 23477 29055 23480
rect 28997 23471 29055 23477
rect 29178 23468 29184 23480
rect 29236 23468 29242 23520
rect 30190 23508 30196 23520
rect 30151 23480 30196 23508
rect 30190 23468 30196 23480
rect 30248 23468 30254 23520
rect 30834 23508 30840 23520
rect 30795 23480 30840 23508
rect 30834 23468 30840 23480
rect 30892 23468 30898 23520
rect 33045 23511 33103 23517
rect 33045 23477 33057 23511
rect 33091 23508 33103 23511
rect 34422 23508 34428 23520
rect 33091 23480 34428 23508
rect 33091 23477 33103 23480
rect 33045 23471 33103 23477
rect 34422 23468 34428 23480
rect 34480 23468 34486 23520
rect 34532 23508 34560 23616
rect 35345 23613 35357 23647
rect 35391 23644 35403 23647
rect 35618 23644 35624 23656
rect 35391 23616 35624 23644
rect 35391 23613 35403 23616
rect 35345 23607 35403 23613
rect 35618 23604 35624 23616
rect 35676 23644 35682 23656
rect 37461 23647 37519 23653
rect 35676 23616 36308 23644
rect 35676 23604 35682 23616
rect 35526 23536 35532 23588
rect 35584 23576 35590 23588
rect 36173 23579 36231 23585
rect 36173 23576 36185 23579
rect 35584 23548 36185 23576
rect 35584 23536 35590 23548
rect 36173 23545 36185 23548
rect 36219 23545 36231 23579
rect 36280 23576 36308 23616
rect 37461 23613 37473 23647
rect 37507 23644 37519 23647
rect 38396 23644 38424 23684
rect 40034 23672 40040 23724
rect 40092 23712 40098 23724
rect 40678 23712 40684 23724
rect 40092 23684 40684 23712
rect 40092 23672 40098 23684
rect 40678 23672 40684 23684
rect 40736 23672 40742 23724
rect 42794 23712 42800 23724
rect 40788 23684 42800 23712
rect 40788 23644 40816 23684
rect 42794 23672 42800 23684
rect 42852 23712 42858 23724
rect 44082 23712 44088 23724
rect 42852 23684 44088 23712
rect 42852 23672 42858 23684
rect 44082 23672 44088 23684
rect 44140 23672 44146 23724
rect 53469 23715 53527 23721
rect 53469 23681 53481 23715
rect 53515 23712 53527 23715
rect 53558 23712 53564 23724
rect 53515 23684 53564 23712
rect 53515 23681 53527 23684
rect 53469 23675 53527 23681
rect 53558 23672 53564 23684
rect 53616 23672 53622 23724
rect 54220 23712 54248 23740
rect 53668 23684 54248 23712
rect 37507 23616 38424 23644
rect 39684 23616 40816 23644
rect 37507 23613 37519 23616
rect 37461 23607 37519 23613
rect 37826 23576 37832 23588
rect 36280 23548 37832 23576
rect 36173 23539 36231 23545
rect 37826 23536 37832 23548
rect 37884 23536 37890 23588
rect 37274 23508 37280 23520
rect 34532 23480 37280 23508
rect 37274 23468 37280 23480
rect 37332 23468 37338 23520
rect 38930 23468 38936 23520
rect 38988 23508 38994 23520
rect 39684 23517 39712 23616
rect 42058 23576 42064 23588
rect 42019 23548 42064 23576
rect 42058 23536 42064 23548
rect 42116 23536 42122 23588
rect 53282 23576 53288 23588
rect 53243 23548 53288 23576
rect 53282 23536 53288 23548
rect 53340 23536 53346 23588
rect 53466 23536 53472 23588
rect 53524 23576 53530 23588
rect 53668 23576 53696 23684
rect 54018 23644 54024 23656
rect 53979 23616 54024 23644
rect 54018 23604 54024 23616
rect 54076 23604 54082 23656
rect 53524 23548 53696 23576
rect 53524 23536 53530 23548
rect 39669 23511 39727 23517
rect 39669 23508 39681 23511
rect 38988 23480 39681 23508
rect 38988 23468 38994 23480
rect 39669 23477 39681 23480
rect 39715 23477 39727 23511
rect 39669 23471 39727 23477
rect 40310 23468 40316 23520
rect 40368 23508 40374 23520
rect 42076 23508 42104 23536
rect 40368 23480 42104 23508
rect 40368 23468 40374 23480
rect 1104 23418 54832 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 54832 23418
rect 1104 23344 54832 23366
rect 22557 23307 22615 23313
rect 22557 23273 22569 23307
rect 22603 23304 22615 23307
rect 22922 23304 22928 23316
rect 22603 23276 22928 23304
rect 22603 23273 22615 23276
rect 22557 23267 22615 23273
rect 22922 23264 22928 23276
rect 22980 23304 22986 23316
rect 23382 23304 23388 23316
rect 22980 23276 23388 23304
rect 22980 23264 22986 23276
rect 23382 23264 23388 23276
rect 23440 23304 23446 23316
rect 24029 23307 24087 23313
rect 24029 23304 24041 23307
rect 23440 23276 24041 23304
rect 23440 23264 23446 23276
rect 24029 23273 24041 23276
rect 24075 23304 24087 23307
rect 24765 23307 24823 23313
rect 24765 23304 24777 23307
rect 24075 23276 24777 23304
rect 24075 23273 24087 23276
rect 24029 23267 24087 23273
rect 24765 23273 24777 23276
rect 24811 23273 24823 23307
rect 24765 23267 24823 23273
rect 25774 23264 25780 23316
rect 25832 23304 25838 23316
rect 25869 23307 25927 23313
rect 25869 23304 25881 23307
rect 25832 23276 25881 23304
rect 25832 23264 25838 23276
rect 25869 23273 25881 23276
rect 25915 23273 25927 23307
rect 25869 23267 25927 23273
rect 27065 23307 27123 23313
rect 27065 23273 27077 23307
rect 27111 23304 27123 23307
rect 27154 23304 27160 23316
rect 27111 23276 27160 23304
rect 27111 23273 27123 23276
rect 27065 23267 27123 23273
rect 27154 23264 27160 23276
rect 27212 23264 27218 23316
rect 28902 23264 28908 23316
rect 28960 23304 28966 23316
rect 29086 23304 29092 23316
rect 28960 23276 29092 23304
rect 28960 23264 28966 23276
rect 29086 23264 29092 23276
rect 29144 23264 29150 23316
rect 30834 23264 30840 23316
rect 30892 23304 30898 23316
rect 32398 23304 32404 23316
rect 30892 23276 32404 23304
rect 30892 23264 30898 23276
rect 32398 23264 32404 23276
rect 32456 23264 32462 23316
rect 33778 23264 33784 23316
rect 33836 23304 33842 23316
rect 34054 23304 34060 23316
rect 33836 23276 34060 23304
rect 33836 23264 33842 23276
rect 34054 23264 34060 23276
rect 34112 23264 34118 23316
rect 34422 23264 34428 23316
rect 34480 23304 34486 23316
rect 34480 23276 37596 23304
rect 34480 23264 34486 23276
rect 35621 23239 35679 23245
rect 35621 23205 35633 23239
rect 35667 23236 35679 23239
rect 37568 23236 37596 23276
rect 37642 23264 37648 23316
rect 37700 23304 37706 23316
rect 38105 23307 38163 23313
rect 38105 23304 38117 23307
rect 37700 23276 38117 23304
rect 37700 23264 37706 23276
rect 38105 23273 38117 23276
rect 38151 23273 38163 23307
rect 38105 23267 38163 23273
rect 38194 23264 38200 23316
rect 38252 23304 38258 23316
rect 40402 23304 40408 23316
rect 38252 23276 39068 23304
rect 40363 23276 40408 23304
rect 38252 23264 38258 23276
rect 38654 23236 38660 23248
rect 35667 23208 35848 23236
rect 37568 23208 38660 23236
rect 35667 23205 35679 23208
rect 35621 23199 35679 23205
rect 23937 23171 23995 23177
rect 23937 23137 23949 23171
rect 23983 23168 23995 23171
rect 24578 23168 24584 23180
rect 23983 23140 24584 23168
rect 23983 23137 23995 23140
rect 23937 23131 23995 23137
rect 24578 23128 24584 23140
rect 24636 23128 24642 23180
rect 24857 23171 24915 23177
rect 24857 23137 24869 23171
rect 24903 23168 24915 23171
rect 25498 23168 25504 23180
rect 24903 23140 25504 23168
rect 24903 23137 24915 23140
rect 24857 23131 24915 23137
rect 25498 23128 25504 23140
rect 25556 23128 25562 23180
rect 26326 23128 26332 23180
rect 26384 23168 26390 23180
rect 26421 23171 26479 23177
rect 26421 23168 26433 23171
rect 26384 23140 26433 23168
rect 26384 23128 26390 23140
rect 26421 23137 26433 23140
rect 26467 23168 26479 23171
rect 27706 23168 27712 23180
rect 26467 23140 27712 23168
rect 26467 23137 26479 23140
rect 26421 23131 26479 23137
rect 27706 23128 27712 23140
rect 27764 23168 27770 23180
rect 28353 23171 28411 23177
rect 28353 23168 28365 23171
rect 27764 23140 28365 23168
rect 27764 23128 27770 23140
rect 28353 23137 28365 23140
rect 28399 23168 28411 23171
rect 28718 23168 28724 23180
rect 28399 23140 28724 23168
rect 28399 23137 28411 23140
rect 28353 23131 28411 23137
rect 28718 23128 28724 23140
rect 28776 23128 28782 23180
rect 33778 23168 33784 23180
rect 33739 23140 33784 23168
rect 33778 23128 33784 23140
rect 33836 23128 33842 23180
rect 34057 23171 34115 23177
rect 34057 23137 34069 23171
rect 34103 23137 34115 23171
rect 34974 23168 34980 23180
rect 34935 23140 34980 23168
rect 34057 23131 34115 23137
rect 1857 23103 1915 23109
rect 1857 23069 1869 23103
rect 1903 23100 1915 23103
rect 2314 23100 2320 23112
rect 1903 23072 2320 23100
rect 1903 23069 1915 23072
rect 1857 23063 1915 23069
rect 2314 23060 2320 23072
rect 2372 23060 2378 23112
rect 23201 23103 23259 23109
rect 23201 23069 23213 23103
rect 23247 23100 23259 23103
rect 23566 23100 23572 23112
rect 23247 23072 23572 23100
rect 23247 23069 23259 23072
rect 23201 23063 23259 23069
rect 23566 23060 23572 23072
rect 23624 23060 23630 23112
rect 24029 23103 24087 23109
rect 24029 23069 24041 23103
rect 24075 23069 24087 23103
rect 24029 23063 24087 23069
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23100 25007 23103
rect 25866 23100 25872 23112
rect 24995 23072 25872 23100
rect 24995 23069 25007 23072
rect 24949 23063 25007 23069
rect 24044 23032 24072 23063
rect 24964 23032 24992 23063
rect 25866 23060 25872 23072
rect 25924 23060 25930 23112
rect 26234 23100 26240 23112
rect 26195 23072 26240 23100
rect 26234 23060 26240 23072
rect 26292 23060 26298 23112
rect 27246 23100 27252 23112
rect 27207 23072 27252 23100
rect 27246 23060 27252 23072
rect 27304 23060 27310 23112
rect 29825 23103 29883 23109
rect 29825 23069 29837 23103
rect 29871 23100 29883 23103
rect 30374 23100 30380 23112
rect 29871 23072 30380 23100
rect 29871 23069 29883 23072
rect 29825 23063 29883 23069
rect 30374 23060 30380 23072
rect 30432 23100 30438 23112
rect 31665 23103 31723 23109
rect 31665 23100 31677 23103
rect 30432 23072 31677 23100
rect 30432 23060 30438 23072
rect 31665 23069 31677 23072
rect 31711 23100 31723 23103
rect 33594 23100 33600 23112
rect 31711 23072 33600 23100
rect 31711 23069 31723 23072
rect 31665 23063 31723 23069
rect 33594 23060 33600 23072
rect 33652 23060 33658 23112
rect 24044 23004 24992 23032
rect 30092 23035 30150 23041
rect 30092 23001 30104 23035
rect 30138 23032 30150 23035
rect 30190 23032 30196 23044
rect 30138 23004 30196 23032
rect 30138 23001 30150 23004
rect 30092 22995 30150 23001
rect 30190 22992 30196 23004
rect 30248 22992 30254 23044
rect 31294 22992 31300 23044
rect 31352 23032 31358 23044
rect 31910 23035 31968 23041
rect 31910 23032 31922 23035
rect 31352 23004 31922 23032
rect 31352 22992 31358 23004
rect 31910 23001 31922 23004
rect 31956 23001 31968 23035
rect 34072 23032 34100 23131
rect 34974 23128 34980 23140
rect 35032 23128 35038 23180
rect 35820 23168 35848 23208
rect 38654 23196 38660 23208
rect 38712 23196 38718 23248
rect 39040 23236 39068 23276
rect 40402 23264 40408 23276
rect 40460 23264 40466 23316
rect 43254 23304 43260 23316
rect 40512 23276 43260 23304
rect 40512 23236 40540 23276
rect 43254 23264 43260 23276
rect 43312 23264 43318 23316
rect 54202 23304 54208 23316
rect 54163 23276 54208 23304
rect 54202 23264 54208 23276
rect 54260 23264 54266 23316
rect 42334 23236 42340 23248
rect 39040 23208 40540 23236
rect 42247 23208 42340 23236
rect 35820 23140 37596 23168
rect 34149 23103 34207 23109
rect 34149 23069 34161 23103
rect 34195 23100 34207 23103
rect 36449 23103 36507 23109
rect 36449 23100 36461 23103
rect 34195 23072 36461 23100
rect 34195 23069 34207 23072
rect 34149 23063 34207 23069
rect 36449 23069 36461 23072
rect 36495 23069 36507 23103
rect 36449 23063 36507 23069
rect 37093 23103 37151 23109
rect 37093 23069 37105 23103
rect 37139 23100 37151 23103
rect 37458 23100 37464 23112
rect 37139 23072 37464 23100
rect 37139 23069 37151 23072
rect 37093 23063 37151 23069
rect 37458 23060 37464 23072
rect 37516 23060 37522 23112
rect 37568 23109 37596 23140
rect 37752 23140 38792 23168
rect 37752 23112 37780 23140
rect 37553 23103 37611 23109
rect 37553 23069 37565 23103
rect 37599 23069 37611 23103
rect 37734 23100 37740 23112
rect 37695 23072 37740 23100
rect 37553 23063 37611 23069
rect 37734 23060 37740 23072
rect 37792 23060 37798 23112
rect 37921 23103 37979 23109
rect 37921 23069 37933 23103
rect 37967 23100 37979 23103
rect 38010 23100 38016 23112
rect 37967 23072 38016 23100
rect 37967 23069 37979 23072
rect 37921 23063 37979 23069
rect 38010 23060 38016 23072
rect 38068 23060 38074 23112
rect 38562 23100 38568 23112
rect 38523 23072 38568 23100
rect 38562 23060 38568 23072
rect 38620 23060 38626 23112
rect 38764 23109 38792 23140
rect 38749 23103 38807 23109
rect 38749 23069 38761 23103
rect 38795 23069 38807 23103
rect 38749 23063 38807 23069
rect 38933 23103 38991 23109
rect 38933 23069 38945 23103
rect 38979 23100 38991 23103
rect 39040 23100 39068 23208
rect 42334 23196 42340 23208
rect 42392 23236 42398 23248
rect 53558 23236 53564 23248
rect 42392 23208 51074 23236
rect 53519 23208 53564 23236
rect 42392 23196 42398 23208
rect 40037 23171 40095 23177
rect 40037 23137 40049 23171
rect 40083 23168 40095 23171
rect 40126 23168 40132 23180
rect 40083 23140 40132 23168
rect 40083 23137 40095 23140
rect 40037 23131 40095 23137
rect 40126 23128 40132 23140
rect 40184 23128 40190 23180
rect 40678 23128 40684 23180
rect 40736 23168 40742 23180
rect 40957 23171 41015 23177
rect 40957 23168 40969 23171
rect 40736 23140 40969 23168
rect 40736 23128 40742 23140
rect 40957 23137 40969 23140
rect 41003 23137 41015 23171
rect 40957 23131 41015 23137
rect 40218 23100 40224 23112
rect 38979 23072 39068 23100
rect 40179 23072 40224 23100
rect 38979 23069 38991 23072
rect 38933 23063 38991 23069
rect 40218 23060 40224 23072
rect 40276 23060 40282 23112
rect 41506 23060 41512 23112
rect 41564 23100 41570 23112
rect 42981 23103 43039 23109
rect 42981 23100 42993 23103
rect 41564 23072 42993 23100
rect 41564 23060 41570 23072
rect 42981 23069 42993 23072
rect 43027 23069 43039 23103
rect 51046 23100 51074 23208
rect 53558 23196 53564 23208
rect 53616 23196 53622 23248
rect 54021 23103 54079 23109
rect 54021 23100 54033 23103
rect 51046 23072 54033 23100
rect 42981 23063 43039 23069
rect 54021 23069 54033 23072
rect 54067 23069 54079 23103
rect 54021 23063 54079 23069
rect 35986 23032 35992 23044
rect 34072 23004 35992 23032
rect 31910 22995 31968 23001
rect 35986 22992 35992 23004
rect 36044 22992 36050 23044
rect 37829 23035 37887 23041
rect 37829 23001 37841 23035
rect 37875 23001 37887 23035
rect 37829 22995 37887 23001
rect 38841 23035 38899 23041
rect 38841 23001 38853 23035
rect 38887 23032 38899 23035
rect 41224 23035 41282 23041
rect 38887 23004 40172 23032
rect 38887 23001 38899 23004
rect 38841 22995 38899 23001
rect 1670 22964 1676 22976
rect 1631 22936 1676 22964
rect 1670 22924 1676 22936
rect 1728 22924 1734 22976
rect 14642 22964 14648 22976
rect 14603 22936 14648 22964
rect 14642 22924 14648 22936
rect 14700 22924 14706 22976
rect 23014 22964 23020 22976
rect 22975 22936 23020 22964
rect 23014 22924 23020 22936
rect 23072 22924 23078 22976
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 23661 22967 23719 22973
rect 23661 22964 23673 22967
rect 23532 22936 23673 22964
rect 23532 22924 23538 22936
rect 23661 22933 23673 22936
rect 23707 22933 23719 22967
rect 23661 22927 23719 22933
rect 23750 22924 23756 22976
rect 23808 22964 23814 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 23808 22936 24593 22964
rect 23808 22924 23814 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 26329 22967 26387 22973
rect 26329 22933 26341 22967
rect 26375 22964 26387 22967
rect 26418 22964 26424 22976
rect 26375 22936 26424 22964
rect 26375 22933 26387 22936
rect 26329 22927 26387 22933
rect 26418 22924 26424 22936
rect 26476 22924 26482 22976
rect 27338 22924 27344 22976
rect 27396 22964 27402 22976
rect 27801 22967 27859 22973
rect 27801 22964 27813 22967
rect 27396 22936 27813 22964
rect 27396 22924 27402 22936
rect 27801 22933 27813 22936
rect 27847 22933 27859 22967
rect 31202 22964 31208 22976
rect 31163 22936 31208 22964
rect 27801 22927 27859 22933
rect 31202 22924 31208 22936
rect 31260 22924 31266 22976
rect 33045 22967 33103 22973
rect 33045 22933 33057 22967
rect 33091 22964 33103 22967
rect 33134 22964 33140 22976
rect 33091 22936 33140 22964
rect 33091 22933 33103 22936
rect 33045 22927 33103 22933
rect 33134 22924 33140 22936
rect 33192 22924 33198 22976
rect 35158 22964 35164 22976
rect 35119 22936 35164 22964
rect 35158 22924 35164 22936
rect 35216 22924 35222 22976
rect 35253 22967 35311 22973
rect 35253 22933 35265 22967
rect 35299 22964 35311 22967
rect 35802 22964 35808 22976
rect 35299 22936 35808 22964
rect 35299 22933 35311 22936
rect 35253 22927 35311 22933
rect 35802 22924 35808 22936
rect 35860 22924 35866 22976
rect 37844 22964 37872 22995
rect 39022 22964 39028 22976
rect 37844 22936 39028 22964
rect 39022 22924 39028 22936
rect 39080 22924 39086 22976
rect 39117 22967 39175 22973
rect 39117 22933 39129 22967
rect 39163 22964 39175 22967
rect 39942 22964 39948 22976
rect 39163 22936 39948 22964
rect 39163 22933 39175 22936
rect 39117 22927 39175 22933
rect 39942 22924 39948 22936
rect 40000 22924 40006 22976
rect 40144 22964 40172 23004
rect 41224 23001 41236 23035
rect 41270 23032 41282 23035
rect 41270 23004 42840 23032
rect 41270 23001 41282 23004
rect 41224 22995 41282 23001
rect 41414 22964 41420 22976
rect 40144 22936 41420 22964
rect 41414 22924 41420 22936
rect 41472 22924 41478 22976
rect 42812 22973 42840 23004
rect 42797 22967 42855 22973
rect 42797 22933 42809 22967
rect 42843 22933 42855 22967
rect 42797 22927 42855 22933
rect 1104 22874 54832 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 54832 22874
rect 1104 22800 54832 22822
rect 2314 22760 2320 22772
rect 2275 22732 2320 22760
rect 2314 22720 2320 22732
rect 2372 22720 2378 22772
rect 14921 22763 14979 22769
rect 14921 22760 14933 22763
rect 6886 22732 14933 22760
rect 1854 22624 1860 22636
rect 1815 22596 1860 22624
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 2501 22627 2559 22633
rect 2501 22593 2513 22627
rect 2547 22624 2559 22627
rect 6886 22624 6914 22732
rect 14921 22729 14933 22732
rect 14967 22729 14979 22763
rect 17218 22760 17224 22772
rect 14921 22723 14979 22729
rect 16546 22732 17224 22760
rect 14550 22652 14556 22704
rect 14608 22692 14614 22704
rect 14608 22664 15424 22692
rect 14608 22652 14614 22664
rect 2547 22596 6914 22624
rect 14461 22627 14519 22633
rect 2547 22593 2559 22596
rect 2501 22587 2559 22593
rect 14461 22593 14473 22627
rect 14507 22624 14519 22627
rect 14734 22624 14740 22636
rect 14507 22596 14740 22624
rect 14507 22593 14519 22596
rect 14461 22587 14519 22593
rect 14734 22584 14740 22596
rect 14792 22584 14798 22636
rect 15396 22633 15424 22664
rect 15381 22627 15439 22633
rect 15381 22593 15393 22627
rect 15427 22624 15439 22627
rect 15841 22627 15899 22633
rect 15841 22624 15853 22627
rect 15427 22596 15853 22624
rect 15427 22593 15439 22596
rect 15381 22587 15439 22593
rect 15841 22593 15853 22596
rect 15887 22624 15899 22627
rect 16546 22624 16574 22732
rect 17218 22720 17224 22732
rect 17276 22720 17282 22772
rect 22922 22760 22928 22772
rect 22883 22732 22928 22760
rect 22922 22720 22928 22732
rect 22980 22720 22986 22772
rect 24302 22720 24308 22772
rect 24360 22760 24366 22772
rect 24765 22763 24823 22769
rect 24765 22760 24777 22763
rect 24360 22732 24777 22760
rect 24360 22720 24366 22732
rect 24765 22729 24777 22732
rect 24811 22729 24823 22763
rect 24765 22723 24823 22729
rect 18782 22652 18788 22704
rect 18840 22692 18846 22704
rect 24780 22692 24808 22723
rect 24854 22720 24860 22772
rect 24912 22760 24918 22772
rect 25317 22763 25375 22769
rect 25317 22760 25329 22763
rect 24912 22732 25329 22760
rect 24912 22720 24918 22732
rect 25317 22729 25329 22732
rect 25363 22729 25375 22763
rect 25682 22760 25688 22772
rect 25643 22732 25688 22760
rect 25317 22723 25375 22729
rect 25682 22720 25688 22732
rect 25740 22720 25746 22772
rect 29917 22763 29975 22769
rect 29917 22729 29929 22763
rect 29963 22760 29975 22763
rect 30006 22760 30012 22772
rect 29963 22732 30012 22760
rect 29963 22729 29975 22732
rect 29917 22723 29975 22729
rect 30006 22720 30012 22732
rect 30064 22720 30070 22772
rect 31754 22720 31760 22772
rect 31812 22760 31818 22772
rect 32306 22760 32312 22772
rect 31812 22732 31857 22760
rect 32267 22732 32312 22760
rect 31812 22720 31818 22732
rect 32306 22720 32312 22732
rect 32364 22720 32370 22772
rect 32677 22763 32735 22769
rect 32677 22729 32689 22763
rect 32723 22760 32735 22763
rect 33134 22760 33140 22772
rect 32723 22732 33140 22760
rect 32723 22729 32735 22732
rect 32677 22723 32735 22729
rect 33134 22720 33140 22732
rect 33192 22760 33198 22772
rect 33318 22760 33324 22772
rect 33192 22732 33324 22760
rect 33192 22720 33198 22732
rect 33318 22720 33324 22732
rect 33376 22760 33382 22772
rect 33873 22763 33931 22769
rect 33873 22760 33885 22763
rect 33376 22732 33885 22760
rect 33376 22720 33382 22732
rect 33873 22729 33885 22732
rect 33919 22729 33931 22763
rect 35526 22760 35532 22772
rect 35487 22732 35532 22760
rect 33873 22723 33931 22729
rect 35526 22720 35532 22732
rect 35584 22720 35590 22772
rect 35989 22763 36047 22769
rect 35989 22729 36001 22763
rect 36035 22760 36047 22763
rect 36722 22760 36728 22772
rect 36035 22732 36728 22760
rect 36035 22729 36047 22732
rect 35989 22723 36047 22729
rect 36722 22720 36728 22732
rect 36780 22720 36786 22772
rect 37458 22720 37464 22772
rect 37516 22720 37522 22772
rect 37734 22760 37740 22772
rect 37660 22732 37740 22760
rect 26326 22692 26332 22704
rect 18840 22664 24624 22692
rect 24780 22664 26332 22692
rect 18840 22652 18846 22664
rect 23474 22624 23480 22636
rect 15887 22596 16574 22624
rect 23435 22596 23480 22624
rect 15887 22593 15899 22596
rect 15841 22587 15899 22593
rect 23474 22584 23480 22596
rect 23532 22584 23538 22636
rect 2590 22516 2596 22568
rect 2648 22556 2654 22568
rect 23753 22559 23811 22565
rect 23753 22556 23765 22559
rect 2648 22528 23765 22556
rect 2648 22516 2654 22528
rect 23753 22525 23765 22528
rect 23799 22525 23811 22559
rect 23753 22519 23811 22525
rect 1670 22420 1676 22432
rect 1631 22392 1676 22420
rect 1670 22380 1676 22392
rect 1728 22380 1734 22432
rect 14001 22423 14059 22429
rect 14001 22389 14013 22423
rect 14047 22420 14059 22423
rect 14090 22420 14096 22432
rect 14047 22392 14096 22420
rect 14047 22389 14059 22392
rect 14001 22383 14059 22389
rect 14090 22380 14096 22392
rect 14148 22380 14154 22432
rect 14369 22423 14427 22429
rect 14369 22389 14381 22423
rect 14415 22420 14427 22423
rect 14642 22420 14648 22432
rect 14415 22392 14648 22420
rect 14415 22389 14427 22392
rect 14369 22383 14427 22389
rect 14642 22380 14648 22392
rect 14700 22420 14706 22432
rect 15286 22420 15292 22432
rect 14700 22392 15292 22420
rect 14700 22380 14706 22392
rect 15286 22380 15292 22392
rect 15344 22380 15350 22432
rect 22465 22423 22523 22429
rect 22465 22389 22477 22423
rect 22511 22420 22523 22423
rect 23474 22420 23480 22432
rect 22511 22392 23480 22420
rect 22511 22389 22523 22392
rect 22465 22383 22523 22389
rect 23474 22380 23480 22392
rect 23532 22380 23538 22432
rect 24596 22420 24624 22664
rect 25884 22565 25912 22664
rect 26326 22652 26332 22664
rect 26384 22652 26390 22704
rect 30926 22692 30932 22704
rect 29748 22664 30932 22692
rect 27522 22624 27528 22636
rect 27483 22596 27528 22624
rect 27522 22584 27528 22596
rect 27580 22584 27586 22636
rect 27709 22627 27767 22633
rect 27709 22593 27721 22627
rect 27755 22624 27767 22627
rect 28353 22627 28411 22633
rect 28353 22624 28365 22627
rect 27755 22596 28365 22624
rect 27755 22593 27767 22596
rect 27709 22587 27767 22593
rect 28353 22593 28365 22596
rect 28399 22593 28411 22627
rect 29089 22627 29147 22633
rect 29089 22624 29101 22627
rect 28353 22587 28411 22593
rect 28966 22596 29101 22624
rect 25777 22559 25835 22565
rect 25777 22556 25789 22559
rect 25700 22528 25789 22556
rect 25700 22500 25728 22528
rect 25777 22525 25789 22528
rect 25823 22525 25835 22559
rect 25777 22519 25835 22525
rect 25869 22559 25927 22565
rect 25869 22525 25881 22559
rect 25915 22525 25927 22559
rect 27338 22556 27344 22568
rect 27299 22528 27344 22556
rect 25869 22519 25927 22525
rect 27338 22516 27344 22528
rect 27396 22556 27402 22568
rect 28966 22556 28994 22596
rect 29089 22593 29101 22596
rect 29135 22624 29147 22627
rect 29638 22624 29644 22636
rect 29135 22596 29644 22624
rect 29135 22593 29147 22596
rect 29089 22587 29147 22593
rect 29638 22584 29644 22596
rect 29696 22584 29702 22636
rect 29748 22633 29776 22664
rect 30926 22652 30932 22664
rect 30984 22652 30990 22704
rect 33410 22652 33416 22704
rect 33468 22692 33474 22704
rect 33781 22695 33839 22701
rect 33781 22692 33793 22695
rect 33468 22664 33793 22692
rect 33468 22652 33474 22664
rect 33781 22661 33793 22664
rect 33827 22692 33839 22695
rect 34238 22692 34244 22704
rect 33827 22664 34244 22692
rect 33827 22661 33839 22664
rect 33781 22655 33839 22661
rect 34238 22652 34244 22664
rect 34296 22652 34302 22704
rect 34514 22652 34520 22704
rect 34572 22692 34578 22704
rect 35069 22695 35127 22701
rect 35069 22692 35081 22695
rect 34572 22664 35081 22692
rect 34572 22652 34578 22664
rect 35069 22661 35081 22664
rect 35115 22692 35127 22695
rect 35710 22692 35716 22704
rect 35115 22664 35716 22692
rect 35115 22661 35127 22664
rect 35069 22655 35127 22661
rect 35710 22652 35716 22664
rect 35768 22652 35774 22704
rect 36170 22692 36176 22704
rect 35820 22664 36176 22692
rect 29733 22627 29791 22633
rect 29733 22593 29745 22627
rect 29779 22593 29791 22627
rect 30374 22624 30380 22636
rect 30335 22596 30380 22624
rect 29733 22587 29791 22593
rect 30374 22584 30380 22596
rect 30432 22584 30438 22636
rect 30644 22627 30702 22633
rect 30644 22593 30656 22627
rect 30690 22624 30702 22627
rect 32214 22624 32220 22636
rect 30690 22596 32220 22624
rect 30690 22593 30702 22596
rect 30644 22587 30702 22593
rect 32214 22584 32220 22596
rect 32272 22584 32278 22636
rect 32398 22584 32404 22636
rect 32456 22624 32462 22636
rect 32456 22596 33640 22624
rect 32456 22584 32462 22596
rect 27396 22528 28994 22556
rect 27396 22516 27402 22528
rect 32122 22516 32128 22568
rect 32180 22556 32186 22568
rect 32766 22556 32772 22568
rect 32180 22528 32772 22556
rect 32180 22516 32186 22528
rect 32766 22516 32772 22528
rect 32824 22516 32830 22568
rect 32858 22516 32864 22568
rect 32916 22556 32922 22568
rect 33612 22565 33640 22596
rect 34698 22584 34704 22636
rect 34756 22624 34762 22636
rect 35161 22627 35219 22633
rect 35161 22624 35173 22627
rect 34756 22596 35173 22624
rect 34756 22584 34762 22596
rect 35161 22593 35173 22596
rect 35207 22593 35219 22627
rect 35161 22587 35219 22593
rect 35250 22584 35256 22636
rect 35308 22624 35314 22636
rect 35526 22624 35532 22636
rect 35308 22596 35532 22624
rect 35308 22584 35314 22596
rect 35526 22584 35532 22596
rect 35584 22624 35590 22636
rect 35820 22624 35848 22664
rect 36170 22652 36176 22664
rect 36228 22652 36234 22704
rect 36357 22695 36415 22701
rect 36357 22661 36369 22695
rect 36403 22692 36415 22695
rect 37476 22692 37504 22720
rect 37660 22701 37688 22732
rect 37734 22720 37740 22732
rect 37792 22720 37798 22772
rect 38013 22763 38071 22769
rect 38013 22729 38025 22763
rect 38059 22760 38071 22763
rect 38746 22760 38752 22772
rect 38059 22732 38752 22760
rect 38059 22729 38071 22732
rect 38013 22723 38071 22729
rect 38746 22720 38752 22732
rect 38804 22720 38810 22772
rect 39301 22763 39359 22769
rect 39301 22729 39313 22763
rect 39347 22760 39359 22763
rect 40218 22760 40224 22772
rect 39347 22732 40224 22760
rect 39347 22729 39359 22732
rect 39301 22723 39359 22729
rect 40218 22720 40224 22732
rect 40276 22720 40282 22772
rect 40402 22720 40408 22772
rect 40460 22760 40466 22772
rect 53282 22760 53288 22772
rect 40460 22732 53288 22760
rect 40460 22720 40466 22732
rect 53282 22720 53288 22732
rect 53340 22720 53346 22772
rect 53466 22760 53472 22772
rect 53427 22732 53472 22760
rect 53466 22720 53472 22732
rect 53524 22720 53530 22772
rect 54202 22760 54208 22772
rect 54163 22732 54208 22760
rect 54202 22720 54208 22732
rect 54260 22720 54266 22772
rect 36403 22664 37504 22692
rect 37645 22695 37703 22701
rect 36403 22661 36415 22664
rect 36357 22655 36415 22661
rect 37645 22661 37657 22695
rect 37691 22692 37703 22695
rect 38378 22692 38384 22704
rect 37691 22664 38384 22692
rect 37691 22661 37703 22664
rect 37645 22655 37703 22661
rect 38378 22652 38384 22664
rect 38436 22692 38442 22704
rect 38933 22695 38991 22701
rect 38933 22692 38945 22695
rect 38436 22664 38945 22692
rect 38436 22652 38442 22664
rect 38933 22661 38945 22664
rect 38979 22661 38991 22695
rect 39758 22692 39764 22704
rect 39719 22664 39764 22692
rect 38933 22655 38991 22661
rect 39758 22652 39764 22664
rect 39816 22652 39822 22704
rect 43254 22692 43260 22704
rect 43215 22664 43260 22692
rect 43254 22652 43260 22664
rect 43312 22652 43318 22704
rect 35584 22596 35848 22624
rect 35584 22584 35590 22596
rect 36078 22584 36084 22636
rect 36136 22624 36142 22636
rect 36446 22624 36452 22636
rect 36136 22596 36452 22624
rect 36136 22584 36142 22596
rect 36446 22584 36452 22596
rect 36504 22584 36510 22636
rect 37461 22627 37519 22633
rect 37461 22593 37473 22627
rect 37507 22593 37519 22627
rect 37461 22587 37519 22593
rect 37737 22627 37795 22633
rect 37737 22593 37749 22627
rect 37783 22593 37795 22627
rect 37737 22587 37795 22593
rect 37829 22627 37887 22633
rect 37829 22593 37841 22627
rect 37875 22624 37887 22627
rect 38010 22624 38016 22636
rect 37875 22596 38016 22624
rect 37875 22593 37887 22596
rect 37829 22587 37887 22593
rect 33597 22559 33655 22565
rect 32916 22528 32961 22556
rect 32916 22516 32922 22528
rect 33597 22525 33609 22559
rect 33643 22556 33655 22559
rect 34790 22556 34796 22568
rect 33643 22528 34796 22556
rect 33643 22525 33655 22528
rect 33597 22519 33655 22525
rect 34790 22516 34796 22528
rect 34848 22556 34854 22568
rect 34885 22559 34943 22565
rect 34885 22556 34897 22559
rect 34848 22528 34897 22556
rect 34848 22516 34854 22528
rect 34885 22525 34897 22528
rect 34931 22556 34943 22559
rect 34974 22556 34980 22568
rect 34931 22528 34980 22556
rect 34931 22525 34943 22528
rect 34885 22519 34943 22525
rect 34974 22516 34980 22528
rect 35032 22556 35038 22568
rect 36541 22559 36599 22565
rect 36541 22556 36553 22559
rect 35032 22528 36553 22556
rect 35032 22516 35038 22528
rect 36541 22525 36553 22528
rect 36587 22525 36599 22559
rect 36541 22519 36599 22525
rect 25682 22448 25688 22500
rect 25740 22448 25746 22500
rect 27430 22488 27436 22500
rect 26344 22460 27436 22488
rect 26344 22420 26372 22460
rect 27430 22448 27436 22460
rect 27488 22448 27494 22500
rect 32582 22448 32588 22500
rect 32640 22488 32646 22500
rect 35618 22488 35624 22500
rect 32640 22460 35624 22488
rect 32640 22448 32646 22460
rect 35618 22448 35624 22460
rect 35676 22448 35682 22500
rect 36078 22448 36084 22500
rect 36136 22488 36142 22500
rect 37476 22488 37504 22587
rect 37752 22556 37780 22587
rect 38010 22584 38016 22596
rect 38068 22584 38074 22636
rect 38654 22584 38660 22636
rect 38712 22624 38718 22636
rect 38749 22627 38807 22633
rect 38749 22624 38761 22627
rect 38712 22596 38761 22624
rect 38712 22584 38718 22596
rect 38749 22593 38761 22596
rect 38795 22593 38807 22627
rect 38749 22587 38807 22593
rect 39025 22627 39083 22633
rect 39025 22593 39037 22627
rect 39071 22593 39083 22627
rect 39025 22587 39083 22593
rect 39117 22627 39175 22633
rect 39117 22593 39129 22627
rect 39163 22624 39175 22627
rect 39206 22624 39212 22636
rect 39163 22596 39212 22624
rect 39163 22593 39175 22596
rect 39117 22587 39175 22593
rect 38930 22556 38936 22568
rect 37752 22528 38936 22556
rect 38930 22516 38936 22528
rect 38988 22516 38994 22568
rect 39040 22556 39068 22587
rect 39206 22584 39212 22596
rect 39264 22584 39270 22636
rect 39942 22624 39948 22636
rect 39903 22596 39948 22624
rect 39942 22584 39948 22596
rect 40000 22584 40006 22636
rect 40310 22624 40316 22636
rect 40052 22596 40316 22624
rect 40052 22556 40080 22596
rect 40310 22584 40316 22596
rect 40368 22584 40374 22636
rect 40678 22624 40684 22636
rect 40639 22596 40684 22624
rect 40678 22584 40684 22596
rect 40736 22584 40742 22636
rect 40948 22627 41006 22633
rect 40948 22593 40960 22627
rect 40994 22624 41006 22627
rect 40994 22596 42656 22624
rect 40994 22593 41006 22596
rect 40948 22587 41006 22593
rect 39040 22528 40080 22556
rect 40126 22516 40132 22568
rect 40184 22556 40190 22568
rect 40586 22556 40592 22568
rect 40184 22528 40592 22556
rect 40184 22516 40190 22528
rect 40586 22516 40592 22528
rect 40644 22516 40650 22568
rect 40034 22488 40040 22500
rect 36136 22460 37504 22488
rect 39684 22460 40040 22488
rect 36136 22448 36142 22460
rect 26510 22420 26516 22432
rect 24596 22392 26372 22420
rect 26471 22392 26516 22420
rect 26510 22380 26516 22392
rect 26568 22380 26574 22432
rect 28166 22420 28172 22432
rect 28127 22392 28172 22420
rect 28166 22380 28172 22392
rect 28224 22380 28230 22432
rect 29638 22380 29644 22432
rect 29696 22420 29702 22432
rect 31294 22420 31300 22432
rect 29696 22392 31300 22420
rect 29696 22380 29702 22392
rect 31294 22380 31300 22392
rect 31352 22380 31358 22432
rect 34241 22423 34299 22429
rect 34241 22389 34253 22423
rect 34287 22420 34299 22423
rect 39684 22420 39712 22460
rect 40034 22448 40040 22460
rect 40092 22448 40098 22500
rect 42628 22497 42656 22596
rect 42702 22584 42708 22636
rect 42760 22624 42766 22636
rect 42797 22627 42855 22633
rect 42797 22624 42809 22627
rect 42760 22596 42809 22624
rect 42760 22584 42766 22596
rect 42797 22593 42809 22596
rect 42843 22593 42855 22627
rect 54021 22627 54079 22633
rect 54021 22624 54033 22627
rect 42797 22587 42855 22593
rect 51046 22596 54033 22624
rect 42613 22491 42671 22497
rect 42613 22457 42625 22491
rect 42659 22457 42671 22491
rect 51046 22488 51074 22596
rect 54021 22593 54033 22596
rect 54067 22593 54079 22627
rect 54021 22587 54079 22593
rect 42613 22451 42671 22457
rect 43180 22460 51074 22488
rect 34287 22392 39712 22420
rect 34287 22389 34299 22392
rect 34241 22383 34299 22389
rect 39758 22380 39764 22432
rect 39816 22420 39822 22432
rect 42061 22423 42119 22429
rect 42061 22420 42073 22423
rect 39816 22392 42073 22420
rect 39816 22380 39822 22392
rect 42061 22389 42073 22392
rect 42107 22420 42119 22423
rect 43180 22420 43208 22460
rect 42107 22392 43208 22420
rect 42107 22389 42119 22392
rect 42061 22383 42119 22389
rect 1104 22330 54832 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 54832 22330
rect 1104 22256 54832 22278
rect 14734 22216 14740 22228
rect 14695 22188 14740 22216
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 22741 22219 22799 22225
rect 22741 22185 22753 22219
rect 22787 22216 22799 22219
rect 22922 22216 22928 22228
rect 22787 22188 22928 22216
rect 22787 22185 22799 22188
rect 22741 22179 22799 22185
rect 22922 22176 22928 22188
rect 22980 22176 22986 22228
rect 24302 22176 24308 22228
rect 24360 22216 24366 22228
rect 24762 22216 24768 22228
rect 24360 22188 24768 22216
rect 24360 22176 24366 22188
rect 24762 22176 24768 22188
rect 24820 22176 24826 22228
rect 25038 22176 25044 22228
rect 25096 22216 25102 22228
rect 26878 22216 26884 22228
rect 25096 22188 26884 22216
rect 25096 22176 25102 22188
rect 26878 22176 26884 22188
rect 26936 22216 26942 22228
rect 27430 22216 27436 22228
rect 26936 22188 27436 22216
rect 26936 22176 26942 22188
rect 27430 22176 27436 22188
rect 27488 22176 27494 22228
rect 30926 22216 30932 22228
rect 30887 22188 30932 22216
rect 30926 22176 30932 22188
rect 30984 22176 30990 22228
rect 32766 22176 32772 22228
rect 32824 22216 32830 22228
rect 40402 22216 40408 22228
rect 32824 22188 40408 22216
rect 32824 22176 32830 22188
rect 40402 22176 40408 22188
rect 40460 22176 40466 22228
rect 40589 22219 40647 22225
rect 40589 22185 40601 22219
rect 40635 22216 40647 22219
rect 43346 22216 43352 22228
rect 40635 22188 41276 22216
rect 43307 22188 43352 22216
rect 40635 22185 40647 22188
rect 40589 22179 40647 22185
rect 1854 22108 1860 22160
rect 1912 22148 1918 22160
rect 2409 22151 2467 22157
rect 2409 22148 2421 22151
rect 1912 22120 2421 22148
rect 1912 22108 1918 22120
rect 2409 22117 2421 22120
rect 2455 22148 2467 22151
rect 23014 22148 23020 22160
rect 2455 22120 23020 22148
rect 2455 22117 2467 22120
rect 2409 22111 2467 22117
rect 23014 22108 23020 22120
rect 23072 22108 23078 22160
rect 23474 22108 23480 22160
rect 23532 22148 23538 22160
rect 27338 22148 27344 22160
rect 23532 22120 27344 22148
rect 23532 22108 23538 22120
rect 15286 22040 15292 22092
rect 15344 22080 15350 22092
rect 15473 22083 15531 22089
rect 15473 22080 15485 22083
rect 15344 22052 15485 22080
rect 15344 22040 15350 22052
rect 15473 22049 15485 22052
rect 15519 22080 15531 22083
rect 20717 22083 20775 22089
rect 20717 22080 20729 22083
rect 15519 22052 20729 22080
rect 15519 22049 15531 22052
rect 15473 22043 15531 22049
rect 20717 22049 20729 22052
rect 20763 22080 20775 22083
rect 21269 22083 21327 22089
rect 21269 22080 21281 22083
rect 20763 22052 21281 22080
rect 20763 22049 20775 22052
rect 20717 22043 20775 22049
rect 21269 22049 21281 22052
rect 21315 22049 21327 22083
rect 21269 22043 21327 22049
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 2406 22012 2412 22024
rect 1903 21984 2412 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 2406 21972 2412 21984
rect 2464 22012 2470 22024
rect 21174 22012 21180 22024
rect 2464 21984 21180 22012
rect 2464 21972 2470 21984
rect 21174 21972 21180 21984
rect 21232 21972 21238 22024
rect 1670 21876 1676 21888
rect 1631 21848 1676 21876
rect 1670 21836 1676 21848
rect 1728 21836 1734 21888
rect 21284 21876 21312 22043
rect 21913 22015 21971 22021
rect 21913 21981 21925 22015
rect 21959 22012 21971 22015
rect 22554 22012 22560 22024
rect 21959 21984 22560 22012
rect 21959 21981 21971 21984
rect 21913 21975 21971 21981
rect 22554 21972 22560 21984
rect 22612 22012 22618 22024
rect 22833 22015 22891 22021
rect 22833 22012 22845 22015
rect 22612 21984 22845 22012
rect 22612 21972 22618 21984
rect 22833 21981 22845 21984
rect 22879 21981 22891 22015
rect 23750 22012 23756 22024
rect 23711 21984 23756 22012
rect 22833 21975 22891 21981
rect 23750 21972 23756 21984
rect 23808 21972 23814 22024
rect 24762 22012 24768 22024
rect 24723 21984 24768 22012
rect 24762 21972 24768 21984
rect 24820 21972 24826 22024
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 22012 25007 22015
rect 25148 22012 25176 22120
rect 27338 22108 27344 22120
rect 27396 22108 27402 22160
rect 30282 22108 30288 22160
rect 30340 22148 30346 22160
rect 32858 22148 32864 22160
rect 30340 22120 32864 22148
rect 30340 22108 30346 22120
rect 27430 22080 27436 22092
rect 27391 22052 27436 22080
rect 27430 22040 27436 22052
rect 27488 22040 27494 22092
rect 28534 22040 28540 22092
rect 28592 22080 28598 22092
rect 29825 22083 29883 22089
rect 29825 22080 29837 22083
rect 28592 22052 29837 22080
rect 28592 22040 28598 22052
rect 29825 22049 29837 22052
rect 29871 22080 29883 22083
rect 30834 22080 30840 22092
rect 29871 22052 30840 22080
rect 29871 22049 29883 22052
rect 29825 22043 29883 22049
rect 30834 22040 30840 22052
rect 30892 22040 30898 22092
rect 31496 22089 31524 22120
rect 31481 22083 31539 22089
rect 31481 22049 31493 22083
rect 31527 22080 31539 22083
rect 32692 22080 32720 22120
rect 32858 22108 32864 22120
rect 32916 22108 32922 22160
rect 36354 22148 36360 22160
rect 36280 22120 36360 22148
rect 36280 22089 36308 22120
rect 36354 22108 36360 22120
rect 36412 22108 36418 22160
rect 36630 22148 36636 22160
rect 36464 22120 36636 22148
rect 32769 22083 32827 22089
rect 32769 22080 32781 22083
rect 31527 22052 31561 22080
rect 32692 22052 32781 22080
rect 31527 22049 31539 22052
rect 31481 22043 31539 22049
rect 32769 22049 32781 22052
rect 32815 22049 32827 22083
rect 32769 22043 32827 22049
rect 36265 22083 36323 22089
rect 36265 22049 36277 22083
rect 36311 22049 36323 22083
rect 36464 22080 36492 22120
rect 36630 22108 36636 22120
rect 36688 22108 36694 22160
rect 36725 22151 36783 22157
rect 36725 22117 36737 22151
rect 36771 22117 36783 22151
rect 36725 22111 36783 22117
rect 36740 22080 36768 22111
rect 36814 22108 36820 22160
rect 36872 22148 36878 22160
rect 36872 22120 37780 22148
rect 36872 22108 36878 22120
rect 37550 22080 37556 22092
rect 36265 22043 36323 22049
rect 36372 22052 36492 22080
rect 36556 22052 36768 22080
rect 37511 22052 37556 22080
rect 24995 21984 25176 22012
rect 25777 22015 25835 22021
rect 24995 21981 25007 21984
rect 24949 21975 25007 21981
rect 25777 21981 25789 22015
rect 25823 21981 25835 22015
rect 25777 21975 25835 21981
rect 25961 22015 26019 22021
rect 25961 21981 25973 22015
rect 26007 22012 26019 22015
rect 27154 22012 27160 22024
rect 26007 21984 27160 22012
rect 26007 21981 26019 21984
rect 25961 21975 26019 21981
rect 22278 21904 22284 21956
rect 22336 21944 22342 21956
rect 25498 21944 25504 21956
rect 22336 21916 25504 21944
rect 22336 21904 22342 21916
rect 25498 21904 25504 21916
rect 25556 21904 25562 21956
rect 25792 21944 25820 21975
rect 27154 21972 27160 21984
rect 27212 21972 27218 22024
rect 27700 22015 27758 22021
rect 27700 21981 27712 22015
rect 27746 22012 27758 22015
rect 28166 22012 28172 22024
rect 27746 21984 28172 22012
rect 27746 21981 27758 21984
rect 27700 21975 27758 21981
rect 28166 21972 28172 21984
rect 28224 21972 28230 22024
rect 28276 21984 31156 22012
rect 26421 21947 26479 21953
rect 26421 21944 26433 21947
rect 25792 21916 26433 21944
rect 26421 21913 26433 21916
rect 26467 21913 26479 21947
rect 26602 21944 26608 21956
rect 26563 21916 26608 21944
rect 26421 21907 26479 21913
rect 26602 21904 26608 21916
rect 26660 21904 26666 21956
rect 26786 21944 26792 21956
rect 26747 21916 26792 21944
rect 26786 21904 26792 21916
rect 26844 21904 26850 21956
rect 28276 21944 28304 21984
rect 30101 21947 30159 21953
rect 30101 21944 30113 21947
rect 26896 21916 28304 21944
rect 28828 21916 30113 21944
rect 22094 21876 22100 21888
rect 21284 21848 22100 21876
rect 22094 21836 22100 21848
rect 22152 21836 22158 21888
rect 22186 21836 22192 21888
rect 22244 21876 22250 21888
rect 22373 21879 22431 21885
rect 22373 21876 22385 21879
rect 22244 21848 22385 21876
rect 22244 21836 22250 21848
rect 22373 21845 22385 21848
rect 22419 21845 22431 21879
rect 23566 21876 23572 21888
rect 23527 21848 23572 21876
rect 22373 21839 22431 21845
rect 23566 21836 23572 21848
rect 23624 21836 23630 21888
rect 23658 21836 23664 21888
rect 23716 21876 23722 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 23716 21848 24593 21876
rect 23716 21836 23722 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 24670 21836 24676 21888
rect 24728 21876 24734 21888
rect 25593 21879 25651 21885
rect 25593 21876 25605 21879
rect 24728 21848 25605 21876
rect 24728 21836 24734 21848
rect 25593 21845 25605 21848
rect 25639 21845 25651 21879
rect 25593 21839 25651 21845
rect 26326 21836 26332 21888
rect 26384 21876 26390 21888
rect 26896 21876 26924 21916
rect 28828 21888 28856 21916
rect 30101 21913 30113 21916
rect 30147 21913 30159 21947
rect 31128 21944 31156 21984
rect 31202 21972 31208 22024
rect 31260 22012 31266 22024
rect 31297 22015 31355 22021
rect 31297 22012 31309 22015
rect 31260 21984 31309 22012
rect 31260 21972 31266 21984
rect 31297 21981 31309 21984
rect 31343 21981 31355 22015
rect 31297 21975 31355 21981
rect 31754 21972 31760 22024
rect 31812 22012 31818 22024
rect 32306 22012 32312 22024
rect 31812 21984 32312 22012
rect 31812 21972 31818 21984
rect 32306 21972 32312 21984
rect 32364 22012 32370 22024
rect 32493 22015 32551 22021
rect 32493 22012 32505 22015
rect 32364 21984 32505 22012
rect 32364 21972 32370 21984
rect 32493 21981 32505 21984
rect 32539 21981 32551 22015
rect 32493 21975 32551 21981
rect 33134 21972 33140 22024
rect 33192 22012 33198 22024
rect 33318 22012 33324 22024
rect 33192 21984 33324 22012
rect 33192 21972 33198 21984
rect 33318 21972 33324 21984
rect 33376 22012 33382 22024
rect 33873 22015 33931 22021
rect 33873 22012 33885 22015
rect 33376 21984 33885 22012
rect 33376 21972 33382 21984
rect 33873 21981 33885 21984
rect 33919 21981 33931 22015
rect 36372 22012 36400 22052
rect 33873 21975 33931 21981
rect 35084 21984 36400 22012
rect 35084 21944 35112 21984
rect 31128 21916 35112 21944
rect 36020 21947 36078 21953
rect 30101 21907 30159 21913
rect 36020 21913 36032 21947
rect 36066 21944 36078 21947
rect 36556 21944 36584 22052
rect 37550 22040 37556 22052
rect 37608 22040 37614 22092
rect 37752 22089 37780 22120
rect 38654 22108 38660 22160
rect 38712 22108 38718 22160
rect 38746 22108 38752 22160
rect 38804 22148 38810 22160
rect 41046 22148 41052 22160
rect 38804 22120 41052 22148
rect 38804 22108 38810 22120
rect 41046 22108 41052 22120
rect 41104 22108 41110 22160
rect 37737 22083 37795 22089
rect 37737 22049 37749 22083
rect 37783 22080 37795 22083
rect 38672 22080 38700 22108
rect 37783 22052 38700 22080
rect 37783 22049 37795 22052
rect 37737 22043 37795 22049
rect 36906 22012 36912 22024
rect 36867 21984 36912 22012
rect 36906 21972 36912 21984
rect 36964 21972 36970 22024
rect 37090 21972 37096 22024
rect 37148 22012 37154 22024
rect 38608 22012 38614 22024
rect 37148 21984 38614 22012
rect 37148 21972 37154 21984
rect 38608 21972 38614 21984
rect 38666 22021 38672 22024
rect 38666 22015 38715 22021
rect 38666 21981 38669 22015
rect 38703 21981 38715 22015
rect 38666 21975 38715 21981
rect 38827 22015 38885 22021
rect 38827 21981 38839 22015
rect 38873 22012 38885 22015
rect 39022 22012 39028 22024
rect 38873 21984 39028 22012
rect 38873 21981 38885 21984
rect 38827 21975 38885 21981
rect 38666 21972 38672 21975
rect 39022 21972 39028 21984
rect 39080 21972 39086 22024
rect 40034 22012 40040 22024
rect 39995 21984 40040 22012
rect 40034 21972 40040 21984
rect 40092 21972 40098 22024
rect 40402 22012 40408 22024
rect 40363 21984 40408 22012
rect 40402 21972 40408 21984
rect 40460 21972 40466 22024
rect 40586 21972 40592 22024
rect 40644 22012 40650 22024
rect 40954 22012 40960 22024
rect 40644 21984 40960 22012
rect 40644 21972 40650 21984
rect 40954 21972 40960 21984
rect 41012 22012 41018 22024
rect 41049 22015 41107 22021
rect 41049 22012 41061 22015
rect 41012 21984 41061 22012
rect 41012 21972 41018 21984
rect 41049 21981 41061 21984
rect 41095 22012 41107 22015
rect 41138 22012 41144 22024
rect 41095 21984 41144 22012
rect 41095 21981 41107 21984
rect 41049 21975 41107 21981
rect 41138 21972 41144 21984
rect 41196 21972 41202 22024
rect 41248 22021 41276 22188
rect 43346 22176 43352 22188
rect 43404 22176 43410 22228
rect 41417 22083 41475 22089
rect 41417 22049 41429 22083
rect 41463 22080 41475 22083
rect 41506 22080 41512 22092
rect 41463 22052 41512 22080
rect 41463 22049 41475 22052
rect 41417 22043 41475 22049
rect 41506 22040 41512 22052
rect 41564 22040 41570 22092
rect 42794 22080 42800 22092
rect 42755 22052 42800 22080
rect 42794 22040 42800 22052
rect 42852 22040 42858 22092
rect 41233 22015 41291 22021
rect 41233 21981 41245 22015
rect 41279 21981 41291 22015
rect 41233 21975 41291 21981
rect 41322 21972 41328 22024
rect 41380 22012 41386 22024
rect 41877 22015 41935 22021
rect 41877 22012 41889 22015
rect 41380 21984 41889 22012
rect 41380 21972 41386 21984
rect 41877 21981 41889 21984
rect 41923 21981 41935 22015
rect 42058 22012 42064 22024
rect 42019 21984 42064 22012
rect 41877 21975 41935 21981
rect 42058 21972 42064 21984
rect 42116 21972 42122 22024
rect 42242 22012 42248 22024
rect 42203 21984 42248 22012
rect 42242 21972 42248 21984
rect 42300 21972 42306 22024
rect 53558 21972 53564 22024
rect 53616 22012 53622 22024
rect 54202 22012 54208 22024
rect 53616 21984 54208 22012
rect 53616 21972 53622 21984
rect 54202 21972 54208 21984
rect 54260 21972 54266 22024
rect 39942 21944 39948 21956
rect 36066 21916 36584 21944
rect 36648 21916 39948 21944
rect 36066 21913 36078 21916
rect 36020 21907 36078 21913
rect 26384 21848 26924 21876
rect 26384 21836 26390 21848
rect 27798 21836 27804 21888
rect 27856 21876 27862 21888
rect 28810 21876 28816 21888
rect 27856 21848 28816 21876
rect 27856 21836 27862 21848
rect 28810 21836 28816 21848
rect 28868 21836 28874 21888
rect 29822 21836 29828 21888
rect 29880 21876 29886 21888
rect 30009 21879 30067 21885
rect 30009 21876 30021 21879
rect 29880 21848 30021 21876
rect 29880 21836 29886 21848
rect 30009 21845 30021 21848
rect 30055 21845 30067 21879
rect 30466 21876 30472 21888
rect 30427 21848 30472 21876
rect 30009 21839 30067 21845
rect 30466 21836 30472 21848
rect 30524 21836 30530 21888
rect 31386 21876 31392 21888
rect 31347 21848 31392 21876
rect 31386 21836 31392 21848
rect 31444 21836 31450 21888
rect 31570 21836 31576 21888
rect 31628 21876 31634 21888
rect 32125 21879 32183 21885
rect 32125 21876 32137 21879
rect 31628 21848 32137 21876
rect 31628 21836 31634 21848
rect 32125 21845 32137 21848
rect 32171 21845 32183 21879
rect 32582 21876 32588 21888
rect 32543 21848 32588 21876
rect 32125 21839 32183 21845
rect 32582 21836 32588 21848
rect 32640 21836 32646 21888
rect 33321 21879 33379 21885
rect 33321 21845 33333 21879
rect 33367 21876 33379 21879
rect 33686 21876 33692 21888
rect 33367 21848 33692 21876
rect 33367 21845 33379 21848
rect 33321 21839 33379 21845
rect 33686 21836 33692 21848
rect 33744 21836 33750 21888
rect 34698 21836 34704 21888
rect 34756 21876 34762 21888
rect 34885 21879 34943 21885
rect 34885 21876 34897 21879
rect 34756 21848 34897 21876
rect 34756 21836 34762 21848
rect 34885 21845 34897 21848
rect 34931 21845 34943 21879
rect 34885 21839 34943 21845
rect 35434 21836 35440 21888
rect 35492 21876 35498 21888
rect 36648 21876 36676 21916
rect 39942 21904 39948 21916
rect 40000 21904 40006 21956
rect 40218 21944 40224 21956
rect 40179 21916 40224 21944
rect 40218 21904 40224 21916
rect 40276 21904 40282 21956
rect 40313 21947 40371 21953
rect 40313 21913 40325 21947
rect 40359 21944 40371 21947
rect 42334 21944 42340 21956
rect 40359 21916 42340 21944
rect 40359 21913 40371 21916
rect 40313 21907 40371 21913
rect 42334 21904 42340 21916
rect 42392 21904 42398 21956
rect 53282 21944 53288 21956
rect 53243 21916 53288 21944
rect 53282 21904 53288 21916
rect 53340 21904 53346 21956
rect 53466 21944 53472 21956
rect 53427 21916 53472 21944
rect 53466 21904 53472 21916
rect 53524 21904 53530 21956
rect 54018 21944 54024 21956
rect 53979 21916 54024 21944
rect 54018 21904 54024 21916
rect 54076 21904 54082 21956
rect 35492 21848 36676 21876
rect 35492 21836 35498 21848
rect 37458 21836 37464 21888
rect 37516 21876 37522 21888
rect 37829 21879 37887 21885
rect 37829 21876 37841 21879
rect 37516 21848 37841 21876
rect 37516 21836 37522 21848
rect 37829 21845 37841 21848
rect 37875 21845 37887 21879
rect 37829 21839 37887 21845
rect 38197 21879 38255 21885
rect 38197 21845 38209 21879
rect 38243 21876 38255 21879
rect 38654 21876 38660 21888
rect 38243 21848 38660 21876
rect 38243 21845 38255 21848
rect 38197 21839 38255 21845
rect 38654 21836 38660 21848
rect 38712 21836 38718 21888
rect 39025 21879 39083 21885
rect 39025 21845 39037 21879
rect 39071 21876 39083 21879
rect 40126 21876 40132 21888
rect 39071 21848 40132 21876
rect 39071 21845 39083 21848
rect 39025 21839 39083 21845
rect 40126 21836 40132 21848
rect 40184 21836 40190 21888
rect 41046 21836 41052 21888
rect 41104 21876 41110 21888
rect 43714 21876 43720 21888
rect 41104 21848 43720 21876
rect 41104 21836 41110 21848
rect 43714 21836 43720 21848
rect 43772 21876 43778 21888
rect 43809 21879 43867 21885
rect 43809 21876 43821 21879
rect 43772 21848 43821 21876
rect 43772 21836 43778 21848
rect 43809 21845 43821 21848
rect 43855 21845 43867 21879
rect 43809 21839 43867 21845
rect 52825 21879 52883 21885
rect 52825 21845 52837 21879
rect 52871 21876 52883 21879
rect 53484 21876 53512 21904
rect 52871 21848 53512 21876
rect 52871 21845 52883 21848
rect 52825 21839 52883 21845
rect 1104 21786 54832 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 54832 21786
rect 1104 21712 54832 21734
rect 2406 21672 2412 21684
rect 2367 21644 2412 21672
rect 2406 21632 2412 21644
rect 2464 21632 2470 21684
rect 2498 21632 2504 21684
rect 2556 21672 2562 21684
rect 23566 21672 23572 21684
rect 2556 21644 23572 21672
rect 2556 21632 2562 21644
rect 23566 21632 23572 21644
rect 23624 21632 23630 21684
rect 25317 21675 25375 21681
rect 25317 21641 25329 21675
rect 25363 21641 25375 21675
rect 25317 21635 25375 21641
rect 27157 21675 27215 21681
rect 27157 21641 27169 21675
rect 27203 21672 27215 21675
rect 27522 21672 27528 21684
rect 27203 21644 27528 21672
rect 27203 21641 27215 21644
rect 27157 21635 27215 21641
rect 20809 21607 20867 21613
rect 20809 21573 20821 21607
rect 20855 21604 20867 21607
rect 22278 21604 22284 21616
rect 20855 21576 22284 21604
rect 20855 21573 20867 21576
rect 20809 21567 20867 21573
rect 22278 21564 22284 21576
rect 22336 21564 22342 21616
rect 24578 21604 24584 21616
rect 23952 21576 24584 21604
rect 1857 21539 1915 21545
rect 1857 21505 1869 21539
rect 1903 21536 1915 21539
rect 2406 21536 2412 21548
rect 1903 21508 2412 21536
rect 1903 21505 1915 21508
rect 1857 21499 1915 21505
rect 2406 21496 2412 21508
rect 2464 21536 2470 21548
rect 14090 21536 14096 21548
rect 2464 21508 6914 21536
rect 14051 21508 14096 21536
rect 2464 21496 2470 21508
rect 6886 21468 6914 21508
rect 14090 21496 14096 21508
rect 14148 21496 14154 21548
rect 21453 21539 21511 21545
rect 21453 21505 21465 21539
rect 21499 21505 21511 21539
rect 22296 21536 22324 21564
rect 22465 21539 22523 21545
rect 22465 21536 22477 21539
rect 22296 21508 22477 21536
rect 21453 21499 21511 21505
rect 22465 21505 22477 21508
rect 22511 21505 22523 21539
rect 22465 21499 22523 21505
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21536 23351 21539
rect 23658 21536 23664 21548
rect 23339 21508 23664 21536
rect 23339 21505 23351 21508
rect 23293 21499 23351 21505
rect 21358 21468 21364 21480
rect 6886 21440 21364 21468
rect 21358 21428 21364 21440
rect 21416 21428 21422 21480
rect 21468 21468 21496 21499
rect 23658 21496 23664 21508
rect 23716 21496 23722 21548
rect 23952 21545 23980 21576
rect 24578 21564 24584 21576
rect 24636 21604 24642 21616
rect 25038 21604 25044 21616
rect 24636 21576 25044 21604
rect 24636 21564 24642 21576
rect 25038 21564 25044 21576
rect 25096 21564 25102 21616
rect 25332 21604 25360 21635
rect 27522 21632 27528 21644
rect 27580 21632 27586 21684
rect 29822 21632 29828 21684
rect 29880 21672 29886 21684
rect 31662 21672 31668 21684
rect 29880 21644 31668 21672
rect 29880 21632 29886 21644
rect 31662 21632 31668 21644
rect 31720 21672 31726 21684
rect 33505 21675 33563 21681
rect 33505 21672 33517 21675
rect 31720 21644 33517 21672
rect 31720 21632 31726 21644
rect 33505 21641 33517 21644
rect 33551 21641 33563 21675
rect 35434 21672 35440 21684
rect 35395 21644 35440 21672
rect 33505 21635 33563 21641
rect 35434 21632 35440 21644
rect 35492 21632 35498 21684
rect 35897 21675 35955 21681
rect 35897 21641 35909 21675
rect 35943 21672 35955 21675
rect 36078 21672 36084 21684
rect 35943 21644 36084 21672
rect 35943 21641 35955 21644
rect 35897 21635 35955 21641
rect 36078 21632 36084 21644
rect 36136 21632 36142 21684
rect 36280 21644 38976 21672
rect 26142 21604 26148 21616
rect 25332 21576 26148 21604
rect 25884 21545 25912 21576
rect 26142 21564 26148 21576
rect 26200 21604 26206 21616
rect 28721 21607 28779 21613
rect 28721 21604 28733 21607
rect 26200 21576 28733 21604
rect 26200 21564 26206 21576
rect 28721 21573 28733 21576
rect 28767 21573 28779 21607
rect 36280 21604 36308 21644
rect 28721 21567 28779 21573
rect 33060 21576 36308 21604
rect 23937 21539 23995 21545
rect 23937 21505 23949 21539
rect 23983 21505 23995 21539
rect 24193 21539 24251 21545
rect 24193 21536 24205 21539
rect 23937 21499 23995 21505
rect 24044 21508 24205 21536
rect 22005 21471 22063 21477
rect 22005 21468 22017 21471
rect 21468 21440 22017 21468
rect 22005 21437 22017 21440
rect 22051 21437 22063 21471
rect 24044 21468 24072 21508
rect 24193 21505 24205 21508
rect 24239 21505 24251 21539
rect 24193 21499 24251 21505
rect 25869 21539 25927 21545
rect 25869 21505 25881 21539
rect 25915 21505 25927 21539
rect 25869 21499 25927 21505
rect 27525 21539 27583 21545
rect 27525 21505 27537 21539
rect 27571 21536 27583 21539
rect 27798 21536 27804 21548
rect 27571 21508 27804 21536
rect 27571 21505 27583 21508
rect 27525 21499 27583 21505
rect 27798 21496 27804 21508
rect 27856 21496 27862 21548
rect 29362 21536 29368 21548
rect 27908 21508 29368 21536
rect 22005 21431 22063 21437
rect 23492 21440 24072 21468
rect 21174 21360 21180 21412
rect 21232 21400 21238 21412
rect 23492 21409 23520 21440
rect 26510 21428 26516 21480
rect 26568 21468 26574 21480
rect 27430 21468 27436 21480
rect 26568 21440 27436 21468
rect 26568 21428 26574 21440
rect 27430 21428 27436 21440
rect 27488 21468 27494 21480
rect 27617 21471 27675 21477
rect 27617 21468 27629 21471
rect 27488 21440 27629 21468
rect 27488 21428 27494 21440
rect 27617 21437 27629 21440
rect 27663 21437 27675 21471
rect 27617 21431 27675 21437
rect 27709 21471 27767 21477
rect 27709 21437 27721 21471
rect 27755 21468 27767 21471
rect 27908 21468 27936 21508
rect 29362 21496 29368 21508
rect 29420 21536 29426 21548
rect 30282 21536 30288 21548
rect 29420 21508 30288 21536
rect 29420 21496 29426 21508
rect 30282 21496 30288 21508
rect 30340 21496 30346 21548
rect 31202 21496 31208 21548
rect 31260 21536 31266 21548
rect 31389 21539 31447 21545
rect 31389 21536 31401 21539
rect 31260 21508 31401 21536
rect 31260 21496 31266 21508
rect 31389 21505 31401 21508
rect 31435 21536 31447 21539
rect 32490 21536 32496 21548
rect 31435 21508 32496 21536
rect 31435 21505 31447 21508
rect 31389 21499 31447 21505
rect 32490 21496 32496 21508
rect 32548 21536 32554 21548
rect 32677 21539 32735 21545
rect 32677 21536 32689 21539
rect 32548 21508 32689 21536
rect 32548 21496 32554 21508
rect 32677 21505 32689 21508
rect 32723 21505 32735 21539
rect 32677 21499 32735 21505
rect 28534 21468 28540 21480
rect 27755 21440 27936 21468
rect 28495 21440 28540 21468
rect 27755 21437 27767 21440
rect 27709 21431 27767 21437
rect 28534 21428 28540 21440
rect 28592 21428 28598 21480
rect 28626 21428 28632 21480
rect 28684 21468 28690 21480
rect 28684 21440 28729 21468
rect 28684 21428 28690 21440
rect 28810 21428 28816 21480
rect 28868 21468 28874 21480
rect 29641 21471 29699 21477
rect 29641 21468 29653 21471
rect 28868 21440 29653 21468
rect 28868 21428 28874 21440
rect 29641 21437 29653 21440
rect 29687 21437 29699 21471
rect 32398 21468 32404 21480
rect 32359 21440 32404 21468
rect 29641 21431 29699 21437
rect 32398 21428 32404 21440
rect 32456 21428 32462 21480
rect 32585 21471 32643 21477
rect 32585 21437 32597 21471
rect 32631 21437 32643 21471
rect 32585 21431 32643 21437
rect 21269 21403 21327 21409
rect 21269 21400 21281 21403
rect 21232 21372 21281 21400
rect 21232 21360 21238 21372
rect 21269 21369 21281 21372
rect 21315 21369 21327 21403
rect 23477 21403 23535 21409
rect 21269 21363 21327 21369
rect 21376 21372 23428 21400
rect 1670 21332 1676 21344
rect 1631 21304 1676 21332
rect 1670 21292 1676 21304
rect 1728 21292 1734 21344
rect 13906 21332 13912 21344
rect 13867 21304 13912 21332
rect 13906 21292 13912 21304
rect 13964 21292 13970 21344
rect 18138 21292 18144 21344
rect 18196 21332 18202 21344
rect 21376 21332 21404 21372
rect 18196 21304 21404 21332
rect 18196 21292 18202 21304
rect 22094 21292 22100 21344
rect 22152 21332 22158 21344
rect 22370 21332 22376 21344
rect 22152 21304 22376 21332
rect 22152 21292 22158 21304
rect 22370 21292 22376 21304
rect 22428 21332 22434 21344
rect 22830 21332 22836 21344
rect 22428 21304 22836 21332
rect 22428 21292 22434 21304
rect 22830 21292 22836 21304
rect 22888 21332 22894 21344
rect 23290 21332 23296 21344
rect 22888 21304 23296 21332
rect 22888 21292 22894 21304
rect 23290 21292 23296 21304
rect 23348 21292 23354 21344
rect 23400 21332 23428 21372
rect 23477 21369 23489 21403
rect 23523 21369 23535 21403
rect 26878 21400 26884 21412
rect 23477 21363 23535 21369
rect 24872 21372 26884 21400
rect 24872 21332 24900 21372
rect 26878 21360 26884 21372
rect 26936 21360 26942 21412
rect 28718 21360 28724 21412
rect 28776 21400 28782 21412
rect 28776 21372 31754 21400
rect 28776 21360 28782 21372
rect 23400 21304 24900 21332
rect 25130 21292 25136 21344
rect 25188 21332 25194 21344
rect 25498 21332 25504 21344
rect 25188 21304 25504 21332
rect 25188 21292 25194 21304
rect 25498 21292 25504 21304
rect 25556 21292 25562 21344
rect 26421 21335 26479 21341
rect 26421 21301 26433 21335
rect 26467 21332 26479 21335
rect 27614 21332 27620 21344
rect 26467 21304 27620 21332
rect 26467 21301 26479 21304
rect 26421 21295 26479 21301
rect 27614 21292 27620 21304
rect 27672 21292 27678 21344
rect 29086 21332 29092 21344
rect 29047 21304 29092 21332
rect 29086 21292 29092 21304
rect 29144 21292 29150 21344
rect 30098 21292 30104 21344
rect 30156 21332 30162 21344
rect 30193 21335 30251 21341
rect 30193 21332 30205 21335
rect 30156 21304 30205 21332
rect 30156 21292 30162 21304
rect 30193 21301 30205 21304
rect 30239 21301 30251 21335
rect 30193 21295 30251 21301
rect 30837 21335 30895 21341
rect 30837 21301 30849 21335
rect 30883 21332 30895 21335
rect 30926 21332 30932 21344
rect 30883 21304 30932 21332
rect 30883 21301 30895 21304
rect 30837 21295 30895 21301
rect 30926 21292 30932 21304
rect 30984 21292 30990 21344
rect 31726 21332 31754 21372
rect 31846 21360 31852 21412
rect 31904 21400 31910 21412
rect 32030 21400 32036 21412
rect 31904 21372 32036 21400
rect 31904 21360 31910 21372
rect 32030 21360 32036 21372
rect 32088 21400 32094 21412
rect 32600 21400 32628 21431
rect 33060 21409 33088 21576
rect 36354 21564 36360 21616
rect 36412 21604 36418 21616
rect 36412 21576 38884 21604
rect 36412 21564 36418 21576
rect 38856 21548 38884 21576
rect 35526 21536 35532 21548
rect 35487 21508 35532 21536
rect 35526 21496 35532 21508
rect 35584 21496 35590 21548
rect 36170 21496 36176 21548
rect 36228 21536 36234 21548
rect 36541 21539 36599 21545
rect 36541 21536 36553 21539
rect 36228 21508 36553 21536
rect 36228 21496 36234 21508
rect 36541 21505 36553 21508
rect 36587 21505 36599 21539
rect 36541 21499 36599 21505
rect 36633 21539 36691 21545
rect 36633 21505 36645 21539
rect 36679 21505 36691 21539
rect 36633 21499 36691 21505
rect 34698 21468 34704 21480
rect 34659 21440 34704 21468
rect 34698 21428 34704 21440
rect 34756 21428 34762 21480
rect 34790 21428 34796 21480
rect 34848 21468 34854 21480
rect 35253 21471 35311 21477
rect 35253 21468 35265 21471
rect 34848 21440 35265 21468
rect 34848 21428 34854 21440
rect 35253 21437 35265 21440
rect 35299 21437 35311 21471
rect 35253 21431 35311 21437
rect 36648 21468 36676 21499
rect 36722 21496 36728 21548
rect 36780 21536 36786 21548
rect 38562 21536 38568 21548
rect 38620 21545 38626 21548
rect 36780 21508 36825 21536
rect 38532 21508 38568 21536
rect 36780 21496 36786 21508
rect 38562 21496 38568 21508
rect 38620 21499 38632 21545
rect 38838 21536 38844 21548
rect 38751 21508 38844 21536
rect 38620 21496 38626 21499
rect 38838 21496 38844 21508
rect 38896 21496 38902 21548
rect 38948 21536 38976 21644
rect 39206 21632 39212 21684
rect 39264 21672 39270 21684
rect 40037 21675 40095 21681
rect 39264 21644 39896 21672
rect 39264 21632 39270 21644
rect 39758 21604 39764 21616
rect 39719 21576 39764 21604
rect 39758 21564 39764 21576
rect 39816 21564 39822 21616
rect 39868 21545 39896 21644
rect 40037 21641 40049 21675
rect 40083 21672 40095 21675
rect 42058 21672 42064 21684
rect 40083 21644 42064 21672
rect 40083 21641 40095 21644
rect 40037 21635 40095 21641
rect 42058 21632 42064 21644
rect 42116 21632 42122 21684
rect 42242 21632 42248 21684
rect 42300 21672 42306 21684
rect 42702 21672 42708 21684
rect 42300 21644 42708 21672
rect 42300 21632 42306 21644
rect 42702 21632 42708 21644
rect 42760 21632 42766 21684
rect 53558 21672 53564 21684
rect 53519 21644 53564 21672
rect 53558 21632 53564 21644
rect 53616 21632 53622 21684
rect 54202 21672 54208 21684
rect 54163 21644 54208 21672
rect 54202 21632 54208 21644
rect 54260 21632 54266 21684
rect 39942 21564 39948 21616
rect 40000 21604 40006 21616
rect 42613 21607 42671 21613
rect 42613 21604 42625 21607
rect 40000 21576 42625 21604
rect 40000 21564 40006 21576
rect 42613 21573 42625 21576
rect 42659 21573 42671 21607
rect 42613 21567 42671 21573
rect 39485 21539 39543 21545
rect 39485 21536 39497 21539
rect 38948 21508 39497 21536
rect 39485 21505 39497 21508
rect 39531 21505 39543 21539
rect 39485 21499 39543 21505
rect 39669 21539 39727 21545
rect 39669 21505 39681 21539
rect 39715 21505 39727 21539
rect 39669 21499 39727 21505
rect 39853 21539 39911 21545
rect 39853 21505 39865 21539
rect 39899 21536 39911 21539
rect 40402 21536 40408 21548
rect 39899 21508 40408 21536
rect 39899 21505 39911 21508
rect 39853 21499 39911 21505
rect 37366 21468 37372 21480
rect 36648 21440 37372 21468
rect 32088 21372 32628 21400
rect 33045 21403 33103 21409
rect 32088 21360 32094 21372
rect 33045 21369 33057 21403
rect 33091 21369 33103 21403
rect 33045 21363 33103 21369
rect 34057 21403 34115 21409
rect 34057 21369 34069 21403
rect 34103 21400 34115 21403
rect 36648 21400 36676 21440
rect 37366 21428 37372 21440
rect 37424 21428 37430 21480
rect 39114 21428 39120 21480
rect 39172 21468 39178 21480
rect 39684 21468 39712 21499
rect 40402 21496 40408 21508
rect 40460 21496 40466 21548
rect 40948 21539 41006 21545
rect 40948 21505 40960 21539
rect 40994 21536 41006 21539
rect 42702 21536 42708 21548
rect 40994 21508 42708 21536
rect 40994 21505 41006 21508
rect 40948 21499 41006 21505
rect 42702 21496 42708 21508
rect 42760 21496 42766 21548
rect 54021 21539 54079 21545
rect 54021 21536 54033 21539
rect 51046 21508 54033 21536
rect 40218 21468 40224 21480
rect 39172 21440 40224 21468
rect 39172 21428 39178 21440
rect 40218 21428 40224 21440
rect 40276 21428 40282 21480
rect 40678 21468 40684 21480
rect 40639 21440 40684 21468
rect 40678 21428 40684 21440
rect 40736 21428 40742 21480
rect 36906 21400 36912 21412
rect 34103 21372 36676 21400
rect 36867 21372 36912 21400
rect 34103 21369 34115 21372
rect 34057 21363 34115 21369
rect 36906 21360 36912 21372
rect 36964 21360 36970 21412
rect 41690 21360 41696 21412
rect 41748 21400 41754 21412
rect 42061 21403 42119 21409
rect 42061 21400 42073 21403
rect 41748 21372 42073 21400
rect 41748 21360 41754 21372
rect 42061 21369 42073 21372
rect 42107 21400 42119 21403
rect 51046 21400 51074 21508
rect 54021 21505 54033 21508
rect 54067 21505 54079 21539
rect 54021 21499 54079 21505
rect 42107 21372 51074 21400
rect 42107 21369 42119 21372
rect 42061 21363 42119 21369
rect 32858 21332 32864 21344
rect 31726 21304 32864 21332
rect 32858 21292 32864 21304
rect 32916 21292 32922 21344
rect 35894 21292 35900 21344
rect 35952 21332 35958 21344
rect 36357 21335 36415 21341
rect 36357 21332 36369 21335
rect 35952 21304 36369 21332
rect 35952 21292 35958 21304
rect 36357 21301 36369 21304
rect 36403 21332 36415 21335
rect 36538 21332 36544 21344
rect 36403 21304 36544 21332
rect 36403 21301 36415 21304
rect 36357 21295 36415 21301
rect 36538 21292 36544 21304
rect 36596 21292 36602 21344
rect 37458 21332 37464 21344
rect 37419 21304 37464 21332
rect 37458 21292 37464 21304
rect 37516 21292 37522 21344
rect 37642 21292 37648 21344
rect 37700 21332 37706 21344
rect 41782 21332 41788 21344
rect 37700 21304 41788 21332
rect 37700 21292 37706 21304
rect 41782 21292 41788 21304
rect 41840 21292 41846 21344
rect 1104 21242 54832 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 54832 21242
rect 1104 21168 54832 21190
rect 2406 21128 2412 21140
rect 2367 21100 2412 21128
rect 2406 21088 2412 21100
rect 2464 21088 2470 21140
rect 21358 21088 21364 21140
rect 21416 21128 21422 21140
rect 22005 21131 22063 21137
rect 22005 21128 22017 21131
rect 21416 21100 22017 21128
rect 21416 21088 21422 21100
rect 22005 21097 22017 21100
rect 22051 21097 22063 21131
rect 22005 21091 22063 21097
rect 23017 21131 23075 21137
rect 23017 21097 23029 21131
rect 23063 21128 23075 21131
rect 23290 21128 23296 21140
rect 23063 21100 23296 21128
rect 23063 21097 23075 21100
rect 23017 21091 23075 21097
rect 23290 21088 23296 21100
rect 23348 21088 23354 21140
rect 26326 21128 26332 21140
rect 24596 21100 26332 21128
rect 19889 21063 19947 21069
rect 19889 21029 19901 21063
rect 19935 21060 19947 21063
rect 19978 21060 19984 21072
rect 19935 21032 19984 21060
rect 19935 21029 19947 21032
rect 19889 21023 19947 21029
rect 19978 21020 19984 21032
rect 20036 21060 20042 21072
rect 24596 21060 24624 21100
rect 26326 21088 26332 21100
rect 26384 21088 26390 21140
rect 26602 21128 26608 21140
rect 26563 21100 26608 21128
rect 26602 21088 26608 21100
rect 26660 21088 26666 21140
rect 26878 21088 26884 21140
rect 26936 21128 26942 21140
rect 32582 21128 32588 21140
rect 26936 21100 32588 21128
rect 26936 21088 26942 21100
rect 32582 21088 32588 21100
rect 32640 21088 32646 21140
rect 34606 21088 34612 21140
rect 34664 21128 34670 21140
rect 34885 21131 34943 21137
rect 34885 21128 34897 21131
rect 34664 21100 34897 21128
rect 34664 21088 34670 21100
rect 34885 21097 34897 21100
rect 34931 21097 34943 21131
rect 34885 21091 34943 21097
rect 35544 21100 35747 21128
rect 20036 21032 24624 21060
rect 27893 21063 27951 21069
rect 20036 21020 20042 21032
rect 27893 21029 27905 21063
rect 27939 21060 27951 21063
rect 28626 21060 28632 21072
rect 27939 21032 28632 21060
rect 27939 21029 27951 21032
rect 27893 21023 27951 21029
rect 28626 21020 28632 21032
rect 28684 21020 28690 21072
rect 29086 21020 29092 21072
rect 29144 21060 29150 21072
rect 35544 21060 35572 21100
rect 29144 21032 35572 21060
rect 35719 21060 35747 21100
rect 35894 21088 35900 21140
rect 35952 21128 35958 21140
rect 37550 21128 37556 21140
rect 35952 21100 37556 21128
rect 35952 21088 35958 21100
rect 37550 21088 37556 21100
rect 37608 21088 37614 21140
rect 38562 21088 38568 21140
rect 38620 21128 38626 21140
rect 40037 21131 40095 21137
rect 40037 21128 40049 21131
rect 38620 21100 40049 21128
rect 38620 21088 38626 21100
rect 40037 21097 40049 21100
rect 40083 21097 40095 21131
rect 43990 21128 43996 21140
rect 40037 21091 40095 21097
rect 40144 21100 42196 21128
rect 43951 21100 43996 21128
rect 35719 21032 38976 21060
rect 29144 21020 29150 21032
rect 20441 20995 20499 21001
rect 20441 20961 20453 20995
rect 20487 20992 20499 20995
rect 22370 20992 22376 21004
rect 20487 20964 22376 20992
rect 20487 20961 20499 20964
rect 20441 20955 20499 20961
rect 22370 20952 22376 20964
rect 22428 20952 22434 21004
rect 22649 20995 22707 21001
rect 22649 20961 22661 20995
rect 22695 20961 22707 20995
rect 27062 20992 27068 21004
rect 22649 20955 22707 20961
rect 23124 20964 24716 20992
rect 1857 20927 1915 20933
rect 1857 20893 1869 20927
rect 1903 20924 1915 20927
rect 13906 20924 13912 20936
rect 1903 20896 13912 20924
rect 1903 20893 1915 20896
rect 1857 20887 1915 20893
rect 13906 20884 13912 20896
rect 13964 20884 13970 20936
rect 22189 20927 22247 20933
rect 22189 20893 22201 20927
rect 22235 20924 22247 20927
rect 22664 20924 22692 20955
rect 23124 20933 23152 20964
rect 22235 20896 22692 20924
rect 23109 20927 23167 20933
rect 22235 20893 22247 20896
rect 22189 20887 22247 20893
rect 23109 20893 23121 20927
rect 23155 20893 23167 20927
rect 23842 20924 23848 20936
rect 23803 20896 23848 20924
rect 23109 20887 23167 20893
rect 20993 20859 21051 20865
rect 20993 20825 21005 20859
rect 21039 20856 21051 20859
rect 23124 20856 23152 20887
rect 23842 20884 23848 20896
rect 23900 20884 23906 20936
rect 24394 20924 24400 20936
rect 23952 20896 24400 20924
rect 21039 20828 23152 20856
rect 21039 20825 21051 20828
rect 20993 20819 21051 20825
rect 1670 20788 1676 20800
rect 1631 20760 1676 20788
rect 1670 20748 1676 20760
rect 1728 20748 1734 20800
rect 21450 20788 21456 20800
rect 21411 20760 21456 20788
rect 21450 20748 21456 20760
rect 21508 20788 21514 20800
rect 23952 20788 23980 20896
rect 24394 20884 24400 20896
rect 24452 20884 24458 20936
rect 24578 20924 24584 20936
rect 24539 20896 24584 20924
rect 24578 20884 24584 20896
rect 24636 20884 24642 20936
rect 24688 20924 24716 20964
rect 25976 20964 27068 20992
rect 25976 20924 26004 20964
rect 27062 20952 27068 20964
rect 27120 20992 27126 21004
rect 28534 20992 28540 21004
rect 27120 20964 27292 20992
rect 28495 20964 28540 20992
rect 27120 20952 27126 20964
rect 27157 20927 27215 20933
rect 27157 20924 27169 20927
rect 24688 20896 26004 20924
rect 26528 20896 27169 20924
rect 24826 20859 24884 20865
rect 24826 20825 24838 20859
rect 24872 20825 24884 20859
rect 24826 20819 24884 20825
rect 21508 20760 23980 20788
rect 24029 20791 24087 20797
rect 21508 20748 21514 20760
rect 24029 20757 24041 20791
rect 24075 20788 24087 20791
rect 24841 20788 24869 20819
rect 26528 20800 26556 20896
rect 27157 20893 27169 20896
rect 27203 20893 27215 20927
rect 27264 20924 27292 20964
rect 28534 20952 28540 20964
rect 28592 20952 28598 21004
rect 31294 20992 31300 21004
rect 28644 20964 31300 20992
rect 28644 20924 28672 20964
rect 31294 20952 31300 20964
rect 31352 20952 31358 21004
rect 32306 20992 32312 21004
rect 32267 20964 32312 20992
rect 32306 20952 32312 20964
rect 32364 20952 32370 21004
rect 33778 20992 33784 21004
rect 33739 20964 33784 20992
rect 33778 20952 33784 20964
rect 33836 20952 33842 21004
rect 35342 20992 35348 21004
rect 33888 20964 35348 20992
rect 30006 20924 30012 20936
rect 27264 20896 28672 20924
rect 28920 20896 30012 20924
rect 27157 20887 27215 20893
rect 24075 20760 24869 20788
rect 24075 20757 24087 20760
rect 24029 20751 24087 20757
rect 25130 20748 25136 20800
rect 25188 20788 25194 20800
rect 25961 20791 26019 20797
rect 25961 20788 25973 20791
rect 25188 20760 25973 20788
rect 25188 20748 25194 20760
rect 25961 20757 25973 20760
rect 26007 20788 26019 20791
rect 26510 20788 26516 20800
rect 26007 20760 26516 20788
rect 26007 20757 26019 20760
rect 25961 20751 26019 20757
rect 26510 20748 26516 20760
rect 26568 20748 26574 20800
rect 27172 20788 27200 20887
rect 28626 20856 28632 20868
rect 28587 20828 28632 20856
rect 28626 20816 28632 20828
rect 28684 20816 28690 20868
rect 28920 20856 28948 20896
rect 30006 20884 30012 20896
rect 30064 20884 30070 20936
rect 30282 20924 30288 20936
rect 30243 20896 30288 20924
rect 30282 20884 30288 20896
rect 30340 20884 30346 20936
rect 31849 20927 31907 20933
rect 31849 20893 31861 20927
rect 31895 20924 31907 20927
rect 32030 20924 32036 20936
rect 31895 20896 32036 20924
rect 31895 20893 31907 20896
rect 31849 20887 31907 20893
rect 32030 20884 32036 20896
rect 32088 20884 32094 20936
rect 32858 20884 32864 20936
rect 32916 20924 32922 20936
rect 33888 20924 33916 20964
rect 35342 20952 35348 20964
rect 35400 20952 35406 21004
rect 35529 20995 35587 21001
rect 35529 20961 35541 20995
rect 35575 20992 35587 20995
rect 35894 20992 35900 21004
rect 35575 20964 35900 20992
rect 35575 20961 35587 20964
rect 35529 20955 35587 20961
rect 35894 20952 35900 20964
rect 35952 20952 35958 21004
rect 36354 20952 36360 21004
rect 36412 20992 36418 21004
rect 36449 20995 36507 21001
rect 36449 20992 36461 20995
rect 36412 20964 36461 20992
rect 36412 20952 36418 20964
rect 36449 20961 36461 20964
rect 36495 20961 36507 20995
rect 36449 20955 36507 20961
rect 36998 20924 37004 20936
rect 32916 20896 33916 20924
rect 34624 20896 37004 20924
rect 32916 20884 32922 20896
rect 34624 20856 34652 20896
rect 36998 20884 37004 20896
rect 37056 20884 37062 20936
rect 38948 20933 38976 21032
rect 40144 20992 40172 21100
rect 42168 21069 42196 21100
rect 43990 21088 43996 21100
rect 44048 21088 44054 21140
rect 42153 21063 42211 21069
rect 42153 21029 42165 21063
rect 42199 21060 42211 21063
rect 54202 21060 54208 21072
rect 42199 21032 51074 21060
rect 54163 21032 54208 21060
rect 42199 21029 42211 21032
rect 42153 21023 42211 21029
rect 39224 20964 40172 20992
rect 39224 20933 39252 20964
rect 38933 20927 38991 20933
rect 38028 20896 38654 20924
rect 28736 20828 28948 20856
rect 29104 20828 34652 20856
rect 28736 20797 28764 20828
rect 29104 20797 29132 20828
rect 34698 20816 34704 20868
rect 34756 20856 34762 20868
rect 35253 20859 35311 20865
rect 35253 20856 35265 20859
rect 34756 20828 35265 20856
rect 34756 20816 34762 20828
rect 35253 20825 35265 20828
rect 35299 20856 35311 20859
rect 35710 20856 35716 20868
rect 35299 20828 35716 20856
rect 35299 20825 35311 20828
rect 35253 20819 35311 20825
rect 35710 20816 35716 20828
rect 35768 20816 35774 20868
rect 38028 20856 38056 20896
rect 38194 20856 38200 20868
rect 35820 20828 38056 20856
rect 38155 20828 38200 20856
rect 28721 20791 28779 20797
rect 28721 20788 28733 20791
rect 27172 20760 28733 20788
rect 28721 20757 28733 20760
rect 28767 20757 28779 20791
rect 28721 20751 28779 20757
rect 29089 20791 29147 20797
rect 29089 20757 29101 20791
rect 29135 20757 29147 20791
rect 29730 20788 29736 20800
rect 29691 20760 29736 20788
rect 29089 20751 29147 20757
rect 29730 20748 29736 20760
rect 29788 20748 29794 20800
rect 30190 20748 30196 20800
rect 30248 20788 30254 20800
rect 31205 20791 31263 20797
rect 31205 20788 31217 20791
rect 30248 20760 31217 20788
rect 30248 20748 30254 20760
rect 31205 20757 31217 20760
rect 31251 20757 31263 20791
rect 31205 20751 31263 20757
rect 32858 20748 32864 20800
rect 32916 20788 32922 20800
rect 32953 20791 33011 20797
rect 32953 20788 32965 20791
rect 32916 20760 32965 20788
rect 32916 20748 32922 20760
rect 32953 20757 32965 20760
rect 32999 20757 33011 20791
rect 32953 20751 33011 20757
rect 34333 20791 34391 20797
rect 34333 20757 34345 20791
rect 34379 20788 34391 20791
rect 34606 20788 34612 20800
rect 34379 20760 34612 20788
rect 34379 20757 34391 20760
rect 34333 20751 34391 20757
rect 34606 20748 34612 20760
rect 34664 20748 34670 20800
rect 34790 20748 34796 20800
rect 34848 20788 34854 20800
rect 35345 20791 35403 20797
rect 35345 20788 35357 20791
rect 34848 20760 35357 20788
rect 34848 20748 34854 20760
rect 35345 20757 35357 20760
rect 35391 20788 35403 20791
rect 35820 20788 35848 20828
rect 38194 20816 38200 20828
rect 38252 20816 38258 20868
rect 38626 20856 38654 20896
rect 38933 20893 38945 20927
rect 38979 20893 38991 20927
rect 38933 20887 38991 20893
rect 39209 20927 39267 20933
rect 39209 20893 39221 20927
rect 39255 20893 39267 20927
rect 39301 20927 39359 20933
rect 39301 20912 39313 20927
rect 39347 20912 39359 20927
rect 39209 20887 39267 20893
rect 38746 20856 38752 20868
rect 38626 20828 38752 20856
rect 38746 20816 38752 20828
rect 38804 20816 38810 20868
rect 39114 20856 39120 20868
rect 39075 20828 39120 20856
rect 39114 20816 39120 20828
rect 39172 20816 39178 20868
rect 39298 20860 39304 20912
rect 39356 20860 39362 20912
rect 40126 20884 40132 20936
rect 40184 20924 40190 20936
rect 40221 20927 40279 20933
rect 40221 20924 40233 20927
rect 40184 20896 40233 20924
rect 40184 20884 40190 20896
rect 40221 20893 40233 20896
rect 40267 20893 40279 20927
rect 40221 20887 40279 20893
rect 40678 20884 40684 20936
rect 40736 20924 40742 20936
rect 40773 20927 40831 20933
rect 40773 20924 40785 20927
rect 40736 20896 40785 20924
rect 40736 20884 40742 20896
rect 40773 20893 40785 20896
rect 40819 20893 40831 20927
rect 40773 20887 40831 20893
rect 42334 20884 42340 20936
rect 42392 20924 42398 20936
rect 42797 20927 42855 20933
rect 42797 20924 42809 20927
rect 42392 20896 42809 20924
rect 42392 20884 42398 20896
rect 42797 20893 42809 20896
rect 42843 20893 42855 20927
rect 43438 20924 43444 20936
rect 43399 20896 43444 20924
rect 42797 20887 42855 20893
rect 43438 20884 43444 20896
rect 43496 20884 43502 20936
rect 51046 20924 51074 21032
rect 54202 21020 54208 21032
rect 54260 21020 54266 21072
rect 54021 20927 54079 20933
rect 54021 20924 54033 20927
rect 51046 20896 54033 20924
rect 54021 20893 54033 20896
rect 54067 20893 54079 20927
rect 54021 20887 54079 20893
rect 41040 20859 41098 20865
rect 41040 20825 41052 20859
rect 41086 20856 41098 20859
rect 41086 20828 43300 20856
rect 41086 20825 41098 20828
rect 41040 20819 41098 20825
rect 35391 20760 35848 20788
rect 35391 20757 35403 20760
rect 35345 20751 35403 20757
rect 36538 20748 36544 20800
rect 36596 20788 36602 20800
rect 39298 20788 39304 20800
rect 36596 20760 39304 20788
rect 36596 20748 36602 20760
rect 39298 20748 39304 20760
rect 39356 20748 39362 20800
rect 39485 20791 39543 20797
rect 39485 20757 39497 20791
rect 39531 20788 39543 20791
rect 42242 20788 42248 20800
rect 39531 20760 42248 20788
rect 39531 20757 39543 20760
rect 39485 20751 39543 20757
rect 42242 20748 42248 20760
rect 42300 20748 42306 20800
rect 42613 20791 42671 20797
rect 42613 20757 42625 20791
rect 42659 20788 42671 20791
rect 42702 20788 42708 20800
rect 42659 20760 42708 20788
rect 42659 20757 42671 20760
rect 42613 20751 42671 20757
rect 42702 20748 42708 20760
rect 42760 20748 42766 20800
rect 43272 20797 43300 20828
rect 43257 20791 43315 20797
rect 43257 20757 43269 20791
rect 43303 20757 43315 20791
rect 53558 20788 53564 20800
rect 53519 20760 53564 20788
rect 43257 20751 43315 20757
rect 53558 20748 53564 20760
rect 53616 20748 53622 20800
rect 1104 20698 54832 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 54832 20698
rect 1104 20624 54832 20646
rect 22005 20587 22063 20593
rect 22005 20584 22017 20587
rect 6886 20556 22017 20584
rect 1857 20451 1915 20457
rect 1857 20417 1869 20451
rect 1903 20448 1915 20451
rect 2409 20451 2467 20457
rect 2409 20448 2421 20451
rect 1903 20420 2421 20448
rect 1903 20417 1915 20420
rect 1857 20411 1915 20417
rect 2409 20417 2421 20420
rect 2455 20448 2467 20451
rect 6886 20448 6914 20556
rect 22005 20553 22017 20556
rect 22051 20553 22063 20587
rect 22005 20547 22063 20553
rect 23569 20587 23627 20593
rect 23569 20553 23581 20587
rect 23615 20584 23627 20587
rect 23842 20584 23848 20596
rect 23615 20556 23848 20584
rect 23615 20553 23627 20556
rect 23569 20547 23627 20553
rect 23842 20544 23848 20556
rect 23900 20544 23906 20596
rect 24029 20587 24087 20593
rect 24029 20553 24041 20587
rect 24075 20553 24087 20587
rect 24029 20547 24087 20553
rect 20349 20519 20407 20525
rect 20349 20485 20361 20519
rect 20395 20516 20407 20519
rect 20901 20519 20959 20525
rect 20901 20516 20913 20519
rect 20395 20488 20913 20516
rect 20395 20485 20407 20488
rect 20349 20479 20407 20485
rect 20901 20485 20913 20488
rect 20947 20516 20959 20519
rect 20947 20488 22094 20516
rect 20947 20485 20959 20488
rect 20901 20479 20959 20485
rect 2455 20420 6914 20448
rect 19429 20451 19487 20457
rect 2455 20417 2467 20420
rect 2409 20411 2467 20417
rect 19429 20417 19441 20451
rect 19475 20448 19487 20451
rect 19610 20448 19616 20460
rect 19475 20420 19616 20448
rect 19475 20417 19487 20420
rect 19429 20411 19487 20417
rect 19610 20408 19616 20420
rect 19668 20408 19674 20460
rect 18966 20340 18972 20392
rect 19024 20380 19030 20392
rect 21450 20380 21456 20392
rect 19024 20352 21456 20380
rect 19024 20340 19030 20352
rect 21450 20340 21456 20352
rect 21508 20340 21514 20392
rect 22066 20380 22094 20488
rect 22186 20448 22192 20460
rect 22147 20420 22192 20448
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 23385 20451 23443 20457
rect 23385 20417 23397 20451
rect 23431 20448 23443 20451
rect 24044 20448 24072 20547
rect 24394 20544 24400 20596
rect 24452 20584 24458 20596
rect 24489 20587 24547 20593
rect 24489 20584 24501 20587
rect 24452 20556 24501 20584
rect 24452 20544 24458 20556
rect 24489 20553 24501 20556
rect 24535 20553 24547 20587
rect 24489 20547 24547 20553
rect 26510 20544 26516 20596
rect 26568 20584 26574 20596
rect 26605 20587 26663 20593
rect 26605 20584 26617 20587
rect 26568 20556 26617 20584
rect 26568 20544 26574 20556
rect 26605 20553 26617 20556
rect 26651 20553 26663 20587
rect 27154 20584 27160 20596
rect 27115 20556 27160 20584
rect 26605 20547 26663 20553
rect 27154 20544 27160 20556
rect 27212 20544 27218 20596
rect 27798 20584 27804 20596
rect 27759 20556 27804 20584
rect 27798 20544 27804 20556
rect 27856 20544 27862 20596
rect 28810 20544 28816 20596
rect 28868 20584 28874 20596
rect 29638 20584 29644 20596
rect 28868 20556 29644 20584
rect 28868 20544 28874 20556
rect 29638 20544 29644 20556
rect 29696 20544 29702 20596
rect 29733 20587 29791 20593
rect 29733 20553 29745 20587
rect 29779 20584 29791 20587
rect 30282 20584 30288 20596
rect 29779 20556 30288 20584
rect 29779 20553 29791 20556
rect 29733 20547 29791 20553
rect 30282 20544 30288 20556
rect 30340 20544 30346 20596
rect 36081 20587 36139 20593
rect 36081 20553 36093 20587
rect 36127 20584 36139 20587
rect 37458 20584 37464 20596
rect 36127 20556 37464 20584
rect 36127 20553 36139 20556
rect 36081 20547 36139 20553
rect 37458 20544 37464 20556
rect 37516 20544 37522 20596
rect 39485 20587 39543 20593
rect 39485 20553 39497 20587
rect 39531 20584 39543 20587
rect 40678 20584 40684 20596
rect 39531 20556 40684 20584
rect 39531 20553 39543 20556
rect 39485 20547 39543 20553
rect 40678 20544 40684 20556
rect 40736 20544 40742 20596
rect 42794 20584 42800 20596
rect 40788 20556 42800 20584
rect 24854 20476 24860 20528
rect 24912 20516 24918 20528
rect 25774 20516 25780 20528
rect 24912 20488 25780 20516
rect 24912 20476 24918 20488
rect 23431 20420 24072 20448
rect 24397 20451 24455 20457
rect 23431 20417 23443 20420
rect 23385 20411 23443 20417
rect 24397 20417 24409 20451
rect 24443 20448 24455 20451
rect 25130 20448 25136 20460
rect 24443 20420 25136 20448
rect 24443 20417 24455 20420
rect 24397 20411 24455 20417
rect 25130 20408 25136 20420
rect 25188 20408 25194 20460
rect 25240 20457 25268 20488
rect 25774 20476 25780 20488
rect 25832 20516 25838 20528
rect 25832 20488 27456 20516
rect 25832 20476 25838 20488
rect 25225 20451 25283 20457
rect 25225 20417 25237 20451
rect 25271 20417 25283 20451
rect 25225 20411 25283 20417
rect 25314 20408 25320 20460
rect 25372 20448 25378 20460
rect 25481 20451 25539 20457
rect 25481 20448 25493 20451
rect 25372 20420 25493 20448
rect 25372 20408 25378 20420
rect 25481 20417 25493 20420
rect 25527 20417 25539 20451
rect 25481 20411 25539 20417
rect 26602 20408 26608 20460
rect 26660 20448 26666 20460
rect 27157 20451 27215 20457
rect 27157 20448 27169 20451
rect 26660 20420 27169 20448
rect 26660 20408 26666 20420
rect 27157 20417 27169 20420
rect 27203 20417 27215 20451
rect 27157 20411 27215 20417
rect 27341 20451 27399 20457
rect 27341 20417 27353 20451
rect 27387 20417 27399 20451
rect 27428 20448 27456 20488
rect 28828 20488 29224 20516
rect 28828 20448 28856 20488
rect 29196 20460 29224 20488
rect 29822 20476 29828 20528
rect 29880 20516 29886 20528
rect 30098 20516 30104 20528
rect 29880 20488 30104 20516
rect 29880 20476 29886 20488
rect 30098 20476 30104 20488
rect 30156 20516 30162 20528
rect 40788 20525 40816 20556
rect 42794 20544 42800 20556
rect 42852 20584 42858 20596
rect 43165 20587 43223 20593
rect 43165 20584 43177 20587
rect 42852 20556 43177 20584
rect 42852 20544 42858 20556
rect 43165 20553 43177 20556
rect 43211 20584 43223 20587
rect 44269 20587 44327 20593
rect 44269 20584 44281 20587
rect 43211 20556 44281 20584
rect 43211 20553 43223 20556
rect 43165 20547 43223 20553
rect 44269 20553 44281 20556
rect 44315 20553 44327 20587
rect 44269 20547 44327 20553
rect 40773 20519 40831 20525
rect 30156 20488 30236 20516
rect 30156 20476 30162 20488
rect 27428 20420 28856 20448
rect 28925 20451 28983 20457
rect 27341 20411 27399 20417
rect 28925 20417 28937 20451
rect 28971 20448 28983 20451
rect 29086 20448 29092 20460
rect 28971 20420 29092 20448
rect 28971 20417 28983 20420
rect 28925 20411 28983 20417
rect 23201 20383 23259 20389
rect 23201 20380 23213 20383
rect 22066 20352 23213 20380
rect 23201 20349 23213 20352
rect 23247 20380 23259 20383
rect 23474 20380 23480 20392
rect 23247 20352 23480 20380
rect 23247 20349 23259 20352
rect 23201 20343 23259 20349
rect 23474 20340 23480 20352
rect 23532 20380 23538 20392
rect 24210 20380 24216 20392
rect 23532 20352 24216 20380
rect 23532 20340 23538 20352
rect 24210 20340 24216 20352
rect 24268 20340 24274 20392
rect 24673 20383 24731 20389
rect 24673 20349 24685 20383
rect 24719 20380 24731 20383
rect 25038 20380 25044 20392
rect 24719 20352 25044 20380
rect 24719 20349 24731 20352
rect 24673 20343 24731 20349
rect 25038 20340 25044 20352
rect 25096 20340 25102 20392
rect 26786 20340 26792 20392
rect 26844 20380 26850 20392
rect 27356 20380 27384 20411
rect 29086 20408 29092 20420
rect 29144 20408 29150 20460
rect 29178 20408 29184 20460
rect 29236 20448 29242 20460
rect 29236 20420 29281 20448
rect 29236 20408 29242 20420
rect 29638 20408 29644 20460
rect 29696 20448 29702 20460
rect 29917 20451 29975 20457
rect 29917 20448 29929 20451
rect 29696 20420 29929 20448
rect 29696 20408 29702 20420
rect 29917 20417 29929 20420
rect 29963 20417 29975 20451
rect 29917 20411 29975 20417
rect 30006 20408 30012 20460
rect 30064 20448 30070 20460
rect 30208 20457 30236 20488
rect 40773 20485 40785 20519
rect 40819 20485 40831 20519
rect 54021 20519 54079 20525
rect 54021 20516 54033 20519
rect 40773 20479 40831 20485
rect 40880 20488 54033 20516
rect 30193 20451 30251 20457
rect 30064 20420 30109 20448
rect 30064 20408 30070 20420
rect 30193 20417 30205 20451
rect 30239 20417 30251 20451
rect 30193 20411 30251 20417
rect 34146 20408 34152 20460
rect 34204 20448 34210 20460
rect 34422 20448 34428 20460
rect 34204 20420 34428 20448
rect 34204 20408 34210 20420
rect 34422 20408 34428 20420
rect 34480 20408 34486 20460
rect 34606 20408 34612 20460
rect 34664 20448 34670 20460
rect 34957 20451 35015 20457
rect 34957 20448 34969 20451
rect 34664 20420 34969 20448
rect 34664 20408 34670 20420
rect 34957 20417 34969 20420
rect 35003 20417 35015 20451
rect 34957 20411 35015 20417
rect 35342 20408 35348 20460
rect 35400 20448 35406 20460
rect 36722 20448 36728 20460
rect 35400 20420 35894 20448
rect 36683 20420 36728 20448
rect 35400 20408 35406 20420
rect 27522 20380 27528 20392
rect 26844 20352 27528 20380
rect 26844 20340 26850 20352
rect 27522 20340 27528 20352
rect 27580 20340 27586 20392
rect 30101 20383 30159 20389
rect 30101 20380 30113 20383
rect 30024 20352 30113 20380
rect 30024 20324 30052 20352
rect 30101 20349 30113 20352
rect 30147 20349 30159 20383
rect 30101 20343 30159 20349
rect 31481 20383 31539 20389
rect 31481 20349 31493 20383
rect 31527 20380 31539 20383
rect 32214 20380 32220 20392
rect 31527 20352 32220 20380
rect 31527 20349 31539 20352
rect 31481 20343 31539 20349
rect 32214 20340 32220 20352
rect 32272 20340 32278 20392
rect 32309 20383 32367 20389
rect 32309 20349 32321 20383
rect 32355 20349 32367 20383
rect 33594 20380 33600 20392
rect 33555 20352 33600 20380
rect 32309 20343 32367 20349
rect 20530 20272 20536 20324
rect 20588 20312 20594 20324
rect 21361 20315 21419 20321
rect 21361 20312 21373 20315
rect 20588 20284 21373 20312
rect 20588 20272 20594 20284
rect 21361 20281 21373 20284
rect 21407 20312 21419 20315
rect 22741 20315 22799 20321
rect 22741 20312 22753 20315
rect 21407 20284 22753 20312
rect 21407 20281 21419 20284
rect 21361 20275 21419 20281
rect 22741 20281 22753 20284
rect 22787 20312 22799 20315
rect 22830 20312 22836 20324
rect 22787 20284 22836 20312
rect 22787 20281 22799 20284
rect 22741 20275 22799 20281
rect 22830 20272 22836 20284
rect 22888 20272 22894 20324
rect 30006 20272 30012 20324
rect 30064 20272 30070 20324
rect 30466 20272 30472 20324
rect 30524 20312 30530 20324
rect 32324 20312 32352 20343
rect 33594 20340 33600 20352
rect 33652 20340 33658 20392
rect 34330 20340 34336 20392
rect 34388 20380 34394 20392
rect 34701 20383 34759 20389
rect 34701 20380 34713 20383
rect 34388 20352 34713 20380
rect 34388 20340 34394 20352
rect 34701 20349 34713 20352
rect 34747 20349 34759 20383
rect 35866 20380 35894 20420
rect 36722 20408 36728 20420
rect 36780 20408 36786 20460
rect 37182 20408 37188 20460
rect 37240 20448 37246 20460
rect 40880 20448 40908 20488
rect 54021 20485 54033 20488
rect 54067 20485 54079 20519
rect 54202 20516 54208 20528
rect 54163 20488 54208 20516
rect 54021 20479 54079 20485
rect 54202 20476 54208 20488
rect 54260 20476 54266 20528
rect 37240 20420 40908 20448
rect 41371 20451 41429 20457
rect 37240 20408 37246 20420
rect 41371 20417 41383 20451
rect 41417 20417 41429 20451
rect 41506 20448 41512 20460
rect 41467 20420 41512 20448
rect 41371 20411 41429 20417
rect 36541 20383 36599 20389
rect 36541 20380 36553 20383
rect 35866 20352 36553 20380
rect 34701 20343 34759 20349
rect 36541 20349 36553 20352
rect 36587 20380 36599 20383
rect 37090 20380 37096 20392
rect 36587 20352 37096 20380
rect 36587 20349 36599 20352
rect 36541 20343 36599 20349
rect 37090 20340 37096 20352
rect 37148 20340 37154 20392
rect 37553 20383 37611 20389
rect 37553 20349 37565 20383
rect 37599 20380 37611 20383
rect 38746 20380 38752 20392
rect 37599 20352 38752 20380
rect 37599 20349 37611 20352
rect 37553 20343 37611 20349
rect 38746 20340 38752 20352
rect 38804 20340 38810 20392
rect 38930 20340 38936 20392
rect 38988 20380 38994 20392
rect 38988 20352 39620 20380
rect 38988 20340 38994 20352
rect 30524 20284 32352 20312
rect 32953 20315 33011 20321
rect 30524 20272 30530 20284
rect 32953 20281 32965 20315
rect 32999 20312 33011 20315
rect 36814 20312 36820 20324
rect 32999 20284 34744 20312
rect 32999 20281 33011 20284
rect 32953 20275 33011 20281
rect 1670 20244 1676 20256
rect 1631 20216 1676 20244
rect 1670 20204 1676 20216
rect 1728 20204 1734 20256
rect 19242 20244 19248 20256
rect 19203 20216 19248 20244
rect 19242 20204 19248 20216
rect 19300 20204 19306 20256
rect 20622 20204 20628 20256
rect 20680 20244 20686 20256
rect 29454 20244 29460 20256
rect 20680 20216 29460 20244
rect 20680 20204 20686 20216
rect 29454 20204 29460 20216
rect 29512 20204 29518 20256
rect 29638 20204 29644 20256
rect 29696 20244 29702 20256
rect 30837 20247 30895 20253
rect 30837 20244 30849 20247
rect 29696 20216 30849 20244
rect 29696 20204 29702 20216
rect 30837 20213 30849 20216
rect 30883 20213 30895 20247
rect 34238 20244 34244 20256
rect 34199 20216 34244 20244
rect 30837 20207 30895 20213
rect 34238 20204 34244 20216
rect 34296 20204 34302 20256
rect 34716 20244 34744 20284
rect 36004 20284 36820 20312
rect 36004 20244 36032 20284
rect 36814 20272 36820 20284
rect 36872 20272 36878 20324
rect 36909 20315 36967 20321
rect 36909 20281 36921 20315
rect 36955 20312 36967 20315
rect 39390 20312 39396 20324
rect 36955 20284 39396 20312
rect 36955 20281 36967 20284
rect 36909 20275 36967 20281
rect 39390 20272 39396 20284
rect 39448 20272 39454 20324
rect 34716 20216 36032 20244
rect 38105 20247 38163 20253
rect 38105 20213 38117 20247
rect 38151 20244 38163 20247
rect 39482 20244 39488 20256
rect 38151 20216 39488 20244
rect 38151 20213 38163 20216
rect 38105 20207 38163 20213
rect 39482 20204 39488 20216
rect 39540 20204 39546 20256
rect 39592 20244 39620 20352
rect 40494 20340 40500 20392
rect 40552 20380 40558 20392
rect 41386 20380 41414 20411
rect 41506 20408 41512 20420
rect 41564 20408 41570 20460
rect 41601 20451 41659 20457
rect 41601 20417 41613 20451
rect 41647 20417 41659 20451
rect 41782 20448 41788 20460
rect 41743 20420 41788 20448
rect 41601 20411 41659 20417
rect 40552 20352 41414 20380
rect 40552 20340 40558 20352
rect 41322 20272 41328 20324
rect 41380 20312 41386 20324
rect 41616 20312 41644 20411
rect 41782 20408 41788 20420
rect 41840 20408 41846 20460
rect 43714 20448 43720 20460
rect 43675 20420 43720 20448
rect 43714 20408 43720 20420
rect 43772 20408 43778 20460
rect 53282 20448 53288 20460
rect 53243 20420 53288 20448
rect 53282 20408 53288 20420
rect 53340 20408 53346 20460
rect 53469 20451 53527 20457
rect 53469 20417 53481 20451
rect 53515 20448 53527 20451
rect 53558 20448 53564 20460
rect 53515 20420 53564 20448
rect 53515 20417 53527 20420
rect 53469 20411 53527 20417
rect 53558 20408 53564 20420
rect 53616 20408 53622 20460
rect 41380 20284 41644 20312
rect 41380 20272 41386 20284
rect 41233 20247 41291 20253
rect 41233 20244 41245 20247
rect 39592 20216 41245 20244
rect 41233 20213 41245 20216
rect 41279 20213 41291 20247
rect 42610 20244 42616 20256
rect 42571 20216 42616 20244
rect 41233 20207 41291 20213
rect 42610 20204 42616 20216
rect 42668 20204 42674 20256
rect 1104 20154 54832 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 54832 20154
rect 1104 20080 54832 20102
rect 2409 20043 2467 20049
rect 2409 20009 2421 20043
rect 2455 20040 2467 20043
rect 2498 20040 2504 20052
rect 2455 20012 2504 20040
rect 2455 20009 2467 20012
rect 2409 20003 2467 20009
rect 1857 19839 1915 19845
rect 1857 19805 1869 19839
rect 1903 19836 1915 19839
rect 2424 19836 2452 20003
rect 2498 20000 2504 20012
rect 2556 20000 2562 20052
rect 19610 20040 19616 20052
rect 19571 20012 19616 20040
rect 19610 20000 19616 20012
rect 19668 20000 19674 20052
rect 21266 20000 21272 20052
rect 21324 20040 21330 20052
rect 24581 20043 24639 20049
rect 21324 20012 22600 20040
rect 21324 20000 21330 20012
rect 20806 19932 20812 19984
rect 20864 19972 20870 19984
rect 21910 19972 21916 19984
rect 20864 19944 21916 19972
rect 20864 19932 20870 19944
rect 21910 19932 21916 19944
rect 21968 19932 21974 19984
rect 22005 19975 22063 19981
rect 22005 19941 22017 19975
rect 22051 19941 22063 19975
rect 22005 19935 22063 19941
rect 15838 19864 15844 19916
rect 15896 19904 15902 19916
rect 20162 19904 20168 19916
rect 15896 19876 20168 19904
rect 15896 19864 15902 19876
rect 20162 19864 20168 19876
rect 20220 19864 20226 19916
rect 20257 19907 20315 19913
rect 20257 19873 20269 19907
rect 20303 19904 20315 19907
rect 21266 19904 21272 19916
rect 20303 19876 21272 19904
rect 20303 19873 20315 19876
rect 20257 19867 20315 19873
rect 21266 19864 21272 19876
rect 21324 19864 21330 19916
rect 14458 19836 14464 19848
rect 1903 19808 2452 19836
rect 14419 19808 14464 19836
rect 1903 19805 1915 19808
rect 1857 19799 1915 19805
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 19978 19836 19984 19848
rect 19939 19808 19984 19836
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 21361 19839 21419 19845
rect 21361 19805 21373 19839
rect 21407 19836 21419 19839
rect 22020 19836 22048 19935
rect 22572 19913 22600 20012
rect 24581 20009 24593 20043
rect 24627 20040 24639 20043
rect 24762 20040 24768 20052
rect 24627 20012 24768 20040
rect 24627 20009 24639 20012
rect 24581 20003 24639 20009
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 26142 20000 26148 20052
rect 26200 20040 26206 20052
rect 27157 20043 27215 20049
rect 27157 20040 27169 20043
rect 26200 20012 27169 20040
rect 26200 20000 26206 20012
rect 27157 20009 27169 20012
rect 27203 20009 27215 20043
rect 27157 20003 27215 20009
rect 27614 20000 27620 20052
rect 27672 20040 27678 20052
rect 30006 20040 30012 20052
rect 27672 20012 30012 20040
rect 27672 20000 27678 20012
rect 30006 20000 30012 20012
rect 30064 20000 30070 20052
rect 30852 20012 32168 20040
rect 27985 19975 28043 19981
rect 27985 19941 27997 19975
rect 28031 19972 28043 19975
rect 29730 19972 29736 19984
rect 28031 19944 29736 19972
rect 28031 19941 28043 19944
rect 27985 19935 28043 19941
rect 29730 19932 29736 19944
rect 29788 19932 29794 19984
rect 30852 19972 30880 20012
rect 30024 19944 30880 19972
rect 22557 19907 22615 19913
rect 22557 19873 22569 19907
rect 22603 19873 22615 19907
rect 22557 19867 22615 19873
rect 22830 19864 22836 19916
rect 22888 19904 22894 19916
rect 23477 19907 23535 19913
rect 23477 19904 23489 19907
rect 22888 19876 23489 19904
rect 22888 19864 22894 19876
rect 23477 19873 23489 19876
rect 23523 19904 23535 19907
rect 24029 19907 24087 19913
rect 24029 19904 24041 19907
rect 23523 19876 24041 19904
rect 23523 19873 23535 19876
rect 23477 19867 23535 19873
rect 24029 19873 24041 19876
rect 24075 19904 24087 19907
rect 24854 19904 24860 19916
rect 24075 19876 24860 19904
rect 24075 19873 24087 19876
rect 24029 19867 24087 19873
rect 24854 19864 24860 19876
rect 24912 19864 24918 19916
rect 25130 19904 25136 19916
rect 25091 19876 25136 19904
rect 25130 19864 25136 19876
rect 25188 19864 25194 19916
rect 25774 19904 25780 19916
rect 25735 19876 25780 19904
rect 25774 19864 25780 19876
rect 25832 19864 25838 19916
rect 28077 19907 28135 19913
rect 28077 19873 28089 19907
rect 28123 19904 28135 19907
rect 28537 19907 28595 19913
rect 28537 19904 28549 19907
rect 28123 19876 28549 19904
rect 28123 19873 28135 19876
rect 28077 19867 28135 19873
rect 28537 19873 28549 19876
rect 28583 19873 28595 19907
rect 28537 19867 28595 19873
rect 29178 19864 29184 19916
rect 29236 19904 29242 19916
rect 30024 19904 30052 19944
rect 30852 19916 30880 19944
rect 29236 19876 30052 19904
rect 30101 19907 30159 19913
rect 29236 19864 29242 19876
rect 30101 19873 30113 19907
rect 30147 19904 30159 19907
rect 30282 19904 30288 19916
rect 30147 19876 30288 19904
rect 30147 19873 30159 19876
rect 30101 19867 30159 19873
rect 30282 19864 30288 19876
rect 30340 19864 30346 19916
rect 30834 19904 30840 19916
rect 30747 19876 30840 19904
rect 30834 19864 30840 19876
rect 30892 19864 30898 19916
rect 22373 19839 22431 19845
rect 22373 19836 22385 19839
rect 21407 19808 22048 19836
rect 22204 19808 22385 19836
rect 21407 19805 21419 19808
rect 21361 19799 21419 19805
rect 18877 19771 18935 19777
rect 18877 19737 18889 19771
rect 18923 19768 18935 19771
rect 22204 19768 22232 19808
rect 22373 19805 22385 19808
rect 22419 19836 22431 19839
rect 27617 19839 27675 19845
rect 22419 19808 26234 19836
rect 22419 19805 22431 19808
rect 22373 19799 22431 19805
rect 18923 19740 22232 19768
rect 18923 19737 18935 19740
rect 18877 19731 18935 19737
rect 22278 19728 22284 19780
rect 22336 19768 22342 19780
rect 26050 19777 26056 19780
rect 22465 19771 22523 19777
rect 22465 19768 22477 19771
rect 22336 19740 22477 19768
rect 22336 19728 22342 19740
rect 22465 19737 22477 19740
rect 22511 19737 22523 19771
rect 22465 19731 22523 19737
rect 24949 19771 25007 19777
rect 24949 19737 24961 19771
rect 24995 19768 25007 19771
rect 24995 19740 26004 19768
rect 24995 19737 25007 19740
rect 24949 19731 25007 19737
rect 1670 19700 1676 19712
rect 1631 19672 1676 19700
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 14274 19700 14280 19712
rect 14235 19672 14280 19700
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 20070 19700 20076 19712
rect 20031 19672 20076 19700
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 20806 19700 20812 19712
rect 20767 19672 20812 19700
rect 20806 19660 20812 19672
rect 20864 19660 20870 19712
rect 21542 19700 21548 19712
rect 21503 19672 21548 19700
rect 21542 19660 21548 19672
rect 21600 19660 21606 19712
rect 22094 19660 22100 19712
rect 22152 19700 22158 19712
rect 25038 19700 25044 19712
rect 22152 19672 25044 19700
rect 22152 19660 22158 19672
rect 25038 19660 25044 19672
rect 25096 19660 25102 19712
rect 25976 19700 26004 19740
rect 26044 19731 26056 19777
rect 26108 19768 26114 19780
rect 26206 19768 26234 19808
rect 27617 19805 27629 19839
rect 27663 19836 27675 19839
rect 27798 19836 27804 19848
rect 27663 19808 27804 19836
rect 27663 19805 27675 19808
rect 27617 19799 27675 19805
rect 27798 19796 27804 19808
rect 27856 19796 27862 19848
rect 28442 19796 28448 19848
rect 28500 19836 28506 19848
rect 29822 19836 29828 19848
rect 28500 19808 29828 19836
rect 28500 19796 28506 19808
rect 29822 19796 29828 19808
rect 29880 19796 29886 19848
rect 30009 19839 30067 19845
rect 30009 19805 30021 19839
rect 30055 19836 30067 19839
rect 30742 19836 30748 19848
rect 30055 19808 30748 19836
rect 30055 19805 30067 19808
rect 30009 19799 30067 19805
rect 30742 19796 30748 19808
rect 30800 19796 30806 19848
rect 31110 19845 31116 19848
rect 31104 19799 31116 19845
rect 31168 19836 31174 19848
rect 32140 19836 32168 20012
rect 32306 20000 32312 20052
rect 32364 20040 32370 20052
rect 32677 20043 32735 20049
rect 32677 20040 32689 20043
rect 32364 20012 32689 20040
rect 32364 20000 32370 20012
rect 32677 20009 32689 20012
rect 32723 20009 32735 20043
rect 32677 20003 32735 20009
rect 34885 20043 34943 20049
rect 34885 20009 34897 20043
rect 34931 20040 34943 20043
rect 35526 20040 35532 20052
rect 34931 20012 35532 20040
rect 34931 20009 34943 20012
rect 34885 20003 34943 20009
rect 35526 20000 35532 20012
rect 35584 20000 35590 20052
rect 39301 20043 39359 20049
rect 39301 20040 39313 20043
rect 37292 20012 39313 20040
rect 32217 19975 32275 19981
rect 32217 19941 32229 19975
rect 32263 19972 32275 19975
rect 32490 19972 32496 19984
rect 32263 19944 32496 19972
rect 32263 19941 32275 19944
rect 32217 19935 32275 19941
rect 32490 19932 32496 19944
rect 32548 19932 32554 19984
rect 37292 19904 37320 20012
rect 39301 20009 39313 20012
rect 39347 20009 39359 20043
rect 39301 20003 39359 20009
rect 39390 20000 39396 20052
rect 39448 20040 39454 20052
rect 42058 20040 42064 20052
rect 39448 20012 42064 20040
rect 39448 20000 39454 20012
rect 42058 20000 42064 20012
rect 42116 20000 42122 20052
rect 42429 20043 42487 20049
rect 42429 20009 42441 20043
rect 42475 20040 42487 20043
rect 43438 20040 43444 20052
rect 42475 20012 43444 20040
rect 42475 20009 42487 20012
rect 42429 20003 42487 20009
rect 43438 20000 43444 20012
rect 43496 20000 43502 20052
rect 54202 20040 54208 20052
rect 54163 20012 54208 20040
rect 54202 20000 54208 20012
rect 54260 20000 54266 20052
rect 37458 19972 37464 19984
rect 37419 19944 37464 19972
rect 37458 19932 37464 19944
rect 37516 19972 37522 19984
rect 37826 19972 37832 19984
rect 37516 19944 37832 19972
rect 37516 19932 37522 19944
rect 37826 19932 37832 19944
rect 37884 19932 37890 19984
rect 53558 19972 53564 19984
rect 53519 19944 53564 19972
rect 53558 19932 53564 19944
rect 53616 19932 53622 19984
rect 38838 19904 38844 19916
rect 36740 19876 37320 19904
rect 38799 19876 38844 19904
rect 34057 19839 34115 19845
rect 34057 19836 34069 19839
rect 31168 19808 31204 19836
rect 32140 19808 34069 19836
rect 31110 19796 31116 19799
rect 31168 19796 31174 19808
rect 34057 19805 34069 19808
rect 34103 19836 34115 19839
rect 34330 19836 34336 19848
rect 34103 19808 34336 19836
rect 34103 19805 34115 19808
rect 34057 19799 34115 19805
rect 34330 19796 34336 19808
rect 34388 19836 34394 19848
rect 36262 19836 36268 19848
rect 34388 19808 36268 19836
rect 34388 19796 34394 19808
rect 36262 19796 36268 19808
rect 36320 19796 36326 19848
rect 33812 19771 33870 19777
rect 26108 19740 26144 19768
rect 26206 19740 31064 19768
rect 26050 19728 26056 19731
rect 26108 19728 26114 19740
rect 26142 19700 26148 19712
rect 25976 19672 26148 19700
rect 26142 19660 26148 19672
rect 26200 19660 26206 19712
rect 29181 19703 29239 19709
rect 29181 19669 29193 19703
rect 29227 19700 29239 19703
rect 29546 19700 29552 19712
rect 29227 19672 29552 19700
rect 29227 19669 29239 19672
rect 29181 19663 29239 19669
rect 29546 19660 29552 19672
rect 29604 19660 29610 19712
rect 30282 19660 30288 19712
rect 30340 19700 30346 19712
rect 30377 19703 30435 19709
rect 30377 19700 30389 19703
rect 30340 19672 30389 19700
rect 30340 19660 30346 19672
rect 30377 19669 30389 19672
rect 30423 19669 30435 19703
rect 31036 19700 31064 19740
rect 33812 19737 33824 19771
rect 33858 19768 33870 19771
rect 36020 19771 36078 19777
rect 33858 19740 35296 19768
rect 33858 19737 33870 19740
rect 33812 19731 33870 19737
rect 34790 19700 34796 19712
rect 31036 19672 34796 19700
rect 30377 19663 30435 19669
rect 34790 19660 34796 19672
rect 34848 19660 34854 19712
rect 35268 19700 35296 19740
rect 36020 19737 36032 19771
rect 36066 19768 36078 19771
rect 36740 19768 36768 19876
rect 38838 19864 38844 19876
rect 38896 19864 38902 19916
rect 42061 19907 42119 19913
rect 42061 19904 42073 19907
rect 39316 19876 40632 19904
rect 36814 19796 36820 19848
rect 36872 19836 36878 19848
rect 36909 19839 36967 19845
rect 36909 19836 36921 19839
rect 36872 19808 36921 19836
rect 36872 19796 36878 19808
rect 36909 19805 36921 19808
rect 36955 19805 36967 19839
rect 36909 19799 36967 19805
rect 36998 19796 37004 19848
rect 37056 19836 37062 19848
rect 39316 19836 39344 19876
rect 39482 19836 39488 19848
rect 37056 19808 39344 19836
rect 39443 19808 39488 19836
rect 37056 19796 37062 19808
rect 39482 19796 39488 19808
rect 39540 19796 39546 19848
rect 36066 19740 36768 19768
rect 38596 19771 38654 19777
rect 36066 19737 36078 19740
rect 36020 19731 36078 19737
rect 38596 19737 38608 19771
rect 38642 19768 38654 19771
rect 40310 19768 40316 19780
rect 38642 19740 40316 19768
rect 38642 19737 38654 19740
rect 38596 19731 38654 19737
rect 40310 19728 40316 19740
rect 40368 19728 40374 19780
rect 40604 19768 40632 19876
rect 41524 19876 42073 19904
rect 41138 19768 41144 19780
rect 40604 19740 41144 19768
rect 41138 19728 41144 19740
rect 41196 19728 41202 19780
rect 41414 19777 41420 19780
rect 41356 19771 41420 19777
rect 41356 19737 41368 19771
rect 41402 19737 41420 19771
rect 41356 19731 41420 19737
rect 41414 19728 41420 19731
rect 41472 19728 41478 19780
rect 36725 19703 36783 19709
rect 36725 19700 36737 19703
rect 35268 19672 36737 19700
rect 36725 19669 36737 19672
rect 36771 19669 36783 19703
rect 36725 19663 36783 19669
rect 38102 19660 38108 19712
rect 38160 19700 38166 19712
rect 40126 19700 40132 19712
rect 38160 19672 40132 19700
rect 38160 19660 38166 19672
rect 40126 19660 40132 19672
rect 40184 19660 40190 19712
rect 40221 19703 40279 19709
rect 40221 19669 40233 19703
rect 40267 19700 40279 19703
rect 40770 19700 40776 19712
rect 40267 19672 40776 19700
rect 40267 19669 40279 19672
rect 40221 19663 40279 19669
rect 40770 19660 40776 19672
rect 40828 19660 40834 19712
rect 40954 19660 40960 19712
rect 41012 19700 41018 19712
rect 41524 19700 41552 19876
rect 42061 19873 42073 19876
rect 42107 19873 42119 19907
rect 42061 19867 42119 19873
rect 41601 19839 41659 19845
rect 41601 19805 41613 19839
rect 41647 19805 41659 19839
rect 42242 19836 42248 19848
rect 42203 19808 42248 19836
rect 41601 19799 41659 19805
rect 41616 19768 41644 19799
rect 42242 19796 42248 19808
rect 42300 19796 42306 19848
rect 44726 19796 44732 19848
rect 44784 19836 44790 19848
rect 54021 19839 54079 19845
rect 54021 19836 54033 19839
rect 44784 19808 54033 19836
rect 44784 19796 44790 19808
rect 54021 19805 54033 19808
rect 54067 19805 54079 19839
rect 54021 19799 54079 19805
rect 42702 19768 42708 19780
rect 41616 19740 42708 19768
rect 42702 19728 42708 19740
rect 42760 19768 42766 19780
rect 43441 19771 43499 19777
rect 43441 19768 43453 19771
rect 42760 19740 43453 19768
rect 42760 19728 42766 19740
rect 43441 19737 43453 19740
rect 43487 19737 43499 19771
rect 43441 19731 43499 19737
rect 41012 19672 41552 19700
rect 41012 19660 41018 19672
rect 42610 19660 42616 19712
rect 42668 19700 42674 19712
rect 42889 19703 42947 19709
rect 42889 19700 42901 19703
rect 42668 19672 42901 19700
rect 42668 19660 42674 19672
rect 42889 19669 42901 19672
rect 42935 19669 42947 19703
rect 42889 19663 42947 19669
rect 1104 19610 54832 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 54832 19610
rect 1104 19536 54832 19558
rect 17034 19456 17040 19508
rect 17092 19496 17098 19508
rect 20070 19496 20076 19508
rect 17092 19468 20076 19496
rect 17092 19456 17098 19468
rect 20070 19456 20076 19468
rect 20128 19456 20134 19508
rect 20162 19456 20168 19508
rect 20220 19496 20226 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 20220 19468 22017 19496
rect 20220 19456 20226 19468
rect 22005 19465 22017 19468
rect 22051 19496 22063 19499
rect 22278 19496 22284 19508
rect 22051 19468 22284 19496
rect 22051 19465 22063 19468
rect 22005 19459 22063 19465
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 22554 19456 22560 19508
rect 22612 19496 22618 19508
rect 23937 19499 23995 19505
rect 23937 19496 23949 19499
rect 22612 19468 23949 19496
rect 22612 19456 22618 19468
rect 23937 19465 23949 19468
rect 23983 19465 23995 19499
rect 23937 19459 23995 19465
rect 25961 19499 26019 19505
rect 25961 19465 25973 19499
rect 26007 19496 26019 19499
rect 26050 19496 26056 19508
rect 26007 19468 26056 19496
rect 26007 19465 26019 19468
rect 25961 19459 26019 19465
rect 26050 19456 26056 19468
rect 26108 19456 26114 19508
rect 26510 19456 26516 19508
rect 26568 19496 26574 19508
rect 27617 19499 27675 19505
rect 27617 19496 27629 19499
rect 26568 19468 27629 19496
rect 26568 19456 26574 19468
rect 27617 19465 27629 19468
rect 27663 19465 27675 19499
rect 27617 19459 27675 19465
rect 28074 19456 28080 19508
rect 28132 19496 28138 19508
rect 28132 19468 28580 19496
rect 28132 19456 28138 19468
rect 19334 19428 19340 19440
rect 18708 19400 19340 19428
rect 1857 19363 1915 19369
rect 1857 19329 1869 19363
rect 1903 19360 1915 19363
rect 14274 19360 14280 19372
rect 1903 19332 14280 19360
rect 1903 19329 1915 19332
rect 1857 19323 1915 19329
rect 14274 19320 14280 19332
rect 14332 19320 14338 19372
rect 18708 19369 18736 19400
rect 19334 19388 19340 19400
rect 19392 19428 19398 19440
rect 22462 19428 22468 19440
rect 19392 19400 22468 19428
rect 19392 19388 19398 19400
rect 22462 19388 22468 19400
rect 22520 19428 22526 19440
rect 23474 19428 23480 19440
rect 22520 19400 23480 19428
rect 22520 19388 22526 19400
rect 18693 19363 18751 19369
rect 18693 19329 18705 19363
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 18960 19363 19018 19369
rect 18960 19329 18972 19363
rect 19006 19360 19018 19363
rect 19242 19360 19248 19372
rect 19006 19332 19248 19360
rect 19006 19329 19018 19332
rect 18960 19323 19018 19329
rect 19242 19320 19248 19332
rect 19300 19320 19306 19372
rect 20622 19360 20628 19372
rect 19996 19332 20628 19360
rect 1670 19156 1676 19168
rect 1631 19128 1676 19156
rect 1670 19116 1676 19128
rect 1728 19116 1734 19168
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 19996 19156 20024 19332
rect 20622 19320 20628 19332
rect 20680 19360 20686 19372
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20680 19332 21097 19360
rect 20680 19320 20686 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 21542 19320 21548 19372
rect 21600 19360 21606 19372
rect 23400 19369 23428 19400
rect 23474 19388 23480 19400
rect 23532 19428 23538 19440
rect 24578 19428 24584 19440
rect 23532 19400 24584 19428
rect 23532 19388 23538 19400
rect 24578 19388 24584 19400
rect 24636 19388 24642 19440
rect 25038 19388 25044 19440
rect 25096 19428 25102 19440
rect 28350 19428 28356 19440
rect 25096 19400 28356 19428
rect 25096 19388 25102 19400
rect 28350 19388 28356 19400
rect 28408 19388 28414 19440
rect 23118 19363 23176 19369
rect 23118 19360 23130 19363
rect 21600 19332 23130 19360
rect 21600 19320 21606 19332
rect 23118 19329 23130 19332
rect 23164 19329 23176 19363
rect 23118 19323 23176 19329
rect 23385 19363 23443 19369
rect 23385 19329 23397 19363
rect 23431 19329 23443 19363
rect 24118 19360 24124 19372
rect 24079 19332 24124 19360
rect 23385 19323 23443 19329
rect 24118 19320 24124 19332
rect 24176 19320 24182 19372
rect 24210 19320 24216 19372
rect 24268 19360 24274 19372
rect 27522 19360 27528 19372
rect 24268 19332 24313 19360
rect 27483 19332 27528 19360
rect 24268 19320 24274 19332
rect 27522 19320 27528 19332
rect 27580 19320 27586 19372
rect 27614 19320 27620 19372
rect 27672 19360 27678 19372
rect 27709 19363 27767 19369
rect 27709 19360 27721 19363
rect 27672 19332 27721 19360
rect 27672 19320 27678 19332
rect 27709 19329 27721 19332
rect 27755 19329 27767 19363
rect 27709 19323 27767 19329
rect 27893 19363 27951 19369
rect 27893 19329 27905 19363
rect 27939 19360 27951 19363
rect 28442 19360 28448 19372
rect 27939 19332 28448 19360
rect 27939 19329 27951 19332
rect 27893 19323 27951 19329
rect 28442 19320 28448 19332
rect 28500 19320 28506 19372
rect 28552 19369 28580 19468
rect 29086 19456 29092 19508
rect 29144 19496 29150 19508
rect 29365 19499 29423 19505
rect 29365 19496 29377 19499
rect 29144 19468 29377 19496
rect 29144 19456 29150 19468
rect 29365 19465 29377 19468
rect 29411 19465 29423 19499
rect 30466 19496 30472 19508
rect 30427 19468 30472 19496
rect 29365 19459 29423 19465
rect 30466 19456 30472 19468
rect 30524 19456 30530 19508
rect 31202 19496 31208 19508
rect 30576 19468 31208 19496
rect 29914 19388 29920 19440
rect 29972 19428 29978 19440
rect 30576 19428 30604 19468
rect 31202 19456 31208 19468
rect 31260 19456 31266 19508
rect 32214 19456 32220 19508
rect 32272 19496 32278 19508
rect 33413 19499 33471 19505
rect 33413 19496 33425 19499
rect 32272 19468 33425 19496
rect 32272 19456 32278 19468
rect 33413 19465 33425 19468
rect 33459 19465 33471 19499
rect 35710 19496 35716 19508
rect 35671 19468 35716 19496
rect 33413 19459 33471 19465
rect 35710 19456 35716 19468
rect 35768 19456 35774 19508
rect 36722 19456 36728 19508
rect 36780 19496 36786 19508
rect 37645 19499 37703 19505
rect 37645 19496 37657 19499
rect 36780 19468 37657 19496
rect 36780 19456 36786 19468
rect 37645 19465 37657 19468
rect 37691 19465 37703 19499
rect 37645 19459 37703 19465
rect 37826 19456 37832 19508
rect 37884 19496 37890 19508
rect 38013 19499 38071 19505
rect 38013 19496 38025 19499
rect 37884 19468 38025 19496
rect 37884 19456 37890 19468
rect 38013 19465 38025 19468
rect 38059 19465 38071 19499
rect 38013 19459 38071 19465
rect 38102 19456 38108 19508
rect 38160 19496 38166 19508
rect 38160 19468 38205 19496
rect 38160 19456 38166 19468
rect 38746 19456 38752 19508
rect 38804 19496 38810 19508
rect 38841 19499 38899 19505
rect 38841 19496 38853 19499
rect 38804 19468 38853 19496
rect 38804 19456 38810 19468
rect 38841 19465 38853 19468
rect 38887 19465 38899 19499
rect 38841 19459 38899 19465
rect 39761 19499 39819 19505
rect 39761 19465 39773 19499
rect 39807 19465 39819 19499
rect 39761 19459 39819 19465
rect 29972 19400 30604 19428
rect 29972 19388 29978 19400
rect 30742 19388 30748 19440
rect 30800 19428 30806 19440
rect 31573 19431 31631 19437
rect 30800 19400 31524 19428
rect 30800 19388 30806 19400
rect 28537 19363 28595 19369
rect 28537 19329 28549 19363
rect 28583 19329 28595 19363
rect 28537 19323 28595 19329
rect 28721 19363 28779 19369
rect 28721 19329 28733 19363
rect 28767 19360 28779 19363
rect 29086 19360 29092 19372
rect 28767 19332 29092 19360
rect 28767 19329 28779 19332
rect 28721 19323 28779 19329
rect 29086 19320 29092 19332
rect 29144 19320 29150 19372
rect 29546 19360 29552 19372
rect 29507 19332 29552 19360
rect 29546 19320 29552 19332
rect 29604 19320 29610 19372
rect 30009 19363 30067 19369
rect 30009 19329 30021 19363
rect 30055 19360 30067 19363
rect 30055 19332 30880 19360
rect 30055 19329 30067 19332
rect 30009 19323 30067 19329
rect 21174 19292 21180 19304
rect 21135 19264 21180 19292
rect 21174 19252 21180 19264
rect 21232 19252 21238 19304
rect 21266 19252 21272 19304
rect 21324 19292 21330 19304
rect 21324 19264 21369 19292
rect 21324 19252 21330 19264
rect 24946 19252 24952 19304
rect 25004 19292 25010 19304
rect 25317 19295 25375 19301
rect 25317 19292 25329 19295
rect 25004 19264 25329 19292
rect 25004 19252 25010 19264
rect 25317 19261 25329 19264
rect 25363 19261 25375 19295
rect 26510 19292 26516 19304
rect 26471 19264 26516 19292
rect 25317 19255 25375 19261
rect 26510 19252 26516 19264
rect 26568 19252 26574 19304
rect 27341 19295 27399 19301
rect 27341 19261 27353 19295
rect 27387 19292 27399 19295
rect 27798 19292 27804 19304
rect 27387 19264 27804 19292
rect 27387 19261 27399 19264
rect 27341 19255 27399 19261
rect 27798 19252 27804 19264
rect 27856 19252 27862 19304
rect 28629 19295 28687 19301
rect 28629 19261 28641 19295
rect 28675 19261 28687 19295
rect 28629 19255 28687 19261
rect 28813 19295 28871 19301
rect 28813 19261 28825 19295
rect 28859 19292 28871 19295
rect 29178 19292 29184 19304
rect 28859 19264 29184 19292
rect 28859 19261 28871 19264
rect 28813 19255 28871 19261
rect 21450 19184 21456 19236
rect 21508 19224 21514 19236
rect 21508 19196 22094 19224
rect 21508 19184 21514 19196
rect 20714 19156 20720 19168
rect 18279 19128 20024 19156
rect 20675 19128 20720 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 22066 19156 22094 19196
rect 28258 19184 28264 19236
rect 28316 19224 28322 19236
rect 28644 19224 28672 19255
rect 29178 19252 29184 19264
rect 29236 19252 29242 19304
rect 28316 19196 28672 19224
rect 28316 19184 28322 19196
rect 30190 19184 30196 19236
rect 30248 19224 30254 19236
rect 30285 19227 30343 19233
rect 30285 19224 30297 19227
rect 30248 19196 30297 19224
rect 30248 19184 30254 19196
rect 30285 19193 30297 19196
rect 30331 19193 30343 19227
rect 30285 19187 30343 19193
rect 23566 19156 23572 19168
rect 22066 19128 23572 19156
rect 23566 19116 23572 19128
rect 23624 19116 23630 19168
rect 23658 19116 23664 19168
rect 23716 19156 23722 19168
rect 24765 19159 24823 19165
rect 24765 19156 24777 19159
rect 23716 19128 24777 19156
rect 23716 19116 23722 19128
rect 24765 19125 24777 19128
rect 24811 19156 24823 19159
rect 28276 19156 28304 19184
rect 24811 19128 28304 19156
rect 28353 19159 28411 19165
rect 24811 19125 24823 19128
rect 24765 19119 24823 19125
rect 28353 19125 28365 19159
rect 28399 19156 28411 19159
rect 28442 19156 28448 19168
rect 28399 19128 28448 19156
rect 28399 19125 28411 19128
rect 28353 19119 28411 19125
rect 28442 19116 28448 19128
rect 28500 19116 28506 19168
rect 30852 19156 30880 19332
rect 31110 19320 31116 19372
rect 31168 19360 31174 19372
rect 31386 19360 31392 19372
rect 31168 19332 31392 19360
rect 31168 19320 31174 19332
rect 31386 19320 31392 19332
rect 31444 19320 31450 19372
rect 31496 19360 31524 19400
rect 31573 19397 31585 19431
rect 31619 19428 31631 19431
rect 31619 19400 33088 19428
rect 31619 19397 31631 19400
rect 31573 19391 31631 19397
rect 31496 19332 31616 19360
rect 31018 19292 31024 19304
rect 30979 19264 31024 19292
rect 31018 19252 31024 19264
rect 31076 19252 31082 19304
rect 31588 19292 31616 19332
rect 31662 19320 31668 19372
rect 31720 19360 31726 19372
rect 32309 19363 32367 19369
rect 32309 19360 32321 19363
rect 31720 19332 32321 19360
rect 31720 19320 31726 19332
rect 32309 19329 32321 19332
rect 32355 19329 32367 19363
rect 32309 19323 32367 19329
rect 31588 19264 31754 19292
rect 31726 19224 31754 19264
rect 32122 19252 32128 19304
rect 32180 19292 32186 19304
rect 32861 19295 32919 19301
rect 32861 19292 32873 19295
rect 32180 19264 32873 19292
rect 32180 19252 32186 19264
rect 32861 19261 32873 19264
rect 32907 19261 32919 19295
rect 33060 19292 33088 19400
rect 34238 19388 34244 19440
rect 34296 19428 34302 19440
rect 34578 19431 34636 19437
rect 34578 19428 34590 19431
rect 34296 19400 34590 19428
rect 34296 19388 34302 19400
rect 34578 19397 34590 19400
rect 34624 19397 34636 19431
rect 34578 19391 34636 19397
rect 37274 19388 37280 19440
rect 37332 19428 37338 19440
rect 39776 19428 39804 19459
rect 39850 19456 39856 19508
rect 39908 19496 39914 19508
rect 40497 19499 40555 19505
rect 40497 19496 40509 19499
rect 39908 19468 40509 19496
rect 39908 19456 39914 19468
rect 40497 19465 40509 19468
rect 40543 19465 40555 19499
rect 40497 19459 40555 19465
rect 41414 19456 41420 19508
rect 41472 19496 41478 19508
rect 41509 19499 41567 19505
rect 41509 19496 41521 19499
rect 41472 19468 41521 19496
rect 41472 19456 41478 19468
rect 41509 19465 41521 19468
rect 41555 19465 41567 19499
rect 54202 19496 54208 19508
rect 54163 19468 54208 19496
rect 41509 19459 41567 19465
rect 54202 19456 54208 19468
rect 54260 19456 54266 19508
rect 40770 19428 40776 19440
rect 37332 19400 39804 19428
rect 39868 19400 40336 19428
rect 40731 19400 40776 19428
rect 37332 19388 37338 19400
rect 33134 19320 33140 19372
rect 33192 19360 33198 19372
rect 33597 19363 33655 19369
rect 33597 19360 33609 19363
rect 33192 19332 33609 19360
rect 33192 19320 33198 19332
rect 33597 19329 33609 19332
rect 33643 19329 33655 19363
rect 39298 19360 39304 19372
rect 33597 19323 33655 19329
rect 38212 19332 39160 19360
rect 39259 19332 39304 19360
rect 33781 19295 33839 19301
rect 33781 19292 33793 19295
rect 33060 19264 33793 19292
rect 32861 19255 32919 19261
rect 33781 19261 33793 19264
rect 33827 19261 33839 19295
rect 34330 19292 34336 19304
rect 34291 19264 34336 19292
rect 33781 19255 33839 19261
rect 34330 19252 34336 19264
rect 34388 19252 34394 19304
rect 35986 19252 35992 19304
rect 36044 19292 36050 19304
rect 36173 19295 36231 19301
rect 36173 19292 36185 19295
rect 36044 19264 36185 19292
rect 36044 19252 36050 19264
rect 36173 19261 36185 19264
rect 36219 19261 36231 19295
rect 36173 19255 36231 19261
rect 36262 19252 36268 19304
rect 36320 19292 36326 19304
rect 37366 19292 37372 19304
rect 36320 19264 37372 19292
rect 36320 19252 36326 19264
rect 37366 19252 37372 19264
rect 37424 19292 37430 19304
rect 38212 19292 38240 19332
rect 37424 19264 38240 19292
rect 37424 19252 37430 19264
rect 38286 19252 38292 19304
rect 38344 19292 38350 19304
rect 39132 19292 39160 19332
rect 39298 19320 39304 19332
rect 39356 19320 39362 19372
rect 39761 19363 39819 19369
rect 39761 19360 39773 19363
rect 39408 19332 39773 19360
rect 39408 19292 39436 19332
rect 39761 19329 39773 19332
rect 39807 19329 39819 19363
rect 39761 19323 39819 19329
rect 38344 19264 38389 19292
rect 39132 19264 39436 19292
rect 38344 19252 38350 19264
rect 33686 19224 33692 19236
rect 31726 19196 33692 19224
rect 33686 19184 33692 19196
rect 33744 19184 33750 19236
rect 37090 19224 37096 19236
rect 35268 19196 37096 19224
rect 32306 19156 32312 19168
rect 30852 19128 32312 19156
rect 32306 19116 32312 19128
rect 32364 19116 32370 19168
rect 33410 19116 33416 19168
rect 33468 19156 33474 19168
rect 35268 19156 35296 19196
rect 37090 19184 37096 19196
rect 37148 19184 37154 19236
rect 38933 19227 38991 19233
rect 38933 19224 38945 19227
rect 37476 19196 38945 19224
rect 33468 19128 35296 19156
rect 36817 19159 36875 19165
rect 33468 19116 33474 19128
rect 36817 19125 36829 19159
rect 36863 19156 36875 19159
rect 37476 19156 37504 19196
rect 38933 19193 38945 19196
rect 38979 19193 38991 19227
rect 38933 19187 38991 19193
rect 39206 19184 39212 19236
rect 39264 19224 39270 19236
rect 39868 19224 39896 19400
rect 39945 19363 40003 19369
rect 39945 19329 39957 19363
rect 39991 19329 40003 19363
rect 40308 19360 40336 19400
rect 40770 19388 40776 19400
rect 40828 19428 40834 19440
rect 44726 19428 44732 19440
rect 40828 19400 41399 19428
rect 40828 19388 40834 19400
rect 40681 19363 40739 19369
rect 40681 19360 40693 19363
rect 40308 19332 40693 19360
rect 39945 19323 40003 19329
rect 40681 19329 40693 19332
rect 40727 19329 40739 19363
rect 40681 19323 40739 19329
rect 40865 19363 40923 19369
rect 40865 19329 40877 19363
rect 40911 19360 40923 19363
rect 41049 19363 41107 19369
rect 40911 19332 40945 19360
rect 40911 19329 40923 19332
rect 40865 19323 40923 19329
rect 41049 19329 41061 19363
rect 41095 19360 41107 19363
rect 41138 19360 41144 19372
rect 41095 19332 41144 19360
rect 41095 19329 41107 19332
rect 41049 19323 41107 19329
rect 39264 19196 39896 19224
rect 39264 19184 39270 19196
rect 36863 19128 37504 19156
rect 36863 19125 36875 19128
rect 36817 19119 36875 19125
rect 38654 19116 38660 19168
rect 38712 19156 38718 19168
rect 39960 19156 39988 19323
rect 40402 19252 40408 19304
rect 40460 19292 40466 19304
rect 40880 19292 40908 19323
rect 41138 19320 41144 19332
rect 41196 19320 41202 19372
rect 41371 19360 41399 19400
rect 41340 19306 41399 19360
rect 41230 19292 41236 19304
rect 40460 19264 41236 19292
rect 40460 19252 40466 19264
rect 41230 19252 41236 19264
rect 41288 19252 41294 19304
rect 41371 19292 41399 19306
rect 41432 19400 44732 19428
rect 41432 19292 41460 19400
rect 44726 19388 44732 19400
rect 44784 19388 44790 19440
rect 41598 19320 41604 19372
rect 41656 19360 41662 19372
rect 41693 19363 41751 19369
rect 41693 19360 41705 19363
rect 41656 19332 41705 19360
rect 41656 19320 41662 19332
rect 41693 19329 41705 19332
rect 41739 19329 41751 19363
rect 41693 19323 41751 19329
rect 54021 19363 54079 19369
rect 54021 19329 54033 19363
rect 54067 19329 54079 19363
rect 54021 19323 54079 19329
rect 41371 19264 41460 19292
rect 40034 19184 40040 19236
rect 40092 19224 40098 19236
rect 54036 19224 54064 19323
rect 40092 19196 54064 19224
rect 40092 19184 40098 19196
rect 38712 19128 39988 19156
rect 38712 19116 38718 19128
rect 40126 19116 40132 19168
rect 40184 19156 40190 19168
rect 42334 19156 42340 19168
rect 40184 19128 42340 19156
rect 40184 19116 40190 19128
rect 42334 19116 42340 19128
rect 42392 19116 42398 19168
rect 42610 19156 42616 19168
rect 42571 19128 42616 19156
rect 42610 19116 42616 19128
rect 42668 19116 42674 19168
rect 53561 19159 53619 19165
rect 53561 19125 53573 19159
rect 53607 19156 53619 19159
rect 54202 19156 54208 19168
rect 53607 19128 54208 19156
rect 53607 19125 53619 19128
rect 53561 19119 53619 19125
rect 54202 19116 54208 19128
rect 54260 19116 54266 19168
rect 1104 19066 54832 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 54832 19066
rect 1104 18992 54832 19014
rect 2409 18955 2467 18961
rect 2409 18921 2421 18955
rect 2455 18952 2467 18955
rect 2590 18952 2596 18964
rect 2455 18924 2596 18952
rect 2455 18921 2467 18924
rect 2409 18915 2467 18921
rect 1857 18751 1915 18757
rect 1857 18717 1869 18751
rect 1903 18748 1915 18751
rect 2424 18748 2452 18915
rect 2590 18912 2596 18924
rect 2648 18912 2654 18964
rect 24857 18955 24915 18961
rect 24857 18921 24869 18955
rect 24903 18952 24915 18955
rect 25314 18952 25320 18964
rect 24903 18924 25320 18952
rect 24903 18921 24915 18924
rect 24857 18915 24915 18921
rect 25314 18912 25320 18924
rect 25372 18912 25378 18964
rect 26510 18952 26516 18964
rect 26471 18924 26516 18952
rect 26510 18912 26516 18924
rect 26568 18912 26574 18964
rect 28626 18912 28632 18964
rect 28684 18952 28690 18964
rect 29178 18952 29184 18964
rect 28684 18924 29184 18952
rect 28684 18912 28690 18924
rect 29178 18912 29184 18924
rect 29236 18952 29242 18964
rect 29733 18955 29791 18961
rect 29733 18952 29745 18955
rect 29236 18924 29745 18952
rect 29236 18912 29242 18924
rect 29733 18921 29745 18924
rect 29779 18921 29791 18955
rect 29733 18915 29791 18921
rect 32030 18912 32036 18964
rect 32088 18952 32094 18964
rect 33229 18955 33287 18961
rect 33229 18952 33241 18955
rect 32088 18924 33241 18952
rect 32088 18912 32094 18924
rect 33229 18921 33241 18924
rect 33275 18921 33287 18955
rect 34330 18952 34336 18964
rect 34291 18924 34336 18952
rect 33229 18915 33287 18921
rect 34330 18912 34336 18924
rect 34388 18912 34394 18964
rect 35986 18952 35992 18964
rect 35947 18924 35992 18952
rect 35986 18912 35992 18924
rect 36044 18912 36050 18964
rect 36906 18912 36912 18964
rect 36964 18952 36970 18964
rect 37001 18955 37059 18961
rect 37001 18952 37013 18955
rect 36964 18924 37013 18952
rect 36964 18912 36970 18924
rect 37001 18921 37013 18924
rect 37047 18921 37059 18955
rect 37001 18915 37059 18921
rect 37090 18912 37096 18964
rect 37148 18952 37154 18964
rect 40034 18952 40040 18964
rect 37148 18924 39436 18952
rect 39995 18924 40040 18952
rect 37148 18912 37154 18924
rect 15470 18844 15476 18896
rect 15528 18884 15534 18896
rect 21085 18887 21143 18893
rect 21085 18884 21097 18887
rect 15528 18856 21097 18884
rect 15528 18844 15534 18856
rect 21085 18853 21097 18856
rect 21131 18884 21143 18887
rect 21174 18884 21180 18896
rect 21131 18856 21180 18884
rect 21131 18853 21143 18856
rect 21085 18847 21143 18853
rect 21174 18844 21180 18856
rect 21232 18844 21238 18896
rect 27709 18887 27767 18893
rect 27709 18853 27721 18887
rect 27755 18884 27767 18887
rect 28442 18884 28448 18896
rect 27755 18856 28448 18884
rect 27755 18853 27767 18856
rect 27709 18847 27767 18853
rect 28442 18844 28448 18856
rect 28500 18844 28506 18896
rect 32769 18887 32827 18893
rect 32769 18853 32781 18887
rect 32815 18884 32827 18887
rect 33042 18884 33048 18896
rect 32815 18856 33048 18884
rect 32815 18853 32827 18856
rect 32769 18847 32827 18853
rect 33042 18844 33048 18856
rect 33100 18844 33106 18896
rect 34882 18884 34888 18896
rect 33428 18856 33732 18884
rect 34843 18856 34888 18884
rect 22462 18816 22468 18828
rect 22423 18788 22468 18816
rect 22462 18776 22468 18788
rect 22520 18776 22526 18828
rect 23753 18819 23811 18825
rect 23753 18785 23765 18819
rect 23799 18816 23811 18819
rect 23934 18816 23940 18828
rect 23799 18788 23940 18816
rect 23799 18785 23811 18788
rect 23753 18779 23811 18785
rect 23934 18776 23940 18788
rect 23992 18776 23998 18828
rect 24029 18819 24087 18825
rect 24029 18785 24041 18819
rect 24075 18816 24087 18819
rect 25869 18819 25927 18825
rect 25869 18816 25881 18819
rect 24075 18788 25881 18816
rect 24075 18785 24087 18788
rect 24029 18779 24087 18785
rect 25869 18785 25881 18788
rect 25915 18785 25927 18819
rect 25869 18779 25927 18785
rect 26881 18819 26939 18825
rect 26881 18785 26893 18819
rect 26927 18816 26939 18819
rect 27154 18816 27160 18828
rect 26927 18788 27160 18816
rect 26927 18785 26939 18788
rect 26881 18779 26939 18785
rect 27154 18776 27160 18788
rect 27212 18776 27218 18828
rect 27614 18816 27620 18828
rect 27448 18788 27620 18816
rect 1903 18720 2452 18748
rect 19429 18751 19487 18757
rect 1903 18717 1915 18720
rect 1857 18711 1915 18717
rect 19429 18717 19441 18751
rect 19475 18748 19487 18751
rect 20346 18748 20352 18760
rect 19475 18720 20352 18748
rect 19475 18717 19487 18720
rect 19429 18711 19487 18717
rect 20346 18708 20352 18720
rect 20404 18708 20410 18760
rect 20441 18751 20499 18757
rect 20441 18717 20453 18751
rect 20487 18748 20499 18751
rect 20714 18748 20720 18760
rect 20487 18720 20720 18748
rect 20487 18717 20499 18720
rect 20441 18711 20499 18717
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 23658 18748 23664 18760
rect 23619 18720 23664 18748
rect 23658 18708 23664 18720
rect 23716 18708 23722 18760
rect 24670 18748 24676 18760
rect 24631 18720 24676 18748
rect 24670 18708 24676 18720
rect 24728 18708 24734 18760
rect 26789 18751 26847 18757
rect 26789 18717 26801 18751
rect 26835 18748 26847 18751
rect 27448 18748 27476 18788
rect 27614 18776 27620 18788
rect 27672 18776 27678 18828
rect 27798 18776 27804 18828
rect 27856 18816 27862 18828
rect 27856 18788 28313 18816
rect 27856 18776 27862 18788
rect 26835 18720 27476 18748
rect 27525 18751 27583 18757
rect 26835 18717 26847 18720
rect 26789 18711 26847 18717
rect 27525 18717 27537 18751
rect 27571 18748 27583 18751
rect 28166 18748 28172 18760
rect 27571 18720 28172 18748
rect 27571 18717 27583 18720
rect 27525 18711 27583 18717
rect 28166 18708 28172 18720
rect 28224 18708 28230 18760
rect 28285 18748 28313 18788
rect 28350 18776 28356 18828
rect 28408 18816 28414 18828
rect 28721 18819 28779 18825
rect 28721 18816 28733 18819
rect 28408 18788 28733 18816
rect 28408 18776 28414 18788
rect 28721 18785 28733 18788
rect 28767 18785 28779 18819
rect 28721 18779 28779 18785
rect 30834 18776 30840 18828
rect 30892 18816 30898 18828
rect 31389 18819 31447 18825
rect 31389 18816 31401 18819
rect 30892 18788 31401 18816
rect 30892 18776 30898 18788
rect 31389 18785 31401 18788
rect 31435 18785 31447 18819
rect 31389 18779 31447 18785
rect 32858 18776 32864 18828
rect 32916 18816 32922 18828
rect 33428 18816 33456 18856
rect 32916 18788 33456 18816
rect 32916 18776 32922 18788
rect 33502 18776 33508 18828
rect 33560 18816 33566 18828
rect 33704 18825 33732 18856
rect 34882 18844 34888 18856
rect 34940 18844 34946 18896
rect 35342 18844 35348 18896
rect 35400 18884 35406 18896
rect 39298 18884 39304 18896
rect 35400 18856 39304 18884
rect 35400 18844 35406 18856
rect 39298 18844 39304 18856
rect 39356 18844 39362 18896
rect 39408 18884 39436 18924
rect 40034 18912 40040 18924
rect 40092 18912 40098 18964
rect 54113 18955 54171 18961
rect 54113 18952 54125 18955
rect 40144 18924 54125 18952
rect 40144 18884 40172 18924
rect 54113 18921 54125 18924
rect 54159 18921 54171 18955
rect 54113 18915 54171 18921
rect 39408 18856 40172 18884
rect 41506 18844 41512 18896
rect 41564 18884 41570 18896
rect 42518 18884 42524 18896
rect 41564 18856 42524 18884
rect 41564 18844 41570 18856
rect 42518 18844 42524 18856
rect 42576 18844 42582 18896
rect 33689 18819 33747 18825
rect 33560 18788 33605 18816
rect 33560 18776 33566 18788
rect 33689 18785 33701 18819
rect 33735 18785 33747 18819
rect 33689 18779 33747 18785
rect 33870 18776 33876 18828
rect 33928 18816 33934 18828
rect 36262 18816 36268 18828
rect 33928 18788 36268 18816
rect 33928 18776 33934 18788
rect 36262 18776 36268 18788
rect 36320 18776 36326 18828
rect 36449 18819 36507 18825
rect 36449 18785 36461 18819
rect 36495 18816 36507 18819
rect 36906 18816 36912 18828
rect 36495 18788 36912 18816
rect 36495 18785 36507 18788
rect 36449 18779 36507 18785
rect 36906 18776 36912 18788
rect 36964 18776 36970 18828
rect 37645 18819 37703 18825
rect 37645 18785 37657 18819
rect 37691 18816 37703 18819
rect 37826 18816 37832 18828
rect 37691 18788 37832 18816
rect 37691 18785 37703 18788
rect 37645 18779 37703 18785
rect 37826 18776 37832 18788
rect 37884 18776 37890 18828
rect 38654 18776 38660 18828
rect 38712 18776 38718 18828
rect 40034 18816 40040 18828
rect 39040 18788 40040 18816
rect 30098 18748 30104 18760
rect 28285 18720 30104 18748
rect 30098 18708 30104 18720
rect 30156 18708 30162 18760
rect 30282 18748 30288 18760
rect 30243 18720 30288 18748
rect 30282 18708 30288 18720
rect 30340 18708 30346 18760
rect 31662 18757 31668 18760
rect 31656 18748 31668 18757
rect 31623 18720 31668 18748
rect 31656 18711 31668 18720
rect 31662 18708 31668 18711
rect 31720 18708 31726 18760
rect 32490 18708 32496 18760
rect 32548 18748 32554 18760
rect 33413 18751 33471 18757
rect 33413 18748 33425 18751
rect 32548 18720 33425 18748
rect 32548 18708 32554 18720
rect 33413 18717 33425 18720
rect 33459 18717 33471 18751
rect 33413 18711 33471 18717
rect 33597 18751 33655 18757
rect 33597 18717 33609 18751
rect 33643 18748 33655 18751
rect 33778 18748 33784 18760
rect 33643 18720 33784 18748
rect 33643 18717 33655 18720
rect 33597 18711 33655 18717
rect 33778 18708 33784 18720
rect 33836 18708 33842 18760
rect 34514 18708 34520 18760
rect 34572 18748 34578 18760
rect 35437 18751 35495 18757
rect 35437 18748 35449 18751
rect 34572 18720 35449 18748
rect 34572 18708 34578 18720
rect 35437 18717 35449 18720
rect 35483 18717 35495 18751
rect 36170 18748 36176 18760
rect 36131 18720 36176 18748
rect 35437 18711 35495 18717
rect 36170 18708 36176 18720
rect 36228 18708 36234 18760
rect 36354 18708 36360 18760
rect 36412 18748 36418 18760
rect 36630 18748 36636 18760
rect 36412 18720 36636 18748
rect 36412 18708 36418 18720
rect 36630 18708 36636 18720
rect 36688 18708 36694 18760
rect 38286 18748 38292 18760
rect 38247 18720 38292 18748
rect 38286 18708 38292 18720
rect 38344 18708 38350 18760
rect 38672 18748 38700 18776
rect 38396 18720 38700 18748
rect 38749 18751 38807 18757
rect 17218 18640 17224 18692
rect 17276 18680 17282 18692
rect 18785 18683 18843 18689
rect 18785 18680 18797 18683
rect 17276 18652 18797 18680
rect 17276 18640 17282 18652
rect 18785 18649 18797 18652
rect 18831 18680 18843 18683
rect 20530 18680 20536 18692
rect 18831 18652 20536 18680
rect 18831 18649 18843 18652
rect 18785 18643 18843 18649
rect 20530 18640 20536 18652
rect 20588 18640 20594 18692
rect 22198 18683 22256 18689
rect 22198 18680 22210 18683
rect 20640 18652 22210 18680
rect 1670 18612 1676 18624
rect 1631 18584 1676 18612
rect 1670 18572 1676 18584
rect 1728 18572 1734 18624
rect 18322 18612 18328 18624
rect 18283 18584 18328 18612
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 19426 18572 19432 18624
rect 19484 18612 19490 18624
rect 20640 18621 20668 18652
rect 22198 18649 22210 18652
rect 22244 18649 22256 18683
rect 22198 18643 22256 18649
rect 23017 18683 23075 18689
rect 23017 18649 23029 18683
rect 23063 18680 23075 18683
rect 27614 18680 27620 18692
rect 23063 18652 27620 18680
rect 23063 18649 23075 18652
rect 23017 18643 23075 18649
rect 27614 18640 27620 18652
rect 27672 18640 27678 18692
rect 28350 18640 28356 18692
rect 28408 18680 28414 18692
rect 28534 18680 28540 18692
rect 28408 18652 28540 18680
rect 28408 18640 28414 18652
rect 28534 18640 28540 18652
rect 28592 18640 28598 18692
rect 36188 18680 36216 18708
rect 38396 18680 38424 18720
rect 38749 18717 38761 18751
rect 38795 18748 38807 18751
rect 38838 18748 38844 18760
rect 38795 18720 38844 18748
rect 38795 18717 38807 18720
rect 38749 18711 38807 18717
rect 38838 18708 38844 18720
rect 38896 18708 38902 18760
rect 39040 18757 39068 18788
rect 40034 18776 40040 18788
rect 40092 18776 40098 18828
rect 41417 18819 41475 18825
rect 41417 18785 41429 18819
rect 41463 18816 41475 18819
rect 42702 18816 42708 18828
rect 41463 18788 42708 18816
rect 41463 18785 41475 18788
rect 41417 18779 41475 18785
rect 42702 18776 42708 18788
rect 42760 18776 42766 18828
rect 39206 18757 39212 18760
rect 39025 18751 39083 18757
rect 39025 18717 39037 18751
rect 39071 18717 39083 18751
rect 39025 18711 39083 18717
rect 39163 18751 39212 18757
rect 39163 18717 39175 18751
rect 39209 18717 39212 18751
rect 39163 18711 39212 18717
rect 39206 18708 39212 18711
rect 39264 18708 39270 18760
rect 39298 18708 39304 18760
rect 39356 18748 39362 18760
rect 41874 18748 41880 18760
rect 39356 18720 41880 18748
rect 39356 18708 39362 18720
rect 41874 18708 41880 18720
rect 41932 18708 41938 18760
rect 42058 18748 42064 18760
rect 42019 18720 42064 18748
rect 42058 18708 42064 18720
rect 42116 18708 42122 18760
rect 54202 18748 54208 18760
rect 54163 18720 54208 18748
rect 54202 18708 54208 18720
rect 54260 18708 54266 18760
rect 36188 18652 38424 18680
rect 38654 18640 38660 18692
rect 38712 18680 38718 18692
rect 38933 18683 38991 18689
rect 38933 18680 38945 18683
rect 38712 18652 38945 18680
rect 38712 18640 38718 18652
rect 38933 18649 38945 18652
rect 38979 18649 38991 18683
rect 40218 18680 40224 18692
rect 38933 18643 38991 18649
rect 39224 18652 40224 18680
rect 19613 18615 19671 18621
rect 19613 18612 19625 18615
rect 19484 18584 19625 18612
rect 19484 18572 19490 18584
rect 19613 18581 19625 18584
rect 19659 18581 19671 18615
rect 19613 18575 19671 18581
rect 20625 18615 20683 18621
rect 20625 18581 20637 18615
rect 20671 18581 20683 18615
rect 25314 18612 25320 18624
rect 25275 18584 25320 18612
rect 20625 18575 20683 18581
rect 25314 18572 25320 18584
rect 25372 18572 25378 18624
rect 28169 18615 28227 18621
rect 28169 18581 28181 18615
rect 28215 18612 28227 18615
rect 28258 18612 28264 18624
rect 28215 18584 28264 18612
rect 28215 18581 28227 18584
rect 28169 18575 28227 18581
rect 28258 18572 28264 18584
rect 28316 18572 28322 18624
rect 30834 18612 30840 18624
rect 30795 18584 30840 18612
rect 30834 18572 30840 18584
rect 30892 18612 30898 18624
rect 31846 18612 31852 18624
rect 30892 18584 31852 18612
rect 30892 18572 30898 18584
rect 31846 18572 31852 18584
rect 31904 18572 31910 18624
rect 32674 18572 32680 18624
rect 32732 18612 32738 18624
rect 33686 18612 33692 18624
rect 32732 18584 33692 18612
rect 32732 18572 32738 18584
rect 33686 18572 33692 18584
rect 33744 18572 33750 18624
rect 38102 18572 38108 18624
rect 38160 18612 38166 18624
rect 38160 18584 38205 18612
rect 38160 18572 38166 18584
rect 38286 18572 38292 18624
rect 38344 18612 38350 18624
rect 39224 18612 39252 18652
rect 40218 18640 40224 18652
rect 40276 18640 40282 18692
rect 40494 18640 40500 18692
rect 40552 18680 40558 18692
rect 40954 18680 40960 18692
rect 40552 18652 40960 18680
rect 40552 18640 40558 18652
rect 40954 18640 40960 18652
rect 41012 18640 41018 18692
rect 41172 18683 41230 18689
rect 41172 18649 41184 18683
rect 41218 18680 41230 18683
rect 41414 18680 41420 18692
rect 41218 18652 41420 18680
rect 41218 18649 41230 18652
rect 41172 18643 41230 18649
rect 41414 18640 41420 18652
rect 41472 18640 41478 18692
rect 49694 18640 49700 18692
rect 49752 18680 49758 18692
rect 53285 18683 53343 18689
rect 53285 18680 53297 18683
rect 49752 18652 53297 18680
rect 49752 18640 49758 18652
rect 53285 18649 53297 18652
rect 53331 18649 53343 18683
rect 53466 18680 53472 18692
rect 53427 18652 53472 18680
rect 53285 18643 53343 18649
rect 53466 18640 53472 18652
rect 53524 18640 53530 18692
rect 38344 18584 39252 18612
rect 39301 18615 39359 18621
rect 38344 18572 38350 18584
rect 39301 18581 39313 18615
rect 39347 18612 39359 18615
rect 39942 18612 39948 18624
rect 39347 18584 39948 18612
rect 39347 18581 39359 18584
rect 39301 18575 39359 18581
rect 39942 18572 39948 18584
rect 40000 18572 40006 18624
rect 40310 18572 40316 18624
rect 40368 18612 40374 18624
rect 41877 18615 41935 18621
rect 41877 18612 41889 18615
rect 40368 18584 41889 18612
rect 40368 18572 40374 18584
rect 41877 18581 41889 18584
rect 41923 18581 41935 18615
rect 41877 18575 41935 18581
rect 42702 18572 42708 18624
rect 42760 18612 42766 18624
rect 43165 18615 43223 18621
rect 43165 18612 43177 18615
rect 42760 18584 43177 18612
rect 42760 18572 42766 18584
rect 43165 18581 43177 18584
rect 43211 18612 43223 18615
rect 44082 18612 44088 18624
rect 43211 18584 44088 18612
rect 43211 18581 43223 18584
rect 43165 18575 43223 18581
rect 44082 18572 44088 18584
rect 44140 18572 44146 18624
rect 52825 18615 52883 18621
rect 52825 18581 52837 18615
rect 52871 18612 52883 18615
rect 53484 18612 53512 18640
rect 52871 18584 53512 18612
rect 52871 18581 52883 18584
rect 52825 18575 52883 18581
rect 1104 18522 54832 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 54832 18522
rect 1104 18448 54832 18470
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 18380 18380 20300 18408
rect 18380 18368 18386 18380
rect 19334 18340 19340 18352
rect 18800 18312 19340 18340
rect 18800 18281 18828 18312
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 20272 18340 20300 18380
rect 20346 18368 20352 18420
rect 20404 18408 20410 18420
rect 20625 18411 20683 18417
rect 20625 18408 20637 18411
rect 20404 18380 20637 18408
rect 20404 18368 20410 18380
rect 20625 18377 20637 18380
rect 20671 18377 20683 18411
rect 31386 18408 31392 18420
rect 20625 18371 20683 18377
rect 22066 18380 31392 18408
rect 20993 18343 21051 18349
rect 20993 18340 21005 18343
rect 20272 18312 21005 18340
rect 20993 18309 21005 18312
rect 21039 18340 21051 18343
rect 22066 18340 22094 18380
rect 31386 18368 31392 18380
rect 31444 18368 31450 18420
rect 31573 18411 31631 18417
rect 31573 18377 31585 18411
rect 31619 18377 31631 18411
rect 31573 18371 31631 18377
rect 23474 18340 23480 18352
rect 21039 18312 22094 18340
rect 23124 18312 23480 18340
rect 21039 18309 21051 18312
rect 20993 18303 21051 18309
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 18785 18275 18843 18281
rect 1811 18244 2360 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 2332 18077 2360 18244
rect 18785 18241 18797 18275
rect 18831 18241 18843 18275
rect 19041 18275 19099 18281
rect 19041 18272 19053 18275
rect 18785 18235 18843 18241
rect 18892 18244 19053 18272
rect 17954 18164 17960 18216
rect 18012 18204 18018 18216
rect 18892 18204 18920 18244
rect 19041 18241 19053 18244
rect 19087 18241 19099 18275
rect 22462 18272 22468 18284
rect 22423 18244 22468 18272
rect 19041 18235 19099 18241
rect 22462 18232 22468 18244
rect 22520 18232 22526 18284
rect 23124 18281 23152 18312
rect 23474 18300 23480 18312
rect 23532 18300 23538 18352
rect 26510 18340 26516 18352
rect 24964 18312 26516 18340
rect 23109 18275 23167 18281
rect 23109 18241 23121 18275
rect 23155 18241 23167 18275
rect 23109 18235 23167 18241
rect 23198 18232 23204 18284
rect 23256 18272 23262 18284
rect 23365 18275 23423 18281
rect 23365 18272 23377 18275
rect 23256 18244 23377 18272
rect 23256 18232 23262 18244
rect 23365 18241 23377 18244
rect 23411 18241 23423 18275
rect 23365 18235 23423 18241
rect 24854 18232 24860 18284
rect 24912 18272 24918 18284
rect 24964 18281 24992 18312
rect 26510 18300 26516 18312
rect 26568 18300 26574 18352
rect 27430 18300 27436 18352
rect 27488 18340 27494 18352
rect 28074 18340 28080 18352
rect 27488 18312 28080 18340
rect 27488 18300 27494 18312
rect 28074 18300 28080 18312
rect 28132 18300 28138 18352
rect 28261 18343 28319 18349
rect 28261 18309 28273 18343
rect 28307 18340 28319 18343
rect 28350 18340 28356 18352
rect 28307 18312 28356 18340
rect 28307 18309 28319 18312
rect 28261 18303 28319 18309
rect 28350 18300 28356 18312
rect 28408 18300 28414 18352
rect 28445 18343 28503 18349
rect 28445 18309 28457 18343
rect 28491 18340 28503 18343
rect 28626 18340 28632 18352
rect 28491 18312 28632 18340
rect 28491 18309 28503 18312
rect 28445 18303 28503 18309
rect 28626 18300 28632 18312
rect 28684 18300 28690 18352
rect 30098 18300 30104 18352
rect 30156 18340 30162 18352
rect 30742 18340 30748 18352
rect 30156 18312 30748 18340
rect 30156 18300 30162 18312
rect 30742 18300 30748 18312
rect 30800 18300 30806 18352
rect 30926 18340 30932 18352
rect 30887 18312 30932 18340
rect 30926 18300 30932 18312
rect 30984 18300 30990 18352
rect 31018 18300 31024 18352
rect 31076 18340 31082 18352
rect 31588 18340 31616 18371
rect 37826 18368 37832 18420
rect 37884 18408 37890 18420
rect 38286 18408 38292 18420
rect 37884 18380 38292 18408
rect 37884 18368 37890 18380
rect 38286 18368 38292 18380
rect 38344 18368 38350 18420
rect 38565 18411 38623 18417
rect 38565 18377 38577 18411
rect 38611 18408 38623 18411
rect 40126 18408 40132 18420
rect 38611 18380 40132 18408
rect 38611 18377 38623 18380
rect 38565 18371 38623 18377
rect 40126 18368 40132 18380
rect 40184 18368 40190 18420
rect 40218 18368 40224 18420
rect 40276 18408 40282 18420
rect 41506 18408 41512 18420
rect 40276 18380 41512 18408
rect 40276 18368 40282 18380
rect 41506 18368 41512 18380
rect 41564 18368 41570 18420
rect 41690 18368 41696 18420
rect 41748 18408 41754 18420
rect 41969 18411 42027 18417
rect 41969 18408 41981 18411
rect 41748 18380 41981 18408
rect 41748 18368 41754 18380
rect 41969 18377 41981 18380
rect 42015 18408 42027 18411
rect 42610 18408 42616 18420
rect 42015 18380 42616 18408
rect 42015 18377 42027 18380
rect 41969 18371 42027 18377
rect 42610 18368 42616 18380
rect 42668 18368 42674 18420
rect 43254 18408 43260 18420
rect 43215 18380 43260 18408
rect 43254 18368 43260 18380
rect 43312 18368 43318 18420
rect 54202 18408 54208 18420
rect 54163 18380 54208 18408
rect 54202 18368 54208 18380
rect 54260 18368 54266 18420
rect 32585 18343 32643 18349
rect 32585 18340 32597 18343
rect 31076 18312 31616 18340
rect 31680 18312 32597 18340
rect 31076 18300 31082 18312
rect 25222 18281 25228 18284
rect 24949 18275 25007 18281
rect 24949 18272 24961 18275
rect 24912 18244 24961 18272
rect 24912 18232 24918 18244
rect 24949 18241 24961 18244
rect 24995 18241 25007 18275
rect 25216 18272 25228 18281
rect 25183 18244 25228 18272
rect 24949 18235 25007 18241
rect 25216 18235 25228 18244
rect 25222 18232 25228 18235
rect 25280 18232 25286 18284
rect 27249 18275 27307 18281
rect 27249 18241 27261 18275
rect 27295 18272 27307 18275
rect 27982 18272 27988 18284
rect 27295 18244 27988 18272
rect 27295 18241 27307 18244
rect 27249 18235 27307 18241
rect 27982 18232 27988 18244
rect 28040 18232 28046 18284
rect 28169 18275 28227 18281
rect 28169 18241 28181 18275
rect 28215 18272 28227 18275
rect 28534 18272 28540 18284
rect 28215 18244 28540 18272
rect 28215 18241 28227 18244
rect 28169 18235 28227 18241
rect 28534 18232 28540 18244
rect 28592 18232 28598 18284
rect 30018 18275 30076 18281
rect 30018 18272 30030 18275
rect 28736 18244 30030 18272
rect 18012 18176 18920 18204
rect 18012 18164 18018 18176
rect 20714 18164 20720 18216
rect 20772 18204 20778 18216
rect 21085 18207 21143 18213
rect 21085 18204 21097 18207
rect 20772 18176 21097 18204
rect 20772 18164 20778 18176
rect 21085 18173 21097 18176
rect 21131 18173 21143 18207
rect 21085 18167 21143 18173
rect 21266 18164 21272 18216
rect 21324 18204 21330 18216
rect 22002 18204 22008 18216
rect 21324 18176 22008 18204
rect 21324 18164 21330 18176
rect 22002 18164 22008 18176
rect 22060 18164 22066 18216
rect 28736 18204 28764 18244
rect 30018 18241 30030 18244
rect 30064 18241 30076 18275
rect 30944 18272 30972 18300
rect 31573 18278 31631 18281
rect 31680 18278 31708 18312
rect 32585 18309 32597 18312
rect 32631 18340 32643 18343
rect 33502 18340 33508 18352
rect 32631 18312 33508 18340
rect 32631 18309 32643 18312
rect 32585 18303 32643 18309
rect 33502 18300 33508 18312
rect 33560 18300 33566 18352
rect 34692 18343 34750 18349
rect 34692 18309 34704 18343
rect 34738 18340 34750 18343
rect 34882 18340 34888 18352
rect 34738 18312 34888 18340
rect 34738 18309 34750 18312
rect 34692 18303 34750 18309
rect 34882 18300 34888 18312
rect 34940 18300 34946 18352
rect 34974 18300 34980 18352
rect 35032 18340 35038 18352
rect 53190 18340 53196 18352
rect 35032 18312 53196 18340
rect 35032 18300 35038 18312
rect 53190 18300 53196 18312
rect 53248 18300 53254 18352
rect 31573 18275 31708 18278
rect 31573 18272 31585 18275
rect 30944 18244 31585 18272
rect 30018 18235 30076 18241
rect 31573 18241 31585 18244
rect 31619 18250 31708 18275
rect 31619 18241 31631 18250
rect 31573 18235 31631 18241
rect 31754 18232 31760 18284
rect 31812 18272 31818 18284
rect 32490 18272 32496 18284
rect 31812 18244 32496 18272
rect 31812 18232 31818 18244
rect 32490 18232 32496 18244
rect 32548 18232 32554 18284
rect 32674 18272 32680 18284
rect 32635 18244 32680 18272
rect 32674 18232 32680 18244
rect 32732 18232 32738 18284
rect 32858 18272 32864 18284
rect 32819 18244 32864 18272
rect 32858 18232 32864 18244
rect 32916 18232 32922 18284
rect 33781 18275 33839 18281
rect 33781 18241 33793 18275
rect 33827 18272 33839 18275
rect 33870 18272 33876 18284
rect 33827 18244 33876 18272
rect 33827 18241 33839 18244
rect 33781 18235 33839 18241
rect 33870 18232 33876 18244
rect 33928 18232 33934 18284
rect 34330 18232 34336 18284
rect 34388 18272 34394 18284
rect 34425 18275 34483 18281
rect 34425 18272 34437 18275
rect 34388 18244 34437 18272
rect 34388 18232 34394 18244
rect 34425 18241 34437 18244
rect 34471 18241 34483 18275
rect 36170 18272 36176 18284
rect 34425 18235 34483 18241
rect 34532 18244 36176 18272
rect 27448 18176 28764 18204
rect 30285 18207 30343 18213
rect 17773 18139 17831 18145
rect 17773 18105 17785 18139
rect 17819 18136 17831 18139
rect 21634 18136 21640 18148
rect 17819 18108 18828 18136
rect 17819 18105 17831 18108
rect 17773 18099 17831 18105
rect 2317 18071 2375 18077
rect 2317 18037 2329 18071
rect 2363 18068 2375 18071
rect 17218 18068 17224 18080
rect 2363 18040 17224 18068
rect 2363 18037 2375 18040
rect 2317 18031 2375 18037
rect 17218 18028 17224 18040
rect 17276 18028 17282 18080
rect 18325 18071 18383 18077
rect 18325 18037 18337 18071
rect 18371 18068 18383 18071
rect 18414 18068 18420 18080
rect 18371 18040 18420 18068
rect 18371 18037 18383 18040
rect 18325 18031 18383 18037
rect 18414 18028 18420 18040
rect 18472 18028 18478 18080
rect 18800 18068 18828 18108
rect 19996 18108 21640 18136
rect 19996 18068 20024 18108
rect 21634 18096 21640 18108
rect 21692 18096 21698 18148
rect 27448 18145 27476 18176
rect 30285 18173 30297 18207
rect 30331 18204 30343 18207
rect 33226 18204 33232 18216
rect 30331 18176 33232 18204
rect 30331 18173 30343 18176
rect 30285 18167 30343 18173
rect 33226 18164 33232 18176
rect 33284 18164 33290 18216
rect 33413 18207 33471 18213
rect 33413 18173 33425 18207
rect 33459 18204 33471 18207
rect 33594 18204 33600 18216
rect 33459 18176 33600 18204
rect 33459 18173 33471 18176
rect 33413 18167 33471 18173
rect 33594 18164 33600 18176
rect 33652 18164 33658 18216
rect 33689 18207 33747 18213
rect 33689 18173 33701 18207
rect 33735 18204 33747 18207
rect 34532 18204 34560 18244
rect 36170 18232 36176 18244
rect 36228 18232 36234 18284
rect 37642 18272 37648 18284
rect 37603 18244 37648 18272
rect 37642 18232 37648 18244
rect 37700 18232 37706 18284
rect 38381 18275 38439 18281
rect 37752 18244 38312 18272
rect 36265 18207 36323 18213
rect 36265 18204 36277 18207
rect 33735 18176 34560 18204
rect 35820 18176 36277 18204
rect 33735 18173 33747 18176
rect 33689 18167 33747 18173
rect 27433 18139 27491 18145
rect 27433 18105 27445 18139
rect 27479 18105 27491 18139
rect 27433 18099 27491 18105
rect 27522 18096 27528 18148
rect 27580 18136 27586 18148
rect 27893 18139 27951 18145
rect 27893 18136 27905 18139
rect 27580 18108 27905 18136
rect 27580 18096 27586 18108
rect 27893 18105 27905 18108
rect 27939 18136 27951 18139
rect 28626 18136 28632 18148
rect 27939 18108 28632 18136
rect 27939 18105 27951 18108
rect 27893 18099 27951 18105
rect 28626 18096 28632 18108
rect 28684 18096 28690 18148
rect 29270 18136 29276 18148
rect 28736 18108 29276 18136
rect 18800 18040 20024 18068
rect 20165 18071 20223 18077
rect 20165 18037 20177 18071
rect 20211 18068 20223 18071
rect 20622 18068 20628 18080
rect 20211 18040 20628 18068
rect 20211 18037 20223 18040
rect 20165 18031 20223 18037
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 22646 18068 22652 18080
rect 22607 18040 22652 18068
rect 22646 18028 22652 18040
rect 22704 18028 22710 18080
rect 24489 18071 24547 18077
rect 24489 18037 24501 18071
rect 24535 18068 24547 18071
rect 24946 18068 24952 18080
rect 24535 18040 24952 18068
rect 24535 18037 24547 18040
rect 24489 18031 24547 18037
rect 24946 18028 24952 18040
rect 25004 18068 25010 18080
rect 26329 18071 26387 18077
rect 26329 18068 26341 18071
rect 25004 18040 26341 18068
rect 25004 18028 25010 18040
rect 26329 18037 26341 18040
rect 26375 18068 26387 18071
rect 28736 18068 28764 18108
rect 29270 18096 29276 18108
rect 29328 18096 29334 18148
rect 31113 18139 31171 18145
rect 31113 18105 31125 18139
rect 31159 18136 31171 18139
rect 33134 18136 33140 18148
rect 31159 18108 33140 18136
rect 31159 18105 31171 18108
rect 31113 18099 31171 18105
rect 33134 18096 33140 18108
rect 33192 18096 33198 18148
rect 33704 18136 33732 18167
rect 35820 18148 35848 18176
rect 36265 18173 36277 18176
rect 36311 18173 36323 18207
rect 36265 18167 36323 18173
rect 36538 18164 36544 18216
rect 36596 18204 36602 18216
rect 37752 18204 37780 18244
rect 36596 18176 37780 18204
rect 36596 18164 36602 18176
rect 38102 18164 38108 18216
rect 38160 18204 38166 18216
rect 38197 18207 38255 18213
rect 38197 18204 38209 18207
rect 38160 18176 38209 18204
rect 38160 18164 38166 18176
rect 38197 18173 38209 18176
rect 38243 18173 38255 18207
rect 38284 18204 38312 18244
rect 38381 18241 38393 18275
rect 38427 18270 38439 18275
rect 38930 18272 38936 18284
rect 38626 18270 38936 18272
rect 38427 18244 38936 18270
rect 38427 18242 38654 18244
rect 38427 18241 38439 18242
rect 38381 18235 38439 18241
rect 38930 18232 38936 18244
rect 38988 18232 38994 18284
rect 39209 18275 39267 18281
rect 39209 18241 39221 18275
rect 39255 18241 39267 18275
rect 39850 18272 39856 18284
rect 39811 18244 39856 18272
rect 39209 18235 39267 18241
rect 39224 18204 39252 18235
rect 39850 18232 39856 18244
rect 39908 18232 39914 18284
rect 39942 18232 39948 18284
rect 40000 18272 40006 18284
rect 40681 18275 40739 18281
rect 40681 18272 40693 18275
rect 40000 18244 40693 18272
rect 40000 18232 40006 18244
rect 40681 18241 40693 18244
rect 40727 18241 40739 18275
rect 40681 18235 40739 18241
rect 41322 18232 41328 18284
rect 41380 18272 41386 18284
rect 41509 18275 41567 18281
rect 41509 18272 41521 18275
rect 41380 18244 41521 18272
rect 41380 18232 41386 18244
rect 41509 18241 41521 18244
rect 41555 18241 41567 18275
rect 41509 18235 41567 18241
rect 41598 18232 41604 18284
rect 41656 18232 41662 18284
rect 41874 18232 41880 18284
rect 41932 18272 41938 18284
rect 42705 18275 42763 18281
rect 42705 18272 42717 18275
rect 41932 18244 42717 18272
rect 41932 18232 41938 18244
rect 42705 18241 42717 18244
rect 42751 18272 42763 18275
rect 49878 18272 49884 18284
rect 42751 18244 49884 18272
rect 42751 18241 42763 18244
rect 42705 18235 42763 18241
rect 49878 18232 49884 18244
rect 49936 18232 49942 18284
rect 54021 18275 54079 18281
rect 54021 18272 54033 18275
rect 53484 18244 54033 18272
rect 38284 18176 39252 18204
rect 38197 18167 38255 18173
rect 39298 18164 39304 18216
rect 39356 18204 39362 18216
rect 39669 18207 39727 18213
rect 39669 18204 39681 18207
rect 39356 18176 39681 18204
rect 39356 18164 39362 18176
rect 39669 18173 39681 18176
rect 39715 18173 39727 18207
rect 39669 18167 39727 18173
rect 39758 18164 39764 18216
rect 39816 18204 39822 18216
rect 40402 18204 40408 18216
rect 39816 18176 40408 18204
rect 39816 18164 39822 18176
rect 40402 18164 40408 18176
rect 40460 18164 40466 18216
rect 40494 18164 40500 18216
rect 40552 18204 40558 18216
rect 41616 18204 41644 18232
rect 40552 18176 40597 18204
rect 40696 18176 41644 18204
rect 40552 18164 40558 18176
rect 35802 18136 35808 18148
rect 33612 18108 33732 18136
rect 35763 18108 35808 18136
rect 26375 18040 28764 18068
rect 26375 18037 26387 18040
rect 26329 18031 26387 18037
rect 28810 18028 28816 18080
rect 28868 18068 28874 18080
rect 28905 18071 28963 18077
rect 28905 18068 28917 18071
rect 28868 18040 28917 18068
rect 28868 18028 28874 18040
rect 28905 18037 28917 18040
rect 28951 18068 28963 18071
rect 30282 18068 30288 18080
rect 28951 18040 30288 18068
rect 28951 18037 28963 18040
rect 28905 18031 28963 18037
rect 30282 18028 30288 18040
rect 30340 18028 30346 18080
rect 32306 18068 32312 18080
rect 32267 18040 32312 18068
rect 32306 18028 32312 18040
rect 32364 18068 32370 18080
rect 33612 18068 33640 18108
rect 35802 18096 35808 18108
rect 35860 18096 35866 18148
rect 36814 18096 36820 18148
rect 36872 18136 36878 18148
rect 36872 18108 38424 18136
rect 36872 18096 36878 18108
rect 32364 18040 33640 18068
rect 32364 18028 32370 18040
rect 34422 18028 34428 18080
rect 34480 18068 34486 18080
rect 36354 18068 36360 18080
rect 34480 18040 36360 18068
rect 34480 18028 34486 18040
rect 36354 18028 36360 18040
rect 36412 18068 36418 18080
rect 36909 18071 36967 18077
rect 36909 18068 36921 18071
rect 36412 18040 36921 18068
rect 36412 18028 36418 18040
rect 36909 18037 36921 18040
rect 36955 18037 36967 18071
rect 36909 18031 36967 18037
rect 37553 18071 37611 18077
rect 37553 18037 37565 18071
rect 37599 18068 37611 18071
rect 37826 18068 37832 18080
rect 37599 18040 37832 18068
rect 37599 18037 37611 18040
rect 37553 18031 37611 18037
rect 37826 18028 37832 18040
rect 37884 18028 37890 18080
rect 38102 18028 38108 18080
rect 38160 18068 38166 18080
rect 38286 18068 38292 18080
rect 38160 18040 38292 18068
rect 38160 18028 38166 18040
rect 38286 18028 38292 18040
rect 38344 18028 38350 18080
rect 38396 18068 38424 18108
rect 38470 18096 38476 18148
rect 38528 18136 38534 18148
rect 40037 18139 40095 18145
rect 38528 18108 39160 18136
rect 38528 18096 38534 18108
rect 39025 18071 39083 18077
rect 39025 18068 39037 18071
rect 38396 18040 39037 18068
rect 39025 18037 39037 18040
rect 39071 18037 39083 18071
rect 39132 18068 39160 18108
rect 40037 18105 40049 18139
rect 40083 18136 40095 18139
rect 40696 18136 40724 18176
rect 40083 18108 40724 18136
rect 40865 18139 40923 18145
rect 40083 18105 40095 18108
rect 40037 18099 40095 18105
rect 40865 18105 40877 18139
rect 40911 18136 40923 18139
rect 41690 18136 41696 18148
rect 40911 18108 41696 18136
rect 40911 18105 40923 18108
rect 40865 18099 40923 18105
rect 41690 18096 41696 18108
rect 41748 18096 41754 18148
rect 53484 18080 53512 18244
rect 54021 18241 54033 18244
rect 54067 18241 54079 18275
rect 54021 18235 54079 18241
rect 41325 18071 41383 18077
rect 41325 18068 41337 18071
rect 39132 18040 41337 18068
rect 39025 18031 39083 18037
rect 41325 18037 41337 18040
rect 41371 18037 41383 18071
rect 41325 18031 41383 18037
rect 41506 18028 41512 18080
rect 41564 18068 41570 18080
rect 43254 18068 43260 18080
rect 41564 18040 43260 18068
rect 41564 18028 41570 18040
rect 43254 18028 43260 18040
rect 43312 18028 43318 18080
rect 53466 18068 53472 18080
rect 53427 18040 53472 18068
rect 53466 18028 53472 18040
rect 53524 18028 53530 18080
rect 1104 17978 54832 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 54832 17978
rect 1104 17904 54832 17926
rect 22462 17824 22468 17876
rect 22520 17864 22526 17876
rect 23109 17867 23167 17873
rect 23109 17864 23121 17867
rect 22520 17836 23121 17864
rect 22520 17824 22526 17836
rect 23109 17833 23121 17836
rect 23155 17833 23167 17867
rect 23109 17827 23167 17833
rect 24118 17824 24124 17876
rect 24176 17864 24182 17876
rect 24581 17867 24639 17873
rect 24581 17864 24593 17867
rect 24176 17836 24593 17864
rect 24176 17824 24182 17836
rect 24581 17833 24593 17836
rect 24627 17833 24639 17867
rect 24581 17827 24639 17833
rect 25038 17824 25044 17876
rect 25096 17864 25102 17876
rect 25096 17836 27016 17864
rect 25096 17824 25102 17836
rect 21269 17799 21327 17805
rect 21269 17765 21281 17799
rect 21315 17765 21327 17799
rect 21269 17759 21327 17765
rect 22649 17799 22707 17805
rect 22649 17765 22661 17799
rect 22695 17796 22707 17799
rect 23198 17796 23204 17808
rect 22695 17768 23204 17796
rect 22695 17765 22707 17768
rect 22649 17759 22707 17765
rect 18230 17728 18236 17740
rect 18191 17700 18236 17728
rect 18230 17688 18236 17700
rect 18288 17688 18294 17740
rect 19334 17688 19340 17740
rect 19392 17728 19398 17740
rect 19429 17731 19487 17737
rect 19429 17728 19441 17731
rect 19392 17700 19441 17728
rect 19392 17688 19398 17700
rect 19429 17697 19441 17700
rect 19475 17697 19487 17731
rect 19429 17691 19487 17697
rect 1857 17663 1915 17669
rect 1857 17629 1869 17663
rect 1903 17660 1915 17663
rect 15378 17660 15384 17672
rect 1903 17632 15384 17660
rect 1903 17629 1915 17632
rect 1857 17623 1915 17629
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17660 18751 17663
rect 21284 17660 21312 17759
rect 23198 17756 23204 17768
rect 23256 17756 23262 17808
rect 23842 17756 23848 17808
rect 23900 17796 23906 17808
rect 26878 17796 26884 17808
rect 23900 17768 26884 17796
rect 23900 17756 23906 17768
rect 26878 17756 26884 17768
rect 26936 17756 26942 17808
rect 26988 17796 27016 17836
rect 27982 17824 27988 17876
rect 28040 17864 28046 17876
rect 30929 17867 30987 17873
rect 30929 17864 30941 17867
rect 28040 17836 30941 17864
rect 28040 17824 28046 17836
rect 30929 17833 30941 17836
rect 30975 17833 30987 17867
rect 54110 17864 54116 17876
rect 30929 17827 30987 17833
rect 31726 17836 54116 17864
rect 31726 17796 31754 17836
rect 54110 17824 54116 17836
rect 54168 17824 54174 17876
rect 26988 17768 31754 17796
rect 33965 17799 34023 17805
rect 33965 17765 33977 17799
rect 34011 17796 34023 17799
rect 34514 17796 34520 17808
rect 34011 17768 34520 17796
rect 34011 17765 34023 17768
rect 33965 17759 34023 17765
rect 34514 17756 34520 17768
rect 34572 17756 34578 17808
rect 36998 17796 37004 17808
rect 35360 17768 37004 17796
rect 21913 17731 21971 17737
rect 21913 17697 21925 17731
rect 21959 17728 21971 17731
rect 22002 17728 22008 17740
rect 21959 17700 22008 17728
rect 21959 17697 21971 17700
rect 21913 17691 21971 17697
rect 22002 17688 22008 17700
rect 22060 17688 22066 17740
rect 24026 17728 24032 17740
rect 23032 17700 24032 17728
rect 21634 17660 21640 17672
rect 18739 17632 21312 17660
rect 21595 17632 21640 17660
rect 18739 17629 18751 17632
rect 18693 17623 18751 17629
rect 21634 17620 21640 17632
rect 21692 17620 21698 17672
rect 22465 17663 22523 17669
rect 22465 17629 22477 17663
rect 22511 17660 22523 17663
rect 22554 17660 22560 17672
rect 22511 17632 22560 17660
rect 22511 17629 22523 17632
rect 22465 17623 22523 17629
rect 22554 17620 22560 17632
rect 22612 17620 22618 17672
rect 18230 17552 18236 17604
rect 18288 17592 18294 17604
rect 18288 17564 19380 17592
rect 18288 17552 18294 17564
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 17126 17524 17132 17536
rect 17087 17496 17132 17524
rect 17126 17484 17132 17496
rect 17184 17484 17190 17536
rect 17678 17524 17684 17536
rect 17639 17496 17684 17524
rect 17678 17484 17684 17496
rect 17736 17484 17742 17536
rect 18877 17527 18935 17533
rect 18877 17493 18889 17527
rect 18923 17524 18935 17527
rect 19242 17524 19248 17536
rect 18923 17496 19248 17524
rect 18923 17493 18935 17496
rect 18877 17487 18935 17493
rect 19242 17484 19248 17496
rect 19300 17484 19306 17536
rect 19352 17524 19380 17564
rect 19426 17552 19432 17604
rect 19484 17592 19490 17604
rect 19674 17595 19732 17601
rect 19674 17592 19686 17595
rect 19484 17564 19686 17592
rect 19484 17552 19490 17564
rect 19674 17561 19686 17564
rect 19720 17561 19732 17595
rect 23032 17592 23060 17700
rect 24026 17688 24032 17700
rect 24084 17688 24090 17740
rect 25130 17728 25136 17740
rect 25091 17700 25136 17728
rect 25130 17688 25136 17700
rect 25188 17688 25194 17740
rect 27522 17728 27528 17740
rect 27483 17700 27528 17728
rect 27522 17688 27528 17700
rect 27580 17688 27586 17740
rect 27706 17688 27712 17740
rect 27764 17728 27770 17740
rect 27764 17700 27809 17728
rect 27764 17688 27770 17700
rect 28350 17688 28356 17740
rect 28408 17728 28414 17740
rect 28537 17731 28595 17737
rect 28537 17728 28549 17731
rect 28408 17700 28549 17728
rect 28408 17688 28414 17700
rect 28537 17697 28549 17700
rect 28583 17697 28595 17731
rect 28537 17691 28595 17697
rect 28902 17688 28908 17740
rect 28960 17728 28966 17740
rect 29362 17728 29368 17740
rect 28960 17700 29368 17728
rect 28960 17688 28966 17700
rect 29362 17688 29368 17700
rect 29420 17728 29426 17740
rect 29917 17731 29975 17737
rect 29917 17728 29929 17731
rect 29420 17700 29929 17728
rect 29420 17688 29426 17700
rect 29917 17697 29929 17700
rect 29963 17728 29975 17731
rect 30098 17728 30104 17740
rect 29963 17700 30104 17728
rect 29963 17697 29975 17700
rect 29917 17691 29975 17697
rect 30098 17688 30104 17700
rect 30156 17688 30162 17740
rect 30282 17688 30288 17740
rect 30340 17688 30346 17740
rect 30374 17688 30380 17740
rect 30432 17728 30438 17740
rect 32493 17731 32551 17737
rect 32493 17728 32505 17731
rect 30432 17700 32505 17728
rect 30432 17688 30438 17700
rect 32493 17697 32505 17700
rect 32539 17728 32551 17731
rect 33134 17728 33140 17740
rect 32539 17700 33140 17728
rect 32539 17697 32551 17700
rect 32493 17691 32551 17697
rect 33134 17688 33140 17700
rect 33192 17688 33198 17740
rect 33689 17731 33747 17737
rect 33689 17697 33701 17731
rect 33735 17728 33747 17731
rect 35360 17728 35388 17768
rect 36998 17756 37004 17768
rect 37056 17756 37062 17808
rect 38010 17756 38016 17808
rect 38068 17796 38074 17808
rect 41322 17796 41328 17808
rect 38068 17768 41328 17796
rect 38068 17756 38074 17768
rect 41322 17756 41328 17768
rect 41380 17756 41386 17808
rect 41414 17756 41420 17808
rect 41472 17796 41478 17808
rect 41509 17799 41567 17805
rect 41509 17796 41521 17799
rect 41472 17768 41521 17796
rect 41472 17756 41478 17768
rect 41509 17765 41521 17768
rect 41555 17765 41567 17799
rect 41509 17759 41567 17765
rect 41598 17756 41604 17808
rect 41656 17796 41662 17808
rect 42153 17799 42211 17805
rect 42153 17796 42165 17799
rect 41656 17768 42165 17796
rect 41656 17756 41662 17768
rect 42153 17765 42165 17768
rect 42199 17765 42211 17799
rect 42153 17759 42211 17765
rect 42797 17799 42855 17805
rect 42797 17765 42809 17799
rect 42843 17796 42855 17799
rect 49694 17796 49700 17808
rect 42843 17768 49700 17796
rect 42843 17765 42855 17768
rect 42797 17759 42855 17765
rect 33735 17700 35388 17728
rect 33735 17697 33747 17700
rect 33689 17691 33747 17697
rect 35526 17688 35532 17740
rect 35584 17728 35590 17740
rect 35584 17700 36308 17728
rect 35584 17688 35590 17700
rect 23293 17663 23351 17669
rect 23293 17629 23305 17663
rect 23339 17629 23351 17663
rect 23293 17623 23351 17629
rect 19674 17555 19732 17561
rect 19812 17564 23060 17592
rect 23308 17592 23336 17623
rect 23382 17620 23388 17672
rect 23440 17660 23446 17672
rect 23440 17632 23485 17660
rect 23440 17620 23446 17632
rect 24670 17620 24676 17672
rect 24728 17660 24734 17672
rect 25777 17663 25835 17669
rect 25777 17660 25789 17663
rect 24728 17632 25789 17660
rect 24728 17620 24734 17632
rect 25777 17629 25789 17632
rect 25823 17629 25835 17663
rect 25777 17623 25835 17629
rect 27433 17663 27491 17669
rect 27433 17629 27445 17663
rect 27479 17629 27491 17663
rect 27433 17623 27491 17629
rect 27617 17663 27675 17669
rect 27617 17629 27629 17663
rect 27663 17629 27675 17663
rect 28810 17660 28816 17672
rect 28771 17632 28816 17660
rect 27617 17623 27675 17629
rect 24578 17592 24584 17604
rect 23308 17564 24584 17592
rect 19812 17524 19840 17564
rect 24578 17552 24584 17564
rect 24636 17552 24642 17604
rect 27448 17592 27476 17623
rect 24688 17564 27476 17592
rect 27632 17592 27660 17623
rect 28810 17620 28816 17632
rect 28868 17620 28874 17672
rect 29454 17660 29460 17672
rect 28966 17632 29460 17660
rect 28966 17592 28994 17632
rect 29454 17620 29460 17632
rect 29512 17620 29518 17672
rect 27632 17564 28994 17592
rect 30101 17595 30159 17601
rect 19352 17496 19840 17524
rect 20714 17484 20720 17536
rect 20772 17524 20778 17536
rect 20809 17527 20867 17533
rect 20809 17524 20821 17527
rect 20772 17496 20821 17524
rect 20772 17484 20778 17496
rect 20809 17493 20821 17496
rect 20855 17493 20867 17527
rect 21726 17524 21732 17536
rect 21687 17496 21732 17524
rect 20809 17487 20867 17493
rect 21726 17484 21732 17496
rect 21784 17484 21790 17536
rect 21818 17484 21824 17536
rect 21876 17524 21882 17536
rect 23842 17524 23848 17536
rect 21876 17496 23848 17524
rect 21876 17484 21882 17496
rect 23842 17484 23848 17496
rect 23900 17484 23906 17536
rect 24026 17524 24032 17536
rect 23987 17496 24032 17524
rect 24026 17484 24032 17496
rect 24084 17484 24090 17536
rect 24118 17484 24124 17536
rect 24176 17524 24182 17536
rect 24688 17524 24716 17564
rect 30101 17561 30113 17595
rect 30147 17592 30159 17595
rect 30300 17592 30328 17688
rect 31113 17663 31171 17669
rect 31113 17660 31125 17663
rect 30147 17564 30328 17592
rect 30484 17632 31125 17660
rect 30147 17561 30159 17564
rect 30101 17555 30159 17561
rect 24946 17524 24952 17536
rect 24176 17496 24716 17524
rect 24907 17496 24952 17524
rect 24176 17484 24182 17496
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 25038 17484 25044 17536
rect 25096 17524 25102 17536
rect 25096 17496 25141 17524
rect 25096 17484 25102 17496
rect 26142 17484 26148 17536
rect 26200 17524 26206 17536
rect 26421 17527 26479 17533
rect 26421 17524 26433 17527
rect 26200 17496 26433 17524
rect 26200 17484 26206 17496
rect 26421 17493 26433 17496
rect 26467 17493 26479 17527
rect 27890 17524 27896 17536
rect 27851 17496 27896 17524
rect 26421 17487 26479 17493
rect 27890 17484 27896 17496
rect 27948 17484 27954 17536
rect 27982 17484 27988 17536
rect 28040 17524 28046 17536
rect 28721 17527 28779 17533
rect 28721 17524 28733 17527
rect 28040 17496 28733 17524
rect 28040 17484 28046 17496
rect 28721 17493 28733 17496
rect 28767 17524 28779 17527
rect 29086 17524 29092 17536
rect 28767 17496 29092 17524
rect 28767 17493 28779 17496
rect 28721 17487 28779 17493
rect 29086 17484 29092 17496
rect 29144 17484 29150 17536
rect 29181 17527 29239 17533
rect 29181 17493 29193 17527
rect 29227 17524 29239 17527
rect 29822 17524 29828 17536
rect 29227 17496 29828 17524
rect 29227 17493 29239 17496
rect 29181 17487 29239 17493
rect 29822 17484 29828 17496
rect 29880 17484 29886 17536
rect 30009 17527 30067 17533
rect 30009 17493 30021 17527
rect 30055 17524 30067 17527
rect 30374 17524 30380 17536
rect 30055 17496 30380 17524
rect 30055 17493 30067 17496
rect 30009 17487 30067 17493
rect 30374 17484 30380 17496
rect 30432 17484 30438 17536
rect 30484 17533 30512 17632
rect 31113 17629 31125 17632
rect 31159 17629 31171 17663
rect 31113 17623 31171 17629
rect 31297 17663 31355 17669
rect 31297 17629 31309 17663
rect 31343 17660 31355 17663
rect 31386 17660 31392 17672
rect 31343 17632 31392 17660
rect 31343 17629 31355 17632
rect 31297 17623 31355 17629
rect 31386 17620 31392 17632
rect 31444 17620 31450 17672
rect 32217 17663 32275 17669
rect 32217 17629 32229 17663
rect 32263 17660 32275 17663
rect 32306 17660 32312 17672
rect 32263 17632 32312 17660
rect 32263 17629 32275 17632
rect 32217 17623 32275 17629
rect 32306 17620 32312 17632
rect 32364 17620 32370 17672
rect 33597 17663 33655 17669
rect 33597 17629 33609 17663
rect 33643 17660 33655 17663
rect 34422 17660 34428 17672
rect 33643 17632 34428 17660
rect 33643 17629 33655 17632
rect 33597 17623 33655 17629
rect 34422 17620 34428 17632
rect 34480 17620 34486 17672
rect 34514 17620 34520 17672
rect 34572 17660 34578 17672
rect 35253 17663 35311 17669
rect 35253 17660 35265 17663
rect 34572 17632 35265 17660
rect 34572 17620 34578 17632
rect 35253 17629 35265 17632
rect 35299 17660 35311 17663
rect 35802 17660 35808 17672
rect 35299 17632 35808 17660
rect 35299 17629 35311 17632
rect 35253 17623 35311 17629
rect 35802 17620 35808 17632
rect 35860 17620 35866 17672
rect 36280 17660 36308 17700
rect 38102 17688 38108 17740
rect 38160 17728 38166 17740
rect 40126 17728 40132 17740
rect 38160 17700 40132 17728
rect 38160 17688 38166 17700
rect 40126 17688 40132 17700
rect 40184 17688 40190 17740
rect 40218 17688 40224 17740
rect 40276 17728 40282 17740
rect 42812 17728 42840 17759
rect 49694 17756 49700 17768
rect 49752 17756 49758 17808
rect 54202 17796 54208 17808
rect 54163 17768 54208 17796
rect 54202 17756 54208 17768
rect 54260 17756 54266 17808
rect 40276 17700 42840 17728
rect 40276 17688 40282 17700
rect 37458 17660 37464 17672
rect 36280 17632 37464 17660
rect 37458 17620 37464 17632
rect 37516 17620 37522 17672
rect 37918 17620 37924 17672
rect 37976 17660 37982 17672
rect 38013 17663 38071 17669
rect 38013 17660 38025 17663
rect 37976 17632 38025 17660
rect 37976 17620 37982 17632
rect 38013 17629 38025 17632
rect 38059 17629 38071 17663
rect 38654 17660 38660 17672
rect 38615 17632 38660 17660
rect 38013 17623 38071 17629
rect 38654 17620 38660 17632
rect 38712 17620 38718 17672
rect 38838 17660 38844 17672
rect 38799 17632 38844 17660
rect 38838 17620 38844 17632
rect 38896 17620 38902 17672
rect 39025 17663 39083 17669
rect 39025 17629 39037 17663
rect 39071 17660 39083 17663
rect 39298 17660 39304 17672
rect 39071 17632 39304 17660
rect 39071 17629 39083 17632
rect 39025 17623 39083 17629
rect 39298 17620 39304 17632
rect 39356 17620 39362 17672
rect 39684 17632 40264 17660
rect 30742 17552 30748 17604
rect 30800 17592 30806 17604
rect 37768 17595 37826 17601
rect 30800 17564 36768 17592
rect 30800 17552 30806 17564
rect 30469 17527 30527 17533
rect 30469 17493 30481 17527
rect 30515 17493 30527 17527
rect 31846 17524 31852 17536
rect 31807 17496 31852 17524
rect 30469 17487 30527 17493
rect 31846 17484 31852 17496
rect 31904 17484 31910 17536
rect 32309 17527 32367 17533
rect 32309 17493 32321 17527
rect 32355 17524 32367 17527
rect 32398 17524 32404 17536
rect 32355 17496 32404 17524
rect 32355 17493 32367 17496
rect 32309 17487 32367 17493
rect 32398 17484 32404 17496
rect 32456 17484 32462 17536
rect 34790 17484 34796 17536
rect 34848 17524 34854 17536
rect 34885 17527 34943 17533
rect 34885 17524 34897 17527
rect 34848 17496 34897 17524
rect 34848 17484 34854 17496
rect 34885 17493 34897 17496
rect 34931 17493 34943 17527
rect 34885 17487 34943 17493
rect 35158 17484 35164 17536
rect 35216 17524 35222 17536
rect 35342 17524 35348 17536
rect 35216 17496 35348 17524
rect 35216 17484 35222 17496
rect 35342 17484 35348 17496
rect 35400 17484 35406 17536
rect 36078 17524 36084 17536
rect 36039 17496 36084 17524
rect 36078 17484 36084 17496
rect 36136 17484 36142 17536
rect 36630 17524 36636 17536
rect 36591 17496 36636 17524
rect 36630 17484 36636 17496
rect 36688 17484 36694 17536
rect 36740 17524 36768 17564
rect 37768 17561 37780 17595
rect 37814 17592 37826 17595
rect 38470 17592 38476 17604
rect 37814 17564 38476 17592
rect 37814 17561 37826 17564
rect 37768 17555 37826 17561
rect 38470 17552 38476 17564
rect 38528 17552 38534 17604
rect 38930 17592 38936 17604
rect 38843 17564 38936 17592
rect 38930 17552 38936 17564
rect 38988 17592 38994 17604
rect 39684 17592 39712 17632
rect 40126 17592 40132 17604
rect 38988 17564 39712 17592
rect 40087 17564 40132 17592
rect 38988 17552 38994 17564
rect 40126 17552 40132 17564
rect 40184 17552 40190 17604
rect 40236 17592 40264 17632
rect 40310 17620 40316 17672
rect 40368 17660 40374 17672
rect 40773 17663 40831 17669
rect 40368 17632 40413 17660
rect 40368 17620 40374 17632
rect 40773 17629 40785 17663
rect 40819 17660 40831 17663
rect 41138 17660 41144 17672
rect 40819 17632 41144 17660
rect 40819 17629 40831 17632
rect 40773 17623 40831 17629
rect 41138 17620 41144 17632
rect 41196 17660 41202 17672
rect 41322 17660 41328 17672
rect 41196 17632 41328 17660
rect 41196 17620 41202 17632
rect 41322 17620 41328 17632
rect 41380 17620 41386 17672
rect 41690 17660 41696 17672
rect 41651 17632 41696 17660
rect 41690 17620 41696 17632
rect 41748 17620 41754 17672
rect 54021 17663 54079 17669
rect 54021 17660 54033 17663
rect 51046 17632 54033 17660
rect 51046 17592 51074 17632
rect 54021 17629 54033 17632
rect 54067 17629 54079 17663
rect 54021 17623 54079 17629
rect 40236 17564 51074 17592
rect 39022 17524 39028 17536
rect 36740 17496 39028 17524
rect 39022 17484 39028 17496
rect 39080 17484 39086 17536
rect 39114 17484 39120 17536
rect 39172 17524 39178 17536
rect 39209 17527 39267 17533
rect 39209 17524 39221 17527
rect 39172 17496 39221 17524
rect 39172 17484 39178 17496
rect 39209 17493 39221 17496
rect 39255 17493 39267 17527
rect 39209 17487 39267 17493
rect 39298 17484 39304 17536
rect 39356 17524 39362 17536
rect 40957 17527 41015 17533
rect 40957 17524 40969 17527
rect 39356 17496 40969 17524
rect 39356 17484 39362 17496
rect 40957 17493 40969 17496
rect 41003 17493 41015 17527
rect 43254 17524 43260 17536
rect 43215 17496 43260 17524
rect 40957 17487 41015 17493
rect 43254 17484 43260 17496
rect 43312 17484 43318 17536
rect 53561 17527 53619 17533
rect 53561 17493 53573 17527
rect 53607 17524 53619 17527
rect 54202 17524 54208 17536
rect 53607 17496 54208 17524
rect 53607 17493 53619 17496
rect 53561 17487 53619 17493
rect 54202 17484 54208 17496
rect 54260 17484 54266 17536
rect 1104 17434 54832 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 54832 17434
rect 1104 17360 54832 17382
rect 17218 17320 17224 17332
rect 17179 17292 17224 17320
rect 17218 17280 17224 17292
rect 17276 17320 17282 17332
rect 19334 17320 19340 17332
rect 17276 17292 19340 17320
rect 17276 17280 17282 17292
rect 19334 17280 19340 17292
rect 19392 17280 19398 17332
rect 24394 17320 24400 17332
rect 22112 17292 24400 17320
rect 16301 17255 16359 17261
rect 16301 17221 16313 17255
rect 16347 17252 16359 17255
rect 18138 17252 18144 17264
rect 16347 17224 18144 17252
rect 16347 17221 16359 17224
rect 16301 17215 16359 17221
rect 18138 17212 18144 17224
rect 18196 17212 18202 17264
rect 20073 17255 20131 17261
rect 20073 17221 20085 17255
rect 20119 17252 20131 17255
rect 21358 17252 21364 17264
rect 20119 17224 21364 17252
rect 20119 17221 20131 17224
rect 20073 17215 20131 17221
rect 21358 17212 21364 17224
rect 21416 17212 21422 17264
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 16482 17184 16488 17196
rect 1903 17156 16488 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 16482 17144 16488 17156
rect 16540 17144 16546 17196
rect 17126 17144 17132 17196
rect 17184 17184 17190 17196
rect 21085 17187 21143 17193
rect 21085 17184 21097 17187
rect 17184 17156 21097 17184
rect 17184 17144 17190 17156
rect 21085 17153 21097 17156
rect 21131 17184 21143 17187
rect 21818 17184 21824 17196
rect 21131 17156 21824 17184
rect 21131 17153 21143 17156
rect 21085 17147 21143 17153
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 22112 17193 22140 17292
rect 24394 17280 24400 17292
rect 24452 17280 24458 17332
rect 24670 17320 24676 17332
rect 24631 17292 24676 17320
rect 24670 17280 24676 17292
rect 24728 17280 24734 17332
rect 27157 17323 27215 17329
rect 27157 17320 27169 17323
rect 24780 17292 27169 17320
rect 22646 17212 22652 17264
rect 22704 17252 22710 17264
rect 22986 17255 23044 17261
rect 22986 17252 22998 17255
rect 22704 17224 22998 17252
rect 22704 17212 22710 17224
rect 22986 17221 22998 17224
rect 23032 17221 23044 17255
rect 22986 17215 23044 17221
rect 22097 17187 22155 17193
rect 22097 17153 22109 17187
rect 22143 17153 22155 17187
rect 22097 17147 22155 17153
rect 22370 17144 22376 17196
rect 22428 17184 22434 17196
rect 22428 17156 23796 17184
rect 22428 17144 22434 17156
rect 18322 17116 18328 17128
rect 18283 17088 18328 17116
rect 18322 17076 18328 17088
rect 18380 17076 18386 17128
rect 20898 17116 20904 17128
rect 20859 17088 20904 17116
rect 20898 17076 20904 17088
rect 20956 17076 20962 17128
rect 20993 17119 21051 17125
rect 20993 17085 21005 17119
rect 21039 17085 21051 17119
rect 20993 17079 21051 17085
rect 20070 17008 20076 17060
rect 20128 17048 20134 17060
rect 21008 17048 21036 17079
rect 22186 17076 22192 17128
rect 22244 17116 22250 17128
rect 22741 17119 22799 17125
rect 22741 17116 22753 17119
rect 22244 17088 22753 17116
rect 22244 17076 22250 17088
rect 22741 17085 22753 17088
rect 22787 17085 22799 17119
rect 23768 17116 23796 17156
rect 23934 17144 23940 17196
rect 23992 17184 23998 17196
rect 24581 17187 24639 17193
rect 24581 17184 24593 17187
rect 23992 17156 24593 17184
rect 23992 17144 23998 17156
rect 24581 17153 24593 17156
rect 24627 17184 24639 17187
rect 24670 17184 24676 17196
rect 24627 17156 24676 17184
rect 24627 17153 24639 17156
rect 24581 17147 24639 17153
rect 24670 17144 24676 17156
rect 24728 17144 24734 17196
rect 24780 17193 24808 17292
rect 27157 17289 27169 17292
rect 27203 17289 27215 17323
rect 27157 17283 27215 17289
rect 27890 17280 27896 17332
rect 27948 17320 27954 17332
rect 36725 17323 36783 17329
rect 27948 17292 36216 17320
rect 27948 17280 27954 17292
rect 25406 17212 25412 17264
rect 25464 17252 25470 17264
rect 25958 17252 25964 17264
rect 25464 17224 25964 17252
rect 25464 17212 25470 17224
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 26142 17212 26148 17264
rect 26200 17252 26206 17264
rect 26338 17255 26396 17261
rect 26338 17252 26350 17255
rect 26200 17224 26350 17252
rect 26200 17212 26206 17224
rect 26338 17221 26350 17224
rect 26384 17221 26396 17255
rect 26338 17215 26396 17221
rect 26510 17212 26516 17264
rect 26568 17252 26574 17264
rect 30742 17252 30748 17264
rect 26568 17224 26648 17252
rect 26568 17212 26574 17224
rect 26620 17193 26648 17224
rect 28368 17224 30236 17252
rect 28368 17193 28396 17224
rect 24765 17187 24823 17193
rect 24765 17153 24777 17187
rect 24811 17153 24823 17187
rect 24765 17147 24823 17153
rect 26605 17188 26663 17193
rect 26605 17187 26924 17188
rect 26605 17153 26617 17187
rect 26651 17184 26924 17187
rect 28353 17187 28411 17193
rect 28353 17184 28365 17187
rect 26651 17160 28365 17184
rect 26651 17153 26663 17160
rect 26896 17156 28365 17160
rect 26605 17147 26663 17153
rect 28353 17153 28365 17156
rect 28399 17153 28411 17187
rect 28353 17147 28411 17153
rect 28442 17144 28448 17196
rect 28500 17184 28506 17196
rect 28609 17187 28667 17193
rect 28609 17184 28621 17187
rect 28500 17156 28621 17184
rect 28500 17144 28506 17156
rect 28609 17153 28621 17156
rect 28655 17153 28667 17187
rect 28609 17147 28667 17153
rect 28902 17144 28908 17196
rect 28960 17184 28966 17196
rect 30208 17193 30236 17224
rect 30300 17224 30748 17252
rect 30193 17187 30251 17193
rect 28960 17156 29776 17184
rect 28960 17144 28966 17156
rect 23768 17088 25360 17116
rect 22741 17079 22799 17085
rect 22646 17048 22652 17060
rect 20128 17020 21036 17048
rect 21376 17020 22652 17048
rect 20128 17008 20134 17020
rect 1670 16980 1676 16992
rect 1631 16952 1676 16980
rect 1670 16940 1676 16952
rect 1728 16940 1734 16992
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 17678 16980 17684 16992
rect 16724 16952 17684 16980
rect 16724 16940 16730 16952
rect 17678 16940 17684 16952
rect 17736 16980 17742 16992
rect 17773 16983 17831 16989
rect 17773 16980 17785 16983
rect 17736 16952 17785 16980
rect 17736 16940 17742 16952
rect 17773 16949 17785 16952
rect 17819 16980 17831 16983
rect 21376 16980 21404 17020
rect 22646 17008 22652 17020
rect 22704 17008 22710 17060
rect 23750 17008 23756 17060
rect 23808 17048 23814 17060
rect 24670 17048 24676 17060
rect 23808 17020 24676 17048
rect 23808 17008 23814 17020
rect 24670 17008 24676 17020
rect 24728 17008 24734 17060
rect 17819 16952 21404 16980
rect 21453 16983 21511 16989
rect 17819 16949 17831 16952
rect 17773 16943 17831 16949
rect 21453 16949 21465 16983
rect 21499 16980 21511 16983
rect 21818 16980 21824 16992
rect 21499 16952 21824 16980
rect 21499 16949 21511 16952
rect 21453 16943 21511 16949
rect 21818 16940 21824 16952
rect 21876 16940 21882 16992
rect 22281 16983 22339 16989
rect 22281 16949 22293 16983
rect 22327 16980 22339 16983
rect 24026 16980 24032 16992
rect 22327 16952 24032 16980
rect 22327 16949 22339 16952
rect 22281 16943 22339 16949
rect 24026 16940 24032 16952
rect 24084 16940 24090 16992
rect 24121 16983 24179 16989
rect 24121 16949 24133 16983
rect 24167 16980 24179 16983
rect 25222 16980 25228 16992
rect 24167 16952 25228 16980
rect 24167 16949 24179 16952
rect 24121 16943 24179 16949
rect 25222 16940 25228 16952
rect 25280 16940 25286 16992
rect 25332 16980 25360 17088
rect 27706 17076 27712 17128
rect 27764 17116 27770 17128
rect 27764 17088 27809 17116
rect 27764 17076 27770 17088
rect 26878 17008 26884 17060
rect 26936 17048 26942 17060
rect 29748 17057 29776 17156
rect 30193 17153 30205 17187
rect 30239 17153 30251 17187
rect 30193 17147 30251 17153
rect 29822 17076 29828 17128
rect 29880 17116 29886 17128
rect 30300 17116 30328 17224
rect 30742 17212 30748 17224
rect 30800 17212 30806 17264
rect 33226 17212 33232 17264
rect 33284 17252 33290 17264
rect 36078 17252 36084 17264
rect 33284 17224 36084 17252
rect 33284 17212 33290 17224
rect 30460 17187 30518 17193
rect 30460 17153 30472 17187
rect 30506 17184 30518 17187
rect 31018 17184 31024 17196
rect 30506 17156 31024 17184
rect 30506 17153 30518 17156
rect 30460 17147 30518 17153
rect 31018 17144 31024 17156
rect 31076 17144 31082 17196
rect 33704 17193 33732 17224
rect 35820 17193 35848 17224
rect 36078 17212 36084 17224
rect 36136 17212 36142 17264
rect 36188 17252 36216 17292
rect 36725 17289 36737 17323
rect 36771 17320 36783 17323
rect 36906 17320 36912 17332
rect 36771 17292 36912 17320
rect 36771 17289 36783 17292
rect 36725 17283 36783 17289
rect 36906 17280 36912 17292
rect 36964 17280 36970 17332
rect 37550 17320 37556 17332
rect 37463 17292 37556 17320
rect 37550 17280 37556 17292
rect 37608 17320 37614 17332
rect 38562 17320 38568 17332
rect 37608 17292 38568 17320
rect 37608 17280 37614 17292
rect 38562 17280 38568 17292
rect 38620 17280 38626 17332
rect 38841 17323 38899 17329
rect 38841 17289 38853 17323
rect 38887 17320 38899 17323
rect 38930 17320 38936 17332
rect 38887 17292 38936 17320
rect 38887 17289 38899 17292
rect 38841 17283 38899 17289
rect 38930 17280 38936 17292
rect 38988 17280 38994 17332
rect 41509 17323 41567 17329
rect 41509 17320 41521 17323
rect 40880 17292 41521 17320
rect 38654 17252 38660 17264
rect 36188 17224 38660 17252
rect 38654 17212 38660 17224
rect 38712 17212 38718 17264
rect 39022 17212 39028 17264
rect 39080 17252 39086 17264
rect 39758 17252 39764 17264
rect 39080 17224 39764 17252
rect 39080 17212 39086 17224
rect 39758 17212 39764 17224
rect 39816 17212 39822 17264
rect 39976 17255 40034 17261
rect 39976 17221 39988 17255
rect 40022 17252 40034 17255
rect 40880 17252 40908 17292
rect 41509 17289 41521 17292
rect 41555 17289 41567 17323
rect 54110 17320 54116 17332
rect 54071 17292 54116 17320
rect 41509 17283 41567 17289
rect 54110 17280 54116 17292
rect 54168 17280 54174 17332
rect 54202 17252 54208 17264
rect 40022 17224 40908 17252
rect 54163 17224 54208 17252
rect 40022 17221 40034 17224
rect 39976 17215 40034 17221
rect 54202 17212 54208 17224
rect 54260 17212 54266 17264
rect 33433 17187 33491 17193
rect 33433 17153 33445 17187
rect 33479 17184 33491 17187
rect 33689 17187 33747 17193
rect 33479 17156 33640 17184
rect 33479 17153 33491 17156
rect 33433 17147 33491 17153
rect 29880 17088 30328 17116
rect 33612 17116 33640 17156
rect 33689 17153 33701 17187
rect 33735 17153 33747 17187
rect 33689 17147 33747 17153
rect 35549 17187 35607 17193
rect 35549 17153 35561 17187
rect 35595 17184 35607 17187
rect 35805 17187 35863 17193
rect 35595 17156 35756 17184
rect 35595 17153 35607 17156
rect 35549 17147 35607 17153
rect 34698 17116 34704 17128
rect 33612 17088 34704 17116
rect 29880 17076 29886 17088
rect 34698 17076 34704 17088
rect 34756 17076 34762 17128
rect 35728 17116 35756 17156
rect 35805 17153 35817 17187
rect 35851 17153 35863 17187
rect 35805 17147 35863 17153
rect 35986 17144 35992 17196
rect 36044 17184 36050 17196
rect 36449 17187 36507 17193
rect 36449 17184 36461 17187
rect 36044 17156 36461 17184
rect 36044 17144 36050 17156
rect 36449 17153 36461 17156
rect 36495 17153 36507 17187
rect 36449 17147 36507 17153
rect 38197 17187 38255 17193
rect 38197 17153 38209 17187
rect 38243 17184 38255 17187
rect 39114 17184 39120 17196
rect 38243 17156 39120 17184
rect 38243 17153 38255 17156
rect 38197 17147 38255 17153
rect 39114 17144 39120 17156
rect 39172 17144 39178 17196
rect 40221 17187 40279 17193
rect 39224 17156 40172 17184
rect 39224 17128 39252 17156
rect 36814 17116 36820 17128
rect 35728 17088 36820 17116
rect 36814 17076 36820 17088
rect 36872 17076 36878 17128
rect 37274 17076 37280 17128
rect 37332 17116 37338 17128
rect 38013 17119 38071 17125
rect 38013 17116 38025 17119
rect 37332 17088 38025 17116
rect 37332 17076 37338 17088
rect 38013 17085 38025 17088
rect 38059 17116 38071 17119
rect 39206 17116 39212 17128
rect 38059 17088 39212 17116
rect 38059 17085 38071 17088
rect 38013 17079 38071 17085
rect 39206 17076 39212 17088
rect 39264 17076 39270 17128
rect 40144 17116 40172 17156
rect 40221 17153 40233 17187
rect 40267 17184 40279 17187
rect 40267 17156 40816 17184
rect 40267 17153 40279 17156
rect 40221 17147 40279 17153
rect 40310 17116 40316 17128
rect 40144 17088 40316 17116
rect 40310 17076 40316 17088
rect 40368 17116 40374 17128
rect 40681 17119 40739 17125
rect 40681 17116 40693 17119
rect 40368 17088 40693 17116
rect 40368 17076 40374 17088
rect 40681 17085 40693 17088
rect 40727 17085 40739 17119
rect 40788 17116 40816 17156
rect 40862 17144 40868 17196
rect 40920 17184 40926 17196
rect 41693 17187 41751 17193
rect 40920 17156 40965 17184
rect 40920 17144 40926 17156
rect 41693 17153 41705 17187
rect 41739 17184 41751 17187
rect 53469 17187 53527 17193
rect 41739 17156 41828 17184
rect 41739 17153 41751 17156
rect 41693 17147 41751 17153
rect 41414 17116 41420 17128
rect 40788 17088 41420 17116
rect 40681 17079 40739 17085
rect 41414 17076 41420 17088
rect 41472 17076 41478 17128
rect 29733 17051 29791 17057
rect 26936 17020 27844 17048
rect 26936 17008 26942 17020
rect 27706 16980 27712 16992
rect 25332 16952 27712 16980
rect 27706 16940 27712 16952
rect 27764 16940 27770 16992
rect 27816 16980 27844 17020
rect 29733 17017 29745 17051
rect 29779 17017 29791 17051
rect 34425 17051 34483 17057
rect 29733 17011 29791 17017
rect 31496 17020 32812 17048
rect 31496 16980 31524 17020
rect 27816 16952 31524 16980
rect 31573 16983 31631 16989
rect 31573 16949 31585 16983
rect 31619 16980 31631 16983
rect 32306 16980 32312 16992
rect 31619 16952 32312 16980
rect 31619 16949 31631 16952
rect 31573 16943 31631 16949
rect 32306 16940 32312 16952
rect 32364 16940 32370 16992
rect 32784 16980 32812 17020
rect 34425 17017 34437 17051
rect 34471 17048 34483 17051
rect 34514 17048 34520 17060
rect 34471 17020 34520 17048
rect 34471 17017 34483 17020
rect 34425 17011 34483 17017
rect 34514 17008 34520 17020
rect 34572 17008 34578 17060
rect 38381 17051 38439 17057
rect 38381 17017 38393 17051
rect 38427 17048 38439 17051
rect 41800 17048 41828 17156
rect 53469 17153 53481 17187
rect 53515 17184 53527 17187
rect 53558 17184 53564 17196
rect 53515 17156 53564 17184
rect 53515 17153 53527 17156
rect 53469 17147 53527 17153
rect 53558 17144 53564 17156
rect 53616 17144 53622 17196
rect 53282 17048 53288 17060
rect 38427 17020 39344 17048
rect 38427 17017 38439 17020
rect 38381 17011 38439 17017
rect 35158 16980 35164 16992
rect 32784 16952 35164 16980
rect 35158 16940 35164 16952
rect 35216 16940 35222 16992
rect 35894 16940 35900 16992
rect 35952 16980 35958 16992
rect 36906 16980 36912 16992
rect 35952 16952 36912 16980
rect 35952 16940 35958 16952
rect 36906 16940 36912 16952
rect 36964 16940 36970 16992
rect 39316 16980 39344 17020
rect 40236 17020 41828 17048
rect 53243 17020 53288 17048
rect 40236 16980 40264 17020
rect 53282 17008 53288 17020
rect 53340 17008 53346 17060
rect 39316 16952 40264 16980
rect 41049 16983 41107 16989
rect 41049 16949 41061 16983
rect 41095 16980 41107 16983
rect 42058 16980 42064 16992
rect 41095 16952 42064 16980
rect 41095 16949 41107 16952
rect 41049 16943 41107 16949
rect 42058 16940 42064 16952
rect 42116 16940 42122 16992
rect 42702 16980 42708 16992
rect 42663 16952 42708 16980
rect 42702 16940 42708 16952
rect 42760 16980 42766 16992
rect 43165 16983 43223 16989
rect 43165 16980 43177 16983
rect 42760 16952 43177 16980
rect 42760 16940 42766 16952
rect 43165 16949 43177 16952
rect 43211 16980 43223 16983
rect 43254 16980 43260 16992
rect 43211 16952 43260 16980
rect 43211 16949 43223 16952
rect 43165 16943 43223 16949
rect 43254 16940 43260 16952
rect 43312 16940 43318 16992
rect 43809 16983 43867 16989
rect 43809 16949 43821 16983
rect 43855 16980 43867 16983
rect 44174 16980 44180 16992
rect 43855 16952 44180 16980
rect 43855 16949 43867 16952
rect 43809 16943 43867 16949
rect 44174 16940 44180 16952
rect 44232 16980 44238 16992
rect 44361 16983 44419 16989
rect 44361 16980 44373 16983
rect 44232 16952 44373 16980
rect 44232 16940 44238 16952
rect 44361 16949 44373 16952
rect 44407 16980 44419 16983
rect 44450 16980 44456 16992
rect 44407 16952 44456 16980
rect 44407 16949 44419 16952
rect 44361 16943 44419 16949
rect 44450 16940 44456 16952
rect 44508 16940 44514 16992
rect 1104 16890 54832 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 54832 16890
rect 1104 16816 54832 16838
rect 15657 16779 15715 16785
rect 15657 16745 15669 16779
rect 15703 16776 15715 16779
rect 18230 16776 18236 16788
rect 15703 16748 18236 16776
rect 15703 16745 15715 16748
rect 15657 16739 15715 16745
rect 18230 16736 18236 16748
rect 18288 16736 18294 16788
rect 22186 16776 22192 16788
rect 22066 16748 22192 16776
rect 16114 16640 16120 16652
rect 16075 16612 16120 16640
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 16758 16640 16764 16652
rect 16719 16612 16764 16640
rect 16758 16600 16764 16612
rect 16816 16600 16822 16652
rect 16942 16600 16948 16652
rect 17000 16640 17006 16652
rect 17865 16643 17923 16649
rect 17865 16640 17877 16643
rect 17000 16612 17877 16640
rect 17000 16600 17006 16612
rect 17865 16609 17877 16612
rect 17911 16609 17923 16643
rect 17865 16603 17923 16609
rect 21269 16643 21327 16649
rect 21269 16609 21281 16643
rect 21315 16640 21327 16643
rect 22066 16640 22094 16748
rect 22186 16736 22192 16748
rect 22244 16736 22250 16788
rect 22370 16776 22376 16788
rect 22331 16748 22376 16776
rect 22370 16736 22376 16748
rect 22428 16736 22434 16788
rect 23017 16779 23075 16785
rect 23017 16745 23029 16779
rect 23063 16776 23075 16779
rect 23106 16776 23112 16788
rect 23063 16748 23112 16776
rect 23063 16745 23075 16748
rect 23017 16739 23075 16745
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 23201 16779 23259 16785
rect 23201 16745 23213 16779
rect 23247 16776 23259 16779
rect 23750 16776 23756 16788
rect 23247 16748 23756 16776
rect 23247 16745 23259 16748
rect 23201 16739 23259 16745
rect 23750 16736 23756 16748
rect 23808 16736 23814 16788
rect 24029 16779 24087 16785
rect 24029 16745 24041 16779
rect 24075 16776 24087 16779
rect 24118 16776 24124 16788
rect 24075 16748 24124 16776
rect 24075 16745 24087 16748
rect 24029 16739 24087 16745
rect 24118 16736 24124 16748
rect 24176 16736 24182 16788
rect 24578 16776 24584 16788
rect 24539 16748 24584 16776
rect 24578 16736 24584 16748
rect 24636 16736 24642 16788
rect 24670 16736 24676 16788
rect 24728 16776 24734 16788
rect 29546 16776 29552 16788
rect 24728 16748 29552 16776
rect 24728 16736 24734 16748
rect 29546 16736 29552 16748
rect 29604 16736 29610 16788
rect 30374 16736 30380 16788
rect 30432 16736 30438 16788
rect 31018 16776 31024 16788
rect 30979 16748 31024 16776
rect 31018 16736 31024 16748
rect 31076 16736 31082 16788
rect 33134 16776 33140 16788
rect 33095 16748 33140 16776
rect 33134 16736 33140 16748
rect 33192 16736 33198 16788
rect 34149 16779 34207 16785
rect 34149 16745 34161 16779
rect 34195 16745 34207 16779
rect 34149 16739 34207 16745
rect 35253 16779 35311 16785
rect 35253 16745 35265 16779
rect 35299 16776 35311 16779
rect 36446 16776 36452 16788
rect 35299 16748 36452 16776
rect 35299 16745 35311 16748
rect 35253 16739 35311 16745
rect 26421 16711 26479 16717
rect 26421 16708 26433 16711
rect 21315 16612 22094 16640
rect 22204 16680 26433 16708
rect 21315 16609 21327 16612
rect 21269 16603 21327 16609
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16572 1915 16575
rect 16574 16572 16580 16584
rect 1903 16544 16580 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 17218 16572 17224 16584
rect 17179 16544 17224 16572
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 18049 16575 18107 16581
rect 18049 16572 18061 16575
rect 17328 16544 18061 16572
rect 14826 16464 14832 16516
rect 14884 16504 14890 16516
rect 15105 16507 15163 16513
rect 15105 16504 15117 16507
rect 14884 16476 15117 16504
rect 14884 16464 14890 16476
rect 15105 16473 15117 16476
rect 15151 16504 15163 16507
rect 17328 16504 17356 16544
rect 18049 16541 18061 16544
rect 18095 16541 18107 16575
rect 18230 16572 18236 16584
rect 18191 16544 18236 16572
rect 18049 16535 18107 16541
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 18693 16575 18751 16581
rect 18693 16541 18705 16575
rect 18739 16572 18751 16575
rect 22094 16572 22100 16584
rect 18739 16544 22100 16572
rect 18739 16541 18751 16544
rect 18693 16535 18751 16541
rect 22094 16532 22100 16544
rect 22152 16532 22158 16584
rect 22204 16581 22232 16680
rect 26421 16677 26433 16680
rect 26467 16708 26479 16711
rect 26881 16711 26939 16717
rect 26881 16708 26893 16711
rect 26467 16680 26893 16708
rect 26467 16677 26479 16680
rect 26421 16671 26479 16677
rect 26881 16677 26893 16680
rect 26927 16677 26939 16711
rect 27430 16708 27436 16720
rect 27391 16680 27436 16708
rect 26881 16671 26939 16677
rect 27430 16668 27436 16680
rect 27488 16708 27494 16720
rect 29086 16708 29092 16720
rect 27488 16680 29092 16708
rect 27488 16668 27494 16680
rect 29086 16668 29092 16680
rect 29144 16668 29150 16720
rect 30392 16708 30420 16736
rect 31570 16708 31576 16720
rect 30392 16680 31576 16708
rect 31570 16668 31576 16680
rect 31628 16708 31634 16720
rect 31628 16680 32260 16708
rect 31628 16668 31634 16680
rect 23661 16643 23719 16649
rect 23661 16609 23673 16643
rect 23707 16640 23719 16643
rect 25038 16640 25044 16652
rect 23707 16612 24869 16640
rect 24999 16612 25044 16640
rect 23707 16609 23719 16612
rect 23661 16603 23719 16609
rect 22189 16575 22247 16581
rect 22189 16541 22201 16575
rect 22235 16541 22247 16575
rect 22189 16535 22247 16541
rect 22373 16575 22431 16581
rect 22373 16541 22385 16575
rect 22419 16572 22431 16575
rect 23750 16572 23756 16584
rect 22419 16544 23756 16572
rect 22419 16541 22431 16544
rect 22373 16535 22431 16541
rect 23750 16532 23756 16544
rect 23808 16532 23814 16584
rect 23845 16575 23903 16581
rect 23845 16541 23857 16575
rect 23891 16572 23903 16575
rect 24210 16572 24216 16584
rect 23891 16544 24216 16572
rect 23891 16541 23903 16544
rect 23845 16535 23903 16541
rect 24210 16532 24216 16544
rect 24268 16532 24274 16584
rect 24841 16572 24869 16612
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 25130 16600 25136 16652
rect 25188 16640 25194 16652
rect 28353 16643 28411 16649
rect 25188 16612 25233 16640
rect 25188 16600 25194 16612
rect 28353 16609 28365 16643
rect 28399 16609 28411 16643
rect 28353 16606 28411 16609
rect 28296 16603 28411 16606
rect 28445 16643 28503 16649
rect 28445 16609 28457 16643
rect 28491 16640 28503 16643
rect 29454 16640 29460 16652
rect 28491 16612 29460 16640
rect 28491 16609 28503 16612
rect 28445 16603 28503 16609
rect 24949 16575 25007 16581
rect 24949 16572 24961 16575
rect 24841 16544 24961 16572
rect 24949 16541 24961 16544
rect 24995 16572 25007 16575
rect 25222 16572 25228 16584
rect 24995 16544 25228 16572
rect 24995 16541 25007 16544
rect 24949 16535 25007 16541
rect 25222 16532 25228 16544
rect 25280 16572 25286 16584
rect 25777 16575 25835 16581
rect 25777 16572 25789 16575
rect 25280 16544 25789 16572
rect 25280 16532 25286 16544
rect 25777 16541 25789 16544
rect 25823 16541 25835 16575
rect 25777 16535 25835 16541
rect 26234 16532 26240 16584
rect 26292 16572 26298 16584
rect 27062 16572 27068 16584
rect 26292 16544 27068 16572
rect 26292 16532 26298 16544
rect 27062 16532 27068 16544
rect 27120 16572 27126 16584
rect 27157 16575 27215 16581
rect 27157 16572 27169 16575
rect 27120 16544 27169 16572
rect 27120 16532 27126 16544
rect 27157 16541 27169 16544
rect 27203 16541 27215 16575
rect 27157 16535 27215 16541
rect 27798 16532 27804 16584
rect 27856 16572 27862 16584
rect 28296 16578 28396 16603
rect 29454 16600 29460 16612
rect 29512 16600 29518 16652
rect 30282 16600 30288 16652
rect 30340 16640 30346 16652
rect 30377 16643 30435 16649
rect 30377 16640 30389 16643
rect 30340 16612 30389 16640
rect 30340 16600 30346 16612
rect 30377 16609 30389 16612
rect 30423 16609 30435 16643
rect 30377 16603 30435 16609
rect 28296 16572 28324 16578
rect 27856 16544 28324 16572
rect 28537 16575 28595 16581
rect 27856 16532 27862 16544
rect 28537 16541 28549 16575
rect 28583 16541 28595 16575
rect 28537 16535 28595 16541
rect 17954 16504 17960 16516
rect 15151 16476 17356 16504
rect 17420 16476 17960 16504
rect 15151 16473 15163 16476
rect 15105 16467 15163 16473
rect 1670 16436 1676 16448
rect 1631 16408 1676 16436
rect 1670 16396 1676 16408
rect 1728 16396 1734 16448
rect 17420 16445 17448 16476
rect 17954 16464 17960 16476
rect 18012 16464 18018 16516
rect 21024 16507 21082 16513
rect 18892 16476 20484 16504
rect 18892 16445 18920 16476
rect 17405 16439 17463 16445
rect 17405 16405 17417 16439
rect 17451 16405 17463 16439
rect 17405 16399 17463 16405
rect 18877 16439 18935 16445
rect 18877 16405 18889 16439
rect 18923 16405 18935 16439
rect 18877 16399 18935 16405
rect 19889 16439 19947 16445
rect 19889 16405 19901 16439
rect 19935 16436 19947 16439
rect 20070 16436 20076 16448
rect 19935 16408 20076 16436
rect 19935 16405 19947 16408
rect 19889 16399 19947 16405
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20456 16436 20484 16476
rect 21024 16473 21036 16507
rect 21070 16504 21082 16507
rect 21634 16504 21640 16516
rect 21070 16476 21640 16504
rect 21070 16473 21082 16476
rect 21024 16467 21082 16473
rect 21634 16464 21640 16476
rect 21692 16464 21698 16516
rect 22646 16464 22652 16516
rect 22704 16504 22710 16516
rect 22833 16507 22891 16513
rect 22833 16504 22845 16507
rect 22704 16476 22845 16504
rect 22704 16464 22710 16476
rect 22833 16473 22845 16476
rect 22879 16473 22891 16507
rect 22833 16467 22891 16473
rect 23049 16507 23107 16513
rect 23049 16473 23061 16507
rect 23095 16504 23107 16507
rect 24578 16504 24584 16516
rect 23095 16476 24584 16504
rect 23095 16473 23107 16476
rect 23049 16467 23107 16473
rect 22186 16436 22192 16448
rect 20456 16408 22192 16436
rect 22186 16396 22192 16408
rect 22244 16396 22250 16448
rect 22848 16436 22876 16467
rect 24578 16464 24584 16476
rect 24636 16504 24642 16516
rect 27249 16507 27307 16513
rect 27249 16504 27261 16507
rect 24636 16476 27261 16504
rect 24636 16464 24642 16476
rect 27249 16473 27261 16476
rect 27295 16473 27307 16507
rect 27249 16467 27307 16473
rect 27522 16464 27528 16516
rect 27580 16504 27586 16516
rect 27816 16504 27844 16532
rect 28350 16504 28356 16516
rect 27580 16476 27844 16504
rect 28092 16476 28356 16504
rect 27580 16464 27586 16476
rect 27065 16439 27123 16445
rect 27065 16436 27077 16439
rect 22848 16408 27077 16436
rect 27065 16405 27077 16408
rect 27111 16436 27123 16439
rect 27430 16436 27436 16448
rect 27111 16408 27436 16436
rect 27111 16405 27123 16408
rect 27065 16399 27123 16405
rect 27430 16396 27436 16408
rect 27488 16396 27494 16448
rect 27614 16396 27620 16448
rect 27672 16436 27678 16448
rect 28092 16436 28120 16476
rect 28350 16464 28356 16476
rect 28408 16504 28414 16516
rect 28552 16504 28580 16535
rect 28626 16532 28632 16584
rect 28684 16572 28690 16584
rect 28684 16544 28729 16572
rect 28684 16532 28690 16544
rect 29638 16532 29644 16584
rect 29696 16572 29702 16584
rect 29733 16575 29791 16581
rect 29733 16572 29745 16575
rect 29696 16544 29745 16572
rect 29696 16532 29702 16544
rect 29733 16541 29745 16544
rect 29779 16541 29791 16575
rect 32232 16572 32260 16680
rect 32950 16668 32956 16720
rect 33008 16708 33014 16720
rect 34164 16708 34192 16739
rect 36446 16736 36452 16748
rect 36504 16736 36510 16788
rect 37458 16776 37464 16788
rect 36556 16748 37464 16776
rect 35342 16708 35348 16720
rect 33008 16680 35348 16708
rect 33008 16668 33014 16680
rect 35342 16668 35348 16680
rect 35400 16668 35406 16720
rect 36173 16711 36231 16717
rect 36173 16677 36185 16711
rect 36219 16708 36231 16711
rect 36556 16708 36584 16748
rect 37458 16736 37464 16748
rect 37516 16736 37522 16788
rect 37645 16779 37703 16785
rect 37645 16745 37657 16779
rect 37691 16776 37703 16779
rect 38010 16776 38016 16788
rect 37691 16748 38016 16776
rect 37691 16745 37703 16748
rect 37645 16739 37703 16745
rect 38010 16736 38016 16748
rect 38068 16736 38074 16788
rect 38197 16779 38255 16785
rect 38197 16745 38209 16779
rect 38243 16776 38255 16779
rect 38286 16776 38292 16788
rect 38243 16748 38292 16776
rect 38243 16745 38255 16748
rect 38197 16739 38255 16745
rect 38286 16736 38292 16748
rect 38344 16736 38350 16788
rect 39390 16776 39396 16788
rect 39351 16748 39396 16776
rect 39390 16736 39396 16748
rect 39448 16736 39454 16788
rect 41230 16776 41236 16788
rect 39500 16748 41236 16776
rect 39500 16708 39528 16748
rect 41230 16736 41236 16748
rect 41288 16736 41294 16788
rect 41506 16736 41512 16788
rect 41564 16776 41570 16788
rect 44269 16779 44327 16785
rect 44269 16776 44281 16779
rect 41564 16748 44281 16776
rect 41564 16736 41570 16748
rect 44269 16745 44281 16748
rect 44315 16776 44327 16779
rect 53466 16776 53472 16788
rect 44315 16748 53472 16776
rect 44315 16745 44327 16748
rect 44269 16739 44327 16745
rect 53466 16736 53472 16748
rect 53524 16736 53530 16788
rect 54202 16776 54208 16788
rect 54163 16748 54208 16776
rect 54202 16736 54208 16748
rect 54260 16736 54266 16788
rect 41874 16708 41880 16720
rect 36219 16680 36584 16708
rect 36832 16680 39528 16708
rect 41835 16680 41880 16708
rect 36219 16677 36231 16680
rect 36173 16671 36231 16677
rect 32306 16600 32312 16652
rect 32364 16640 32370 16652
rect 32493 16643 32551 16649
rect 32493 16640 32505 16643
rect 32364 16612 32505 16640
rect 32364 16600 32370 16612
rect 32493 16609 32505 16612
rect 32539 16640 32551 16643
rect 33042 16640 33048 16652
rect 32539 16612 33048 16640
rect 32539 16609 32551 16612
rect 32493 16603 32551 16609
rect 33042 16600 33048 16612
rect 33100 16600 33106 16652
rect 33410 16640 33416 16652
rect 33152 16612 33416 16640
rect 33152 16572 33180 16612
rect 33410 16600 33416 16612
rect 33468 16600 33474 16652
rect 33502 16600 33508 16652
rect 33560 16600 33566 16652
rect 34882 16640 34888 16652
rect 34843 16612 34888 16640
rect 34882 16600 34888 16612
rect 34940 16600 34946 16652
rect 35158 16600 35164 16652
rect 35216 16640 35222 16652
rect 35894 16640 35900 16652
rect 35216 16612 35900 16640
rect 35216 16600 35222 16612
rect 35894 16600 35900 16612
rect 35952 16600 35958 16652
rect 36630 16600 36636 16652
rect 36688 16640 36694 16652
rect 36832 16649 36860 16680
rect 41874 16668 41880 16680
rect 41932 16668 41938 16720
rect 42886 16668 42892 16720
rect 42944 16708 42950 16720
rect 43073 16711 43131 16717
rect 43073 16708 43085 16711
rect 42944 16680 43085 16708
rect 42944 16668 42950 16680
rect 43073 16677 43085 16680
rect 43119 16677 43131 16711
rect 53558 16708 53564 16720
rect 53519 16680 53564 16708
rect 43073 16671 43131 16677
rect 53558 16668 53564 16680
rect 53616 16668 53622 16720
rect 36817 16643 36875 16649
rect 36817 16640 36829 16643
rect 36688 16612 36829 16640
rect 36688 16600 36694 16612
rect 36817 16609 36829 16612
rect 36863 16609 36875 16643
rect 36817 16603 36875 16609
rect 37826 16600 37832 16652
rect 37884 16640 37890 16652
rect 40402 16640 40408 16652
rect 37884 16612 40408 16640
rect 37884 16600 37890 16612
rect 40402 16600 40408 16612
rect 40460 16600 40466 16652
rect 41414 16640 41420 16652
rect 41375 16612 41420 16640
rect 41414 16600 41420 16612
rect 41472 16600 41478 16652
rect 43622 16640 43628 16652
rect 43583 16612 43628 16640
rect 43622 16600 43628 16612
rect 43680 16600 43686 16652
rect 32232 16544 33180 16572
rect 29733 16535 29791 16541
rect 33413 16507 33471 16513
rect 28408 16476 28580 16504
rect 28966 16476 33364 16504
rect 28408 16464 28414 16476
rect 27672 16408 28120 16436
rect 28169 16439 28227 16445
rect 27672 16396 27678 16408
rect 28169 16405 28181 16439
rect 28215 16436 28227 16439
rect 28966 16436 28994 16476
rect 29914 16436 29920 16448
rect 28215 16408 28994 16436
rect 29875 16408 29920 16436
rect 28215 16405 28227 16408
rect 28169 16399 28227 16405
rect 29914 16396 29920 16408
rect 29972 16396 29978 16448
rect 30006 16396 30012 16448
rect 30064 16436 30070 16448
rect 31849 16439 31907 16445
rect 31849 16436 31861 16439
rect 30064 16408 31861 16436
rect 30064 16396 30070 16408
rect 31849 16405 31861 16408
rect 31895 16405 31907 16439
rect 33336 16436 33364 16476
rect 33413 16473 33425 16507
rect 33459 16504 33471 16507
rect 33520 16504 33548 16600
rect 33594 16532 33600 16584
rect 33652 16572 33658 16584
rect 33965 16575 34023 16581
rect 33965 16572 33977 16575
rect 33652 16544 33977 16572
rect 33652 16532 33658 16544
rect 33965 16541 33977 16544
rect 34011 16541 34023 16575
rect 33965 16535 34023 16541
rect 34790 16532 34796 16584
rect 34848 16572 34854 16584
rect 35069 16575 35127 16581
rect 35069 16572 35081 16575
rect 34848 16544 35081 16572
rect 34848 16532 34854 16544
rect 35069 16541 35081 16544
rect 35115 16541 35127 16575
rect 36354 16572 36360 16584
rect 36315 16544 36360 16572
rect 35069 16535 35127 16541
rect 36354 16532 36360 16544
rect 36412 16532 36418 16584
rect 37274 16572 37280 16584
rect 37235 16544 37280 16572
rect 37274 16532 37280 16544
rect 37332 16532 37338 16584
rect 37458 16572 37464 16584
rect 37419 16544 37464 16572
rect 37458 16532 37464 16544
rect 37516 16532 37522 16584
rect 38654 16532 38660 16584
rect 38712 16572 38718 16584
rect 38841 16575 38899 16581
rect 38841 16572 38853 16575
rect 38712 16544 38853 16572
rect 38712 16532 38718 16544
rect 38841 16541 38853 16544
rect 38887 16541 38899 16575
rect 38841 16535 38899 16541
rect 39209 16575 39267 16581
rect 39209 16541 39221 16575
rect 39255 16572 39267 16575
rect 39298 16572 39304 16584
rect 39255 16544 39304 16572
rect 39255 16541 39267 16544
rect 39209 16535 39267 16541
rect 39298 16532 39304 16544
rect 39356 16532 39362 16584
rect 41161 16575 41219 16581
rect 41161 16541 41173 16575
rect 41207 16572 41219 16575
rect 41874 16572 41880 16584
rect 41207 16568 41399 16572
rect 41524 16568 41880 16572
rect 41207 16544 41880 16568
rect 41207 16541 41219 16544
rect 41161 16535 41219 16541
rect 41371 16540 41552 16544
rect 41874 16532 41880 16544
rect 41932 16532 41938 16584
rect 42058 16572 42064 16584
rect 42019 16544 42064 16572
rect 42058 16532 42064 16544
rect 42116 16532 42122 16584
rect 42518 16572 42524 16584
rect 42479 16544 42524 16572
rect 42518 16532 42524 16544
rect 42576 16532 42582 16584
rect 54021 16575 54079 16581
rect 54021 16541 54033 16575
rect 54067 16541 54079 16575
rect 54021 16535 54079 16541
rect 33459 16476 33548 16504
rect 33459 16473 33471 16476
rect 33413 16467 33471 16473
rect 33686 16464 33692 16516
rect 33744 16504 33750 16516
rect 36449 16507 36507 16513
rect 36449 16504 36461 16507
rect 33744 16476 36461 16504
rect 33744 16464 33750 16476
rect 36449 16473 36461 16476
rect 36495 16473 36507 16507
rect 36449 16467 36507 16473
rect 36538 16464 36544 16516
rect 36596 16504 36602 16516
rect 36679 16507 36737 16513
rect 36596 16476 36641 16504
rect 36596 16464 36602 16476
rect 36679 16473 36691 16507
rect 36725 16504 36737 16507
rect 37366 16504 37372 16516
rect 36725 16476 37372 16504
rect 36725 16473 36737 16476
rect 36679 16467 36737 16473
rect 37366 16464 37372 16476
rect 37424 16464 37430 16516
rect 37642 16464 37648 16516
rect 37700 16504 37706 16516
rect 38102 16504 38108 16516
rect 37700 16476 38108 16504
rect 37700 16464 37706 16476
rect 38102 16464 38108 16476
rect 38160 16504 38166 16516
rect 38289 16507 38347 16513
rect 38289 16504 38301 16507
rect 38160 16476 38301 16504
rect 38160 16464 38166 16476
rect 38289 16473 38301 16476
rect 38335 16473 38347 16507
rect 39022 16504 39028 16516
rect 38983 16476 39028 16504
rect 38289 16467 38347 16473
rect 39022 16464 39028 16476
rect 39080 16464 39086 16516
rect 39117 16507 39175 16513
rect 39117 16473 39129 16507
rect 39163 16504 39175 16507
rect 39163 16476 48314 16504
rect 39163 16473 39175 16476
rect 39117 16467 39175 16473
rect 38746 16436 38752 16448
rect 33336 16408 38752 16436
rect 31849 16399 31907 16405
rect 38746 16396 38752 16408
rect 38804 16396 38810 16448
rect 40052 16445 40080 16476
rect 40037 16439 40095 16445
rect 40037 16405 40049 16439
rect 40083 16405 40095 16439
rect 48286 16436 48314 16476
rect 54036 16436 54064 16535
rect 48286 16408 54064 16436
rect 40037 16399 40095 16405
rect 1104 16346 54832 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 54832 16346
rect 1104 16272 54832 16294
rect 14550 16232 14556 16244
rect 14511 16204 14556 16232
rect 14550 16192 14556 16204
rect 14608 16192 14614 16244
rect 15378 16192 15384 16244
rect 15436 16232 15442 16244
rect 16853 16235 16911 16241
rect 16853 16232 16865 16235
rect 15436 16204 16865 16232
rect 15436 16192 15442 16204
rect 16853 16201 16865 16204
rect 16899 16201 16911 16235
rect 16853 16195 16911 16201
rect 17310 16192 17316 16244
rect 17368 16232 17374 16244
rect 20533 16235 20591 16241
rect 20533 16232 20545 16235
rect 17368 16204 20545 16232
rect 17368 16192 17374 16204
rect 20533 16201 20545 16204
rect 20579 16201 20591 16235
rect 20533 16195 20591 16201
rect 20622 16192 20628 16244
rect 20680 16232 20686 16244
rect 20993 16235 21051 16241
rect 20993 16232 21005 16235
rect 20680 16204 21005 16232
rect 20680 16192 20686 16204
rect 20993 16201 21005 16204
rect 21039 16201 21051 16235
rect 20993 16195 21051 16201
rect 22094 16192 22100 16244
rect 22152 16232 22158 16244
rect 22557 16235 22615 16241
rect 22557 16232 22569 16235
rect 22152 16204 22569 16232
rect 22152 16192 22158 16204
rect 22557 16201 22569 16204
rect 22603 16201 22615 16235
rect 22557 16195 22615 16201
rect 24394 16192 24400 16244
rect 24452 16232 24458 16244
rect 25593 16235 25651 16241
rect 25593 16232 25605 16235
rect 24452 16204 25605 16232
rect 24452 16192 24458 16204
rect 25593 16201 25605 16204
rect 25639 16201 25651 16235
rect 28166 16232 28172 16244
rect 28127 16204 28172 16232
rect 25593 16195 25651 16201
rect 28166 16192 28172 16204
rect 28224 16192 28230 16244
rect 28534 16192 28540 16244
rect 28592 16232 28598 16244
rect 30282 16232 30288 16244
rect 28592 16204 29316 16232
rect 30243 16204 30288 16232
rect 28592 16192 28598 16204
rect 15102 16164 15108 16176
rect 6886 16136 12434 16164
rect 15063 16136 15108 16164
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 6886 16096 6914 16136
rect 1903 16068 6914 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 12406 16028 12434 16136
rect 15102 16124 15108 16136
rect 15160 16124 15166 16176
rect 17494 16164 17500 16176
rect 17328 16136 17500 16164
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16850 16096 16856 16108
rect 16163 16068 16856 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 16850 16056 16856 16068
rect 16908 16056 16914 16108
rect 17328 16105 17356 16136
rect 17494 16124 17500 16136
rect 17552 16124 17558 16176
rect 18233 16167 18291 16173
rect 18233 16133 18245 16167
rect 18279 16164 18291 16167
rect 18322 16164 18328 16176
rect 18279 16136 18328 16164
rect 18279 16133 18291 16136
rect 18233 16127 18291 16133
rect 18322 16124 18328 16136
rect 18380 16124 18386 16176
rect 22830 16164 22836 16176
rect 22066 16136 22836 16164
rect 17313 16099 17371 16105
rect 17313 16065 17325 16099
rect 17359 16065 17371 16099
rect 17313 16059 17371 16065
rect 17402 16056 17408 16108
rect 17460 16096 17466 16108
rect 18414 16096 18420 16108
rect 17460 16068 18420 16096
rect 17460 16056 17466 16068
rect 18414 16056 18420 16068
rect 18472 16096 18478 16108
rect 20622 16096 20628 16108
rect 18472 16068 20628 16096
rect 18472 16056 18478 16068
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 20898 16096 20904 16108
rect 20859 16068 20904 16096
rect 20898 16056 20904 16068
rect 20956 16096 20962 16108
rect 22066 16096 22094 16136
rect 22830 16124 22836 16136
rect 22888 16124 22894 16176
rect 23474 16164 23480 16176
rect 23435 16136 23480 16164
rect 23474 16124 23480 16136
rect 23532 16124 23538 16176
rect 25133 16167 25191 16173
rect 25133 16133 25145 16167
rect 25179 16164 25191 16167
rect 25866 16164 25872 16176
rect 25179 16136 25872 16164
rect 25179 16133 25191 16136
rect 25133 16127 25191 16133
rect 25866 16124 25872 16136
rect 25924 16164 25930 16176
rect 28994 16164 29000 16176
rect 25924 16136 29000 16164
rect 25924 16124 25930 16136
rect 28994 16124 29000 16136
rect 29052 16124 29058 16176
rect 22738 16096 22744 16108
rect 20956 16068 22094 16096
rect 22699 16068 22744 16096
rect 20956 16056 20962 16068
rect 22738 16056 22744 16068
rect 22796 16056 22802 16108
rect 27154 16096 27160 16108
rect 27115 16068 27160 16096
rect 27154 16056 27160 16068
rect 27212 16056 27218 16108
rect 27338 16096 27344 16108
rect 27299 16068 27344 16096
rect 27338 16056 27344 16068
rect 27396 16056 27402 16108
rect 27433 16099 27491 16105
rect 27433 16065 27445 16099
rect 27479 16065 27491 16099
rect 27433 16059 27491 16065
rect 27525 16099 27583 16105
rect 27525 16065 27537 16099
rect 27571 16065 27583 16099
rect 27525 16059 27583 16065
rect 28629 16099 28687 16105
rect 28629 16065 28641 16099
rect 28675 16096 28687 16099
rect 28810 16096 28816 16108
rect 28675 16068 28816 16096
rect 28675 16065 28687 16068
rect 28629 16059 28687 16065
rect 16758 16028 16764 16040
rect 12406 16000 16764 16028
rect 16758 15988 16764 16000
rect 16816 15988 16822 16040
rect 16942 15988 16948 16040
rect 17000 16028 17006 16040
rect 17037 16031 17095 16037
rect 17037 16028 17049 16031
rect 17000 16000 17049 16028
rect 17000 15988 17006 16000
rect 17037 15997 17049 16000
rect 17083 15997 17095 16031
rect 17037 15991 17095 15997
rect 17129 16031 17187 16037
rect 17129 15997 17141 16031
rect 17175 15997 17187 16031
rect 17129 15991 17187 15997
rect 17144 15960 17172 15991
rect 17218 15988 17224 16040
rect 17276 16028 17282 16040
rect 17276 16000 17321 16028
rect 17276 15988 17282 16000
rect 17586 15988 17592 16040
rect 17644 16028 17650 16040
rect 19978 16028 19984 16040
rect 17644 16000 19984 16028
rect 17644 15988 17650 16000
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 21082 15988 21088 16040
rect 21140 16028 21146 16040
rect 21177 16031 21235 16037
rect 21177 16028 21189 16031
rect 21140 16000 21189 16028
rect 21140 15988 21146 16000
rect 21177 15997 21189 16000
rect 21223 16028 21235 16031
rect 22002 16028 22008 16040
rect 21223 16000 22008 16028
rect 21223 15997 21235 16000
rect 21177 15991 21235 15997
rect 22002 15988 22008 16000
rect 22060 15988 22066 16040
rect 22925 16031 22983 16037
rect 22925 15997 22937 16031
rect 22971 16028 22983 16031
rect 23382 16028 23388 16040
rect 22971 16000 23388 16028
rect 22971 15997 22983 16000
rect 22925 15991 22983 15997
rect 20530 15960 20536 15972
rect 17144 15932 20536 15960
rect 20530 15920 20536 15932
rect 20588 15920 20594 15972
rect 20622 15920 20628 15972
rect 20680 15960 20686 15972
rect 22830 15960 22836 15972
rect 20680 15932 22836 15960
rect 20680 15920 20686 15932
rect 22830 15920 22836 15932
rect 22888 15960 22894 15972
rect 22940 15960 22968 15991
rect 23382 15988 23388 16000
rect 23440 15988 23446 16040
rect 26234 16028 26240 16040
rect 26195 16000 26240 16028
rect 26234 15988 26240 16000
rect 26292 15988 26298 16040
rect 26326 15988 26332 16040
rect 26384 16028 26390 16040
rect 27448 16028 27476 16059
rect 26384 16000 27476 16028
rect 26384 15988 26390 16000
rect 22888 15932 22968 15960
rect 22888 15920 22894 15932
rect 25498 15920 25504 15972
rect 25556 15960 25562 15972
rect 27338 15960 27344 15972
rect 25556 15932 27344 15960
rect 25556 15920 25562 15932
rect 27338 15920 27344 15932
rect 27396 15920 27402 15972
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 14274 15852 14280 15904
rect 14332 15892 14338 15904
rect 15562 15892 15568 15904
rect 14332 15864 15568 15892
rect 14332 15852 14338 15864
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 16301 15895 16359 15901
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 17862 15892 17868 15904
rect 16347 15864 17868 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 20806 15892 20812 15904
rect 18012 15864 20812 15892
rect 18012 15852 18018 15864
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 22097 15895 22155 15901
rect 22097 15861 22109 15895
rect 22143 15892 22155 15895
rect 24118 15892 24124 15904
rect 22143 15864 24124 15892
rect 22143 15861 22155 15864
rect 22097 15855 22155 15861
rect 24118 15852 24124 15864
rect 24176 15852 24182 15904
rect 24210 15852 24216 15904
rect 24268 15892 24274 15904
rect 27540 15892 27568 16059
rect 28810 16056 28816 16068
rect 28868 16056 28874 16108
rect 29086 16056 29092 16108
rect 29144 16096 29150 16108
rect 29288 16105 29316 16204
rect 30282 16192 30288 16204
rect 30340 16192 30346 16244
rect 33321 16235 33379 16241
rect 33321 16201 33333 16235
rect 33367 16232 33379 16235
rect 36354 16232 36360 16244
rect 33367 16204 36360 16232
rect 33367 16201 33379 16204
rect 33321 16195 33379 16201
rect 36354 16192 36360 16204
rect 36412 16192 36418 16244
rect 37274 16192 37280 16244
rect 37332 16232 37338 16244
rect 41506 16232 41512 16244
rect 37332 16204 41512 16232
rect 37332 16192 37338 16204
rect 41506 16192 41512 16204
rect 41564 16192 41570 16244
rect 41598 16192 41604 16244
rect 41656 16232 41662 16244
rect 41969 16235 42027 16241
rect 41969 16232 41981 16235
rect 41656 16204 41981 16232
rect 41656 16192 41662 16204
rect 41969 16201 41981 16204
rect 42015 16201 42027 16235
rect 41969 16195 42027 16201
rect 42886 16192 42892 16244
rect 42944 16232 42950 16244
rect 44821 16235 44879 16241
rect 44821 16232 44833 16235
rect 42944 16204 44833 16232
rect 42944 16192 42950 16204
rect 44821 16201 44833 16204
rect 44867 16201 44879 16235
rect 54202 16232 54208 16244
rect 54163 16204 54208 16232
rect 44821 16195 44879 16201
rect 54202 16192 54208 16204
rect 54260 16192 54266 16244
rect 34241 16167 34299 16173
rect 34241 16133 34253 16167
rect 34287 16164 34299 16167
rect 35158 16164 35164 16176
rect 34287 16136 34369 16164
rect 35119 16136 35164 16164
rect 34287 16133 34299 16136
rect 34241 16127 34299 16133
rect 29273 16099 29331 16105
rect 29144 16068 29189 16096
rect 29144 16056 29150 16068
rect 29273 16065 29285 16099
rect 29319 16065 29331 16099
rect 29273 16059 29331 16065
rect 29917 16099 29975 16105
rect 29917 16065 29929 16099
rect 29963 16096 29975 16099
rect 30006 16096 30012 16108
rect 29963 16068 30012 16096
rect 29963 16065 29975 16068
rect 29917 16059 29975 16065
rect 30006 16056 30012 16068
rect 30064 16056 30070 16108
rect 31110 16096 31116 16108
rect 31071 16068 31116 16096
rect 31110 16056 31116 16068
rect 31168 16056 31174 16108
rect 31205 16099 31263 16105
rect 31205 16065 31217 16099
rect 31251 16096 31263 16099
rect 31846 16096 31852 16108
rect 31251 16068 31852 16096
rect 31251 16065 31263 16068
rect 31205 16059 31263 16065
rect 31846 16056 31852 16068
rect 31904 16056 31910 16108
rect 32306 16096 32312 16108
rect 32267 16068 32312 16096
rect 32306 16056 32312 16068
rect 32364 16056 32370 16108
rect 32490 16096 32496 16108
rect 32451 16068 32496 16096
rect 32490 16056 32496 16068
rect 32548 16056 32554 16108
rect 32950 16096 32956 16108
rect 32911 16068 32956 16096
rect 32950 16056 32956 16068
rect 33008 16056 33014 16108
rect 33042 16056 33048 16108
rect 33100 16096 33106 16108
rect 33137 16099 33195 16105
rect 33137 16096 33149 16099
rect 33100 16068 33149 16096
rect 33100 16056 33106 16068
rect 33137 16065 33149 16068
rect 33183 16065 33195 16099
rect 33137 16059 33195 16065
rect 29181 16031 29239 16037
rect 27724 16000 28580 16028
rect 27724 15969 27752 16000
rect 27709 15963 27767 15969
rect 27709 15929 27721 15963
rect 27755 15929 27767 15963
rect 28258 15960 28264 15972
rect 28219 15932 28264 15960
rect 27709 15923 27767 15929
rect 28258 15920 28264 15932
rect 28316 15920 28322 15972
rect 28442 15892 28448 15904
rect 24268 15864 28448 15892
rect 24268 15852 24274 15864
rect 28442 15852 28448 15864
rect 28500 15852 28506 15904
rect 28552 15892 28580 16000
rect 29181 15997 29193 16031
rect 29227 16028 29239 16031
rect 29825 16031 29883 16037
rect 29825 16028 29837 16031
rect 29227 16000 29837 16028
rect 29227 15997 29239 16000
rect 29181 15991 29239 15997
rect 29825 15997 29837 16000
rect 29871 15997 29883 16031
rect 29825 15991 29883 15997
rect 31389 16031 31447 16037
rect 31389 15997 31401 16031
rect 31435 16028 31447 16031
rect 32030 16028 32036 16040
rect 31435 16000 32036 16028
rect 31435 15997 31447 16000
rect 31389 15991 31447 15997
rect 32030 15988 32036 16000
rect 32088 15988 32094 16040
rect 32401 16031 32459 16037
rect 32401 16028 32413 16031
rect 32140 16000 32413 16028
rect 28810 15920 28816 15972
rect 28868 15960 28874 15972
rect 32140 15960 32168 16000
rect 32401 15997 32413 16000
rect 32447 15997 32459 16031
rect 32401 15991 32459 15997
rect 28868 15932 32168 15960
rect 28868 15920 28874 15932
rect 33134 15892 33140 15904
rect 28552 15864 33140 15892
rect 33134 15852 33140 15864
rect 33192 15852 33198 15904
rect 33318 15852 33324 15904
rect 33376 15892 33382 15904
rect 33965 15895 34023 15901
rect 33965 15892 33977 15895
rect 33376 15864 33977 15892
rect 33376 15852 33382 15864
rect 33965 15861 33977 15864
rect 34011 15861 34023 15895
rect 34341 15892 34369 16136
rect 35158 16124 35164 16136
rect 35216 16164 35222 16176
rect 36446 16164 36452 16176
rect 35216 16136 36452 16164
rect 35216 16124 35222 16136
rect 36446 16124 36452 16136
rect 36504 16164 36510 16176
rect 38194 16164 38200 16176
rect 36504 16136 38200 16164
rect 36504 16124 36510 16136
rect 38194 16124 38200 16136
rect 38252 16164 38258 16176
rect 39025 16167 39083 16173
rect 39025 16164 39037 16167
rect 38252 16136 39037 16164
rect 38252 16124 38258 16136
rect 39025 16133 39037 16136
rect 39071 16164 39083 16167
rect 42794 16164 42800 16176
rect 39071 16136 42800 16164
rect 39071 16133 39083 16136
rect 39025 16127 39083 16133
rect 42794 16124 42800 16136
rect 42852 16124 42858 16176
rect 36906 16096 36912 16108
rect 36867 16068 36912 16096
rect 36906 16056 36912 16068
rect 36964 16056 36970 16108
rect 37645 16099 37703 16105
rect 37645 16065 37657 16099
rect 37691 16065 37703 16099
rect 37645 16059 37703 16065
rect 38473 16099 38531 16105
rect 38473 16065 38485 16099
rect 38519 16065 38531 16099
rect 38473 16059 38531 16065
rect 34698 15988 34704 16040
rect 34756 16028 34762 16040
rect 37660 16028 37688 16059
rect 34756 16000 37688 16028
rect 34756 15988 34762 16000
rect 38102 15960 38108 15972
rect 36004 15932 38108 15960
rect 36004 15904 36032 15932
rect 38102 15920 38108 15932
rect 38160 15920 38166 15972
rect 38488 15960 38516 16059
rect 38562 16056 38568 16108
rect 38620 16096 38626 16108
rect 41233 16099 41291 16105
rect 41233 16096 41245 16099
rect 38620 16068 41245 16096
rect 38620 16056 38626 16068
rect 41233 16065 41245 16068
rect 41279 16065 41291 16099
rect 41233 16059 41291 16065
rect 41322 16056 41328 16108
rect 41380 16096 41386 16108
rect 54018 16096 54024 16108
rect 41380 16068 51074 16096
rect 53979 16068 54024 16096
rect 41380 16056 41386 16068
rect 40773 16031 40831 16037
rect 40773 15997 40785 16031
rect 40819 16028 40831 16031
rect 41414 16028 41420 16040
rect 40819 16000 41420 16028
rect 40819 15997 40831 16000
rect 40773 15991 40831 15997
rect 41414 15988 41420 16000
rect 41472 15988 41478 16040
rect 42518 16028 42524 16040
rect 42168 16000 42524 16028
rect 42168 15960 42196 16000
rect 42518 15988 42524 16000
rect 42576 16028 42582 16040
rect 43806 16028 43812 16040
rect 42576 16000 43812 16028
rect 42576 15988 42582 16000
rect 43806 15988 43812 16000
rect 43864 16028 43870 16040
rect 43864 16000 44404 16028
rect 43864 15988 43870 16000
rect 43714 15960 43720 15972
rect 38488 15932 42196 15960
rect 43675 15932 43720 15960
rect 43714 15920 43720 15932
rect 43772 15920 43778 15972
rect 34422 15892 34428 15904
rect 34341 15864 34428 15892
rect 33965 15855 34023 15861
rect 34422 15852 34428 15864
rect 34480 15852 34486 15904
rect 34514 15852 34520 15904
rect 34572 15892 34578 15904
rect 35986 15892 35992 15904
rect 34572 15864 35992 15892
rect 34572 15852 34578 15864
rect 35986 15852 35992 15864
rect 36044 15852 36050 15904
rect 37458 15892 37464 15904
rect 37419 15864 37464 15892
rect 37458 15852 37464 15864
rect 37516 15852 37522 15904
rect 38194 15892 38200 15904
rect 38155 15864 38200 15892
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 38286 15852 38292 15904
rect 38344 15892 38350 15904
rect 41230 15892 41236 15904
rect 38344 15864 41236 15892
rect 38344 15852 38350 15864
rect 41230 15852 41236 15864
rect 41288 15852 41294 15904
rect 41322 15852 41328 15904
rect 41380 15892 41386 15904
rect 41417 15895 41475 15901
rect 41417 15892 41429 15895
rect 41380 15864 41429 15892
rect 41380 15852 41386 15864
rect 41417 15861 41429 15864
rect 41463 15861 41475 15895
rect 42610 15892 42616 15904
rect 42571 15864 42616 15892
rect 41417 15855 41475 15861
rect 42610 15852 42616 15864
rect 42668 15852 42674 15904
rect 42978 15852 42984 15904
rect 43036 15892 43042 15904
rect 44376 15901 44404 16000
rect 51046 15960 51074 16068
rect 54018 16056 54024 16068
rect 54076 16056 54082 16108
rect 53282 15960 53288 15972
rect 51046 15932 53288 15960
rect 53282 15920 53288 15932
rect 53340 15920 53346 15972
rect 43165 15895 43223 15901
rect 43165 15892 43177 15895
rect 43036 15864 43177 15892
rect 43036 15852 43042 15864
rect 43165 15861 43177 15864
rect 43211 15861 43223 15895
rect 43165 15855 43223 15861
rect 44361 15895 44419 15901
rect 44361 15861 44373 15895
rect 44407 15892 44419 15895
rect 53650 15892 53656 15904
rect 44407 15864 53656 15892
rect 44407 15861 44419 15864
rect 44361 15855 44419 15861
rect 53650 15852 53656 15864
rect 53708 15852 53714 15904
rect 1104 15802 54832 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 54832 15802
rect 1104 15728 54832 15750
rect 16482 15648 16488 15700
rect 16540 15688 16546 15700
rect 16761 15691 16819 15697
rect 16761 15688 16773 15691
rect 16540 15660 16773 15688
rect 16540 15648 16546 15660
rect 16761 15657 16773 15660
rect 16807 15657 16819 15691
rect 16761 15651 16819 15657
rect 16850 15648 16856 15700
rect 16908 15688 16914 15700
rect 17770 15688 17776 15700
rect 16908 15660 17776 15688
rect 16908 15648 16914 15660
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 20622 15688 20628 15700
rect 19444 15660 20628 15688
rect 19444 15620 19472 15660
rect 20622 15648 20628 15660
rect 20680 15648 20686 15700
rect 21634 15688 21640 15700
rect 21595 15660 21640 15688
rect 21634 15648 21640 15660
rect 21692 15648 21698 15700
rect 24762 15648 24768 15700
rect 24820 15688 24826 15700
rect 25961 15691 26019 15697
rect 25961 15688 25973 15691
rect 24820 15660 25973 15688
rect 24820 15648 24826 15660
rect 25961 15657 25973 15660
rect 26007 15688 26019 15691
rect 26326 15688 26332 15700
rect 26007 15660 26332 15688
rect 26007 15657 26019 15660
rect 25961 15651 26019 15657
rect 26326 15648 26332 15660
rect 26384 15648 26390 15700
rect 28626 15648 28632 15700
rect 28684 15688 28690 15700
rect 29733 15691 29791 15697
rect 29733 15688 29745 15691
rect 28684 15660 29745 15688
rect 28684 15648 28690 15660
rect 29733 15657 29745 15660
rect 29779 15657 29791 15691
rect 33686 15688 33692 15700
rect 29733 15651 29791 15657
rect 31726 15660 33692 15688
rect 20806 15620 20812 15632
rect 16132 15592 19472 15620
rect 20719 15592 20812 15620
rect 13725 15555 13783 15561
rect 13725 15521 13737 15555
rect 13771 15552 13783 15555
rect 15930 15552 15936 15564
rect 13771 15524 15936 15552
rect 13771 15521 13783 15524
rect 13725 15515 13783 15521
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 1857 15487 1915 15493
rect 1857 15453 1869 15487
rect 1903 15484 1915 15487
rect 15562 15484 15568 15496
rect 1903 15456 15568 15484
rect 1903 15453 1915 15456
rect 1857 15447 1915 15453
rect 15562 15444 15568 15456
rect 15620 15444 15626 15496
rect 16132 15493 16160 15592
rect 20806 15580 20812 15592
rect 20864 15620 20870 15632
rect 21726 15620 21732 15632
rect 20864 15592 21732 15620
rect 20864 15580 20870 15592
rect 21726 15580 21732 15592
rect 21784 15580 21790 15632
rect 28537 15623 28595 15629
rect 28537 15589 28549 15623
rect 28583 15620 28595 15623
rect 31726 15620 31754 15660
rect 33686 15648 33692 15660
rect 33744 15648 33750 15700
rect 33873 15691 33931 15697
rect 33873 15657 33885 15691
rect 33919 15688 33931 15691
rect 34698 15688 34704 15700
rect 33919 15660 34704 15688
rect 33919 15657 33931 15660
rect 33873 15651 33931 15657
rect 34698 15648 34704 15660
rect 34756 15648 34762 15700
rect 35989 15691 36047 15697
rect 35084 15660 35664 15688
rect 33594 15620 33600 15632
rect 28583 15592 31754 15620
rect 32784 15592 33600 15620
rect 28583 15589 28595 15592
rect 28537 15583 28595 15589
rect 17037 15555 17095 15561
rect 17037 15521 17049 15555
rect 17083 15552 17095 15555
rect 17954 15552 17960 15564
rect 17083 15524 17960 15552
rect 17083 15521 17095 15524
rect 17037 15515 17095 15521
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 18782 15552 18788 15564
rect 18743 15524 18788 15552
rect 18782 15512 18788 15524
rect 18840 15512 18846 15564
rect 22278 15552 22284 15564
rect 22239 15524 22284 15552
rect 22278 15512 22284 15524
rect 22336 15512 22342 15564
rect 26234 15512 26240 15564
rect 26292 15552 26298 15564
rect 28902 15552 28908 15564
rect 26292 15524 28908 15552
rect 26292 15512 26298 15524
rect 28902 15512 28908 15524
rect 28960 15512 28966 15564
rect 29089 15555 29147 15561
rect 29089 15521 29101 15555
rect 29135 15552 29147 15555
rect 29362 15552 29368 15564
rect 29135 15524 29368 15552
rect 29135 15521 29147 15524
rect 29089 15515 29147 15521
rect 29362 15512 29368 15524
rect 29420 15552 29426 15564
rect 32784 15561 32812 15592
rect 33594 15580 33600 15592
rect 33652 15580 33658 15632
rect 32769 15555 32827 15561
rect 29420 15524 31800 15552
rect 29420 15512 29426 15524
rect 16117 15487 16175 15493
rect 16117 15453 16129 15487
rect 16163 15453 16175 15487
rect 16942 15484 16948 15496
rect 16903 15456 16948 15484
rect 16117 15447 16175 15453
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 17126 15484 17132 15496
rect 17087 15456 17132 15484
rect 17126 15444 17132 15456
rect 17184 15444 17190 15496
rect 17218 15444 17224 15496
rect 17276 15484 17282 15496
rect 19426 15484 19432 15496
rect 17276 15456 17321 15484
rect 19387 15456 19432 15484
rect 17276 15444 17282 15456
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 19518 15444 19524 15496
rect 19576 15484 19582 15496
rect 19685 15487 19743 15493
rect 19685 15484 19697 15487
rect 19576 15456 19697 15484
rect 19576 15444 19582 15456
rect 19685 15453 19697 15456
rect 19731 15453 19743 15487
rect 21818 15484 21824 15496
rect 21779 15456 21824 15484
rect 19685 15447 19743 15453
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 22066 15456 24593 15484
rect 14553 15419 14611 15425
rect 14553 15385 14565 15419
rect 14599 15416 14611 15419
rect 14734 15416 14740 15428
rect 14599 15388 14740 15416
rect 14599 15385 14611 15388
rect 14553 15379 14611 15385
rect 14734 15376 14740 15388
rect 14792 15376 14798 15428
rect 15102 15376 15108 15428
rect 15160 15416 15166 15428
rect 15657 15419 15715 15425
rect 15657 15416 15669 15419
rect 15160 15388 15669 15416
rect 15160 15376 15166 15388
rect 15657 15385 15669 15388
rect 15703 15416 15715 15419
rect 17586 15416 17592 15428
rect 15703 15388 17592 15416
rect 15703 15385 15715 15388
rect 15657 15379 15715 15385
rect 17586 15376 17592 15388
rect 17644 15376 17650 15428
rect 20346 15416 20352 15428
rect 17972 15388 20352 15416
rect 1670 15348 1676 15360
rect 1631 15320 1676 15348
rect 1670 15308 1676 15320
rect 1728 15308 1734 15360
rect 15010 15348 15016 15360
rect 14971 15320 15016 15348
rect 15010 15308 15016 15320
rect 15068 15308 15074 15360
rect 16301 15351 16359 15357
rect 16301 15317 16313 15351
rect 16347 15348 16359 15351
rect 17972 15348 18000 15388
rect 20346 15376 20352 15388
rect 20404 15376 20410 15428
rect 18138 15348 18144 15360
rect 16347 15320 18000 15348
rect 18099 15320 18144 15348
rect 16347 15317 16359 15320
rect 16301 15311 16359 15317
rect 18138 15308 18144 15320
rect 18196 15308 18202 15360
rect 18230 15308 18236 15360
rect 18288 15348 18294 15360
rect 18509 15351 18567 15357
rect 18509 15348 18521 15351
rect 18288 15320 18521 15348
rect 18288 15308 18294 15320
rect 18509 15317 18521 15320
rect 18555 15317 18567 15351
rect 18509 15311 18567 15317
rect 18598 15308 18604 15360
rect 18656 15348 18662 15360
rect 18656 15320 18701 15348
rect 18656 15308 18662 15320
rect 19978 15308 19984 15360
rect 20036 15348 20042 15360
rect 22066 15348 22094 15456
rect 24581 15453 24593 15456
rect 24627 15484 24639 15487
rect 24670 15484 24676 15496
rect 24627 15456 24676 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 24670 15444 24676 15456
rect 24728 15444 24734 15496
rect 26510 15484 26516 15496
rect 26471 15456 26516 15484
rect 26510 15444 26516 15456
rect 26568 15444 26574 15496
rect 27890 15444 27896 15496
rect 27948 15484 27954 15496
rect 28074 15484 28080 15496
rect 27948 15456 28080 15484
rect 27948 15444 27954 15456
rect 28074 15444 28080 15456
rect 28132 15444 28138 15496
rect 28353 15487 28411 15493
rect 28353 15453 28365 15487
rect 28399 15484 28411 15487
rect 28534 15484 28540 15496
rect 28399 15456 28540 15484
rect 28399 15453 28411 15456
rect 28353 15447 28411 15453
rect 28534 15444 28540 15456
rect 28592 15444 28598 15496
rect 28997 15487 29055 15493
rect 28997 15453 29009 15487
rect 29043 15484 29055 15487
rect 29454 15484 29460 15496
rect 29043 15456 29460 15484
rect 29043 15453 29055 15456
rect 28997 15447 29055 15453
rect 29454 15444 29460 15456
rect 29512 15444 29518 15496
rect 29914 15484 29920 15496
rect 29875 15456 29920 15484
rect 29914 15444 29920 15456
rect 29972 15444 29978 15496
rect 30009 15487 30067 15493
rect 30009 15453 30021 15487
rect 30055 15453 30067 15487
rect 30009 15447 30067 15453
rect 30745 15487 30803 15493
rect 30745 15453 30757 15487
rect 30791 15484 30803 15487
rect 31294 15484 31300 15496
rect 30791 15456 31300 15484
rect 30791 15453 30803 15456
rect 30745 15447 30803 15453
rect 22186 15376 22192 15428
rect 22244 15416 22250 15428
rect 22526 15419 22584 15425
rect 22526 15416 22538 15419
rect 22244 15388 22538 15416
rect 22244 15376 22250 15388
rect 22526 15385 22538 15388
rect 22572 15385 22584 15419
rect 22526 15379 22584 15385
rect 24026 15376 24032 15428
rect 24084 15416 24090 15428
rect 24826 15419 24884 15425
rect 24826 15416 24838 15419
rect 24084 15388 24838 15416
rect 24084 15376 24090 15388
rect 24826 15385 24838 15388
rect 24872 15385 24884 15419
rect 24826 15379 24884 15385
rect 27065 15419 27123 15425
rect 27065 15385 27077 15419
rect 27111 15416 27123 15419
rect 29178 15416 29184 15428
rect 27111 15388 29184 15416
rect 27111 15385 27123 15388
rect 27065 15379 27123 15385
rect 29178 15376 29184 15388
rect 29236 15376 29242 15428
rect 29270 15376 29276 15428
rect 29328 15416 29334 15428
rect 30024 15416 30052 15447
rect 31294 15444 31300 15456
rect 31352 15444 31358 15496
rect 31772 15484 31800 15524
rect 32769 15521 32781 15555
rect 32815 15521 32827 15555
rect 32769 15515 32827 15521
rect 33134 15512 33140 15564
rect 33192 15552 33198 15564
rect 35084 15552 35112 15660
rect 33192 15524 35112 15552
rect 35253 15555 35311 15561
rect 33192 15512 33198 15524
rect 35253 15521 35265 15555
rect 35299 15552 35311 15555
rect 35526 15552 35532 15564
rect 35299 15524 35532 15552
rect 35299 15521 35311 15524
rect 35253 15515 35311 15521
rect 35526 15512 35532 15524
rect 35584 15512 35590 15564
rect 35636 15552 35664 15660
rect 35989 15657 36001 15691
rect 36035 15688 36047 15691
rect 37550 15688 37556 15700
rect 36035 15660 37556 15688
rect 36035 15657 36047 15660
rect 35989 15651 36047 15657
rect 37550 15648 37556 15660
rect 37608 15648 37614 15700
rect 37918 15688 37924 15700
rect 37879 15660 37924 15688
rect 37918 15648 37924 15660
rect 37976 15648 37982 15700
rect 40037 15691 40095 15697
rect 40037 15657 40049 15691
rect 40083 15688 40095 15691
rect 40083 15660 42748 15688
rect 40083 15657 40095 15660
rect 40037 15651 40095 15657
rect 36538 15580 36544 15632
rect 36596 15620 36602 15632
rect 38378 15620 38384 15632
rect 36596 15592 38384 15620
rect 36596 15580 36602 15592
rect 38378 15580 38384 15592
rect 38436 15580 38442 15632
rect 39022 15580 39028 15632
rect 39080 15620 39086 15632
rect 39666 15620 39672 15632
rect 39080 15592 39672 15620
rect 39080 15580 39086 15592
rect 35636 15524 38976 15552
rect 32214 15484 32220 15496
rect 31772 15456 32220 15484
rect 32214 15444 32220 15456
rect 32272 15444 32278 15496
rect 33229 15487 33287 15493
rect 33229 15484 33241 15487
rect 32324 15456 33241 15484
rect 30926 15416 30932 15428
rect 29328 15388 30052 15416
rect 30887 15388 30932 15416
rect 29328 15376 29334 15388
rect 30926 15376 30932 15388
rect 30984 15376 30990 15428
rect 31110 15376 31116 15428
rect 31168 15416 31174 15428
rect 32324 15416 32352 15456
rect 33229 15453 33241 15456
rect 33275 15453 33287 15487
rect 33229 15447 33287 15453
rect 34514 15444 34520 15496
rect 34572 15484 34578 15496
rect 35069 15487 35127 15493
rect 35069 15484 35081 15487
rect 34572 15456 35081 15484
rect 34572 15444 34578 15456
rect 35069 15453 35081 15456
rect 35115 15453 35127 15487
rect 35069 15447 35127 15453
rect 35158 15444 35164 15496
rect 35216 15484 35222 15496
rect 35345 15487 35403 15493
rect 35216 15456 35261 15484
rect 35216 15444 35222 15456
rect 35345 15453 35357 15487
rect 35391 15484 35403 15487
rect 35710 15484 35716 15496
rect 35391 15456 35716 15484
rect 35391 15453 35403 15456
rect 35345 15447 35403 15453
rect 35710 15444 35716 15456
rect 35768 15444 35774 15496
rect 36446 15484 36452 15496
rect 36407 15456 36452 15484
rect 36446 15444 36452 15456
rect 36504 15444 36510 15496
rect 38948 15493 38976 15524
rect 39132 15493 39160 15592
rect 39666 15580 39672 15592
rect 39724 15580 39730 15632
rect 40052 15552 40080 15651
rect 41506 15580 41512 15632
rect 41564 15620 41570 15632
rect 42720 15620 42748 15660
rect 42794 15648 42800 15700
rect 42852 15688 42858 15700
rect 43162 15688 43168 15700
rect 42852 15660 43168 15688
rect 42852 15648 42858 15660
rect 43162 15648 43168 15660
rect 43220 15688 43226 15700
rect 43809 15691 43867 15697
rect 43809 15688 43821 15691
rect 43220 15660 43821 15688
rect 43220 15648 43226 15660
rect 43809 15657 43821 15660
rect 43855 15657 43867 15691
rect 54018 15688 54024 15700
rect 43809 15651 43867 15657
rect 51046 15660 54024 15688
rect 51046 15620 51074 15660
rect 54018 15648 54024 15660
rect 54076 15648 54082 15700
rect 53282 15620 53288 15632
rect 41564 15592 41828 15620
rect 42720 15592 51074 15620
rect 53243 15592 53288 15620
rect 41564 15580 41570 15592
rect 41414 15552 41420 15564
rect 39224 15524 40080 15552
rect 41375 15524 41420 15552
rect 39224 15493 39252 15524
rect 41414 15512 41420 15524
rect 41472 15512 41478 15564
rect 41800 15552 41828 15592
rect 53282 15580 53288 15592
rect 53340 15580 53346 15632
rect 54021 15555 54079 15561
rect 54021 15552 54033 15555
rect 41800 15524 54033 15552
rect 54021 15521 54033 15524
rect 54067 15521 54079 15555
rect 54021 15515 54079 15521
rect 38933 15487 38991 15493
rect 38933 15453 38945 15487
rect 38979 15453 38991 15487
rect 38933 15447 38991 15453
rect 39117 15487 39175 15493
rect 39117 15453 39129 15487
rect 39163 15453 39175 15487
rect 39117 15447 39175 15453
rect 39209 15487 39267 15493
rect 39209 15453 39221 15487
rect 39255 15453 39267 15487
rect 39209 15447 39267 15453
rect 39298 15444 39304 15496
rect 39356 15484 39362 15496
rect 39356 15456 39401 15484
rect 39356 15444 39362 15456
rect 41506 15444 41512 15496
rect 41564 15484 41570 15496
rect 41877 15487 41935 15493
rect 41877 15484 41889 15487
rect 41564 15456 41889 15484
rect 41564 15444 41570 15456
rect 41877 15453 41889 15456
rect 41923 15453 41935 15487
rect 42058 15484 42064 15496
rect 42019 15456 42064 15484
rect 41877 15447 41935 15453
rect 42058 15444 42064 15456
rect 42116 15444 42122 15496
rect 42518 15484 42524 15496
rect 42479 15456 42524 15484
rect 42518 15444 42524 15456
rect 42576 15444 42582 15496
rect 42705 15487 42763 15493
rect 42705 15453 42717 15487
rect 42751 15484 42763 15487
rect 42886 15484 42892 15496
rect 42751 15456 42892 15484
rect 42751 15453 42763 15456
rect 42705 15447 42763 15453
rect 42886 15444 42892 15456
rect 42944 15444 42950 15496
rect 43346 15484 43352 15496
rect 43307 15456 43352 15484
rect 43346 15444 43352 15456
rect 43404 15444 43410 15496
rect 53558 15444 53564 15496
rect 53616 15484 53622 15496
rect 54202 15484 54208 15496
rect 53616 15456 54208 15484
rect 53616 15444 53622 15456
rect 54202 15444 54208 15456
rect 54260 15444 54266 15496
rect 31168 15388 32352 15416
rect 32524 15419 32582 15425
rect 31168 15376 31174 15388
rect 32524 15385 32536 15419
rect 32570 15416 32582 15419
rect 37458 15416 37464 15428
rect 32570 15388 37464 15416
rect 32570 15385 32582 15388
rect 32524 15379 32582 15385
rect 37458 15376 37464 15388
rect 37516 15376 37522 15428
rect 40494 15416 40500 15428
rect 39500 15388 40500 15416
rect 23658 15348 23664 15360
rect 20036 15320 22094 15348
rect 23619 15320 23664 15348
rect 20036 15308 20042 15320
rect 23658 15308 23664 15320
rect 23716 15308 23722 15360
rect 24118 15308 24124 15360
rect 24176 15348 24182 15360
rect 26786 15348 26792 15360
rect 24176 15320 26792 15348
rect 24176 15308 24182 15320
rect 26786 15308 26792 15320
rect 26844 15348 26850 15360
rect 27525 15351 27583 15357
rect 27525 15348 27537 15351
rect 26844 15320 27537 15348
rect 26844 15308 26850 15320
rect 27525 15317 27537 15320
rect 27571 15348 27583 15351
rect 27614 15348 27620 15360
rect 27571 15320 27620 15348
rect 27571 15317 27583 15320
rect 27525 15311 27583 15317
rect 27614 15308 27620 15320
rect 27672 15308 27678 15360
rect 28169 15351 28227 15357
rect 28169 15317 28181 15351
rect 28215 15348 28227 15351
rect 28626 15348 28632 15360
rect 28215 15320 28632 15348
rect 28215 15317 28227 15320
rect 28169 15311 28227 15317
rect 28626 15308 28632 15320
rect 28684 15348 28690 15360
rect 28810 15348 28816 15360
rect 28684 15320 28816 15348
rect 28684 15308 28690 15320
rect 28810 15308 28816 15320
rect 28868 15308 28874 15360
rect 30374 15308 30380 15360
rect 30432 15348 30438 15360
rect 30561 15351 30619 15357
rect 30561 15348 30573 15351
rect 30432 15320 30573 15348
rect 30432 15308 30438 15320
rect 30561 15317 30573 15320
rect 30607 15317 30619 15351
rect 30561 15311 30619 15317
rect 30834 15308 30840 15360
rect 30892 15348 30898 15360
rect 31389 15351 31447 15357
rect 31389 15348 31401 15351
rect 30892 15320 31401 15348
rect 30892 15308 30898 15320
rect 31389 15317 31401 15320
rect 31435 15317 31447 15351
rect 31389 15311 31447 15317
rect 34790 15308 34796 15360
rect 34848 15348 34854 15360
rect 34885 15351 34943 15357
rect 34885 15348 34897 15351
rect 34848 15320 34897 15348
rect 34848 15308 34854 15320
rect 34885 15317 34897 15320
rect 34931 15317 34943 15351
rect 34885 15311 34943 15317
rect 35342 15308 35348 15360
rect 35400 15348 35406 15360
rect 38838 15348 38844 15360
rect 35400 15320 38844 15348
rect 35400 15308 35406 15320
rect 38838 15308 38844 15320
rect 38896 15348 38902 15360
rect 39390 15348 39396 15360
rect 38896 15320 39396 15348
rect 38896 15308 38902 15320
rect 39390 15308 39396 15320
rect 39448 15308 39454 15360
rect 39500 15357 39528 15388
rect 40494 15376 40500 15388
rect 40552 15376 40558 15428
rect 41172 15419 41230 15425
rect 41172 15385 41184 15419
rect 41218 15416 41230 15419
rect 41218 15388 43208 15416
rect 41218 15385 41230 15388
rect 41172 15379 41230 15385
rect 39485 15351 39543 15357
rect 39485 15317 39497 15351
rect 39531 15317 39543 15351
rect 39485 15311 39543 15317
rect 39666 15308 39672 15360
rect 39724 15348 39730 15360
rect 41322 15348 41328 15360
rect 39724 15320 41328 15348
rect 39724 15308 39730 15320
rect 41322 15308 41328 15320
rect 41380 15308 41386 15360
rect 41690 15308 41696 15360
rect 41748 15348 41754 15360
rect 41969 15351 42027 15357
rect 41969 15348 41981 15351
rect 41748 15320 41981 15348
rect 41748 15308 41754 15320
rect 41969 15317 41981 15320
rect 42015 15317 42027 15351
rect 42610 15348 42616 15360
rect 42571 15320 42616 15348
rect 41969 15311 42027 15317
rect 42610 15308 42616 15320
rect 42668 15308 42674 15360
rect 43180 15357 43208 15388
rect 43438 15376 43444 15428
rect 43496 15416 43502 15428
rect 45189 15419 45247 15425
rect 45189 15416 45201 15419
rect 43496 15388 45201 15416
rect 43496 15376 43502 15388
rect 45189 15385 45201 15388
rect 45235 15385 45247 15419
rect 45189 15379 45247 15385
rect 52825 15419 52883 15425
rect 52825 15385 52837 15419
rect 52871 15416 52883 15419
rect 53466 15416 53472 15428
rect 52871 15388 53472 15416
rect 52871 15385 52883 15388
rect 52825 15379 52883 15385
rect 53466 15376 53472 15388
rect 53524 15376 53530 15428
rect 43165 15351 43223 15357
rect 43165 15317 43177 15351
rect 43211 15317 43223 15351
rect 44450 15348 44456 15360
rect 44411 15320 44456 15348
rect 43165 15311 43223 15317
rect 44450 15308 44456 15320
rect 44508 15308 44514 15360
rect 1104 15258 54832 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 54832 15258
rect 1104 15184 54832 15206
rect 13725 15147 13783 15153
rect 13725 15113 13737 15147
rect 13771 15144 13783 15147
rect 18690 15144 18696 15156
rect 13771 15116 18696 15144
rect 13771 15113 13783 15116
rect 13725 15107 13783 15113
rect 18690 15104 18696 15116
rect 18748 15104 18754 15156
rect 19334 15104 19340 15156
rect 19392 15144 19398 15156
rect 19521 15147 19579 15153
rect 19521 15144 19533 15147
rect 19392 15116 19533 15144
rect 19392 15104 19398 15116
rect 19521 15113 19533 15116
rect 19567 15113 19579 15147
rect 20806 15144 20812 15156
rect 20767 15116 20812 15144
rect 19521 15107 19579 15113
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 22738 15104 22744 15156
rect 22796 15144 22802 15156
rect 23293 15147 23351 15153
rect 23293 15144 23305 15147
rect 22796 15116 23305 15144
rect 22796 15104 22802 15116
rect 23293 15113 23305 15116
rect 23339 15113 23351 15147
rect 26050 15144 26056 15156
rect 23293 15107 23351 15113
rect 23584 15116 26056 15144
rect 14274 15076 14280 15088
rect 14235 15048 14280 15076
rect 14274 15036 14280 15048
rect 14332 15036 14338 15088
rect 15930 15076 15936 15088
rect 15843 15048 15936 15076
rect 15930 15036 15936 15048
rect 15988 15076 15994 15088
rect 17678 15076 17684 15088
rect 15988 15048 17684 15076
rect 15988 15036 15994 15048
rect 17678 15036 17684 15048
rect 17736 15036 17742 15088
rect 18233 15079 18291 15085
rect 18233 15045 18245 15079
rect 18279 15076 18291 15079
rect 18322 15076 18328 15088
rect 18279 15048 18328 15076
rect 18279 15045 18291 15048
rect 18233 15039 18291 15045
rect 18322 15036 18328 15048
rect 18380 15036 18386 15088
rect 18414 15036 18420 15088
rect 18472 15076 18478 15088
rect 23584 15076 23612 15116
rect 26050 15104 26056 15116
rect 26108 15104 26114 15156
rect 26510 15104 26516 15156
rect 26568 15144 26574 15156
rect 27157 15147 27215 15153
rect 27157 15144 27169 15147
rect 26568 15116 27169 15144
rect 26568 15104 26574 15116
rect 27157 15113 27169 15116
rect 27203 15113 27215 15147
rect 27157 15107 27215 15113
rect 27430 15104 27436 15156
rect 27488 15144 27494 15156
rect 28350 15144 28356 15156
rect 27488 15116 28356 15144
rect 27488 15104 27494 15116
rect 23750 15076 23756 15088
rect 18472 15048 23612 15076
rect 23711 15048 23756 15076
rect 18472 15036 18478 15048
rect 23750 15036 23756 15048
rect 23808 15036 23814 15088
rect 25130 15036 25136 15088
rect 25188 15076 25194 15088
rect 28276 15076 28304 15116
rect 28350 15104 28356 15116
rect 28408 15104 28414 15156
rect 28994 15104 29000 15156
rect 29052 15144 29058 15156
rect 41322 15153 41328 15156
rect 29089 15147 29147 15153
rect 29089 15144 29101 15147
rect 29052 15116 29101 15144
rect 29052 15104 29058 15116
rect 29089 15113 29101 15116
rect 29135 15113 29147 15147
rect 41309 15147 41328 15153
rect 29089 15107 29147 15113
rect 29196 15116 39896 15144
rect 25188 15048 27476 15076
rect 28276 15048 28704 15076
rect 25188 15036 25194 15048
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 15008 1915 15011
rect 4614 15008 4620 15020
rect 1903 14980 4620 15008
rect 1903 14977 1915 14980
rect 1857 14971 1915 14977
rect 4614 14968 4620 14980
rect 4672 14968 4678 15020
rect 14734 15008 14740 15020
rect 14695 14980 14740 15008
rect 14734 14968 14740 14980
rect 14792 14968 14798 15020
rect 15378 14968 15384 15020
rect 15436 15008 15442 15020
rect 16666 15008 16672 15020
rect 15436 14980 16672 15008
rect 15436 14968 15442 14980
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 15008 17187 15011
rect 20070 15008 20076 15020
rect 17175 14980 20076 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 20070 14968 20076 14980
rect 20128 14968 20134 15020
rect 22554 15008 22560 15020
rect 20824 14980 22560 15008
rect 11698 14900 11704 14952
rect 11756 14940 11762 14952
rect 16853 14943 16911 14949
rect 16853 14940 16865 14943
rect 11756 14912 16865 14940
rect 11756 14900 11762 14912
rect 16853 14909 16865 14912
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 17037 14943 17095 14949
rect 17037 14909 17049 14943
rect 17083 14909 17095 14943
rect 17037 14903 17095 14909
rect 17221 14943 17279 14949
rect 17221 14909 17233 14943
rect 17267 14909 17279 14943
rect 17221 14903 17279 14909
rect 17052 14872 17080 14903
rect 16500 14844 17080 14872
rect 16500 14816 16528 14844
rect 17126 14832 17132 14884
rect 17184 14872 17190 14884
rect 17236 14872 17264 14903
rect 17310 14900 17316 14952
rect 17368 14940 17374 14952
rect 17368 14912 17413 14940
rect 17368 14900 17374 14912
rect 17586 14900 17592 14952
rect 17644 14940 17650 14952
rect 20530 14940 20536 14952
rect 17644 14912 20536 14940
rect 17644 14900 17650 14912
rect 20530 14900 20536 14912
rect 20588 14940 20594 14952
rect 20824 14940 20852 14980
rect 22554 14968 22560 14980
rect 22612 14968 22618 15020
rect 22649 15011 22707 15017
rect 22649 14977 22661 15011
rect 22695 15008 22707 15011
rect 23382 15008 23388 15020
rect 22695 14980 23388 15008
rect 22695 14977 22707 14980
rect 22649 14971 22707 14977
rect 23382 14968 23388 14980
rect 23440 14968 23446 15020
rect 23658 15008 23664 15020
rect 23571 14980 23664 15008
rect 23658 14968 23664 14980
rect 23716 15008 23722 15020
rect 24762 15008 24768 15020
rect 23716 14980 24768 15008
rect 23716 14968 23722 14980
rect 24762 14968 24768 14980
rect 24820 14968 24826 15020
rect 27448 15008 27476 15048
rect 27525 15011 27583 15017
rect 27525 15008 27537 15011
rect 27448 14980 27537 15008
rect 27525 14977 27537 14980
rect 27571 14977 27583 15011
rect 28169 15011 28227 15017
rect 28169 15008 28181 15011
rect 27525 14971 27583 14977
rect 27724 14980 28181 15008
rect 20588 14912 20852 14940
rect 20901 14943 20959 14949
rect 20588 14900 20594 14912
rect 20901 14909 20913 14943
rect 20947 14909 20959 14943
rect 20901 14903 20959 14909
rect 21085 14943 21143 14949
rect 21085 14909 21097 14943
rect 21131 14940 21143 14943
rect 21174 14940 21180 14952
rect 21131 14912 21180 14940
rect 21131 14909 21143 14912
rect 21085 14903 21143 14909
rect 17184 14844 17264 14872
rect 17184 14832 17190 14844
rect 17770 14832 17776 14884
rect 17828 14872 17834 14884
rect 20441 14875 20499 14881
rect 20441 14872 20453 14875
rect 17828 14844 20453 14872
rect 17828 14832 17834 14844
rect 20441 14841 20453 14844
rect 20487 14841 20499 14875
rect 20441 14835 20499 14841
rect 20806 14832 20812 14884
rect 20864 14872 20870 14884
rect 20916 14872 20944 14903
rect 21174 14900 21180 14912
rect 21232 14900 21238 14952
rect 22830 14940 22836 14952
rect 22791 14912 22836 14940
rect 22830 14900 22836 14912
rect 22888 14900 22894 14952
rect 23842 14940 23848 14952
rect 23803 14912 23848 14940
rect 23842 14900 23848 14912
rect 23900 14900 23906 14952
rect 25314 14940 25320 14952
rect 25275 14912 25320 14940
rect 25314 14900 25320 14912
rect 25372 14900 25378 14952
rect 25774 14940 25780 14952
rect 25735 14912 25780 14940
rect 25774 14900 25780 14912
rect 25832 14900 25838 14952
rect 26326 14940 26332 14952
rect 26287 14912 26332 14940
rect 26326 14900 26332 14912
rect 26384 14900 26390 14952
rect 26878 14900 26884 14952
rect 26936 14940 26942 14952
rect 27062 14940 27068 14952
rect 26936 14912 27068 14940
rect 26936 14900 26942 14912
rect 27062 14900 27068 14912
rect 27120 14940 27126 14952
rect 27333 14943 27391 14949
rect 27333 14940 27345 14943
rect 27120 14912 27345 14940
rect 27120 14900 27126 14912
rect 27333 14909 27345 14912
rect 27379 14909 27391 14943
rect 27333 14903 27391 14909
rect 27430 14900 27436 14952
rect 27488 14940 27494 14952
rect 27614 14940 27620 14952
rect 27488 14912 27533 14940
rect 27575 14912 27620 14940
rect 27488 14900 27494 14912
rect 27614 14900 27620 14912
rect 27672 14900 27678 14952
rect 20864 14844 20944 14872
rect 20864 14832 20870 14844
rect 21634 14832 21640 14884
rect 21692 14872 21698 14884
rect 23198 14872 23204 14884
rect 21692 14844 23204 14872
rect 21692 14832 21698 14844
rect 23198 14832 23204 14844
rect 23256 14832 23262 14884
rect 24762 14832 24768 14884
rect 24820 14872 24826 14884
rect 27154 14872 27160 14884
rect 24820 14844 27160 14872
rect 24820 14832 24826 14844
rect 27154 14832 27160 14844
rect 27212 14872 27218 14884
rect 27724 14872 27752 14980
rect 28169 14977 28181 14980
rect 28215 14977 28227 15011
rect 28169 14971 28227 14977
rect 28258 14968 28264 15020
rect 28316 15008 28322 15020
rect 28353 15011 28411 15017
rect 28353 15008 28365 15011
rect 28316 14980 28365 15008
rect 28316 14968 28322 14980
rect 28353 14977 28365 14980
rect 28399 14977 28411 15011
rect 28353 14971 28411 14977
rect 28445 15011 28503 15017
rect 28445 14977 28457 15011
rect 28491 14977 28503 15011
rect 28445 14971 28503 14977
rect 27798 14900 27804 14952
rect 27856 14940 27862 14952
rect 28460 14940 28488 14971
rect 28534 14968 28540 15020
rect 28592 15017 28598 15020
rect 28592 15008 28600 15017
rect 28676 15008 28704 15048
rect 28902 15036 28908 15088
rect 28960 15076 28966 15088
rect 29196 15076 29224 15116
rect 29546 15076 29552 15088
rect 28960 15048 29224 15076
rect 29507 15048 29552 15076
rect 28960 15036 28966 15048
rect 29546 15036 29552 15048
rect 29604 15036 29610 15088
rect 36725 15079 36783 15085
rect 36725 15045 36737 15079
rect 36771 15076 36783 15079
rect 36771 15048 37964 15076
rect 36771 15045 36783 15048
rect 36725 15039 36783 15045
rect 30561 15011 30619 15017
rect 30561 15008 30573 15011
rect 28592 14980 28637 15008
rect 28676 14998 28764 15008
rect 28920 14998 30573 15008
rect 28676 14980 30573 14998
rect 28592 14971 28600 14980
rect 28592 14968 28598 14971
rect 28736 14970 28948 14980
rect 30561 14977 30573 14980
rect 30607 14977 30619 15011
rect 30561 14971 30619 14977
rect 33433 15011 33491 15017
rect 33433 14977 33445 15011
rect 33479 15008 33491 15011
rect 34149 15011 34207 15017
rect 34149 15008 34161 15011
rect 33479 14980 34161 15008
rect 33479 14977 33491 14980
rect 33433 14971 33491 14977
rect 34149 14977 34161 14980
rect 34195 14977 34207 15011
rect 34149 14971 34207 14977
rect 30466 14940 30472 14952
rect 27856 14912 28488 14940
rect 28966 14912 30472 14940
rect 27856 14900 27862 14912
rect 28966 14872 28994 14912
rect 30466 14900 30472 14912
rect 30524 14900 30530 14952
rect 30576 14940 30604 14971
rect 35158 14968 35164 15020
rect 35216 15008 35222 15020
rect 35434 15008 35440 15020
rect 35216 14980 35440 15008
rect 35216 14968 35222 14980
rect 35434 14968 35440 14980
rect 35492 15008 35498 15020
rect 35621 15011 35679 15017
rect 35621 15008 35633 15011
rect 35492 14980 35633 15008
rect 35492 14968 35498 14980
rect 35621 14977 35633 14980
rect 35667 14977 35679 15011
rect 35621 14971 35679 14977
rect 36909 15011 36967 15017
rect 36909 14977 36921 15011
rect 36955 15008 36967 15011
rect 37826 15008 37832 15020
rect 36955 14980 37832 15008
rect 36955 14977 36967 14980
rect 36909 14971 36967 14977
rect 37826 14968 37832 14980
rect 37884 14968 37890 15020
rect 37936 15008 37964 15048
rect 38010 15036 38016 15088
rect 38068 15076 38074 15088
rect 38470 15076 38476 15088
rect 38068 15048 38476 15076
rect 38068 15036 38074 15048
rect 38470 15036 38476 15048
rect 38528 15076 38534 15088
rect 39666 15076 39672 15088
rect 38528 15048 38884 15076
rect 39627 15048 39672 15076
rect 38528 15036 38534 15048
rect 38194 15008 38200 15020
rect 37936 14980 38200 15008
rect 38194 14968 38200 14980
rect 38252 14968 38258 15020
rect 38856 15017 38884 15048
rect 39666 15036 39672 15048
rect 39724 15036 39730 15088
rect 38585 15011 38643 15017
rect 38585 14977 38597 15011
rect 38631 15008 38643 15011
rect 38841 15011 38899 15017
rect 38631 14980 38792 15008
rect 38631 14977 38643 14980
rect 38585 14971 38643 14977
rect 31662 14940 31668 14952
rect 30576 14912 31156 14940
rect 31623 14912 31668 14940
rect 29178 14872 29184 14884
rect 27212 14844 27752 14872
rect 27816 14844 28994 14872
rect 29139 14844 29184 14872
rect 27212 14832 27218 14844
rect 1670 14804 1676 14816
rect 1631 14776 1676 14804
rect 1670 14764 1676 14776
rect 1728 14764 1734 14816
rect 13170 14804 13176 14816
rect 13131 14776 13176 14804
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 15378 14804 15384 14816
rect 15339 14776 15384 14804
rect 15378 14764 15384 14776
rect 15436 14764 15442 14816
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 16025 14807 16083 14813
rect 16025 14804 16037 14807
rect 15988 14776 16037 14804
rect 15988 14764 15994 14776
rect 16025 14773 16037 14776
rect 16071 14804 16083 14807
rect 16482 14804 16488 14816
rect 16071 14776 16488 14804
rect 16071 14773 16083 14776
rect 16025 14767 16083 14773
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 17402 14764 17408 14816
rect 17460 14804 17466 14816
rect 20714 14804 20720 14816
rect 17460 14776 20720 14804
rect 17460 14764 17466 14776
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 20898 14764 20904 14816
rect 20956 14804 20962 14816
rect 22465 14807 22523 14813
rect 22465 14804 22477 14807
rect 20956 14776 22477 14804
rect 20956 14764 20962 14776
rect 22465 14773 22477 14776
rect 22511 14773 22523 14807
rect 22465 14767 22523 14773
rect 22554 14764 22560 14816
rect 22612 14804 22618 14816
rect 23934 14804 23940 14816
rect 22612 14776 23940 14804
rect 22612 14764 22618 14776
rect 23934 14764 23940 14776
rect 23992 14804 23998 14816
rect 27816 14804 27844 14844
rect 29178 14832 29184 14844
rect 29236 14832 29242 14884
rect 30285 14875 30343 14881
rect 30285 14841 30297 14875
rect 30331 14872 30343 14875
rect 31021 14875 31079 14881
rect 31021 14872 31033 14875
rect 30331 14844 31033 14872
rect 30331 14841 30343 14844
rect 30285 14835 30343 14841
rect 31021 14841 31033 14844
rect 31067 14841 31079 14875
rect 31128 14872 31156 14912
rect 31662 14900 31668 14912
rect 31720 14900 31726 14952
rect 33686 14940 33692 14952
rect 33647 14912 33692 14940
rect 33686 14900 33692 14912
rect 33744 14900 33750 14952
rect 34698 14940 34704 14952
rect 34659 14912 34704 14940
rect 34698 14900 34704 14912
rect 34756 14900 34762 14952
rect 35529 14943 35587 14949
rect 35529 14909 35541 14943
rect 35575 14909 35587 14943
rect 38764 14940 38792 14980
rect 38841 14977 38853 15011
rect 38887 14977 38899 15011
rect 39482 15008 39488 15020
rect 39443 14980 39488 15008
rect 38841 14971 38899 14977
rect 39482 14968 39488 14980
rect 39540 14968 39546 15020
rect 39868 15017 39896 15116
rect 41309 15113 41321 15147
rect 41309 15107 41328 15113
rect 41322 15104 41328 15107
rect 41380 15104 41386 15156
rect 43162 15144 43168 15156
rect 43123 15116 43168 15144
rect 43162 15104 43168 15116
rect 43220 15104 43226 15156
rect 53558 15144 53564 15156
rect 53519 15116 53564 15144
rect 53558 15104 53564 15116
rect 53616 15104 53622 15156
rect 54202 15144 54208 15156
rect 54163 15116 54208 15144
rect 54202 15104 54208 15116
rect 54260 15104 54266 15156
rect 41509 15079 41567 15085
rect 41509 15045 41521 15079
rect 41555 15076 41567 15079
rect 41874 15076 41880 15088
rect 41555 15048 41880 15076
rect 41555 15045 41567 15048
rect 41509 15039 41567 15045
rect 41874 15036 41880 15048
rect 41932 15036 41938 15088
rect 42058 15036 42064 15088
rect 42116 15076 42122 15088
rect 42518 15076 42524 15088
rect 42116 15048 42524 15076
rect 42116 15036 42122 15048
rect 42518 15036 42524 15048
rect 42576 15076 42582 15088
rect 43438 15076 43444 15088
rect 42576 15048 43444 15076
rect 42576 15036 42582 15048
rect 43438 15036 43444 15048
rect 43496 15036 43502 15088
rect 39577 15011 39635 15017
rect 39577 14977 39589 15011
rect 39623 14977 39635 15011
rect 39577 14971 39635 14977
rect 39853 15011 39911 15017
rect 39853 14977 39865 15011
rect 39899 14977 39911 15011
rect 40494 15008 40500 15020
rect 40455 14980 40500 15008
rect 39853 14971 39911 14977
rect 39592 14940 39620 14971
rect 40494 14968 40500 14980
rect 40552 14968 40558 15020
rect 40681 15011 40739 15017
rect 40681 14977 40693 15011
rect 40727 15008 40739 15011
rect 43346 15008 43352 15020
rect 40727 14980 43352 15008
rect 40727 14977 40739 14980
rect 40681 14971 40739 14977
rect 43346 14968 43352 14980
rect 43404 14968 43410 15020
rect 54018 15008 54024 15020
rect 53979 14980 54024 15008
rect 54018 14968 54024 14980
rect 54076 14968 54082 15020
rect 40034 14940 40040 14952
rect 38764 14912 39528 14940
rect 39592 14912 40040 14940
rect 35529 14903 35587 14909
rect 32674 14872 32680 14884
rect 31128 14844 32680 14872
rect 31021 14835 31079 14841
rect 32674 14832 32680 14844
rect 32732 14832 32738 14884
rect 33870 14832 33876 14884
rect 33928 14872 33934 14884
rect 35544 14872 35572 14903
rect 37458 14872 37464 14884
rect 33928 14844 37320 14872
rect 37419 14844 37464 14872
rect 33928 14832 33934 14844
rect 28166 14804 28172 14816
rect 23992 14776 27844 14804
rect 28127 14776 28172 14804
rect 23992 14764 23998 14776
rect 28166 14764 28172 14776
rect 28224 14764 28230 14816
rect 30098 14804 30104 14816
rect 30059 14776 30104 14804
rect 30098 14764 30104 14776
rect 30156 14764 30162 14816
rect 32309 14807 32367 14813
rect 32309 14773 32321 14807
rect 32355 14804 32367 14807
rect 33502 14804 33508 14816
rect 32355 14776 33508 14804
rect 32355 14773 32367 14776
rect 32309 14767 32367 14773
rect 33502 14764 33508 14776
rect 33560 14764 33566 14816
rect 33778 14764 33784 14816
rect 33836 14804 33842 14816
rect 35345 14807 35403 14813
rect 35345 14804 35357 14807
rect 33836 14776 35357 14804
rect 33836 14764 33842 14776
rect 35345 14773 35357 14776
rect 35391 14773 35403 14807
rect 35345 14767 35403 14773
rect 36541 14807 36599 14813
rect 36541 14773 36553 14807
rect 36587 14804 36599 14807
rect 37090 14804 37096 14816
rect 36587 14776 37096 14804
rect 36587 14773 36599 14776
rect 36541 14767 36599 14773
rect 37090 14764 37096 14776
rect 37148 14764 37154 14816
rect 37292 14804 37320 14844
rect 37458 14832 37464 14844
rect 37516 14832 37522 14884
rect 39500 14872 39528 14912
rect 40034 14900 40040 14912
rect 40092 14900 40098 14952
rect 40218 14900 40224 14952
rect 40276 14940 40282 14952
rect 40313 14943 40371 14949
rect 40313 14940 40325 14943
rect 40276 14912 40325 14940
rect 40276 14900 40282 14912
rect 40313 14909 40325 14912
rect 40359 14909 40371 14943
rect 40313 14903 40371 14909
rect 40402 14900 40408 14952
rect 40460 14940 40466 14952
rect 42610 14940 42616 14952
rect 40460 14912 42616 14940
rect 40460 14900 40466 14912
rect 41690 14872 41696 14884
rect 39500 14844 41696 14872
rect 41690 14832 41696 14844
rect 41748 14832 41754 14884
rect 39114 14804 39120 14816
rect 37292 14776 39120 14804
rect 39114 14764 39120 14776
rect 39172 14764 39178 14816
rect 39298 14804 39304 14816
rect 39259 14776 39304 14804
rect 39298 14764 39304 14776
rect 39356 14764 39362 14816
rect 39390 14764 39396 14816
rect 39448 14804 39454 14816
rect 40218 14804 40224 14816
rect 39448 14776 40224 14804
rect 39448 14764 39454 14776
rect 40218 14764 40224 14776
rect 40276 14764 40282 14816
rect 41046 14764 41052 14816
rect 41104 14804 41110 14816
rect 41141 14807 41199 14813
rect 41141 14804 41153 14807
rect 41104 14776 41153 14804
rect 41104 14764 41110 14776
rect 41141 14773 41153 14776
rect 41187 14773 41199 14807
rect 41141 14767 41199 14773
rect 41325 14807 41383 14813
rect 41325 14773 41337 14807
rect 41371 14804 41383 14807
rect 41800 14804 41828 14912
rect 42610 14900 42616 14912
rect 42668 14900 42674 14952
rect 41874 14832 41880 14884
rect 41932 14872 41938 14884
rect 42058 14872 42064 14884
rect 41932 14844 42064 14872
rect 41932 14832 41938 14844
rect 42058 14832 42064 14844
rect 42116 14872 42122 14884
rect 42116 14844 44956 14872
rect 42116 14832 42122 14844
rect 41966 14804 41972 14816
rect 41371 14776 41828 14804
rect 41927 14776 41972 14804
rect 41371 14773 41383 14776
rect 41325 14767 41383 14773
rect 41966 14764 41972 14776
rect 42024 14764 42030 14816
rect 42610 14804 42616 14816
rect 42571 14776 42616 14804
rect 42610 14764 42616 14776
rect 42668 14764 42674 14816
rect 43254 14764 43260 14816
rect 43312 14804 43318 14816
rect 43717 14807 43775 14813
rect 43717 14804 43729 14807
rect 43312 14776 43729 14804
rect 43312 14764 43318 14776
rect 43717 14773 43729 14776
rect 43763 14773 43775 14807
rect 44266 14804 44272 14816
rect 44227 14776 44272 14804
rect 43717 14767 43775 14773
rect 44266 14764 44272 14776
rect 44324 14764 44330 14816
rect 44928 14813 44956 14844
rect 44913 14807 44971 14813
rect 44913 14773 44925 14807
rect 44959 14804 44971 14807
rect 53742 14804 53748 14816
rect 44959 14776 53748 14804
rect 44959 14773 44971 14776
rect 44913 14767 44971 14773
rect 53742 14764 53748 14776
rect 53800 14764 53806 14816
rect 1104 14714 54832 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 54832 14714
rect 1104 14640 54832 14662
rect 15102 14600 15108 14612
rect 15063 14572 15108 14600
rect 15102 14560 15108 14572
rect 15160 14560 15166 14612
rect 15562 14600 15568 14612
rect 15523 14572 15568 14600
rect 15562 14560 15568 14572
rect 15620 14560 15626 14612
rect 16574 14600 16580 14612
rect 15948 14572 16436 14600
rect 16535 14572 16580 14600
rect 13725 14535 13783 14541
rect 13725 14501 13737 14535
rect 13771 14532 13783 14535
rect 15948 14532 15976 14572
rect 13771 14504 15976 14532
rect 16408 14532 16436 14572
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 17681 14603 17739 14609
rect 17681 14569 17693 14603
rect 17727 14600 17739 14603
rect 18414 14600 18420 14612
rect 17727 14572 18420 14600
rect 17727 14569 17739 14572
rect 17681 14563 17739 14569
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 19444 14572 20484 14600
rect 19444 14532 19472 14572
rect 16408 14504 19472 14532
rect 13771 14501 13783 14504
rect 13725 14495 13783 14501
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 11698 14464 11704 14476
rect 4672 14436 11704 14464
rect 4672 14424 4678 14436
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 14553 14467 14611 14473
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 14734 14464 14740 14476
rect 14599 14436 14740 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 14734 14424 14740 14436
rect 14792 14464 14798 14476
rect 15102 14464 15108 14476
rect 14792 14436 15108 14464
rect 14792 14424 14798 14436
rect 15102 14424 15108 14436
rect 15160 14424 15166 14476
rect 15470 14424 15476 14476
rect 15528 14464 15534 14476
rect 15841 14467 15899 14473
rect 15841 14464 15853 14467
rect 15528 14436 15853 14464
rect 15528 14424 15534 14436
rect 15841 14433 15853 14436
rect 15887 14433 15899 14467
rect 15841 14427 15899 14433
rect 15933 14467 15991 14473
rect 15933 14433 15945 14467
rect 15979 14464 15991 14467
rect 15979 14436 16436 14464
rect 15979 14433 15991 14436
rect 15933 14427 15991 14433
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14396 1915 14399
rect 15654 14396 15660 14408
rect 1903 14368 15660 14396
rect 1903 14365 1915 14368
rect 1857 14359 1915 14365
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14365 15807 14399
rect 16022 14396 16028 14408
rect 15983 14368 16028 14396
rect 15749 14359 15807 14365
rect 4338 14288 4344 14340
rect 4396 14328 4402 14340
rect 15562 14328 15568 14340
rect 4396 14300 15568 14328
rect 4396 14288 4402 14300
rect 15562 14288 15568 14300
rect 15620 14288 15626 14340
rect 1670 14260 1676 14272
rect 1631 14232 1676 14260
rect 1670 14220 1676 14232
rect 1728 14220 1734 14272
rect 12621 14263 12679 14269
rect 12621 14229 12633 14263
rect 12667 14260 12679 14263
rect 13170 14260 13176 14272
rect 12667 14232 13176 14260
rect 12667 14229 12679 14232
rect 12621 14223 12679 14229
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 14918 14220 14924 14272
rect 14976 14260 14982 14272
rect 15470 14260 15476 14272
rect 14976 14232 15476 14260
rect 14976 14220 14982 14232
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 15764 14260 15792 14359
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16408 14328 16436 14436
rect 16482 14424 16488 14476
rect 16540 14464 16546 14476
rect 16761 14467 16819 14473
rect 16761 14464 16773 14467
rect 16540 14436 16773 14464
rect 16540 14424 16546 14436
rect 16761 14433 16773 14436
rect 16807 14433 16819 14467
rect 17402 14464 17408 14476
rect 16761 14427 16819 14433
rect 16868 14436 17408 14464
rect 16868 14405 16896 14436
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 18782 14464 18788 14476
rect 18743 14436 18788 14464
rect 18782 14424 18788 14436
rect 18840 14424 18846 14476
rect 16853 14399 16911 14405
rect 16853 14365 16865 14399
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14396 17095 14399
rect 17678 14396 17684 14408
rect 17083 14368 17684 14396
rect 17083 14365 17095 14368
rect 17037 14359 17095 14365
rect 16574 14328 16580 14340
rect 16408 14300 16580 14328
rect 16574 14288 16580 14300
rect 16632 14328 16638 14340
rect 16960 14328 16988 14359
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 17862 14356 17868 14408
rect 17920 14396 17926 14408
rect 19426 14396 19432 14408
rect 17920 14368 18736 14396
rect 19339 14368 19432 14396
rect 17920 14356 17926 14368
rect 17126 14328 17132 14340
rect 16632 14300 17132 14328
rect 16632 14288 16638 14300
rect 17126 14288 17132 14300
rect 17184 14288 17190 14340
rect 17954 14288 17960 14340
rect 18012 14328 18018 14340
rect 18601 14331 18659 14337
rect 18601 14328 18613 14331
rect 18012 14300 18613 14328
rect 18012 14288 18018 14300
rect 18601 14297 18613 14300
rect 18647 14297 18659 14331
rect 18708 14328 18736 14368
rect 19426 14356 19432 14368
rect 19484 14396 19490 14408
rect 20070 14396 20076 14408
rect 19484 14368 20076 14396
rect 19484 14356 19490 14368
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 20456 14396 20484 14572
rect 20714 14560 20720 14612
rect 20772 14600 20778 14612
rect 20772 14572 23704 14600
rect 20772 14560 20778 14572
rect 23676 14532 23704 14572
rect 23750 14560 23756 14612
rect 23808 14600 23814 14612
rect 23937 14603 23995 14609
rect 23937 14600 23949 14603
rect 23808 14572 23949 14600
rect 23808 14560 23814 14572
rect 23937 14569 23949 14572
rect 23983 14600 23995 14603
rect 25225 14603 25283 14609
rect 25225 14600 25237 14603
rect 23983 14572 25237 14600
rect 23983 14569 23995 14572
rect 23937 14563 23995 14569
rect 25225 14569 25237 14572
rect 25271 14600 25283 14603
rect 27798 14600 27804 14612
rect 25271 14572 27804 14600
rect 25271 14569 25283 14572
rect 25225 14563 25283 14569
rect 27798 14560 27804 14572
rect 27856 14560 27862 14612
rect 28166 14560 28172 14612
rect 28224 14600 28230 14612
rect 31662 14600 31668 14612
rect 28224 14572 30788 14600
rect 31623 14572 31668 14600
rect 28224 14560 28230 14572
rect 28077 14535 28135 14541
rect 23676 14504 24164 14532
rect 24136 14476 24164 14504
rect 28077 14501 28089 14535
rect 28123 14532 28135 14535
rect 28902 14532 28908 14544
rect 28123 14504 28908 14532
rect 28123 14501 28135 14504
rect 28077 14495 28135 14501
rect 28902 14492 28908 14504
rect 28960 14492 28966 14544
rect 30760 14532 30788 14572
rect 31662 14560 31668 14572
rect 31720 14560 31726 14612
rect 33137 14603 33195 14609
rect 33137 14569 33149 14603
rect 33183 14600 33195 14603
rect 34698 14600 34704 14612
rect 33183 14572 34704 14600
rect 33183 14569 33195 14572
rect 33137 14563 33195 14569
rect 34698 14560 34704 14572
rect 34756 14560 34762 14612
rect 37001 14603 37059 14609
rect 37001 14600 37013 14603
rect 34808 14572 37013 14600
rect 34808 14532 34836 14572
rect 37001 14569 37013 14572
rect 37047 14569 37059 14603
rect 37001 14563 37059 14569
rect 37553 14603 37611 14609
rect 37553 14569 37565 14603
rect 37599 14600 37611 14603
rect 41506 14600 41512 14612
rect 37599 14572 41512 14600
rect 37599 14569 37611 14572
rect 37553 14563 37611 14569
rect 41506 14560 41512 14572
rect 41564 14560 41570 14612
rect 43073 14603 43131 14609
rect 43073 14569 43085 14603
rect 43119 14600 43131 14603
rect 43438 14600 43444 14612
rect 43119 14572 43444 14600
rect 43119 14569 43131 14572
rect 43073 14563 43131 14569
rect 43438 14560 43444 14572
rect 43496 14560 43502 14612
rect 30760 14504 34836 14532
rect 37826 14492 37832 14544
rect 37884 14532 37890 14544
rect 38930 14532 38936 14544
rect 37884 14504 38936 14532
rect 37884 14492 37890 14504
rect 38930 14492 38936 14504
rect 38988 14492 38994 14544
rect 39206 14492 39212 14544
rect 39264 14492 39270 14544
rect 39298 14492 39304 14544
rect 39356 14492 39362 14544
rect 54202 14532 54208 14544
rect 54163 14504 54208 14532
rect 54202 14492 54208 14504
rect 54260 14492 54266 14544
rect 21174 14424 21180 14476
rect 21232 14464 21238 14476
rect 21821 14467 21879 14473
rect 21821 14464 21833 14467
rect 21232 14436 21833 14464
rect 21232 14424 21238 14436
rect 21821 14433 21833 14436
rect 21867 14433 21879 14467
rect 21821 14427 21879 14433
rect 22278 14424 22284 14476
rect 22336 14464 22342 14476
rect 22557 14467 22615 14473
rect 22557 14464 22569 14467
rect 22336 14436 22569 14464
rect 22336 14424 22342 14436
rect 22557 14433 22569 14436
rect 22603 14433 22615 14467
rect 22557 14427 22615 14433
rect 24118 14424 24124 14476
rect 24176 14464 24182 14476
rect 24302 14464 24308 14476
rect 24176 14436 24308 14464
rect 24176 14424 24182 14436
rect 24302 14424 24308 14436
rect 24360 14464 24366 14476
rect 26605 14467 26663 14473
rect 24360 14436 24808 14464
rect 24360 14424 24366 14436
rect 21634 14396 21640 14408
rect 20456 14368 21640 14396
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 24210 14356 24216 14408
rect 24268 14396 24274 14408
rect 24780 14405 24808 14436
rect 26605 14433 26617 14467
rect 26651 14464 26663 14467
rect 29270 14464 29276 14476
rect 26651 14436 29276 14464
rect 26651 14433 26663 14436
rect 26605 14427 26663 14433
rect 29270 14424 29276 14436
rect 29328 14464 29334 14476
rect 29822 14464 29828 14476
rect 29328 14436 29828 14464
rect 29328 14424 29334 14436
rect 29822 14424 29828 14436
rect 29880 14424 29886 14476
rect 31294 14424 31300 14476
rect 31352 14464 31358 14476
rect 31754 14464 31760 14476
rect 31352 14436 31760 14464
rect 31352 14424 31358 14436
rect 31754 14424 31760 14436
rect 31812 14464 31818 14476
rect 31941 14467 31999 14473
rect 31941 14464 31953 14467
rect 31812 14436 31953 14464
rect 31812 14424 31818 14436
rect 31941 14433 31953 14436
rect 31987 14433 31999 14467
rect 31941 14427 31999 14433
rect 32030 14424 32036 14476
rect 32088 14464 32094 14476
rect 32950 14464 32956 14476
rect 32088 14436 32444 14464
rect 32911 14436 32956 14464
rect 32088 14424 32094 14436
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 24268 14368 24593 14396
rect 24268 14356 24274 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 24765 14399 24823 14405
rect 24765 14365 24777 14399
rect 24811 14365 24823 14399
rect 27246 14396 27252 14408
rect 24765 14359 24823 14365
rect 26160 14368 27252 14396
rect 19674 14331 19732 14337
rect 19674 14328 19686 14331
rect 18708 14300 19686 14328
rect 18601 14291 18659 14297
rect 19674 14297 19686 14300
rect 19720 14297 19732 14331
rect 19674 14291 19732 14297
rect 20714 14288 20720 14340
rect 20772 14328 20778 14340
rect 22802 14331 22860 14337
rect 22802 14328 22814 14331
rect 20772 14300 22814 14328
rect 20772 14288 20778 14300
rect 22802 14297 22814 14300
rect 22848 14297 22860 14331
rect 22802 14291 22860 14297
rect 24673 14331 24731 14337
rect 24673 14297 24685 14331
rect 24719 14328 24731 14331
rect 26160 14328 26188 14368
rect 27246 14356 27252 14368
rect 27304 14396 27310 14408
rect 27525 14399 27583 14405
rect 27525 14396 27537 14399
rect 27304 14368 27537 14396
rect 27304 14356 27310 14368
rect 27525 14365 27537 14368
rect 27571 14365 27583 14399
rect 27706 14396 27712 14408
rect 27667 14368 27712 14396
rect 27525 14359 27583 14365
rect 27706 14356 27712 14368
rect 27764 14356 27770 14408
rect 27893 14399 27951 14405
rect 27893 14365 27905 14399
rect 27939 14396 27951 14399
rect 28534 14396 28540 14408
rect 27939 14368 28540 14396
rect 27939 14365 27951 14368
rect 27893 14359 27951 14365
rect 28534 14356 28540 14368
rect 28592 14356 28598 14408
rect 28905 14399 28963 14405
rect 28905 14365 28917 14399
rect 28951 14396 28963 14399
rect 29086 14396 29092 14408
rect 28951 14368 29092 14396
rect 28951 14365 28963 14368
rect 28905 14359 28963 14365
rect 24719 14300 26188 14328
rect 24719 14297 24731 14300
rect 24673 14291 24731 14297
rect 26234 14288 26240 14340
rect 26292 14328 26298 14340
rect 26338 14331 26396 14337
rect 26338 14328 26350 14331
rect 26292 14300 26350 14328
rect 26292 14288 26298 14300
rect 26338 14297 26350 14300
rect 26384 14297 26396 14331
rect 26338 14291 26396 14297
rect 26602 14288 26608 14340
rect 26660 14328 26666 14340
rect 27801 14331 27859 14337
rect 27801 14328 27813 14331
rect 26660 14300 27813 14328
rect 26660 14288 26666 14300
rect 27801 14297 27813 14300
rect 27847 14297 27859 14331
rect 27801 14291 27859 14297
rect 28442 14288 28448 14340
rect 28500 14328 28506 14340
rect 28920 14328 28948 14359
rect 29086 14356 29092 14368
rect 29144 14396 29150 14408
rect 29914 14396 29920 14408
rect 29144 14368 29920 14396
rect 29144 14356 29150 14368
rect 29914 14356 29920 14368
rect 29972 14356 29978 14408
rect 30926 14356 30932 14408
rect 30984 14396 30990 14408
rect 31849 14399 31907 14405
rect 31849 14396 31861 14399
rect 30984 14368 31861 14396
rect 30984 14356 30990 14368
rect 31849 14365 31861 14368
rect 31895 14365 31907 14399
rect 31849 14359 31907 14365
rect 28500 14300 28948 14328
rect 28500 14288 28506 14300
rect 29178 14288 29184 14340
rect 29236 14328 29242 14340
rect 30070 14331 30128 14337
rect 30070 14328 30082 14331
rect 29236 14300 30082 14328
rect 29236 14288 29242 14300
rect 30070 14297 30082 14300
rect 30116 14297 30128 14331
rect 31864 14328 31892 14359
rect 32122 14356 32128 14408
rect 32180 14396 32186 14408
rect 32416 14396 32444 14436
rect 32950 14424 32956 14436
rect 33008 14424 33014 14476
rect 33778 14464 33784 14476
rect 33739 14436 33784 14464
rect 33778 14424 33784 14436
rect 33836 14424 33842 14476
rect 39022 14464 39028 14476
rect 38212 14436 39028 14464
rect 32858 14396 32864 14408
rect 32180 14368 32225 14396
rect 32416 14368 32864 14396
rect 32180 14356 32186 14368
rect 32858 14356 32864 14368
rect 32916 14356 32922 14408
rect 33594 14356 33600 14408
rect 33652 14396 33658 14408
rect 36262 14396 36268 14408
rect 33652 14368 36124 14396
rect 36223 14368 36268 14396
rect 33652 14356 33658 14368
rect 34238 14328 34244 14340
rect 31864 14300 34244 14328
rect 30070 14291 30128 14297
rect 34238 14288 34244 14300
rect 34296 14288 34302 14340
rect 34606 14288 34612 14340
rect 34664 14328 34670 14340
rect 35250 14328 35256 14340
rect 34664 14300 35256 14328
rect 34664 14288 34670 14300
rect 35250 14288 35256 14300
rect 35308 14288 35314 14340
rect 35894 14288 35900 14340
rect 35952 14328 35958 14340
rect 35998 14331 36056 14337
rect 35998 14328 36010 14331
rect 35952 14300 36010 14328
rect 35952 14288 35958 14300
rect 35998 14297 36010 14300
rect 36044 14297 36056 14331
rect 36096 14328 36124 14368
rect 36262 14356 36268 14368
rect 36320 14356 36326 14408
rect 36909 14399 36967 14405
rect 36909 14365 36921 14399
rect 36955 14396 36967 14399
rect 37090 14396 37096 14408
rect 36955 14368 37096 14396
rect 36955 14365 36967 14368
rect 36909 14359 36967 14365
rect 37090 14356 37096 14368
rect 37148 14356 37154 14408
rect 37458 14405 37464 14408
rect 37428 14399 37464 14405
rect 37428 14365 37440 14399
rect 37428 14359 37464 14365
rect 37458 14356 37464 14359
rect 37516 14356 37522 14408
rect 38212 14405 38240 14436
rect 39022 14424 39028 14436
rect 39080 14424 39086 14476
rect 38197 14399 38255 14405
rect 38197 14365 38209 14399
rect 38243 14365 38255 14399
rect 38197 14359 38255 14365
rect 38286 14356 38292 14408
rect 38344 14396 38350 14408
rect 39117 14399 39175 14405
rect 38344 14368 38389 14396
rect 38344 14356 38350 14368
rect 39117 14365 39129 14399
rect 39163 14396 39175 14399
rect 39224 14396 39252 14492
rect 39163 14368 39252 14396
rect 39316 14405 39344 14492
rect 41340 14436 44404 14464
rect 41340 14408 41368 14436
rect 39316 14399 39379 14405
rect 39316 14368 39333 14399
rect 39163 14365 39175 14368
rect 39117 14359 39175 14365
rect 39321 14365 39333 14368
rect 39367 14365 39379 14399
rect 39321 14359 39379 14365
rect 40218 14356 40224 14408
rect 40276 14396 40282 14408
rect 41322 14396 41328 14408
rect 40276 14368 41328 14396
rect 40276 14356 40282 14368
rect 41322 14356 41328 14368
rect 41380 14356 41386 14408
rect 41414 14356 41420 14408
rect 41472 14396 41478 14408
rect 42702 14396 42708 14408
rect 41472 14368 42708 14396
rect 41472 14356 41478 14368
rect 42702 14356 42708 14368
rect 42760 14396 42766 14408
rect 43533 14399 43591 14405
rect 43533 14396 43545 14399
rect 42760 14368 43545 14396
rect 42760 14356 42766 14368
rect 43533 14365 43545 14368
rect 43579 14396 43591 14399
rect 44266 14396 44272 14408
rect 43579 14368 44272 14396
rect 43579 14365 43591 14368
rect 43533 14359 43591 14365
rect 44266 14356 44272 14368
rect 44324 14356 44330 14408
rect 38746 14328 38752 14340
rect 36096 14300 38752 14328
rect 35998 14291 36056 14297
rect 38746 14288 38752 14300
rect 38804 14288 38810 14340
rect 39485 14331 39543 14337
rect 39485 14297 39497 14331
rect 39531 14328 39543 14331
rect 40678 14328 40684 14340
rect 39531 14300 40684 14328
rect 39531 14297 39543 14300
rect 39485 14291 39543 14297
rect 40678 14288 40684 14300
rect 40736 14288 40742 14340
rect 40770 14288 40776 14340
rect 40828 14328 40834 14340
rect 41150 14331 41208 14337
rect 41150 14328 41162 14331
rect 40828 14300 41162 14328
rect 40828 14288 40834 14300
rect 41150 14297 41162 14300
rect 41196 14297 41208 14331
rect 41150 14291 41208 14297
rect 41506 14288 41512 14340
rect 41564 14328 41570 14340
rect 41877 14331 41935 14337
rect 41877 14328 41889 14331
rect 41564 14300 41889 14328
rect 41564 14288 41570 14300
rect 41877 14297 41889 14300
rect 41923 14328 41935 14331
rect 42429 14331 42487 14337
rect 42429 14328 42441 14331
rect 41923 14300 42441 14328
rect 41923 14297 41935 14300
rect 41877 14291 41935 14297
rect 42429 14297 42441 14300
rect 42475 14328 42487 14331
rect 42610 14328 42616 14340
rect 42475 14300 42616 14328
rect 42475 14297 42487 14300
rect 42429 14291 42487 14297
rect 42610 14288 42616 14300
rect 42668 14288 42674 14340
rect 15930 14260 15936 14272
rect 15764 14232 15936 14260
rect 15930 14220 15936 14232
rect 15988 14220 15994 14272
rect 18138 14260 18144 14272
rect 18099 14232 18144 14260
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 18509 14263 18567 14269
rect 18509 14229 18521 14263
rect 18555 14260 18567 14263
rect 18690 14260 18696 14272
rect 18555 14232 18696 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 20806 14260 20812 14272
rect 20767 14232 20812 14260
rect 20806 14220 20812 14232
rect 20864 14220 20870 14272
rect 21266 14260 21272 14272
rect 21227 14232 21272 14260
rect 21266 14220 21272 14232
rect 21324 14220 21330 14272
rect 21726 14260 21732 14272
rect 21687 14232 21732 14260
rect 21726 14220 21732 14232
rect 21784 14220 21790 14272
rect 21818 14220 21824 14272
rect 21876 14260 21882 14272
rect 25498 14260 25504 14272
rect 21876 14232 25504 14260
rect 21876 14220 21882 14232
rect 25498 14220 25504 14232
rect 25556 14220 25562 14272
rect 28534 14220 28540 14272
rect 28592 14260 28598 14272
rect 29089 14263 29147 14269
rect 29089 14260 29101 14263
rect 28592 14232 29101 14260
rect 28592 14220 28598 14232
rect 29089 14229 29101 14232
rect 29135 14260 29147 14263
rect 30742 14260 30748 14272
rect 29135 14232 30748 14260
rect 29135 14229 29147 14232
rect 29089 14223 29147 14229
rect 30742 14220 30748 14232
rect 30800 14220 30806 14272
rect 31202 14260 31208 14272
rect 31163 14232 31208 14260
rect 31202 14220 31208 14232
rect 31260 14220 31266 14272
rect 32674 14220 32680 14272
rect 32732 14260 32738 14272
rect 33594 14260 33600 14272
rect 32732 14232 33600 14260
rect 32732 14220 32738 14232
rect 33594 14220 33600 14232
rect 33652 14220 33658 14272
rect 34333 14263 34391 14269
rect 34333 14229 34345 14263
rect 34379 14260 34391 14263
rect 34422 14260 34428 14272
rect 34379 14232 34428 14260
rect 34379 14229 34391 14232
rect 34333 14223 34391 14229
rect 34422 14220 34428 14232
rect 34480 14220 34486 14272
rect 34885 14263 34943 14269
rect 34885 14229 34897 14263
rect 34931 14260 34943 14263
rect 35342 14260 35348 14272
rect 34931 14232 35348 14260
rect 34931 14229 34943 14232
rect 34885 14223 34943 14229
rect 35342 14220 35348 14232
rect 35400 14220 35406 14272
rect 37366 14260 37372 14272
rect 37327 14232 37372 14260
rect 37366 14220 37372 14232
rect 37424 14220 37430 14272
rect 38289 14263 38347 14269
rect 38289 14229 38301 14263
rect 38335 14260 38347 14263
rect 38378 14260 38384 14272
rect 38335 14232 38384 14260
rect 38335 14229 38347 14232
rect 38289 14223 38347 14229
rect 38378 14220 38384 14232
rect 38436 14220 38442 14272
rect 39114 14220 39120 14272
rect 39172 14260 39178 14272
rect 39850 14260 39856 14272
rect 39172 14232 39856 14260
rect 39172 14220 39178 14232
rect 39850 14220 39856 14232
rect 39908 14220 39914 14272
rect 40034 14220 40040 14272
rect 40092 14260 40098 14272
rect 43898 14260 43904 14272
rect 40092 14232 43904 14260
rect 40092 14220 40098 14232
rect 43898 14220 43904 14232
rect 43956 14220 43962 14272
rect 44177 14263 44235 14269
rect 44177 14229 44189 14263
rect 44223 14260 44235 14263
rect 44376 14260 44404 14436
rect 54018 14396 54024 14408
rect 53979 14368 54024 14396
rect 54018 14356 54024 14368
rect 54076 14356 54082 14408
rect 49050 14260 49056 14272
rect 44223 14232 49056 14260
rect 44223 14229 44235 14232
rect 44177 14223 44235 14229
rect 49050 14220 49056 14232
rect 49108 14220 49114 14272
rect 53561 14263 53619 14269
rect 53561 14229 53573 14263
rect 53607 14260 53619 14263
rect 54202 14260 54208 14272
rect 53607 14232 54208 14260
rect 53607 14229 53619 14232
rect 53561 14223 53619 14229
rect 54202 14220 54208 14232
rect 54260 14220 54266 14272
rect 1104 14170 54832 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 54832 14170
rect 1104 14096 54832 14118
rect 13909 14059 13967 14065
rect 13909 14025 13921 14059
rect 13955 14056 13967 14059
rect 13998 14056 14004 14068
rect 13955 14028 14004 14056
rect 13955 14025 13967 14028
rect 13909 14019 13967 14025
rect 13998 14016 14004 14028
rect 14056 14056 14062 14068
rect 15010 14056 15016 14068
rect 14056 14028 15016 14056
rect 14056 14016 14062 14028
rect 15010 14016 15016 14028
rect 15068 14016 15074 14068
rect 17586 14056 17592 14068
rect 15764 14028 17592 14056
rect 13357 13991 13415 13997
rect 13357 13957 13369 13991
rect 13403 13988 13415 13991
rect 14458 13988 14464 14000
rect 13403 13960 14464 13988
rect 13403 13957 13415 13960
rect 13357 13951 13415 13957
rect 14458 13948 14464 13960
rect 14516 13948 14522 14000
rect 14550 13948 14556 14000
rect 14608 13988 14614 14000
rect 15102 13988 15108 14000
rect 14608 13960 15108 13988
rect 14608 13948 14614 13960
rect 15102 13948 15108 13960
rect 15160 13948 15166 14000
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 4338 13920 4344 13932
rect 1903 13892 4344 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 14918 13920 14924 13932
rect 12299 13892 14924 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 14461 13855 14519 13861
rect 14461 13821 14473 13855
rect 14507 13852 14519 13855
rect 15764 13852 15792 14028
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 18322 14056 18328 14068
rect 18235 14028 18328 14056
rect 18322 14016 18328 14028
rect 18380 14056 18386 14068
rect 18598 14056 18604 14068
rect 18380 14028 18604 14056
rect 18380 14016 18386 14028
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 20257 14059 20315 14065
rect 20257 14025 20269 14059
rect 20303 14056 20315 14059
rect 21818 14056 21824 14068
rect 20303 14028 21824 14056
rect 20303 14025 20315 14028
rect 20257 14019 20315 14025
rect 21818 14016 21824 14028
rect 21876 14016 21882 14068
rect 23382 14056 23388 14068
rect 23343 14028 23388 14056
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 23750 14056 23756 14068
rect 23711 14028 23756 14056
rect 23750 14016 23756 14028
rect 23808 14016 23814 14068
rect 23845 14059 23903 14065
rect 23845 14025 23857 14059
rect 23891 14056 23903 14059
rect 23934 14056 23940 14068
rect 23891 14028 23940 14056
rect 23891 14025 23903 14028
rect 23845 14019 23903 14025
rect 23934 14016 23940 14028
rect 23992 14016 23998 14068
rect 29365 14059 29423 14065
rect 29365 14056 29377 14059
rect 24596 14028 29377 14056
rect 16868 13960 17246 13988
rect 16868 13932 16896 13960
rect 15838 13880 15844 13932
rect 15896 13920 15902 13932
rect 16117 13923 16175 13929
rect 15896 13892 16068 13920
rect 15896 13880 15902 13892
rect 15930 13852 15936 13864
rect 14507 13824 15792 13852
rect 15891 13824 15936 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 15930 13812 15936 13824
rect 15988 13812 15994 13864
rect 16040 13861 16068 13892
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16574 13920 16580 13932
rect 16163 13892 16580 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16574 13880 16580 13892
rect 16632 13920 16638 13932
rect 16850 13920 16856 13932
rect 16632 13892 16856 13920
rect 16632 13880 16638 13892
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 17218 13929 17246 13960
rect 18230 13948 18236 14000
rect 18288 13988 18294 14000
rect 21726 13988 21732 14000
rect 18288 13960 21732 13988
rect 18288 13948 18294 13960
rect 21726 13948 21732 13960
rect 21784 13948 21790 14000
rect 22094 13948 22100 14000
rect 22152 13988 22158 14000
rect 22465 13991 22523 13997
rect 22465 13988 22477 13991
rect 22152 13960 22477 13988
rect 22152 13948 22158 13960
rect 22465 13957 22477 13960
rect 22511 13957 22523 13991
rect 22465 13951 22523 13957
rect 22833 13991 22891 13997
rect 22833 13957 22845 13991
rect 22879 13988 22891 13991
rect 24596 13988 24624 14028
rect 29365 14025 29377 14028
rect 29411 14025 29423 14059
rect 31294 14056 31300 14068
rect 31255 14028 31300 14056
rect 29365 14019 29423 14025
rect 31294 14016 31300 14028
rect 31352 14016 31358 14068
rect 31389 14059 31447 14065
rect 31389 14025 31401 14059
rect 31435 14056 31447 14059
rect 32030 14056 32036 14068
rect 31435 14028 32036 14056
rect 31435 14025 31447 14028
rect 31389 14019 31447 14025
rect 32030 14016 32036 14028
rect 32088 14016 32094 14068
rect 35529 14059 35587 14065
rect 35529 14025 35541 14059
rect 35575 14056 35587 14059
rect 35802 14056 35808 14068
rect 35575 14028 35808 14056
rect 35575 14025 35587 14028
rect 35529 14019 35587 14025
rect 35802 14016 35808 14028
rect 35860 14016 35866 14068
rect 39942 14056 39948 14068
rect 38600 14028 39948 14056
rect 22879 13960 24624 13988
rect 22879 13957 22891 13960
rect 22833 13951 22891 13957
rect 24670 13948 24676 14000
rect 24728 13988 24734 14000
rect 29270 13988 29276 14000
rect 24728 13960 29276 13988
rect 24728 13948 24734 13960
rect 17212 13923 17270 13929
rect 17212 13889 17224 13923
rect 17258 13889 17270 13923
rect 17212 13883 17270 13889
rect 17586 13880 17592 13932
rect 17644 13920 17650 13932
rect 19438 13923 19496 13929
rect 19438 13920 19450 13923
rect 17644 13892 19450 13920
rect 17644 13880 17650 13892
rect 19438 13889 19450 13892
rect 19484 13889 19496 13923
rect 19438 13883 19496 13889
rect 19610 13880 19616 13932
rect 19668 13920 19674 13932
rect 20990 13920 20996 13932
rect 19668 13892 20996 13920
rect 19668 13880 19674 13892
rect 20990 13880 20996 13892
rect 21048 13920 21054 13932
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 21048 13892 21097 13920
rect 21048 13880 21054 13892
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13920 21235 13923
rect 21450 13920 21456 13932
rect 21223 13892 21456 13920
rect 21223 13889 21235 13892
rect 21177 13883 21235 13889
rect 21450 13880 21456 13892
rect 21508 13880 21514 13932
rect 24210 13880 24216 13932
rect 24268 13920 24274 13932
rect 25240 13929 25268 13960
rect 24581 13923 24639 13929
rect 24581 13920 24593 13923
rect 24268 13892 24593 13920
rect 24268 13880 24274 13892
rect 24581 13889 24593 13892
rect 24627 13889 24639 13923
rect 24581 13883 24639 13889
rect 24765 13923 24823 13929
rect 24765 13889 24777 13923
rect 24811 13889 24823 13923
rect 24765 13883 24823 13889
rect 25225 13923 25283 13929
rect 25225 13889 25237 13923
rect 25271 13889 25283 13923
rect 25225 13883 25283 13889
rect 25492 13923 25550 13929
rect 25492 13889 25504 13923
rect 25538 13920 25550 13923
rect 25774 13920 25780 13932
rect 25538 13892 25780 13920
rect 25538 13889 25550 13892
rect 25492 13883 25550 13889
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13821 16083 13855
rect 16025 13815 16083 13821
rect 16209 13855 16267 13861
rect 16209 13821 16221 13855
rect 16255 13852 16267 13855
rect 16390 13852 16396 13864
rect 16255 13824 16396 13852
rect 16255 13821 16267 13824
rect 16209 13815 16267 13821
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 17037 13855 17095 13861
rect 17037 13821 17049 13855
rect 17083 13821 17095 13855
rect 17037 13815 17095 13821
rect 15948 13784 15976 13812
rect 17052 13784 17080 13815
rect 17126 13812 17132 13864
rect 17184 13852 17190 13864
rect 17313 13855 17371 13861
rect 17184 13824 17229 13852
rect 17184 13812 17190 13824
rect 17313 13821 17325 13855
rect 17359 13852 17371 13855
rect 17402 13852 17408 13864
rect 17359 13824 17408 13852
rect 17359 13821 17371 13824
rect 17313 13815 17371 13821
rect 17402 13812 17408 13824
rect 17460 13812 17466 13864
rect 19705 13855 19763 13861
rect 19705 13821 19717 13855
rect 19751 13852 19763 13855
rect 20070 13852 20076 13864
rect 19751 13824 20076 13852
rect 19751 13821 19763 13824
rect 19705 13815 19763 13821
rect 20070 13812 20076 13824
rect 20128 13812 20134 13864
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13821 21327 13855
rect 21269 13815 21327 13821
rect 15948 13756 17080 13784
rect 19886 13744 19892 13796
rect 19944 13784 19950 13796
rect 20898 13784 20904 13796
rect 19944 13756 20904 13784
rect 19944 13744 19950 13756
rect 20898 13744 20904 13756
rect 20956 13744 20962 13796
rect 21174 13744 21180 13796
rect 21232 13784 21238 13796
rect 21284 13784 21312 13815
rect 23934 13812 23940 13864
rect 23992 13852 23998 13864
rect 23992 13824 24037 13852
rect 23992 13812 23998 13824
rect 24302 13812 24308 13864
rect 24360 13852 24366 13864
rect 24486 13852 24492 13864
rect 24360 13824 24492 13852
rect 24360 13812 24366 13824
rect 24486 13812 24492 13824
rect 24544 13852 24550 13864
rect 24780 13852 24808 13883
rect 25774 13880 25780 13892
rect 25832 13880 25838 13932
rect 26050 13880 26056 13932
rect 26108 13920 26114 13932
rect 26694 13920 26700 13932
rect 26108 13892 26700 13920
rect 26108 13880 26114 13892
rect 26694 13880 26700 13892
rect 26752 13880 26758 13932
rect 27706 13920 27712 13932
rect 27540 13892 27712 13920
rect 24544 13824 24808 13852
rect 24544 13812 24550 13824
rect 24762 13784 24768 13796
rect 21232 13756 21312 13784
rect 24723 13756 24768 13784
rect 21232 13744 21238 13756
rect 24762 13744 24768 13756
rect 24820 13744 24826 13796
rect 26602 13784 26608 13796
rect 26563 13756 26608 13784
rect 26602 13744 26608 13756
rect 26660 13744 26666 13796
rect 27540 13784 27568 13892
rect 27706 13880 27712 13892
rect 27764 13880 27770 13932
rect 27982 13880 27988 13932
rect 28040 13920 28046 13932
rect 28270 13923 28328 13929
rect 28270 13920 28282 13923
rect 28040 13892 28282 13920
rect 28040 13880 28046 13892
rect 28270 13889 28282 13892
rect 28316 13889 28328 13923
rect 28270 13883 28328 13889
rect 28537 13923 28595 13929
rect 28537 13889 28549 13923
rect 28583 13920 28595 13923
rect 28644 13920 28672 13960
rect 29270 13948 29276 13960
rect 29328 13948 29334 14000
rect 30466 13948 30472 14000
rect 30524 13988 30530 14000
rect 32309 13991 32367 13997
rect 32309 13988 32321 13991
rect 30524 13960 32321 13988
rect 30524 13948 30530 13960
rect 32309 13957 32321 13960
rect 32355 13957 32367 13991
rect 32309 13951 32367 13957
rect 33686 13948 33692 14000
rect 33744 13988 33750 14000
rect 38600 13997 38628 14028
rect 39942 14016 39948 14028
rect 40000 14016 40006 14068
rect 43254 14056 43260 14068
rect 43215 14028 43260 14056
rect 43254 14016 43260 14028
rect 43312 14016 43318 14068
rect 43806 14056 43812 14068
rect 43767 14028 43812 14056
rect 43806 14016 43812 14028
rect 43864 14016 43870 14068
rect 43898 14016 43904 14068
rect 43956 14056 43962 14068
rect 54018 14056 54024 14068
rect 43956 14028 54024 14056
rect 43956 14016 43962 14028
rect 54018 14016 54024 14028
rect 54076 14016 54082 14068
rect 38585 13991 38643 13997
rect 33744 13960 36308 13988
rect 33744 13948 33750 13960
rect 28583 13892 28672 13920
rect 28583 13889 28595 13892
rect 28537 13883 28595 13889
rect 29086 13880 29092 13932
rect 29144 13920 29150 13932
rect 29549 13923 29607 13929
rect 29549 13920 29561 13923
rect 29144 13892 29561 13920
rect 29144 13880 29150 13892
rect 29549 13889 29561 13892
rect 29595 13889 29607 13923
rect 30006 13920 30012 13932
rect 29967 13892 30012 13920
rect 29549 13883 29607 13889
rect 30006 13880 30012 13892
rect 30064 13880 30070 13932
rect 30926 13880 30932 13932
rect 30984 13920 30990 13932
rect 31205 13923 31263 13929
rect 31205 13920 31217 13923
rect 30984 13892 31217 13920
rect 30984 13880 30990 13892
rect 31205 13889 31217 13892
rect 31251 13889 31263 13923
rect 31205 13883 31263 13889
rect 31573 13923 31631 13929
rect 31573 13889 31585 13923
rect 31619 13920 31631 13923
rect 32122 13920 32128 13932
rect 31619 13892 32128 13920
rect 31619 13889 31631 13892
rect 31573 13883 31631 13889
rect 32122 13880 32128 13892
rect 32180 13880 32186 13932
rect 34164 13929 34192 13960
rect 36280 13932 36308 13960
rect 38585 13957 38597 13991
rect 38631 13957 38643 13991
rect 43272 13988 43300 14016
rect 54202 13988 54208 14000
rect 38585 13951 38643 13957
rect 41524 13960 43300 13988
rect 54163 13960 54208 13988
rect 34422 13929 34428 13932
rect 33505 13923 33563 13929
rect 33505 13920 33517 13923
rect 32600 13892 33517 13920
rect 29733 13855 29791 13861
rect 29733 13821 29745 13855
rect 29779 13852 29791 13855
rect 31021 13855 31079 13861
rect 29779 13824 30972 13852
rect 29779 13821 29791 13824
rect 29733 13815 29791 13821
rect 30944 13796 30972 13824
rect 31021 13821 31033 13855
rect 31067 13852 31079 13855
rect 32600 13852 32628 13892
rect 33505 13889 33517 13892
rect 33551 13889 33563 13923
rect 33505 13883 33563 13889
rect 34149 13923 34207 13929
rect 34149 13889 34161 13923
rect 34195 13889 34207 13923
rect 34416 13920 34428 13929
rect 34383 13892 34428 13920
rect 34149 13883 34207 13889
rect 34416 13883 34428 13892
rect 34422 13880 34428 13883
rect 34480 13880 34486 13932
rect 36262 13880 36268 13932
rect 36320 13920 36326 13932
rect 38194 13920 38200 13932
rect 36320 13892 38200 13920
rect 36320 13880 36326 13892
rect 38194 13880 38200 13892
rect 38252 13880 38258 13932
rect 38841 13923 38899 13929
rect 38841 13889 38853 13923
rect 38887 13889 38899 13923
rect 38841 13883 38899 13889
rect 32950 13852 32956 13864
rect 31067 13824 32628 13852
rect 32911 13824 32956 13852
rect 31067 13821 31079 13824
rect 31021 13815 31079 13821
rect 32950 13812 32956 13824
rect 33008 13812 33014 13864
rect 33594 13812 33600 13864
rect 33652 13852 33658 13864
rect 33689 13855 33747 13861
rect 33689 13852 33701 13855
rect 33652 13824 33701 13852
rect 33652 13812 33658 13824
rect 33689 13821 33701 13824
rect 33735 13821 33747 13855
rect 36538 13852 36544 13864
rect 36499 13824 36544 13852
rect 33689 13815 33747 13821
rect 36538 13812 36544 13824
rect 36596 13812 36602 13864
rect 38856 13852 38884 13883
rect 38930 13880 38936 13932
rect 38988 13920 38994 13932
rect 39393 13923 39451 13929
rect 39393 13920 39405 13923
rect 38988 13892 39405 13920
rect 38988 13880 38994 13892
rect 39393 13889 39405 13892
rect 39439 13920 39451 13923
rect 39758 13920 39764 13932
rect 39439 13892 39764 13920
rect 39439 13889 39451 13892
rect 39393 13883 39451 13889
rect 39758 13880 39764 13892
rect 39816 13880 39822 13932
rect 39850 13880 39856 13932
rect 39908 13920 39914 13932
rect 40129 13923 40187 13929
rect 40129 13920 40141 13923
rect 39908 13892 40141 13920
rect 39908 13880 39914 13892
rect 40129 13889 40141 13892
rect 40175 13920 40187 13923
rect 40494 13920 40500 13932
rect 40175 13892 40500 13920
rect 40175 13889 40187 13892
rect 40129 13883 40187 13889
rect 40494 13880 40500 13892
rect 40552 13880 40558 13932
rect 41046 13920 41052 13932
rect 41007 13892 41052 13920
rect 41046 13880 41052 13892
rect 41104 13880 41110 13932
rect 41138 13880 41144 13932
rect 41196 13920 41202 13932
rect 41524 13920 41552 13960
rect 54202 13948 54208 13960
rect 54260 13948 54266 14000
rect 41196 13892 41552 13920
rect 53469 13923 53527 13929
rect 41196 13880 41202 13892
rect 53469 13889 53481 13923
rect 53515 13920 53527 13923
rect 53558 13920 53564 13932
rect 53515 13892 53564 13920
rect 53515 13889 53527 13892
rect 53469 13883 53527 13889
rect 53558 13880 53564 13892
rect 53616 13880 53622 13932
rect 39114 13852 39120 13864
rect 38856 13824 39120 13852
rect 39114 13812 39120 13824
rect 39172 13812 39178 13864
rect 41414 13812 41420 13864
rect 41472 13852 41478 13864
rect 42613 13855 42671 13861
rect 42613 13852 42625 13855
rect 41472 13824 42625 13852
rect 41472 13812 41478 13824
rect 42613 13821 42625 13824
rect 42659 13821 42671 13855
rect 42613 13815 42671 13821
rect 53834 13812 53840 13864
rect 53892 13852 53898 13864
rect 54021 13855 54079 13861
rect 54021 13852 54033 13855
rect 53892 13824 54033 13852
rect 53892 13812 53898 13824
rect 54021 13821 54033 13824
rect 54067 13821 54079 13855
rect 54021 13815 54079 13821
rect 30469 13787 30527 13793
rect 30469 13784 30481 13787
rect 26712 13756 27568 13784
rect 29748 13756 30481 13784
rect 1670 13716 1676 13728
rect 1631 13688 1676 13716
rect 1670 13676 1676 13688
rect 1728 13676 1734 13728
rect 12805 13719 12863 13725
rect 12805 13685 12817 13719
rect 12851 13716 12863 13719
rect 13170 13716 13176 13728
rect 12851 13688 13176 13716
rect 12851 13685 12863 13688
rect 12805 13679 12863 13685
rect 13170 13676 13176 13688
rect 13228 13676 13234 13728
rect 15286 13716 15292 13728
rect 15247 13688 15292 13716
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 15749 13719 15807 13725
rect 15749 13716 15761 13719
rect 15712 13688 15761 13716
rect 15712 13676 15718 13688
rect 15749 13685 15761 13688
rect 15795 13685 15807 13719
rect 15749 13679 15807 13685
rect 16758 13676 16764 13728
rect 16816 13716 16822 13728
rect 16853 13719 16911 13725
rect 16853 13716 16865 13719
rect 16816 13688 16865 13716
rect 16816 13676 16822 13688
rect 16853 13685 16865 13688
rect 16899 13685 16911 13719
rect 16853 13679 16911 13685
rect 18414 13676 18420 13728
rect 18472 13716 18478 13728
rect 18966 13716 18972 13728
rect 18472 13688 18972 13716
rect 18472 13676 18478 13688
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 20622 13676 20628 13728
rect 20680 13716 20686 13728
rect 20717 13719 20775 13725
rect 20717 13716 20729 13719
rect 20680 13688 20729 13716
rect 20680 13676 20686 13688
rect 20717 13685 20729 13688
rect 20763 13685 20775 13719
rect 20717 13679 20775 13685
rect 22646 13676 22652 13728
rect 22704 13716 22710 13728
rect 26712 13716 26740 13756
rect 27154 13716 27160 13728
rect 22704 13688 26740 13716
rect 27115 13688 27160 13716
rect 22704 13676 22710 13688
rect 27154 13676 27160 13688
rect 27212 13676 27218 13728
rect 27338 13676 27344 13728
rect 27396 13716 27402 13728
rect 28902 13716 28908 13728
rect 27396 13688 28908 13716
rect 27396 13676 27402 13688
rect 28902 13676 28908 13688
rect 28960 13716 28966 13728
rect 29748 13716 29776 13756
rect 30469 13753 30481 13756
rect 30515 13753 30527 13787
rect 30926 13784 30932 13796
rect 30839 13756 30932 13784
rect 30469 13747 30527 13753
rect 30926 13744 30932 13756
rect 30984 13784 30990 13796
rect 31478 13784 31484 13796
rect 30984 13756 31484 13784
rect 30984 13744 30990 13756
rect 31478 13744 31484 13756
rect 31536 13744 31542 13796
rect 35526 13744 35532 13796
rect 35584 13784 35590 13796
rect 36354 13784 36360 13796
rect 35584 13756 36360 13784
rect 35584 13744 35590 13756
rect 36354 13744 36360 13756
rect 36412 13744 36418 13796
rect 53282 13784 53288 13796
rect 38856 13756 51074 13784
rect 53243 13756 53288 13784
rect 29914 13716 29920 13728
rect 28960 13688 29776 13716
rect 29875 13688 29920 13716
rect 28960 13676 28966 13688
rect 29914 13676 29920 13688
rect 29972 13676 29978 13728
rect 33686 13676 33692 13728
rect 33744 13716 33750 13728
rect 35434 13716 35440 13728
rect 33744 13688 35440 13716
rect 33744 13676 33750 13688
rect 35434 13676 35440 13688
rect 35492 13676 35498 13728
rect 35986 13716 35992 13728
rect 35947 13688 35992 13716
rect 35986 13676 35992 13688
rect 36044 13676 36050 13728
rect 37461 13719 37519 13725
rect 37461 13685 37473 13719
rect 37507 13716 37519 13719
rect 37550 13716 37556 13728
rect 37507 13688 37556 13716
rect 37507 13685 37519 13688
rect 37461 13679 37519 13685
rect 37550 13676 37556 13688
rect 37608 13716 37614 13728
rect 38856 13716 38884 13756
rect 39482 13716 39488 13728
rect 37608 13688 38884 13716
rect 39443 13688 39488 13716
rect 37608 13676 37614 13688
rect 39482 13676 39488 13688
rect 39540 13676 39546 13728
rect 39850 13676 39856 13728
rect 39908 13716 39914 13728
rect 40129 13719 40187 13725
rect 40129 13716 40141 13719
rect 39908 13688 40141 13716
rect 39908 13676 39914 13688
rect 40129 13685 40141 13688
rect 40175 13685 40187 13719
rect 40862 13716 40868 13728
rect 40823 13688 40868 13716
rect 40129 13679 40187 13685
rect 40862 13676 40868 13688
rect 40920 13676 40926 13728
rect 41506 13716 41512 13728
rect 41467 13688 41512 13716
rect 41506 13676 41512 13688
rect 41564 13676 41570 13728
rect 51046 13716 51074 13756
rect 53282 13744 53288 13756
rect 53340 13744 53346 13796
rect 54018 13716 54024 13728
rect 51046 13688 54024 13716
rect 54018 13676 54024 13688
rect 54076 13676 54082 13728
rect 1104 13626 54832 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 54832 13626
rect 1104 13552 54832 13574
rect 14829 13515 14887 13521
rect 14829 13481 14841 13515
rect 14875 13512 14887 13515
rect 14918 13512 14924 13524
rect 14875 13484 14924 13512
rect 14875 13481 14887 13484
rect 14829 13475 14887 13481
rect 14918 13472 14924 13484
rect 14976 13472 14982 13524
rect 15562 13472 15568 13524
rect 15620 13512 15626 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15620 13484 16037 13512
rect 15620 13472 15626 13484
rect 16025 13481 16037 13484
rect 16071 13481 16083 13515
rect 16025 13475 16083 13481
rect 16114 13472 16120 13524
rect 16172 13512 16178 13524
rect 22278 13512 22284 13524
rect 16172 13484 20300 13512
rect 22239 13484 22284 13512
rect 16172 13472 16178 13484
rect 13722 13404 13728 13456
rect 13780 13444 13786 13456
rect 17126 13444 17132 13456
rect 13780 13416 17132 13444
rect 13780 13404 13786 13416
rect 17126 13404 17132 13416
rect 17184 13404 17190 13456
rect 20070 13404 20076 13456
rect 20128 13404 20134 13456
rect 13633 13379 13691 13385
rect 13633 13345 13645 13379
rect 13679 13376 13691 13379
rect 15378 13376 15384 13388
rect 13679 13348 15384 13376
rect 13679 13345 13691 13348
rect 13633 13339 13691 13345
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13376 16359 13379
rect 18877 13379 18935 13385
rect 16347 13348 17816 13376
rect 16347 13345 16359 13348
rect 16301 13339 16359 13345
rect 1854 13308 1860 13320
rect 1815 13280 1860 13308
rect 1854 13268 1860 13280
rect 1912 13268 1918 13320
rect 14642 13308 14648 13320
rect 14603 13280 14648 13308
rect 14642 13268 14648 13280
rect 14700 13268 14706 13320
rect 15286 13308 15292 13320
rect 15247 13280 15292 13308
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 15930 13268 15936 13320
rect 15988 13308 15994 13320
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 15988 13280 16221 13308
rect 15988 13268 15994 13280
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13277 16451 13311
rect 16393 13271 16451 13277
rect 1670 13172 1676 13184
rect 1631 13144 1676 13172
rect 1670 13132 1676 13144
rect 1728 13132 1734 13184
rect 12621 13175 12679 13181
rect 12621 13141 12633 13175
rect 12667 13172 12679 13175
rect 13170 13172 13176 13184
rect 12667 13144 13176 13172
rect 12667 13141 12679 13144
rect 12621 13135 12679 13141
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 14826 13132 14832 13184
rect 14884 13172 14890 13184
rect 15473 13175 15531 13181
rect 15473 13172 15485 13175
rect 14884 13144 15485 13172
rect 14884 13132 14890 13144
rect 15473 13141 15485 13144
rect 15519 13141 15531 13175
rect 15473 13135 15531 13141
rect 16298 13132 16304 13184
rect 16356 13172 16362 13184
rect 16408 13172 16436 13271
rect 16482 13268 16488 13320
rect 16540 13308 16546 13320
rect 16540 13280 16585 13308
rect 16540 13268 16546 13280
rect 16666 13268 16672 13320
rect 16724 13308 16730 13320
rect 17586 13308 17592 13320
rect 16724 13280 17592 13308
rect 16724 13268 16730 13280
rect 17586 13268 17592 13280
rect 17644 13268 17650 13320
rect 17788 13308 17816 13348
rect 18877 13345 18889 13379
rect 18923 13376 18935 13379
rect 20088 13376 20116 13404
rect 18923 13348 20116 13376
rect 20272 13376 20300 13484
rect 22278 13472 22284 13484
rect 22336 13472 22342 13524
rect 23385 13515 23443 13521
rect 23385 13481 23397 13515
rect 23431 13512 23443 13515
rect 23658 13512 23664 13524
rect 23431 13484 23664 13512
rect 23431 13481 23443 13484
rect 23385 13475 23443 13481
rect 23658 13472 23664 13484
rect 23716 13512 23722 13524
rect 24578 13512 24584 13524
rect 23716 13484 24440 13512
rect 24539 13484 24584 13512
rect 23716 13472 23722 13484
rect 20349 13447 20407 13453
rect 20349 13413 20361 13447
rect 20395 13444 20407 13447
rect 24026 13444 24032 13456
rect 20395 13416 24032 13444
rect 20395 13413 20407 13416
rect 20349 13407 20407 13413
rect 24026 13404 24032 13416
rect 24084 13404 24090 13456
rect 24412 13444 24440 13484
rect 24578 13472 24584 13484
rect 24636 13472 24642 13524
rect 26053 13515 26111 13521
rect 26053 13481 26065 13515
rect 26099 13512 26111 13515
rect 26234 13512 26240 13524
rect 26099 13484 26240 13512
rect 26099 13481 26111 13484
rect 26053 13475 26111 13481
rect 26234 13472 26240 13484
rect 26292 13472 26298 13524
rect 26786 13472 26792 13524
rect 26844 13512 26850 13524
rect 26881 13515 26939 13521
rect 26881 13512 26893 13515
rect 26844 13484 26893 13512
rect 26844 13472 26850 13484
rect 26881 13481 26893 13484
rect 26927 13512 26939 13515
rect 27338 13512 27344 13524
rect 26927 13484 27344 13512
rect 26927 13481 26939 13484
rect 26881 13475 26939 13481
rect 27338 13472 27344 13484
rect 27396 13472 27402 13524
rect 29086 13512 29092 13524
rect 29047 13484 29092 13512
rect 29086 13472 29092 13484
rect 29144 13472 29150 13524
rect 30285 13515 30343 13521
rect 30285 13481 30297 13515
rect 30331 13512 30343 13515
rect 31110 13512 31116 13524
rect 30331 13484 31116 13512
rect 30331 13481 30343 13484
rect 30285 13475 30343 13481
rect 31110 13472 31116 13484
rect 31168 13472 31174 13524
rect 32122 13472 32128 13524
rect 32180 13512 32186 13524
rect 32309 13515 32367 13521
rect 32309 13512 32321 13515
rect 32180 13484 32321 13512
rect 32180 13472 32186 13484
rect 32309 13481 32321 13484
rect 32355 13481 32367 13515
rect 32309 13475 32367 13481
rect 32858 13472 32864 13524
rect 32916 13512 32922 13524
rect 32953 13515 33011 13521
rect 32953 13512 32965 13515
rect 32916 13484 32965 13512
rect 32916 13472 32922 13484
rect 32953 13481 32965 13484
rect 32999 13481 33011 13515
rect 37185 13515 37243 13521
rect 37185 13512 37197 13515
rect 32953 13475 33011 13481
rect 33060 13484 37197 13512
rect 27433 13447 27491 13453
rect 24412 13416 24808 13444
rect 20272 13348 20852 13376
rect 18923 13345 18935 13348
rect 18877 13339 18935 13345
rect 18322 13308 18328 13320
rect 17788 13280 18328 13308
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13308 19487 13311
rect 19886 13308 19892 13320
rect 19475 13280 19892 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 19978 13268 19984 13320
rect 20036 13308 20042 13320
rect 20824 13317 20852 13348
rect 23750 13336 23756 13388
rect 23808 13376 23814 13388
rect 23937 13379 23995 13385
rect 23937 13376 23949 13379
rect 23808 13348 23949 13376
rect 23808 13336 23814 13348
rect 23937 13345 23949 13348
rect 23983 13345 23995 13379
rect 23937 13339 23995 13345
rect 20073 13311 20131 13317
rect 20073 13308 20085 13311
rect 20036 13280 20085 13308
rect 20036 13268 20042 13280
rect 20073 13277 20085 13280
rect 20119 13277 20131 13311
rect 20073 13271 20131 13277
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 23382 13308 23388 13320
rect 20855 13280 23388 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 24780 13317 24808 13416
rect 27433 13413 27445 13447
rect 27479 13444 27491 13447
rect 33060 13444 33088 13484
rect 37185 13481 37197 13484
rect 37231 13481 37243 13515
rect 37185 13475 37243 13481
rect 37274 13472 37280 13524
rect 37332 13512 37338 13524
rect 37734 13512 37740 13524
rect 37332 13484 37740 13512
rect 37332 13472 37338 13484
rect 37734 13472 37740 13484
rect 37792 13512 37798 13524
rect 38381 13515 38439 13521
rect 38381 13512 38393 13515
rect 37792 13484 38393 13512
rect 37792 13472 37798 13484
rect 38381 13481 38393 13484
rect 38427 13481 38439 13515
rect 38381 13475 38439 13481
rect 38470 13472 38476 13524
rect 38528 13512 38534 13524
rect 39850 13512 39856 13524
rect 38528 13484 39856 13512
rect 38528 13472 38534 13484
rect 39850 13472 39856 13484
rect 39908 13472 39914 13524
rect 40770 13512 40776 13524
rect 40731 13484 40776 13512
rect 40770 13472 40776 13484
rect 40828 13472 40834 13524
rect 41506 13512 41512 13524
rect 41467 13484 41512 13512
rect 41506 13472 41512 13484
rect 41564 13512 41570 13524
rect 41969 13515 42027 13521
rect 41969 13512 41981 13515
rect 41564 13484 41981 13512
rect 41564 13472 41570 13484
rect 41969 13481 41981 13484
rect 42015 13481 42027 13515
rect 42518 13512 42524 13524
rect 42479 13484 42524 13512
rect 41969 13475 42027 13481
rect 42518 13472 42524 13484
rect 42576 13472 42582 13524
rect 53282 13512 53288 13524
rect 51046 13484 53288 13512
rect 51046 13444 51074 13484
rect 53282 13472 53288 13484
rect 53340 13472 53346 13524
rect 54202 13512 54208 13524
rect 54163 13484 54208 13512
rect 54202 13472 54208 13484
rect 54260 13472 54266 13524
rect 53558 13444 53564 13456
rect 27479 13416 33088 13444
rect 36372 13416 51074 13444
rect 53519 13416 53564 13444
rect 27479 13413 27491 13416
rect 27433 13407 27491 13413
rect 24949 13379 25007 13385
rect 24949 13345 24961 13379
rect 24995 13376 25007 13379
rect 25314 13376 25320 13388
rect 24995 13348 25320 13376
rect 24995 13345 25007 13348
rect 24949 13339 25007 13345
rect 25314 13336 25320 13348
rect 25372 13336 25378 13388
rect 26789 13379 26847 13385
rect 26789 13345 26801 13379
rect 26835 13376 26847 13379
rect 29917 13379 29975 13385
rect 26835 13348 28028 13376
rect 26835 13345 26847 13348
rect 26789 13339 26847 13345
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13308 24823 13311
rect 25130 13308 25136 13320
rect 24811 13280 25136 13308
rect 24811 13277 24823 13280
rect 24765 13271 24823 13277
rect 25130 13268 25136 13280
rect 25188 13268 25194 13320
rect 25406 13308 25412 13320
rect 25367 13280 25412 13308
rect 25406 13268 25412 13280
rect 25464 13268 25470 13320
rect 27062 13268 27068 13320
rect 27120 13308 27126 13320
rect 28000 13317 28028 13348
rect 29917 13345 29929 13379
rect 29963 13376 29975 13379
rect 30466 13376 30472 13388
rect 29963 13348 30472 13376
rect 29963 13345 29975 13348
rect 29917 13339 29975 13345
rect 30466 13336 30472 13348
rect 30524 13336 30530 13388
rect 31202 13336 31208 13388
rect 31260 13376 31266 13388
rect 31665 13379 31723 13385
rect 31665 13376 31677 13379
rect 31260 13348 31677 13376
rect 31260 13336 31266 13348
rect 31665 13345 31677 13348
rect 31711 13345 31723 13379
rect 33134 13376 33140 13388
rect 31665 13339 31723 13345
rect 31772 13348 33140 13376
rect 27308 13311 27366 13317
rect 27308 13308 27320 13311
rect 27120 13280 27320 13308
rect 27120 13268 27126 13280
rect 27308 13277 27320 13280
rect 27354 13308 27366 13311
rect 27985 13311 28043 13317
rect 27354 13280 27936 13308
rect 27354 13277 27366 13280
rect 27308 13271 27366 13277
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 18610 13243 18668 13249
rect 18610 13240 18622 13243
rect 17092 13212 18622 13240
rect 17092 13200 17098 13212
rect 18610 13209 18622 13212
rect 18656 13209 18668 13243
rect 20349 13243 20407 13249
rect 18610 13203 18668 13209
rect 19628 13212 20300 13240
rect 16356 13144 16436 13172
rect 17497 13175 17555 13181
rect 16356 13132 16362 13144
rect 17497 13141 17509 13175
rect 17543 13172 17555 13175
rect 17954 13172 17960 13184
rect 17543 13144 17960 13172
rect 17543 13141 17555 13144
rect 17497 13135 17555 13141
rect 17954 13132 17960 13144
rect 18012 13132 18018 13184
rect 19628 13181 19656 13212
rect 19613 13175 19671 13181
rect 19613 13141 19625 13175
rect 19659 13141 19671 13175
rect 20162 13172 20168 13184
rect 20123 13144 20168 13172
rect 19613 13135 19671 13141
rect 20162 13132 20168 13144
rect 20220 13132 20226 13184
rect 20272 13172 20300 13212
rect 20349 13209 20361 13243
rect 20395 13240 20407 13243
rect 25038 13240 25044 13252
rect 20395 13212 25044 13240
rect 20395 13209 20407 13212
rect 20349 13203 20407 13209
rect 25038 13200 25044 13212
rect 25096 13200 25102 13252
rect 27908 13240 27936 13280
rect 27985 13277 27997 13311
rect 28031 13308 28043 13311
rect 28350 13308 28356 13320
rect 28031 13280 28356 13308
rect 28031 13277 28043 13280
rect 27985 13271 28043 13277
rect 28350 13268 28356 13280
rect 28408 13268 28414 13320
rect 29181 13311 29239 13317
rect 29181 13277 29193 13311
rect 29227 13308 29239 13311
rect 29546 13308 29552 13320
rect 29227 13280 29552 13308
rect 29227 13277 29239 13280
rect 29181 13271 29239 13277
rect 29546 13268 29552 13280
rect 29604 13268 29610 13320
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13308 30159 13311
rect 30374 13308 30380 13320
rect 30147 13280 30380 13308
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 30374 13268 30380 13280
rect 30432 13268 30438 13320
rect 30742 13308 30748 13320
rect 30703 13280 30748 13308
rect 30742 13268 30748 13280
rect 30800 13268 30806 13320
rect 30834 13268 30840 13320
rect 30892 13308 30898 13320
rect 31021 13311 31079 13317
rect 30892 13280 30937 13308
rect 30892 13268 30898 13280
rect 31021 13277 31033 13311
rect 31067 13277 31079 13311
rect 31021 13271 31079 13277
rect 28994 13240 29000 13252
rect 27908 13212 29000 13240
rect 28994 13200 29000 13212
rect 29052 13200 29058 13252
rect 29914 13200 29920 13252
rect 29972 13240 29978 13252
rect 31036 13240 31064 13271
rect 31478 13268 31484 13320
rect 31536 13308 31542 13320
rect 31772 13308 31800 13348
rect 33134 13336 33140 13348
rect 33192 13336 33198 13388
rect 33502 13376 33508 13388
rect 33463 13348 33508 13376
rect 33502 13336 33508 13348
rect 33560 13336 33566 13388
rect 36262 13376 36268 13388
rect 36223 13348 36268 13376
rect 36262 13336 36268 13348
rect 36320 13336 36326 13388
rect 31536 13280 31800 13308
rect 31536 13268 31542 13280
rect 31846 13268 31852 13320
rect 31904 13308 31910 13320
rect 36372 13308 36400 13416
rect 53558 13404 53564 13416
rect 53616 13404 53622 13456
rect 37366 13336 37372 13388
rect 37424 13376 37430 13388
rect 37826 13376 37832 13388
rect 37424 13348 37832 13376
rect 37424 13336 37430 13348
rect 37826 13336 37832 13348
rect 37884 13376 37890 13388
rect 39482 13376 39488 13388
rect 37884 13348 39488 13376
rect 37884 13336 37890 13348
rect 37090 13308 37096 13320
rect 31904 13280 36400 13308
rect 37051 13280 37096 13308
rect 31904 13268 31910 13280
rect 37090 13268 37096 13280
rect 37148 13268 37154 13320
rect 37550 13268 37556 13320
rect 37608 13308 37614 13320
rect 37608 13280 37653 13308
rect 37608 13268 37614 13280
rect 38102 13268 38108 13320
rect 38160 13308 38166 13320
rect 38197 13311 38255 13317
rect 38197 13308 38209 13311
rect 38160 13280 38209 13308
rect 38160 13268 38166 13280
rect 38197 13277 38209 13280
rect 38243 13308 38255 13311
rect 38470 13308 38476 13320
rect 38243 13280 38476 13308
rect 38243 13277 38255 13280
rect 38197 13271 38255 13277
rect 38470 13268 38476 13280
rect 38528 13268 38534 13320
rect 39224 13317 39252 13348
rect 39482 13336 39488 13348
rect 39540 13336 39546 13388
rect 39209 13311 39267 13317
rect 39209 13277 39221 13311
rect 39255 13277 39267 13311
rect 39390 13308 39396 13320
rect 39351 13280 39396 13308
rect 39209 13271 39267 13277
rect 39390 13268 39396 13280
rect 39448 13268 39454 13320
rect 40034 13308 40040 13320
rect 39995 13280 40040 13308
rect 40034 13268 40040 13280
rect 40092 13268 40098 13320
rect 40678 13268 40684 13320
rect 40736 13308 40742 13320
rect 40957 13311 41015 13317
rect 40957 13308 40969 13311
rect 40736 13280 40969 13308
rect 40736 13268 40742 13280
rect 40957 13277 40969 13280
rect 41003 13277 41015 13311
rect 54018 13308 54024 13320
rect 53979 13280 54024 13308
rect 40957 13271 41015 13277
rect 54018 13268 54024 13280
rect 54076 13268 54082 13320
rect 32674 13240 32680 13252
rect 29972 13212 32680 13240
rect 29972 13200 29978 13212
rect 32674 13200 32680 13212
rect 32732 13200 32738 13252
rect 34241 13243 34299 13249
rect 34241 13209 34253 13243
rect 34287 13240 34299 13243
rect 34422 13240 34428 13252
rect 34287 13212 34428 13240
rect 34287 13209 34299 13212
rect 34241 13203 34299 13209
rect 34422 13200 34428 13212
rect 34480 13200 34486 13252
rect 35986 13200 35992 13252
rect 36044 13249 36050 13252
rect 36044 13240 36056 13249
rect 40126 13240 40132 13252
rect 36044 13212 36089 13240
rect 37752 13212 40132 13240
rect 36044 13203 36056 13212
rect 36044 13200 36050 13203
rect 20714 13172 20720 13184
rect 20272 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 24118 13132 24124 13184
rect 24176 13172 24182 13184
rect 24394 13172 24400 13184
rect 24176 13144 24400 13172
rect 24176 13132 24182 13144
rect 24394 13132 24400 13144
rect 24452 13132 24458 13184
rect 27246 13172 27252 13184
rect 27207 13144 27252 13172
rect 27246 13132 27252 13144
rect 27304 13132 27310 13184
rect 28537 13175 28595 13181
rect 28537 13141 28549 13175
rect 28583 13172 28595 13175
rect 28810 13172 28816 13184
rect 28583 13144 28816 13172
rect 28583 13141 28595 13144
rect 28537 13135 28595 13141
rect 28810 13132 28816 13144
rect 28868 13132 28874 13184
rect 28902 13132 28908 13184
rect 28960 13172 28966 13184
rect 30374 13172 30380 13184
rect 28960 13144 30380 13172
rect 28960 13132 28966 13144
rect 30374 13132 30380 13144
rect 30432 13172 30438 13184
rect 30650 13172 30656 13184
rect 30432 13144 30656 13172
rect 30432 13132 30438 13144
rect 30650 13132 30656 13144
rect 30708 13132 30714 13184
rect 31202 13172 31208 13184
rect 31163 13144 31208 13172
rect 31202 13132 31208 13144
rect 31260 13132 31266 13184
rect 33042 13132 33048 13184
rect 33100 13172 33106 13184
rect 34149 13175 34207 13181
rect 34149 13172 34161 13175
rect 33100 13144 34161 13172
rect 33100 13132 33106 13144
rect 34149 13141 34161 13144
rect 34195 13141 34207 13175
rect 34149 13135 34207 13141
rect 34885 13175 34943 13181
rect 34885 13141 34897 13175
rect 34931 13172 34943 13175
rect 35526 13172 35532 13184
rect 34931 13144 35532 13172
rect 34931 13141 34943 13144
rect 34885 13135 34943 13141
rect 35526 13132 35532 13144
rect 35584 13132 35590 13184
rect 37366 13132 37372 13184
rect 37424 13172 37430 13184
rect 37752 13181 37780 13212
rect 40126 13200 40132 13212
rect 40184 13200 40190 13252
rect 37553 13175 37611 13181
rect 37553 13172 37565 13175
rect 37424 13144 37565 13172
rect 37424 13132 37430 13144
rect 37553 13141 37565 13144
rect 37599 13141 37611 13175
rect 37553 13135 37611 13141
rect 37737 13175 37795 13181
rect 37737 13141 37749 13175
rect 37783 13141 37795 13175
rect 39022 13172 39028 13184
rect 38983 13144 39028 13172
rect 37737 13135 37795 13141
rect 39022 13132 39028 13144
rect 39080 13132 39086 13184
rect 39758 13132 39764 13184
rect 39816 13172 39822 13184
rect 40221 13175 40279 13181
rect 40221 13172 40233 13175
rect 39816 13144 40233 13172
rect 39816 13132 39822 13144
rect 40221 13141 40233 13144
rect 40267 13172 40279 13175
rect 41138 13172 41144 13184
rect 40267 13144 41144 13172
rect 40267 13141 40279 13144
rect 40221 13135 40279 13141
rect 41138 13132 41144 13144
rect 41196 13132 41202 13184
rect 1104 13082 54832 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 54832 13082
rect 1104 13008 54832 13030
rect 1854 12928 1860 12980
rect 1912 12968 1918 12980
rect 12437 12971 12495 12977
rect 1912 12940 6914 12968
rect 1912 12928 1918 12940
rect 6886 12900 6914 12940
rect 12437 12937 12449 12971
rect 12483 12968 12495 12971
rect 14182 12968 14188 12980
rect 12483 12940 14188 12968
rect 12483 12937 12495 12940
rect 12437 12931 12495 12937
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 14461 12971 14519 12977
rect 14461 12937 14473 12971
rect 14507 12968 14519 12971
rect 16114 12968 16120 12980
rect 14507 12940 16120 12968
rect 14507 12937 14519 12940
rect 14461 12931 14519 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 17034 12968 17040 12980
rect 16995 12940 17040 12968
rect 17034 12928 17040 12940
rect 17092 12928 17098 12980
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 17681 12971 17739 12977
rect 17681 12968 17693 12971
rect 17184 12940 17693 12968
rect 17184 12928 17190 12940
rect 17681 12937 17693 12940
rect 17727 12937 17739 12971
rect 18230 12968 18236 12980
rect 18191 12940 18236 12968
rect 17681 12931 17739 12937
rect 18230 12928 18236 12940
rect 18288 12928 18294 12980
rect 19978 12968 19984 12980
rect 19306 12940 19984 12968
rect 11885 12903 11943 12909
rect 6886 12872 11376 12900
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 1903 12804 6914 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 6886 12696 6914 12804
rect 11348 12764 11376 12872
rect 11885 12869 11897 12903
rect 11931 12900 11943 12903
rect 15102 12900 15108 12912
rect 11931 12872 15108 12900
rect 11931 12869 11943 12872
rect 11885 12863 11943 12869
rect 15102 12860 15108 12872
rect 15160 12860 15166 12912
rect 15289 12903 15347 12909
rect 15289 12869 15301 12903
rect 15335 12900 15347 12903
rect 15335 12872 17540 12900
rect 15335 12869 15347 12872
rect 15289 12863 15347 12869
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 13170 12832 13176 12844
rect 13035 12804 13176 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 13412 12804 13461 12832
rect 13412 12792 13418 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 13538 12792 13544 12844
rect 13596 12832 13602 12844
rect 13722 12832 13728 12844
rect 13596 12804 13641 12832
rect 13683 12804 13728 12832
rect 13596 12792 13602 12804
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 14182 12792 14188 12844
rect 14240 12832 14246 12844
rect 14734 12832 14740 12844
rect 14240 12804 14740 12832
rect 14240 12792 14246 12804
rect 14734 12792 14740 12804
rect 14792 12832 14798 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14792 12804 14933 12832
rect 14792 12792 14798 12804
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 16114 12832 16120 12844
rect 16027 12804 16120 12832
rect 14921 12795 14979 12801
rect 16114 12792 16120 12804
rect 16172 12832 16178 12844
rect 16298 12832 16304 12844
rect 16172 12804 16304 12832
rect 16172 12792 16178 12804
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 17512 12841 17540 12872
rect 17586 12860 17592 12912
rect 17644 12900 17650 12912
rect 19306 12900 19334 12940
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 20162 12928 20168 12980
rect 20220 12968 20226 12980
rect 24949 12971 25007 12977
rect 20220 12940 24900 12968
rect 20220 12928 20226 12940
rect 22278 12900 22284 12912
rect 17644 12872 19334 12900
rect 20180 12872 22284 12900
rect 17644 12860 17650 12872
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12801 17555 12835
rect 17497 12795 17555 12801
rect 19357 12835 19415 12841
rect 19357 12801 19369 12835
rect 19403 12832 19415 12835
rect 19978 12832 19984 12844
rect 19403 12804 19984 12832
rect 19403 12801 19415 12804
rect 19357 12795 19415 12801
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 11348 12736 15761 12764
rect 15749 12733 15761 12736
rect 15795 12733 15807 12767
rect 15930 12764 15936 12776
rect 15891 12736 15936 12764
rect 15749 12727 15807 12733
rect 15930 12724 15936 12736
rect 15988 12724 15994 12776
rect 16025 12767 16083 12773
rect 16025 12733 16037 12767
rect 16071 12733 16083 12767
rect 16025 12727 16083 12733
rect 15838 12696 15844 12708
rect 6886 12668 15844 12696
rect 15838 12656 15844 12668
rect 15896 12656 15902 12708
rect 16040 12696 16068 12727
rect 16206 12724 16212 12776
rect 16264 12764 16270 12776
rect 16868 12764 16896 12795
rect 19978 12792 19984 12804
rect 20036 12792 20042 12844
rect 20070 12792 20076 12844
rect 20128 12832 20134 12844
rect 20180 12832 20208 12872
rect 22278 12860 22284 12872
rect 22336 12900 22342 12912
rect 22554 12900 22560 12912
rect 22336 12872 22560 12900
rect 22336 12860 22342 12872
rect 22554 12860 22560 12872
rect 22612 12860 22618 12912
rect 23014 12900 23020 12912
rect 22975 12872 23020 12900
rect 23014 12860 23020 12872
rect 23072 12860 23078 12912
rect 24872 12900 24900 12940
rect 24949 12937 24961 12971
rect 24995 12968 25007 12971
rect 26602 12968 26608 12980
rect 24995 12940 26608 12968
rect 24995 12937 25007 12940
rect 24949 12931 25007 12937
rect 26602 12928 26608 12940
rect 26660 12928 26666 12980
rect 27982 12968 27988 12980
rect 27943 12940 27988 12968
rect 27982 12928 27988 12940
rect 28040 12928 28046 12980
rect 29730 12928 29736 12980
rect 29788 12968 29794 12980
rect 29788 12940 29960 12968
rect 29788 12928 29794 12940
rect 26145 12903 26203 12909
rect 26145 12900 26157 12903
rect 24872 12872 26157 12900
rect 26145 12869 26157 12872
rect 26191 12900 26203 12903
rect 26234 12900 26240 12912
rect 26191 12872 26240 12900
rect 26191 12869 26203 12872
rect 26145 12863 26203 12869
rect 26234 12860 26240 12872
rect 26292 12900 26298 12912
rect 27154 12900 27160 12912
rect 26292 12872 27160 12900
rect 26292 12860 26298 12872
rect 27154 12860 27160 12872
rect 27212 12860 27218 12912
rect 27430 12860 27436 12912
rect 27488 12900 27494 12912
rect 28442 12900 28448 12912
rect 27488 12872 28448 12900
rect 27488 12860 27494 12872
rect 28442 12860 28448 12872
rect 28500 12900 28506 12912
rect 29822 12900 29828 12912
rect 28500 12872 28652 12900
rect 28500 12860 28506 12872
rect 20346 12841 20352 12844
rect 20340 12832 20352 12841
rect 20128 12804 20221 12832
rect 20307 12804 20352 12832
rect 20128 12792 20134 12804
rect 20340 12795 20352 12804
rect 20346 12792 20352 12795
rect 20404 12792 20410 12844
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 21450 12832 21456 12844
rect 20772 12804 21456 12832
rect 20772 12792 20778 12804
rect 21450 12792 21456 12804
rect 21508 12792 21514 12844
rect 22094 12792 22100 12844
rect 22152 12832 22158 12844
rect 22373 12835 22431 12841
rect 22373 12832 22385 12835
rect 22152 12804 22385 12832
rect 22152 12792 22158 12804
rect 22373 12801 22385 12804
rect 22419 12801 22431 12835
rect 24026 12832 24032 12844
rect 23987 12804 24032 12832
rect 22373 12795 22431 12801
rect 24026 12792 24032 12804
rect 24084 12792 24090 12844
rect 25041 12835 25099 12841
rect 25041 12801 25053 12835
rect 25087 12832 25099 12835
rect 25314 12832 25320 12844
rect 25087 12804 25320 12832
rect 25087 12801 25099 12804
rect 25041 12795 25099 12801
rect 25314 12792 25320 12804
rect 25372 12832 25378 12844
rect 25372 12804 28580 12832
rect 25372 12792 25378 12804
rect 18138 12764 18144 12776
rect 16264 12736 16309 12764
rect 16868 12736 18144 12764
rect 16264 12724 16270 12736
rect 18138 12724 18144 12736
rect 18196 12724 18202 12776
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12733 19671 12767
rect 23477 12767 23535 12773
rect 23477 12764 23489 12767
rect 19613 12727 19671 12733
rect 21100 12736 23489 12764
rect 17954 12696 17960 12708
rect 16040 12668 17960 12696
rect 17954 12656 17960 12668
rect 18012 12656 18018 12708
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 13906 12628 13912 12640
rect 13867 12600 13912 12628
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 19628 12628 19656 12727
rect 19392 12600 19656 12628
rect 19392 12588 19398 12600
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 21100 12628 21128 12736
rect 23477 12733 23489 12736
rect 23523 12733 23535 12767
rect 23477 12727 23535 12733
rect 23842 12724 23848 12776
rect 23900 12764 23906 12776
rect 25133 12767 25191 12773
rect 23900 12736 24992 12764
rect 23900 12724 23906 12736
rect 21450 12696 21456 12708
rect 21411 12668 21456 12696
rect 21450 12656 21456 12668
rect 21508 12656 21514 12708
rect 22738 12656 22744 12708
rect 22796 12696 22802 12708
rect 24964 12696 24992 12736
rect 25133 12733 25145 12767
rect 25179 12733 25191 12767
rect 26237 12767 26295 12773
rect 26237 12764 26249 12767
rect 25133 12727 25191 12733
rect 26160 12736 26249 12764
rect 25148 12696 25176 12727
rect 26160 12708 26188 12736
rect 26237 12733 26249 12736
rect 26283 12733 26295 12767
rect 26237 12727 26295 12733
rect 26329 12767 26387 12773
rect 26329 12733 26341 12767
rect 26375 12733 26387 12767
rect 26329 12727 26387 12733
rect 27433 12767 27491 12773
rect 27433 12733 27445 12767
rect 27479 12733 27491 12767
rect 27433 12727 27491 12733
rect 22796 12668 23060 12696
rect 24964 12668 26096 12696
rect 22796 12656 22802 12668
rect 20772 12600 21128 12628
rect 20772 12588 20778 12600
rect 21174 12588 21180 12640
rect 21232 12628 21238 12640
rect 22097 12631 22155 12637
rect 22097 12628 22109 12631
rect 21232 12600 22109 12628
rect 21232 12588 21238 12600
rect 22097 12597 22109 12600
rect 22143 12597 22155 12631
rect 23032 12628 23060 12668
rect 24581 12631 24639 12637
rect 24581 12628 24593 12631
rect 23032 12600 24593 12628
rect 22097 12591 22155 12597
rect 24581 12597 24593 12600
rect 24627 12597 24639 12631
rect 24581 12591 24639 12597
rect 24946 12588 24952 12640
rect 25004 12628 25010 12640
rect 25777 12631 25835 12637
rect 25777 12628 25789 12631
rect 25004 12600 25789 12628
rect 25004 12588 25010 12600
rect 25777 12597 25789 12600
rect 25823 12597 25835 12631
rect 26068 12628 26096 12668
rect 26142 12656 26148 12708
rect 26200 12656 26206 12708
rect 26344 12628 26372 12727
rect 27448 12696 27476 12727
rect 28445 12699 28503 12705
rect 28445 12696 28457 12699
rect 27448 12668 28457 12696
rect 28445 12665 28457 12668
rect 28491 12665 28503 12699
rect 28552 12696 28580 12804
rect 28624 12764 28652 12872
rect 29656 12872 29828 12900
rect 28810 12832 28816 12844
rect 28771 12804 28816 12832
rect 28810 12792 28816 12804
rect 28868 12792 28874 12844
rect 29656 12841 29684 12872
rect 29822 12860 29828 12872
rect 29880 12860 29886 12912
rect 29932 12909 29960 12940
rect 30558 12928 30564 12980
rect 30616 12968 30622 12980
rect 30745 12971 30803 12977
rect 30745 12968 30757 12971
rect 30616 12940 30757 12968
rect 30616 12928 30622 12940
rect 30745 12937 30757 12940
rect 30791 12937 30803 12971
rect 30745 12931 30803 12937
rect 32122 12928 32128 12980
rect 32180 12968 32186 12980
rect 35989 12971 36047 12977
rect 32180 12940 35848 12968
rect 32180 12928 32186 12940
rect 29917 12903 29975 12909
rect 29917 12869 29929 12903
rect 29963 12869 29975 12903
rect 29917 12863 29975 12869
rect 29641 12835 29699 12841
rect 29641 12801 29653 12835
rect 29687 12801 29699 12835
rect 29641 12795 29699 12801
rect 29730 12792 29736 12844
rect 29788 12832 29794 12844
rect 29788 12804 29833 12832
rect 29788 12792 29794 12804
rect 28721 12767 28779 12773
rect 28721 12764 28733 12767
rect 28624 12736 28733 12764
rect 28721 12733 28733 12736
rect 28767 12733 28779 12767
rect 29932 12764 29960 12863
rect 30650 12860 30656 12912
rect 30708 12900 30714 12912
rect 31386 12900 31392 12912
rect 30708 12872 30880 12900
rect 30708 12860 30714 12872
rect 30006 12792 30012 12844
rect 30064 12832 30070 12844
rect 30147 12835 30205 12841
rect 30064 12804 30109 12832
rect 30064 12792 30070 12804
rect 30147 12801 30159 12835
rect 30193 12832 30205 12835
rect 30742 12832 30748 12844
rect 30193 12804 30748 12832
rect 30193 12801 30205 12804
rect 30147 12795 30205 12801
rect 30742 12792 30748 12804
rect 30800 12792 30806 12844
rect 30852 12764 30880 12872
rect 30944 12872 31392 12900
rect 30944 12841 30972 12872
rect 31386 12860 31392 12872
rect 31444 12860 31450 12912
rect 32766 12900 32772 12912
rect 32232 12872 32772 12900
rect 30929 12835 30987 12841
rect 30929 12801 30941 12835
rect 30975 12801 30987 12835
rect 30929 12795 30987 12801
rect 31018 12792 31024 12844
rect 31076 12832 31082 12844
rect 31076 12804 31121 12832
rect 31076 12792 31082 12804
rect 31202 12792 31208 12844
rect 31260 12832 31266 12844
rect 31260 12804 31305 12832
rect 31260 12792 31266 12804
rect 31113 12767 31171 12773
rect 31113 12764 31125 12767
rect 29932 12736 30696 12764
rect 30852 12736 31125 12764
rect 28721 12727 28779 12733
rect 30668 12696 30696 12736
rect 31113 12733 31125 12736
rect 31159 12764 31171 12767
rect 32232 12764 32260 12872
rect 32766 12860 32772 12872
rect 32824 12860 32830 12912
rect 34082 12903 34140 12909
rect 34082 12869 34094 12903
rect 34128 12900 34140 12903
rect 34701 12903 34759 12909
rect 34701 12900 34713 12903
rect 34128 12872 34713 12900
rect 34128 12869 34140 12872
rect 34082 12863 34140 12869
rect 34701 12869 34713 12872
rect 34747 12900 34759 12903
rect 35710 12900 35716 12912
rect 34747 12872 35716 12900
rect 34747 12869 34759 12872
rect 34701 12863 34759 12869
rect 35710 12860 35716 12872
rect 35768 12860 35774 12912
rect 35820 12900 35848 12940
rect 35989 12937 36001 12971
rect 36035 12968 36047 12971
rect 36538 12968 36544 12980
rect 36035 12940 36544 12968
rect 36035 12937 36047 12940
rect 35989 12931 36047 12937
rect 36538 12928 36544 12940
rect 36596 12928 36602 12980
rect 38838 12968 38844 12980
rect 37844 12940 38844 12968
rect 37629 12903 37687 12909
rect 35820 12872 36492 12900
rect 32582 12832 32588 12844
rect 32543 12804 32588 12832
rect 32582 12792 32588 12804
rect 32640 12792 32646 12844
rect 32677 12835 32735 12841
rect 32677 12801 32689 12835
rect 32723 12832 32735 12835
rect 32784 12832 32812 12860
rect 32723 12804 32812 12832
rect 32723 12801 32735 12804
rect 32677 12795 32735 12801
rect 33134 12792 33140 12844
rect 33192 12832 33198 12844
rect 33597 12835 33655 12841
rect 33597 12832 33609 12835
rect 33192 12804 33609 12832
rect 33192 12792 33198 12804
rect 33597 12801 33609 12804
rect 33643 12832 33655 12835
rect 33778 12832 33784 12844
rect 33643 12804 33784 12832
rect 33643 12801 33655 12804
rect 33597 12795 33655 12801
rect 33778 12792 33784 12804
rect 33836 12792 33842 12844
rect 35342 12832 35348 12844
rect 35303 12804 35348 12832
rect 35342 12792 35348 12804
rect 35400 12792 35406 12844
rect 36354 12832 36360 12844
rect 35452 12804 36360 12832
rect 31159 12736 32260 12764
rect 31159 12733 31171 12736
rect 31113 12727 31171 12733
rect 32398 12724 32404 12776
rect 32456 12764 32462 12776
rect 32493 12767 32551 12773
rect 32493 12764 32505 12767
rect 32456 12736 32505 12764
rect 32456 12724 32462 12736
rect 32493 12733 32505 12736
rect 32539 12733 32551 12767
rect 32493 12727 32551 12733
rect 31202 12696 31208 12708
rect 28552 12668 30604 12696
rect 30668 12668 31208 12696
rect 28445 12659 28503 12665
rect 26510 12628 26516 12640
rect 26068 12600 26516 12628
rect 25777 12591 25835 12597
rect 26510 12588 26516 12600
rect 26568 12628 26574 12640
rect 27338 12628 27344 12640
rect 26568 12600 27344 12628
rect 26568 12588 26574 12600
rect 27338 12588 27344 12600
rect 27396 12588 27402 12640
rect 30282 12628 30288 12640
rect 30243 12600 30288 12628
rect 30282 12588 30288 12600
rect 30340 12588 30346 12640
rect 30576 12628 30604 12668
rect 31202 12656 31208 12668
rect 31260 12656 31266 12708
rect 31386 12656 31392 12708
rect 31444 12696 31450 12708
rect 32214 12696 32220 12708
rect 31444 12668 32220 12696
rect 31444 12656 31450 12668
rect 32214 12656 32220 12668
rect 32272 12656 32278 12708
rect 32600 12696 32628 12792
rect 32766 12724 32772 12776
rect 32824 12764 32830 12776
rect 32824 12736 32869 12764
rect 32824 12724 32830 12736
rect 33686 12724 33692 12776
rect 33744 12764 33750 12776
rect 33873 12767 33931 12773
rect 33873 12764 33885 12767
rect 33744 12736 33885 12764
rect 33744 12724 33750 12736
rect 33873 12733 33885 12736
rect 33919 12733 33931 12767
rect 33873 12727 33931 12733
rect 33965 12767 34023 12773
rect 33965 12733 33977 12767
rect 34011 12764 34023 12767
rect 35452 12764 35480 12804
rect 36354 12792 36360 12804
rect 36412 12792 36418 12844
rect 36464 12832 36492 12872
rect 37629 12869 37641 12903
rect 37675 12900 37687 12903
rect 37734 12900 37740 12912
rect 37675 12872 37740 12900
rect 37675 12869 37687 12872
rect 37629 12863 37687 12869
rect 37734 12860 37740 12872
rect 37792 12860 37798 12912
rect 37844 12909 37872 12940
rect 38838 12928 38844 12940
rect 38896 12928 38902 12980
rect 39942 12928 39948 12980
rect 40000 12968 40006 12980
rect 40221 12971 40279 12977
rect 40221 12968 40233 12971
rect 40000 12940 40233 12968
rect 40000 12928 40006 12940
rect 40221 12937 40233 12940
rect 40267 12937 40279 12971
rect 40221 12931 40279 12937
rect 41414 12928 41420 12980
rect 41472 12968 41478 12980
rect 41877 12971 41935 12977
rect 41877 12968 41889 12971
rect 41472 12940 41889 12968
rect 41472 12928 41478 12940
rect 41877 12937 41889 12940
rect 41923 12937 41935 12971
rect 53834 12968 53840 12980
rect 41877 12931 41935 12937
rect 48286 12940 53840 12968
rect 37829 12903 37887 12909
rect 37829 12869 37841 12903
rect 37875 12869 37887 12903
rect 48286 12900 48314 12940
rect 53834 12928 53840 12940
rect 53892 12928 53898 12980
rect 54202 12968 54208 12980
rect 54163 12940 54208 12968
rect 54202 12928 54208 12940
rect 54260 12928 54266 12980
rect 37829 12863 37887 12869
rect 37936 12872 39528 12900
rect 37936 12832 37964 12872
rect 36464 12804 37964 12832
rect 38378 12792 38384 12844
rect 38436 12832 38442 12844
rect 38545 12835 38603 12841
rect 38545 12832 38557 12835
rect 38436 12804 38557 12832
rect 38436 12792 38442 12804
rect 38545 12801 38557 12804
rect 38591 12801 38603 12835
rect 39500 12832 39528 12872
rect 39684 12872 48314 12900
rect 39684 12832 39712 12872
rect 40126 12832 40132 12844
rect 39500 12804 39712 12832
rect 40087 12804 40132 12832
rect 38545 12795 38603 12801
rect 40126 12792 40132 12804
rect 40184 12792 40190 12844
rect 40313 12835 40371 12841
rect 40313 12801 40325 12835
rect 40359 12832 40371 12835
rect 40494 12832 40500 12844
rect 40359 12804 40500 12832
rect 40359 12801 40371 12804
rect 40313 12795 40371 12801
rect 40494 12792 40500 12804
rect 40552 12832 40558 12844
rect 41782 12832 41788 12844
rect 40552 12804 41788 12832
rect 40552 12792 40558 12804
rect 41782 12792 41788 12804
rect 41840 12792 41846 12844
rect 54021 12835 54079 12841
rect 54021 12832 54033 12835
rect 51046 12804 54033 12832
rect 36262 12764 36268 12776
rect 34011 12736 35480 12764
rect 36223 12736 36268 12764
rect 34011 12733 34023 12736
rect 33965 12727 34023 12733
rect 36262 12724 36268 12736
rect 36320 12724 36326 12776
rect 38194 12724 38200 12776
rect 38252 12764 38258 12776
rect 38289 12767 38347 12773
rect 38289 12764 38301 12767
rect 38252 12736 38301 12764
rect 38252 12724 38258 12736
rect 38289 12733 38301 12736
rect 38335 12733 38347 12767
rect 38289 12727 38347 12733
rect 32600 12668 37780 12696
rect 32122 12628 32128 12640
rect 30576 12600 32128 12628
rect 32122 12588 32128 12600
rect 32180 12588 32186 12640
rect 32306 12628 32312 12640
rect 32267 12600 32312 12628
rect 32306 12588 32312 12600
rect 32364 12588 32370 12640
rect 34238 12628 34244 12640
rect 34199 12600 34244 12628
rect 34238 12588 34244 12600
rect 34296 12588 34302 12640
rect 34514 12588 34520 12640
rect 34572 12628 34578 12640
rect 37461 12631 37519 12637
rect 37461 12628 37473 12631
rect 34572 12600 37473 12628
rect 34572 12588 34578 12600
rect 37461 12597 37473 12600
rect 37507 12597 37519 12631
rect 37642 12628 37648 12640
rect 37603 12600 37648 12628
rect 37461 12591 37519 12597
rect 37642 12588 37648 12600
rect 37700 12588 37706 12640
rect 37752 12628 37780 12668
rect 39390 12656 39396 12708
rect 39448 12696 39454 12708
rect 39669 12699 39727 12705
rect 39669 12696 39681 12699
rect 39448 12668 39681 12696
rect 39448 12656 39454 12668
rect 39669 12665 39681 12668
rect 39715 12696 39727 12699
rect 51046 12696 51074 12804
rect 54021 12801 54033 12804
rect 54067 12801 54079 12835
rect 54021 12795 54079 12801
rect 39715 12668 51074 12696
rect 39715 12665 39727 12668
rect 39669 12659 39727 12665
rect 40773 12631 40831 12637
rect 40773 12628 40785 12631
rect 37752 12600 40785 12628
rect 40773 12597 40785 12600
rect 40819 12597 40831 12631
rect 40773 12591 40831 12597
rect 41417 12631 41475 12637
rect 41417 12597 41429 12631
rect 41463 12628 41475 12631
rect 41782 12628 41788 12640
rect 41463 12600 41788 12628
rect 41463 12597 41475 12600
rect 41417 12591 41475 12597
rect 41782 12588 41788 12600
rect 41840 12588 41846 12640
rect 1104 12538 54832 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 54832 12538
rect 1104 12464 54832 12486
rect 12069 12427 12127 12433
rect 12069 12393 12081 12427
rect 12115 12424 12127 12427
rect 13538 12424 13544 12436
rect 12115 12396 13544 12424
rect 12115 12393 12127 12396
rect 12069 12387 12127 12393
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 15838 12424 15844 12436
rect 15799 12396 15844 12424
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 17310 12424 17316 12436
rect 17271 12396 17316 12424
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 17586 12384 17592 12436
rect 17644 12424 17650 12436
rect 20806 12424 20812 12436
rect 17644 12396 20812 12424
rect 17644 12384 17650 12396
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 22554 12384 22560 12436
rect 22612 12424 22618 12436
rect 25961 12427 26019 12433
rect 22612 12396 24624 12424
rect 22612 12384 22618 12396
rect 13173 12359 13231 12365
rect 13173 12325 13185 12359
rect 13219 12356 13231 12359
rect 13725 12359 13783 12365
rect 13725 12356 13737 12359
rect 13219 12328 13737 12356
rect 13219 12325 13231 12328
rect 13173 12319 13231 12325
rect 13725 12325 13737 12328
rect 13771 12356 13783 12359
rect 16666 12356 16672 12368
rect 13771 12328 16672 12356
rect 13771 12325 13783 12328
rect 13725 12319 13783 12325
rect 16666 12316 16672 12328
rect 16724 12316 16730 12368
rect 17034 12316 17040 12368
rect 17092 12356 17098 12368
rect 17129 12359 17187 12365
rect 17129 12356 17141 12359
rect 17092 12328 17141 12356
rect 17092 12316 17098 12328
rect 17129 12325 17141 12328
rect 17175 12325 17187 12359
rect 17129 12319 17187 12325
rect 17862 12316 17868 12368
rect 17920 12356 17926 12368
rect 19794 12356 19800 12368
rect 17920 12328 19800 12356
rect 17920 12316 17926 12328
rect 19794 12316 19800 12328
rect 19852 12316 19858 12368
rect 22741 12359 22799 12365
rect 19904 12328 22094 12356
rect 15746 12288 15752 12300
rect 2746 12260 15752 12288
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12220 1915 12223
rect 2746 12220 2774 12260
rect 15746 12248 15752 12260
rect 15804 12248 15810 12300
rect 16117 12291 16175 12297
rect 16117 12257 16129 12291
rect 16163 12288 16175 12291
rect 18230 12288 18236 12300
rect 16163 12260 18236 12288
rect 16163 12257 16175 12260
rect 16117 12251 16175 12257
rect 18230 12248 18236 12260
rect 18288 12248 18294 12300
rect 18785 12291 18843 12297
rect 18785 12257 18797 12291
rect 18831 12288 18843 12291
rect 18874 12288 18880 12300
rect 18831 12260 18880 12288
rect 18831 12257 18843 12260
rect 18785 12251 18843 12257
rect 18874 12248 18880 12260
rect 18932 12248 18938 12300
rect 1903 12192 2774 12220
rect 1903 12189 1915 12192
rect 1857 12183 1915 12189
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 14369 12223 14427 12229
rect 14369 12220 14381 12223
rect 13964 12192 14381 12220
rect 13964 12180 13970 12192
rect 14369 12189 14381 12192
rect 14415 12189 14427 12223
rect 14369 12183 14427 12189
rect 15930 12180 15936 12232
rect 15988 12220 15994 12232
rect 16025 12223 16083 12229
rect 16025 12220 16037 12223
rect 15988 12192 16037 12220
rect 15988 12180 15994 12192
rect 16025 12189 16037 12192
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12189 16267 12223
rect 16209 12183 16267 12189
rect 16301 12223 16359 12229
rect 16301 12189 16313 12223
rect 16347 12220 16359 12223
rect 16574 12220 16580 12232
rect 16347 12192 16580 12220
rect 16347 12189 16359 12192
rect 16301 12183 16359 12189
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 14056 12124 15056 12152
rect 14056 12112 14062 12124
rect 15028 12096 15056 12124
rect 15194 12112 15200 12164
rect 15252 12152 15258 12164
rect 16114 12152 16120 12164
rect 15252 12124 16120 12152
rect 15252 12112 15258 12124
rect 16114 12112 16120 12124
rect 16172 12152 16178 12164
rect 16224 12152 16252 12183
rect 16574 12180 16580 12192
rect 16632 12180 16638 12232
rect 16666 12180 16672 12232
rect 16724 12220 16730 12232
rect 16853 12223 16911 12229
rect 16853 12220 16865 12223
rect 16724 12192 16865 12220
rect 16724 12180 16730 12192
rect 16853 12189 16865 12192
rect 16899 12220 16911 12223
rect 17126 12220 17132 12232
rect 16899 12192 17132 12220
rect 16899 12189 16911 12192
rect 16853 12183 16911 12189
rect 17126 12180 17132 12192
rect 17184 12220 17190 12232
rect 17862 12220 17868 12232
rect 17184 12192 17868 12220
rect 17184 12180 17190 12192
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 18196 12192 18613 12220
rect 18196 12180 18202 12192
rect 18601 12189 18613 12192
rect 18647 12220 18659 12223
rect 19242 12220 19248 12232
rect 18647 12192 19248 12220
rect 18647 12189 18659 12192
rect 18601 12183 18659 12189
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 19904 12229 19932 12328
rect 20622 12288 20628 12300
rect 19996 12260 20628 12288
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12189 19947 12223
rect 19889 12183 19947 12189
rect 19996 12152 20024 12260
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 21174 12288 21180 12300
rect 21135 12260 21180 12288
rect 21174 12248 21180 12260
rect 21232 12248 21238 12300
rect 22066 12288 22094 12328
rect 22741 12325 22753 12359
rect 22787 12356 22799 12359
rect 23198 12356 23204 12368
rect 22787 12328 23204 12356
rect 22787 12325 22799 12328
rect 22741 12319 22799 12325
rect 23198 12316 23204 12328
rect 23256 12316 23262 12368
rect 23753 12291 23811 12297
rect 23753 12288 23765 12291
rect 22066 12260 23765 12288
rect 23753 12257 23765 12260
rect 23799 12288 23811 12291
rect 23934 12288 23940 12300
rect 23799 12260 23940 12288
rect 23799 12257 23811 12260
rect 23753 12251 23811 12257
rect 23934 12248 23940 12260
rect 23992 12248 23998 12300
rect 24596 12297 24624 12396
rect 25961 12393 25973 12427
rect 26007 12424 26019 12427
rect 26602 12424 26608 12436
rect 26007 12396 26608 12424
rect 26007 12393 26019 12396
rect 25961 12387 26019 12393
rect 26602 12384 26608 12396
rect 26660 12384 26666 12436
rect 29086 12384 29092 12436
rect 29144 12424 29150 12436
rect 29730 12424 29736 12436
rect 29144 12396 29736 12424
rect 29144 12384 29150 12396
rect 29730 12384 29736 12396
rect 29788 12384 29794 12436
rect 30006 12384 30012 12436
rect 30064 12424 30070 12436
rect 31110 12424 31116 12436
rect 30064 12396 31116 12424
rect 30064 12384 30070 12396
rect 31110 12384 31116 12396
rect 31168 12384 31174 12436
rect 31478 12384 31484 12436
rect 31536 12424 31542 12436
rect 36173 12427 36231 12433
rect 31536 12396 35204 12424
rect 31536 12384 31542 12396
rect 26528 12328 27376 12356
rect 24029 12291 24087 12297
rect 24029 12257 24041 12291
rect 24075 12257 24087 12291
rect 24029 12251 24087 12257
rect 24581 12291 24639 12297
rect 24581 12257 24593 12291
rect 24627 12257 24639 12291
rect 24581 12251 24639 12257
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12220 20131 12223
rect 20714 12220 20720 12232
rect 20119 12192 20720 12220
rect 20119 12189 20131 12192
rect 20073 12183 20131 12189
rect 20714 12180 20720 12192
rect 20772 12180 20778 12232
rect 23658 12220 23664 12232
rect 23619 12192 23664 12220
rect 23658 12180 23664 12192
rect 23716 12180 23722 12232
rect 24044 12220 24072 12251
rect 25406 12220 25412 12232
rect 24044 12192 25412 12220
rect 25406 12180 25412 12192
rect 25464 12180 25470 12232
rect 26421 12223 26479 12229
rect 26421 12220 26433 12223
rect 25516 12192 26433 12220
rect 22186 12152 22192 12164
rect 16172 12124 16252 12152
rect 17880 12124 20024 12152
rect 22147 12124 22192 12152
rect 16172 12112 16178 12124
rect 1670 12084 1676 12096
rect 1631 12056 1676 12084
rect 1670 12044 1676 12056
rect 1728 12044 1734 12096
rect 12618 12084 12624 12096
rect 12579 12056 12624 12084
rect 12618 12044 12624 12056
rect 12676 12084 12682 12096
rect 13722 12084 13728 12096
rect 12676 12056 13728 12084
rect 12676 12044 12682 12056
rect 13722 12044 13728 12056
rect 13780 12044 13786 12096
rect 14461 12087 14519 12093
rect 14461 12053 14473 12087
rect 14507 12084 14519 12087
rect 14826 12084 14832 12096
rect 14507 12056 14832 12084
rect 14507 12053 14519 12056
rect 14461 12047 14519 12053
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 15010 12044 15016 12096
rect 15068 12084 15074 12096
rect 15289 12087 15347 12093
rect 15289 12084 15301 12087
rect 15068 12056 15301 12084
rect 15068 12044 15074 12056
rect 15289 12053 15301 12056
rect 15335 12053 15347 12087
rect 15289 12047 15347 12053
rect 15838 12044 15844 12096
rect 15896 12084 15902 12096
rect 17880 12084 17908 12124
rect 22186 12112 22192 12124
rect 22244 12112 22250 12164
rect 22462 12152 22468 12164
rect 22423 12124 22468 12152
rect 22462 12112 22468 12124
rect 22520 12112 22526 12164
rect 24026 12112 24032 12164
rect 24084 12152 24090 12164
rect 24826 12155 24884 12161
rect 24826 12152 24838 12155
rect 24084 12124 24838 12152
rect 24084 12112 24090 12124
rect 24826 12121 24838 12124
rect 24872 12121 24884 12155
rect 24826 12115 24884 12121
rect 25038 12112 25044 12164
rect 25096 12152 25102 12164
rect 25516 12152 25544 12192
rect 26421 12189 26433 12192
rect 26467 12189 26479 12223
rect 26421 12183 26479 12189
rect 26528 12152 26556 12328
rect 27154 12248 27160 12300
rect 27212 12288 27218 12300
rect 27249 12291 27307 12297
rect 27249 12288 27261 12291
rect 27212 12260 27261 12288
rect 27212 12248 27218 12260
rect 27249 12257 27261 12260
rect 27295 12257 27307 12291
rect 27348 12288 27376 12328
rect 28994 12316 29000 12368
rect 29052 12356 29058 12368
rect 29181 12359 29239 12365
rect 29181 12356 29193 12359
rect 29052 12328 29193 12356
rect 29052 12316 29058 12328
rect 29181 12325 29193 12328
rect 29227 12325 29239 12359
rect 34054 12356 34060 12368
rect 33967 12328 34060 12356
rect 29181 12319 29239 12325
rect 34054 12316 34060 12328
rect 34112 12356 34118 12368
rect 34238 12356 34244 12368
rect 34112 12328 34244 12356
rect 34112 12316 34118 12328
rect 34238 12316 34244 12328
rect 34296 12316 34302 12368
rect 34514 12316 34520 12368
rect 34572 12356 34578 12368
rect 34698 12356 34704 12368
rect 34572 12328 34704 12356
rect 34572 12316 34578 12328
rect 34698 12316 34704 12328
rect 34756 12316 34762 12368
rect 34790 12316 34796 12368
rect 34848 12356 34854 12368
rect 34977 12359 35035 12365
rect 34977 12356 34989 12359
rect 34848 12328 34989 12356
rect 34848 12316 34854 12328
rect 34977 12325 34989 12328
rect 35023 12325 35035 12359
rect 35176 12356 35204 12396
rect 36173 12393 36185 12427
rect 36219 12424 36231 12427
rect 36354 12424 36360 12436
rect 36219 12396 36360 12424
rect 36219 12393 36231 12396
rect 36173 12387 36231 12393
rect 36354 12384 36360 12396
rect 36412 12384 36418 12436
rect 37550 12384 37556 12436
rect 37608 12424 37614 12436
rect 37645 12427 37703 12433
rect 37645 12424 37657 12427
rect 37608 12396 37657 12424
rect 37608 12384 37614 12396
rect 37645 12393 37657 12396
rect 37691 12424 37703 12427
rect 37734 12424 37740 12436
rect 37691 12396 37740 12424
rect 37691 12393 37703 12396
rect 37645 12387 37703 12393
rect 37734 12384 37740 12396
rect 37792 12384 37798 12436
rect 38289 12427 38347 12433
rect 38289 12393 38301 12427
rect 38335 12424 38347 12427
rect 38378 12424 38384 12436
rect 38335 12396 38384 12424
rect 38335 12393 38347 12396
rect 38289 12387 38347 12393
rect 38378 12384 38384 12396
rect 38436 12384 38442 12436
rect 40034 12424 40040 12436
rect 39995 12396 40040 12424
rect 40034 12384 40040 12396
rect 40092 12384 40098 12436
rect 38657 12359 38715 12365
rect 38657 12356 38669 12359
rect 35176 12328 38669 12356
rect 34977 12319 35035 12325
rect 38657 12325 38669 12328
rect 38703 12325 38715 12359
rect 38657 12319 38715 12325
rect 38838 12316 38844 12368
rect 38896 12356 38902 12368
rect 40589 12359 40647 12365
rect 40589 12356 40601 12359
rect 38896 12328 40601 12356
rect 38896 12316 38902 12328
rect 40589 12325 40601 12328
rect 40635 12356 40647 12359
rect 41141 12359 41199 12365
rect 41141 12356 41153 12359
rect 40635 12328 41153 12356
rect 40635 12325 40647 12328
rect 40589 12319 40647 12325
rect 41141 12325 41153 12328
rect 41187 12325 41199 12359
rect 41141 12319 41199 12325
rect 27348 12260 28028 12288
rect 27249 12251 27307 12257
rect 26605 12223 26663 12229
rect 26605 12189 26617 12223
rect 26651 12220 26663 12223
rect 28000 12220 28028 12260
rect 28534 12248 28540 12300
rect 28592 12288 28598 12300
rect 29733 12291 29791 12297
rect 29733 12288 29745 12291
rect 28592 12260 29745 12288
rect 28592 12248 28598 12260
rect 29733 12257 29745 12260
rect 29779 12257 29791 12291
rect 29733 12251 29791 12257
rect 30834 12248 30840 12300
rect 30892 12288 30898 12300
rect 32122 12288 32128 12300
rect 30892 12260 32128 12288
rect 30892 12248 30898 12260
rect 32122 12248 32128 12260
rect 32180 12248 32186 12300
rect 28813 12223 28871 12229
rect 28813 12220 28825 12223
rect 26651 12192 27936 12220
rect 28000 12192 28825 12220
rect 26651 12189 26663 12192
rect 26605 12183 26663 12189
rect 25096 12124 25544 12152
rect 26252 12124 26556 12152
rect 25096 12112 25102 12124
rect 15896 12056 17908 12084
rect 15896 12044 15902 12056
rect 18046 12044 18052 12096
rect 18104 12084 18110 12096
rect 18141 12087 18199 12093
rect 18141 12084 18153 12087
rect 18104 12056 18153 12084
rect 18104 12044 18110 12056
rect 18141 12053 18153 12056
rect 18187 12053 18199 12087
rect 18506 12084 18512 12096
rect 18467 12056 18512 12084
rect 18141 12047 18199 12053
rect 18506 12044 18512 12056
rect 18564 12044 18570 12096
rect 19981 12087 20039 12093
rect 19981 12053 19993 12087
rect 20027 12084 20039 12087
rect 20070 12084 20076 12096
rect 20027 12056 20076 12084
rect 20027 12053 20039 12056
rect 19981 12047 20039 12053
rect 20070 12044 20076 12056
rect 20128 12044 20134 12096
rect 20162 12044 20168 12096
rect 20220 12084 20226 12096
rect 20533 12087 20591 12093
rect 20533 12084 20545 12087
rect 20220 12056 20545 12084
rect 20220 12044 20226 12056
rect 20533 12053 20545 12056
rect 20579 12053 20591 12087
rect 20898 12084 20904 12096
rect 20859 12056 20904 12084
rect 20533 12047 20591 12053
rect 20898 12044 20904 12056
rect 20956 12044 20962 12096
rect 20990 12044 20996 12096
rect 21048 12084 21054 12096
rect 22281 12087 22339 12093
rect 21048 12056 21093 12084
rect 21048 12044 21054 12056
rect 22281 12053 22293 12087
rect 22327 12084 22339 12087
rect 22370 12084 22376 12096
rect 22327 12056 22376 12084
rect 22327 12053 22339 12056
rect 22281 12047 22339 12053
rect 22370 12044 22376 12056
rect 22428 12044 22434 12096
rect 22830 12044 22836 12096
rect 22888 12084 22894 12096
rect 23014 12084 23020 12096
rect 22888 12056 23020 12084
rect 22888 12044 22894 12056
rect 23014 12044 23020 12056
rect 23072 12084 23078 12096
rect 24210 12084 24216 12096
rect 23072 12056 24216 12084
rect 23072 12044 23078 12056
rect 24210 12044 24216 12056
rect 24268 12084 24274 12096
rect 26252 12084 26280 12124
rect 24268 12056 26280 12084
rect 24268 12044 24274 12056
rect 26326 12044 26332 12096
rect 26384 12084 26390 12096
rect 26789 12087 26847 12093
rect 26789 12084 26801 12087
rect 26384 12056 26801 12084
rect 26384 12044 26390 12056
rect 26789 12053 26801 12056
rect 26835 12084 26847 12087
rect 26878 12084 26884 12096
rect 26835 12056 26884 12084
rect 26835 12053 26847 12056
rect 26789 12047 26847 12053
rect 26878 12044 26884 12056
rect 26936 12044 26942 12096
rect 27908 12093 27936 12192
rect 28813 12189 28825 12192
rect 28859 12189 28871 12223
rect 28813 12183 28871 12189
rect 28997 12223 29055 12229
rect 28997 12189 29009 12223
rect 29043 12220 29055 12223
rect 29638 12220 29644 12232
rect 29043 12192 29644 12220
rect 29043 12189 29055 12192
rect 28997 12183 29055 12189
rect 29638 12180 29644 12192
rect 29696 12180 29702 12232
rect 29822 12180 29828 12232
rect 29880 12220 29886 12232
rect 30742 12220 30748 12232
rect 29880 12192 30748 12220
rect 29880 12180 29886 12192
rect 30742 12180 30748 12192
rect 30800 12220 30806 12232
rect 33134 12220 33140 12232
rect 30800 12192 33140 12220
rect 30800 12180 30806 12192
rect 33134 12180 33140 12192
rect 33192 12220 33198 12232
rect 34072 12229 34100 12316
rect 37090 12288 37096 12300
rect 34341 12260 37096 12288
rect 34341 12229 34369 12260
rect 37090 12248 37096 12260
rect 37148 12248 37154 12300
rect 37734 12288 37740 12300
rect 37695 12260 37740 12288
rect 37734 12248 37740 12260
rect 37792 12248 37798 12300
rect 38286 12248 38292 12300
rect 38344 12288 38350 12300
rect 38749 12291 38807 12297
rect 38344 12260 38654 12288
rect 38344 12248 38350 12260
rect 33827 12223 33885 12229
rect 33827 12220 33839 12223
rect 33192 12192 33839 12220
rect 33192 12180 33198 12192
rect 33827 12189 33839 12192
rect 33873 12189 33885 12223
rect 33827 12183 33885 12189
rect 34057 12223 34115 12229
rect 34057 12189 34069 12223
rect 34103 12189 34115 12223
rect 34057 12183 34115 12189
rect 34240 12223 34298 12229
rect 34240 12189 34252 12223
rect 34286 12189 34298 12223
rect 34240 12183 34298 12189
rect 34333 12223 34391 12229
rect 34333 12189 34345 12223
rect 34379 12189 34391 12223
rect 36538 12220 36544 12232
rect 34333 12183 34391 12189
rect 34431 12192 36544 12220
rect 28902 12112 28908 12164
rect 28960 12152 28966 12164
rect 28960 12124 29224 12152
rect 28960 12112 28966 12124
rect 27893 12087 27951 12093
rect 27893 12053 27905 12087
rect 27939 12084 27951 12087
rect 28258 12084 28264 12096
rect 27939 12056 28264 12084
rect 27939 12053 27951 12056
rect 27893 12047 27951 12053
rect 28258 12044 28264 12056
rect 28316 12044 28322 12096
rect 29196 12084 29224 12124
rect 29270 12112 29276 12164
rect 29328 12152 29334 12164
rect 29978 12155 30036 12161
rect 29978 12152 29990 12155
rect 29328 12124 29990 12152
rect 29328 12112 29334 12124
rect 29978 12121 29990 12124
rect 30024 12121 30036 12155
rect 29978 12115 30036 12121
rect 30650 12112 30656 12164
rect 30708 12152 30714 12164
rect 31662 12152 31668 12164
rect 30708 12124 31668 12152
rect 30708 12112 30714 12124
rect 31662 12112 31668 12124
rect 31720 12112 31726 12164
rect 33502 12112 33508 12164
rect 33560 12152 33566 12164
rect 33965 12155 34023 12161
rect 33965 12152 33977 12155
rect 33560 12124 33977 12152
rect 33560 12112 33566 12124
rect 33965 12121 33977 12124
rect 34011 12121 34023 12155
rect 34255 12152 34283 12183
rect 34431 12152 34459 12192
rect 36538 12180 36544 12192
rect 36596 12180 36602 12232
rect 36722 12180 36728 12232
rect 36780 12220 36786 12232
rect 36817 12223 36875 12229
rect 36817 12220 36829 12223
rect 36780 12192 36829 12220
rect 36780 12180 36786 12192
rect 36817 12189 36829 12192
rect 36863 12220 36875 12223
rect 36906 12220 36912 12232
rect 36863 12192 36912 12220
rect 36863 12189 36875 12192
rect 36817 12183 36875 12189
rect 36906 12180 36912 12192
rect 36964 12180 36970 12232
rect 36998 12180 37004 12232
rect 37056 12220 37062 12232
rect 37461 12223 37519 12229
rect 37461 12220 37473 12223
rect 37056 12192 37473 12220
rect 37056 12180 37062 12192
rect 37461 12189 37473 12192
rect 37507 12189 37519 12223
rect 37461 12183 37519 12189
rect 35342 12152 35348 12164
rect 34255 12124 34459 12152
rect 35303 12124 35348 12152
rect 33965 12115 34023 12121
rect 35342 12112 35348 12124
rect 35400 12112 35406 12164
rect 37182 12112 37188 12164
rect 37240 12152 37246 12164
rect 38304 12152 38332 12248
rect 38470 12220 38476 12232
rect 38383 12192 38476 12220
rect 38470 12180 38476 12192
rect 38528 12180 38534 12232
rect 38626 12220 38654 12260
rect 38749 12257 38761 12291
rect 38795 12288 38807 12291
rect 39022 12288 39028 12300
rect 38795 12260 39028 12288
rect 38795 12257 38807 12260
rect 38749 12251 38807 12257
rect 39022 12248 39028 12260
rect 39080 12248 39086 12300
rect 39209 12223 39267 12229
rect 39209 12220 39221 12223
rect 38626 12192 39221 12220
rect 39209 12189 39221 12192
rect 39255 12189 39267 12223
rect 39209 12183 39267 12189
rect 39298 12180 39304 12232
rect 39356 12180 39362 12232
rect 49694 12180 49700 12232
rect 49752 12220 49758 12232
rect 54021 12223 54079 12229
rect 54021 12220 54033 12223
rect 49752 12192 54033 12220
rect 49752 12180 49758 12192
rect 54021 12189 54033 12192
rect 54067 12189 54079 12223
rect 54202 12220 54208 12232
rect 54163 12192 54208 12220
rect 54021 12183 54079 12189
rect 54202 12180 54208 12192
rect 54260 12180 54266 12232
rect 37240 12124 38332 12152
rect 38479 12152 38507 12180
rect 39316 12152 39344 12180
rect 39758 12152 39764 12164
rect 38479 12124 39764 12152
rect 37240 12112 37246 12124
rect 39758 12112 39764 12124
rect 39816 12112 39822 12164
rect 53190 12112 53196 12164
rect 53248 12152 53254 12164
rect 53285 12155 53343 12161
rect 53285 12152 53297 12155
rect 53248 12124 53297 12152
rect 53248 12112 53254 12124
rect 53285 12121 53297 12124
rect 53331 12121 53343 12155
rect 53466 12152 53472 12164
rect 53427 12124 53472 12152
rect 53285 12115 53343 12121
rect 53466 12112 53472 12124
rect 53524 12112 53530 12164
rect 53558 12112 53564 12164
rect 53616 12152 53622 12164
rect 54220 12152 54248 12180
rect 53616 12124 54248 12152
rect 53616 12112 53622 12124
rect 31570 12084 31576 12096
rect 29196 12056 31576 12084
rect 31570 12044 31576 12056
rect 31628 12044 31634 12096
rect 31754 12044 31760 12096
rect 31812 12084 31818 12096
rect 32769 12087 32827 12093
rect 32769 12084 32781 12087
rect 31812 12056 32781 12084
rect 31812 12044 31818 12056
rect 32769 12053 32781 12056
rect 32815 12084 32827 12087
rect 33594 12084 33600 12096
rect 32815 12056 33600 12084
rect 32815 12053 32827 12056
rect 32769 12047 32827 12053
rect 33594 12044 33600 12056
rect 33652 12044 33658 12096
rect 33689 12087 33747 12093
rect 33689 12053 33701 12087
rect 33735 12084 33747 12087
rect 34698 12084 34704 12096
rect 33735 12056 34704 12084
rect 33735 12053 33747 12056
rect 33689 12047 33747 12053
rect 34698 12044 34704 12056
rect 34756 12044 34762 12096
rect 34790 12044 34796 12096
rect 34848 12084 34854 12096
rect 34885 12087 34943 12093
rect 34885 12084 34897 12087
rect 34848 12056 34897 12084
rect 34848 12044 34854 12056
rect 34885 12053 34897 12056
rect 34931 12053 34943 12087
rect 34885 12047 34943 12053
rect 36630 12044 36636 12096
rect 36688 12084 36694 12096
rect 37277 12087 37335 12093
rect 37277 12084 37289 12087
rect 36688 12056 37289 12084
rect 36688 12044 36694 12056
rect 37277 12053 37289 12056
rect 37323 12053 37335 12087
rect 37277 12047 37335 12053
rect 37366 12044 37372 12096
rect 37424 12084 37430 12096
rect 37642 12084 37648 12096
rect 37424 12056 37648 12084
rect 37424 12044 37430 12056
rect 37642 12044 37648 12056
rect 37700 12084 37706 12096
rect 39301 12087 39359 12093
rect 39301 12084 39313 12087
rect 37700 12056 39313 12084
rect 37700 12044 37706 12056
rect 39301 12053 39313 12056
rect 39347 12053 39359 12087
rect 39301 12047 39359 12053
rect 39390 12044 39396 12096
rect 39448 12084 39454 12096
rect 41230 12084 41236 12096
rect 39448 12056 41236 12084
rect 39448 12044 39454 12056
rect 41230 12044 41236 12056
rect 41288 12044 41294 12096
rect 41782 12084 41788 12096
rect 41695 12056 41788 12084
rect 41782 12044 41788 12056
rect 41840 12084 41846 12096
rect 42518 12084 42524 12096
rect 41840 12056 42524 12084
rect 41840 12044 41846 12056
rect 42518 12044 42524 12056
rect 42576 12044 42582 12096
rect 52825 12087 52883 12093
rect 52825 12053 52837 12087
rect 52871 12084 52883 12087
rect 53484 12084 53512 12112
rect 52871 12056 53512 12084
rect 52871 12053 52883 12056
rect 52825 12047 52883 12053
rect 1104 11994 54832 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 54832 11994
rect 1104 11920 54832 11942
rect 12621 11883 12679 11889
rect 12621 11849 12633 11883
rect 12667 11880 12679 11883
rect 13354 11880 13360 11892
rect 12667 11852 13360 11880
rect 12667 11849 12679 11852
rect 12621 11843 12679 11849
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 15746 11880 15752 11892
rect 15707 11852 15752 11880
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 18506 11880 18512 11892
rect 16868 11852 18512 11880
rect 13725 11815 13783 11821
rect 13725 11781 13737 11815
rect 13771 11812 13783 11815
rect 16868 11812 16896 11852
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 18782 11840 18788 11892
rect 18840 11880 18846 11892
rect 18840 11852 19472 11880
rect 18840 11840 18846 11852
rect 13771 11784 16896 11812
rect 13771 11781 13783 11784
rect 13725 11775 13783 11781
rect 16942 11772 16948 11824
rect 17000 11812 17006 11824
rect 17037 11815 17095 11821
rect 17037 11812 17049 11815
rect 17000 11784 17049 11812
rect 17000 11772 17006 11784
rect 17037 11781 17049 11784
rect 17083 11781 17095 11815
rect 19444 11812 19472 11852
rect 20898 11840 20904 11892
rect 20956 11880 20962 11892
rect 26145 11883 26203 11889
rect 20956 11852 26096 11880
rect 20956 11840 20962 11852
rect 20134 11815 20192 11821
rect 20134 11812 20146 11815
rect 17037 11775 17095 11781
rect 17880 11784 19380 11812
rect 19444 11784 20146 11812
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11744 1915 11747
rect 15013 11747 15071 11753
rect 1903 11716 2774 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 2746 11676 2774 11716
rect 15013 11713 15025 11747
rect 15059 11744 15071 11747
rect 15838 11744 15844 11756
rect 15059 11716 15844 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11744 16083 11747
rect 17586 11744 17592 11756
rect 16071 11716 17592 11744
rect 16071 11713 16083 11716
rect 16025 11707 16083 11713
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 17880 11753 17908 11784
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11713 17923 11747
rect 17865 11707 17923 11713
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18121 11747 18179 11753
rect 18121 11744 18133 11747
rect 18012 11716 18133 11744
rect 18012 11704 18018 11716
rect 18121 11713 18133 11716
rect 18167 11713 18179 11747
rect 18121 11707 18179 11713
rect 19352 11688 19380 11784
rect 20134 11781 20146 11784
rect 20180 11781 20192 11815
rect 20134 11775 20192 11781
rect 22278 11772 22284 11824
rect 22336 11812 22342 11824
rect 22646 11812 22652 11824
rect 22336 11784 22652 11812
rect 22336 11772 22342 11784
rect 22646 11772 22652 11784
rect 22704 11772 22710 11824
rect 22833 11815 22891 11821
rect 22833 11781 22845 11815
rect 22879 11812 22891 11815
rect 23566 11812 23572 11824
rect 22879 11784 23572 11812
rect 22879 11781 22891 11784
rect 22833 11775 22891 11781
rect 23566 11772 23572 11784
rect 23624 11772 23630 11824
rect 23750 11772 23756 11824
rect 23808 11812 23814 11824
rect 25010 11815 25068 11821
rect 25010 11812 25022 11815
rect 23808 11784 25022 11812
rect 23808 11772 23814 11784
rect 25010 11781 25022 11784
rect 25056 11781 25068 11815
rect 26068 11812 26096 11852
rect 26145 11849 26157 11883
rect 26191 11880 26203 11883
rect 26234 11880 26240 11892
rect 26191 11852 26240 11880
rect 26191 11849 26203 11852
rect 26145 11843 26203 11849
rect 26234 11840 26240 11852
rect 26292 11840 26298 11892
rect 27338 11840 27344 11892
rect 27396 11880 27402 11892
rect 29638 11880 29644 11892
rect 27396 11852 29500 11880
rect 29599 11852 29644 11880
rect 27396 11840 27402 11852
rect 28902 11812 28908 11824
rect 26068 11784 28908 11812
rect 25010 11775 25068 11781
rect 28902 11772 28908 11784
rect 28960 11772 28966 11824
rect 29086 11812 29092 11824
rect 29047 11784 29092 11812
rect 29086 11772 29092 11784
rect 29144 11772 29150 11824
rect 19426 11704 19432 11756
rect 19484 11744 19490 11756
rect 20990 11744 20996 11756
rect 19484 11716 20996 11744
rect 19484 11704 19490 11716
rect 14737 11679 14795 11685
rect 14737 11676 14749 11679
rect 2746 11648 14749 11676
rect 14737 11645 14749 11648
rect 14783 11645 14795 11679
rect 14918 11676 14924 11688
rect 14879 11648 14924 11676
rect 14737 11639 14795 11645
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 15102 11676 15108 11688
rect 15063 11648 15108 11676
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 15194 11636 15200 11688
rect 15252 11676 15258 11688
rect 15930 11676 15936 11688
rect 15252 11648 15297 11676
rect 15891 11648 15936 11676
rect 15252 11636 15258 11648
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 16114 11676 16120 11688
rect 16075 11648 16120 11676
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 16209 11679 16267 11685
rect 16209 11645 16221 11679
rect 16255 11645 16267 11679
rect 16209 11639 16267 11645
rect 15286 11568 15292 11620
rect 15344 11608 15350 11620
rect 16224 11608 16252 11639
rect 19334 11636 19340 11688
rect 19392 11676 19398 11688
rect 19889 11679 19947 11685
rect 19889 11676 19901 11679
rect 19392 11648 19901 11676
rect 19392 11636 19398 11648
rect 19889 11645 19901 11648
rect 19935 11645 19947 11679
rect 19889 11639 19947 11645
rect 20916 11608 20944 11716
rect 20990 11704 20996 11716
rect 21048 11704 21054 11756
rect 24121 11747 24179 11753
rect 24121 11713 24133 11747
rect 24167 11744 24179 11747
rect 24854 11744 24860 11756
rect 24167 11716 24860 11744
rect 24167 11713 24179 11716
rect 24121 11707 24179 11713
rect 24854 11704 24860 11716
rect 24912 11704 24918 11756
rect 28281 11747 28339 11753
rect 28281 11713 28293 11747
rect 28327 11744 28339 11747
rect 28997 11747 29055 11753
rect 28327 11716 28948 11744
rect 28327 11713 28339 11716
rect 28281 11707 28339 11713
rect 22278 11636 22284 11688
rect 22336 11676 22342 11688
rect 22830 11676 22836 11688
rect 22336 11648 22836 11676
rect 22336 11636 22342 11648
rect 22830 11636 22836 11648
rect 22888 11636 22894 11688
rect 22925 11679 22983 11685
rect 22925 11645 22937 11679
rect 22971 11676 22983 11679
rect 23658 11676 23664 11688
rect 22971 11648 23664 11676
rect 22971 11645 22983 11648
rect 22925 11639 22983 11645
rect 23658 11636 23664 11648
rect 23716 11636 23722 11688
rect 24210 11636 24216 11688
rect 24268 11676 24274 11688
rect 24305 11679 24363 11685
rect 24305 11676 24317 11679
rect 24268 11648 24317 11676
rect 24268 11636 24274 11648
rect 24305 11645 24317 11648
rect 24351 11645 24363 11679
rect 24762 11676 24768 11688
rect 24723 11648 24768 11676
rect 24305 11639 24363 11645
rect 24762 11636 24768 11648
rect 24820 11636 24826 11688
rect 28534 11636 28540 11688
rect 28592 11676 28598 11688
rect 28592 11648 28685 11676
rect 28592 11636 28598 11648
rect 21269 11611 21327 11617
rect 21269 11608 21281 11611
rect 15344 11580 16252 11608
rect 16868 11580 17908 11608
rect 15344 11568 15350 11580
rect 1670 11540 1676 11552
rect 1631 11512 1676 11540
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 13170 11540 13176 11552
rect 13083 11512 13176 11540
rect 13170 11500 13176 11512
rect 13228 11540 13234 11552
rect 13722 11540 13728 11552
rect 13228 11512 13728 11540
rect 13228 11500 13234 11512
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 14277 11543 14335 11549
rect 14277 11509 14289 11543
rect 14323 11540 14335 11543
rect 16868 11540 16896 11580
rect 14323 11512 16896 11540
rect 16945 11543 17003 11549
rect 14323 11509 14335 11512
rect 14277 11503 14335 11509
rect 16945 11509 16957 11543
rect 16991 11540 17003 11543
rect 17770 11540 17776 11552
rect 16991 11512 17776 11540
rect 16991 11509 17003 11512
rect 16945 11503 17003 11509
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 17880 11540 17908 11580
rect 19168 11580 19932 11608
rect 20916 11580 21281 11608
rect 19168 11540 19196 11580
rect 17880 11512 19196 11540
rect 19242 11500 19248 11552
rect 19300 11540 19306 11552
rect 19904 11540 19932 11580
rect 21269 11577 21281 11580
rect 21315 11577 21327 11611
rect 22370 11608 22376 11620
rect 22331 11580 22376 11608
rect 21269 11571 21327 11577
rect 22370 11568 22376 11580
rect 22428 11568 22434 11620
rect 20898 11540 20904 11552
rect 19300 11512 19345 11540
rect 19904 11512 20904 11540
rect 19300 11500 19306 11512
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 22186 11500 22192 11552
rect 22244 11540 22250 11552
rect 23937 11543 23995 11549
rect 23937 11540 23949 11543
rect 22244 11512 23949 11540
rect 22244 11500 22250 11512
rect 23937 11509 23949 11512
rect 23983 11509 23995 11543
rect 27154 11540 27160 11552
rect 27115 11512 27160 11540
rect 23937 11503 23995 11509
rect 27154 11500 27160 11512
rect 27212 11500 27218 11552
rect 27614 11500 27620 11552
rect 27672 11540 27678 11552
rect 28552 11540 28580 11636
rect 27672 11512 28580 11540
rect 28920 11540 28948 11716
rect 28997 11713 29009 11747
rect 29043 11744 29055 11747
rect 29181 11747 29239 11753
rect 29043 11716 29132 11744
rect 29043 11713 29055 11716
rect 28997 11707 29055 11713
rect 29104 11688 29132 11716
rect 29181 11713 29193 11747
rect 29227 11713 29239 11747
rect 29472 11744 29500 11852
rect 29638 11840 29644 11852
rect 29696 11840 29702 11892
rect 30006 11880 30012 11892
rect 29967 11852 30012 11880
rect 30006 11840 30012 11852
rect 30064 11840 30070 11892
rect 31478 11880 31484 11892
rect 31439 11852 31484 11880
rect 31478 11840 31484 11852
rect 31536 11840 31542 11892
rect 31662 11840 31668 11892
rect 31720 11880 31726 11892
rect 32309 11883 32367 11889
rect 32309 11880 32321 11883
rect 31720 11852 32321 11880
rect 31720 11840 31726 11852
rect 32309 11849 32321 11852
rect 32355 11849 32367 11883
rect 32309 11843 32367 11849
rect 32861 11883 32919 11889
rect 32861 11849 32873 11883
rect 32907 11880 32919 11883
rect 33502 11880 33508 11892
rect 32907 11852 33508 11880
rect 32907 11849 32919 11852
rect 32861 11843 32919 11849
rect 33502 11840 33508 11852
rect 33560 11840 33566 11892
rect 34977 11883 35035 11889
rect 34977 11849 34989 11883
rect 35023 11880 35035 11883
rect 35894 11880 35900 11892
rect 35023 11852 35900 11880
rect 35023 11849 35035 11852
rect 34977 11843 35035 11849
rect 35894 11840 35900 11852
rect 35952 11840 35958 11892
rect 36817 11883 36875 11889
rect 36817 11849 36829 11883
rect 36863 11880 36875 11883
rect 37734 11880 37740 11892
rect 36863 11852 37740 11880
rect 36863 11849 36875 11852
rect 36817 11843 36875 11849
rect 37734 11840 37740 11852
rect 37792 11840 37798 11892
rect 39206 11880 39212 11892
rect 37844 11852 39212 11880
rect 29914 11772 29920 11824
rect 29972 11812 29978 11824
rect 30101 11815 30159 11821
rect 30101 11812 30113 11815
rect 29972 11784 30113 11812
rect 29972 11772 29978 11784
rect 30101 11781 30113 11784
rect 30147 11781 30159 11815
rect 30101 11775 30159 11781
rect 30742 11772 30748 11824
rect 30800 11812 30806 11824
rect 31754 11812 31760 11824
rect 30800 11784 30959 11812
rect 30800 11772 30806 11784
rect 29472 11716 30236 11744
rect 29181 11707 29239 11713
rect 29086 11636 29092 11688
rect 29144 11636 29150 11688
rect 29196 11608 29224 11707
rect 30208 11685 30236 11716
rect 30282 11704 30288 11756
rect 30340 11744 30346 11756
rect 30837 11747 30895 11753
rect 30837 11744 30849 11747
rect 30340 11716 30849 11744
rect 30340 11704 30346 11716
rect 30837 11713 30849 11716
rect 30883 11713 30895 11747
rect 30837 11707 30895 11713
rect 30193 11679 30251 11685
rect 30193 11645 30205 11679
rect 30239 11676 30251 11679
rect 30931 11676 30959 11784
rect 31036 11784 31760 11812
rect 31036 11753 31064 11784
rect 31754 11772 31760 11784
rect 31812 11772 31818 11824
rect 33996 11815 34054 11821
rect 33996 11781 34008 11815
rect 34042 11812 34054 11815
rect 37844 11812 37872 11852
rect 39206 11840 39212 11852
rect 39264 11840 39270 11892
rect 39298 11840 39304 11892
rect 39356 11880 39362 11892
rect 41138 11880 41144 11892
rect 39356 11852 41144 11880
rect 39356 11840 39362 11852
rect 41138 11840 41144 11852
rect 41196 11840 41202 11892
rect 41230 11840 41236 11892
rect 41288 11880 41294 11892
rect 41693 11883 41751 11889
rect 41693 11880 41705 11883
rect 41288 11852 41705 11880
rect 41288 11840 41294 11852
rect 41693 11849 41705 11852
rect 41739 11849 41751 11883
rect 53558 11880 53564 11892
rect 53519 11852 53564 11880
rect 41693 11843 41751 11849
rect 53558 11840 53564 11852
rect 53616 11840 53622 11892
rect 54202 11880 54208 11892
rect 54163 11852 54208 11880
rect 54202 11840 54208 11852
rect 54260 11840 54266 11892
rect 39114 11812 39120 11824
rect 34042 11784 36768 11812
rect 34042 11781 34054 11784
rect 33996 11775 34054 11781
rect 31021 11747 31079 11753
rect 31021 11713 31033 11747
rect 31067 11713 31079 11747
rect 31021 11707 31079 11713
rect 31113 11747 31171 11753
rect 31113 11713 31125 11747
rect 31159 11713 31171 11747
rect 31113 11707 31171 11713
rect 31128 11676 31156 11707
rect 31202 11704 31208 11756
rect 31260 11744 31266 11756
rect 34790 11744 34796 11756
rect 31260 11716 31305 11744
rect 34751 11716 34796 11744
rect 31260 11704 31266 11716
rect 34790 11704 34796 11716
rect 34848 11704 34854 11756
rect 35704 11747 35762 11753
rect 35704 11713 35716 11747
rect 35750 11744 35762 11747
rect 35986 11744 35992 11756
rect 35750 11716 35992 11744
rect 35750 11713 35762 11716
rect 35704 11707 35762 11713
rect 35986 11704 35992 11716
rect 36044 11704 36050 11756
rect 32582 11676 32588 11688
rect 30239 11648 30788 11676
rect 30931 11648 32588 11676
rect 30239 11645 30251 11648
rect 30193 11639 30251 11645
rect 29454 11608 29460 11620
rect 29196 11580 29460 11608
rect 29454 11568 29460 11580
rect 29512 11568 29518 11620
rect 30650 11608 30656 11620
rect 29564 11580 30656 11608
rect 29564 11540 29592 11580
rect 30650 11568 30656 11580
rect 30708 11568 30714 11620
rect 30760 11608 30788 11648
rect 32582 11636 32588 11648
rect 32640 11636 32646 11688
rect 34241 11679 34299 11685
rect 34241 11645 34253 11679
rect 34287 11676 34299 11679
rect 35342 11676 35348 11688
rect 34287 11648 35348 11676
rect 34287 11645 34299 11648
rect 34241 11639 34299 11645
rect 35342 11636 35348 11648
rect 35400 11676 35406 11688
rect 35437 11679 35495 11685
rect 35437 11676 35449 11679
rect 35400 11648 35449 11676
rect 35400 11636 35406 11648
rect 35437 11645 35449 11648
rect 35483 11645 35495 11679
rect 35437 11639 35495 11645
rect 32858 11608 32864 11620
rect 30760 11580 32864 11608
rect 32858 11568 32864 11580
rect 32916 11608 32922 11620
rect 33226 11608 33232 11620
rect 32916 11580 33232 11608
rect 32916 11568 32922 11580
rect 33226 11568 33232 11580
rect 33284 11568 33290 11620
rect 36740 11608 36768 11784
rect 37568 11784 37872 11812
rect 38488 11784 39120 11812
rect 36814 11704 36820 11756
rect 36872 11744 36878 11756
rect 37568 11753 37596 11784
rect 37553 11747 37611 11753
rect 37553 11744 37565 11747
rect 36872 11716 37565 11744
rect 36872 11704 36878 11716
rect 37553 11713 37565 11716
rect 37599 11713 37611 11747
rect 37553 11707 37611 11713
rect 37642 11704 37648 11756
rect 37700 11744 37706 11756
rect 37700 11716 37745 11744
rect 37700 11704 37706 11716
rect 38194 11704 38200 11756
rect 38252 11744 38258 11756
rect 38488 11753 38516 11784
rect 39114 11772 39120 11784
rect 39172 11812 39178 11824
rect 40954 11812 40960 11824
rect 39172 11784 40960 11812
rect 39172 11772 39178 11784
rect 40954 11772 40960 11784
rect 41012 11772 41018 11824
rect 51074 11812 51080 11824
rect 46216 11784 51080 11812
rect 38473 11747 38531 11753
rect 38473 11744 38485 11747
rect 38252 11716 38485 11744
rect 38252 11704 38258 11716
rect 38473 11713 38485 11716
rect 38519 11713 38531 11747
rect 38473 11707 38531 11713
rect 38740 11747 38798 11753
rect 38740 11713 38752 11747
rect 38786 11744 38798 11747
rect 40034 11744 40040 11756
rect 38786 11716 40040 11744
rect 38786 11713 38798 11716
rect 38740 11707 38798 11713
rect 40034 11704 40040 11716
rect 40092 11704 40098 11756
rect 40218 11704 40224 11756
rect 40276 11744 40282 11756
rect 40497 11747 40555 11753
rect 40497 11744 40509 11747
rect 40276 11716 40509 11744
rect 40276 11704 40282 11716
rect 40497 11713 40509 11716
rect 40543 11713 40555 11747
rect 46216 11744 46244 11784
rect 51074 11772 51080 11784
rect 51132 11772 51138 11824
rect 40497 11707 40555 11713
rect 40696 11716 46244 11744
rect 40696 11685 40724 11716
rect 46934 11704 46940 11756
rect 46992 11744 46998 11756
rect 54021 11747 54079 11753
rect 54021 11744 54033 11747
rect 46992 11716 54033 11744
rect 46992 11704 46998 11716
rect 54021 11713 54033 11716
rect 54067 11713 54079 11747
rect 54021 11707 54079 11713
rect 40681 11679 40739 11685
rect 40681 11645 40693 11679
rect 40727 11645 40739 11679
rect 40681 11639 40739 11645
rect 38378 11608 38384 11620
rect 36740 11580 38384 11608
rect 38378 11568 38384 11580
rect 38436 11568 38442 11620
rect 39853 11611 39911 11617
rect 39853 11577 39865 11611
rect 39899 11608 39911 11611
rect 40696 11608 40724 11639
rect 41138 11636 41144 11688
rect 41196 11676 41202 11688
rect 43622 11676 43628 11688
rect 41196 11648 43628 11676
rect 41196 11636 41202 11648
rect 43622 11636 43628 11648
rect 43680 11636 43686 11688
rect 39899 11580 40724 11608
rect 39899 11577 39911 11580
rect 39853 11571 39911 11577
rect 28920 11512 29592 11540
rect 27672 11500 27678 11512
rect 29638 11500 29644 11552
rect 29696 11540 29702 11552
rect 31846 11540 31852 11552
rect 29696 11512 31852 11540
rect 29696 11500 29702 11512
rect 31846 11500 31852 11512
rect 31904 11500 31910 11552
rect 33870 11500 33876 11552
rect 33928 11540 33934 11552
rect 37642 11540 37648 11552
rect 33928 11512 37648 11540
rect 33928 11500 33934 11512
rect 37642 11500 37648 11512
rect 37700 11500 37706 11552
rect 37829 11543 37887 11549
rect 37829 11509 37841 11543
rect 37875 11540 37887 11543
rect 39206 11540 39212 11552
rect 37875 11512 39212 11540
rect 37875 11509 37887 11512
rect 37829 11503 37887 11509
rect 39206 11500 39212 11512
rect 39264 11500 39270 11552
rect 40313 11543 40371 11549
rect 40313 11509 40325 11543
rect 40359 11540 40371 11543
rect 40494 11540 40500 11552
rect 40359 11512 40500 11540
rect 40359 11509 40371 11512
rect 40313 11503 40371 11509
rect 40494 11500 40500 11512
rect 40552 11500 40558 11552
rect 1104 11450 54832 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 54832 11450
rect 1104 11376 54832 11398
rect 15197 11339 15255 11345
rect 15197 11305 15209 11339
rect 15243 11336 15255 11339
rect 15286 11336 15292 11348
rect 15243 11308 15292 11336
rect 15243 11305 15255 11308
rect 15197 11299 15255 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 16117 11339 16175 11345
rect 16117 11305 16129 11339
rect 16163 11336 16175 11339
rect 16206 11336 16212 11348
rect 16163 11308 16212 11336
rect 16163 11305 16175 11308
rect 16117 11299 16175 11305
rect 16206 11296 16212 11308
rect 16264 11296 16270 11348
rect 23842 11336 23848 11348
rect 16960 11308 23848 11336
rect 14458 11228 14464 11280
rect 14516 11268 14522 11280
rect 15013 11271 15071 11277
rect 15013 11268 15025 11271
rect 14516 11240 15025 11268
rect 14516 11228 14522 11240
rect 15013 11237 15025 11240
rect 15059 11237 15071 11271
rect 15930 11268 15936 11280
rect 15891 11240 15936 11268
rect 15013 11231 15071 11237
rect 15930 11228 15936 11240
rect 15988 11228 15994 11280
rect 16853 11271 16911 11277
rect 16853 11237 16865 11271
rect 16899 11237 16911 11271
rect 16853 11231 16911 11237
rect 15286 11160 15292 11212
rect 15344 11200 15350 11212
rect 16114 11200 16120 11212
rect 15344 11172 16120 11200
rect 15344 11160 15350 11172
rect 16114 11160 16120 11172
rect 16172 11200 16178 11212
rect 16868 11200 16896 11231
rect 16172 11172 16896 11200
rect 16172 11160 16178 11172
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 11054 11132 11060 11144
rect 1903 11104 11060 11132
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 15010 11092 15016 11144
rect 15068 11132 15074 11144
rect 16960 11132 16988 11308
rect 23842 11296 23848 11308
rect 23900 11296 23906 11348
rect 25038 11336 25044 11348
rect 24999 11308 25044 11336
rect 25038 11296 25044 11308
rect 25096 11296 25102 11348
rect 27154 11296 27160 11348
rect 27212 11336 27218 11348
rect 35986 11336 35992 11348
rect 27212 11308 34008 11336
rect 35947 11308 35992 11336
rect 27212 11296 27218 11308
rect 18690 11228 18696 11280
rect 18748 11268 18754 11280
rect 20162 11268 20168 11280
rect 18748 11240 20168 11268
rect 18748 11228 18754 11240
rect 20162 11228 20168 11240
rect 20220 11228 20226 11280
rect 23934 11228 23940 11280
rect 23992 11268 23998 11280
rect 26145 11271 26203 11277
rect 26145 11268 26157 11271
rect 23992 11240 26157 11268
rect 23992 11228 23998 11240
rect 26145 11237 26157 11240
rect 26191 11237 26203 11271
rect 26145 11231 26203 11237
rect 25685 11203 25743 11209
rect 21284 11172 22416 11200
rect 15068 11104 16988 11132
rect 17037 11135 17095 11141
rect 15068 11092 15074 11104
rect 17037 11101 17049 11135
rect 17083 11101 17095 11135
rect 17037 11095 17095 11101
rect 17497 11135 17555 11141
rect 17497 11101 17509 11135
rect 17543 11132 17555 11135
rect 19334 11132 19340 11144
rect 17543 11104 19340 11132
rect 17543 11101 17555 11104
rect 17497 11095 17555 11101
rect 13173 11067 13231 11073
rect 13173 11033 13185 11067
rect 13219 11064 13231 11067
rect 13814 11064 13820 11076
rect 13219 11036 13820 11064
rect 13219 11033 13231 11036
rect 13173 11027 13231 11033
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 13998 11024 14004 11076
rect 14056 11064 14062 11076
rect 14737 11067 14795 11073
rect 14737 11064 14749 11067
rect 14056 11036 14749 11064
rect 14056 11024 14062 11036
rect 14737 11033 14749 11036
rect 14783 11064 14795 11067
rect 15657 11067 15715 11073
rect 15657 11064 15669 11067
rect 14783 11036 15669 11064
rect 14783 11033 14795 11036
rect 14737 11027 14795 11033
rect 15657 11033 15669 11036
rect 15703 11064 15715 11067
rect 15703 11036 16574 11064
rect 15703 11033 15715 11036
rect 15657 11027 15715 11033
rect 1670 10996 1676 11008
rect 1631 10968 1676 10996
rect 1670 10956 1676 10968
rect 1728 10956 1734 11008
rect 13722 10996 13728 11008
rect 13635 10968 13728 10996
rect 13722 10956 13728 10968
rect 13780 10996 13786 11008
rect 15838 10996 15844 11008
rect 13780 10968 15844 10996
rect 13780 10956 13786 10968
rect 15838 10956 15844 10968
rect 15896 10956 15902 11008
rect 16546 10996 16574 11036
rect 16666 11024 16672 11076
rect 16724 11064 16730 11076
rect 16850 11064 16856 11076
rect 16724 11036 16856 11064
rect 16724 11024 16730 11036
rect 16850 11024 16856 11036
rect 16908 11064 16914 11076
rect 17052 11064 17080 11095
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11132 19579 11135
rect 21284 11132 21312 11172
rect 19567 11104 21312 11132
rect 21361 11135 21419 11141
rect 19567 11101 19579 11104
rect 19521 11095 19579 11101
rect 21361 11101 21373 11135
rect 21407 11132 21419 11135
rect 22278 11132 22284 11144
rect 21407 11104 22284 11132
rect 21407 11101 21419 11104
rect 21361 11095 21419 11101
rect 22278 11092 22284 11104
rect 22336 11092 22342 11144
rect 22388 11132 22416 11172
rect 25685 11169 25697 11203
rect 25731 11200 25743 11203
rect 26602 11200 26608 11212
rect 25731 11172 26608 11200
rect 25731 11169 25743 11172
rect 25685 11163 25743 11169
rect 26602 11160 26608 11172
rect 26660 11160 26666 11212
rect 27724 11209 27752 11308
rect 29454 11268 29460 11280
rect 27908 11240 29460 11268
rect 27908 11209 27936 11240
rect 29454 11228 29460 11240
rect 29512 11268 29518 11280
rect 29825 11271 29883 11277
rect 29825 11268 29837 11271
rect 29512 11240 29837 11268
rect 29512 11228 29518 11240
rect 29825 11237 29837 11240
rect 29871 11237 29883 11271
rect 29825 11231 29883 11237
rect 31205 11271 31263 11277
rect 31205 11237 31217 11271
rect 31251 11268 31263 11271
rect 32030 11268 32036 11280
rect 31251 11240 32036 11268
rect 31251 11237 31263 11240
rect 31205 11231 31263 11237
rect 32030 11228 32036 11240
rect 32088 11228 32094 11280
rect 32309 11271 32367 11277
rect 32309 11237 32321 11271
rect 32355 11268 32367 11271
rect 33410 11268 33416 11280
rect 32355 11240 33416 11268
rect 32355 11237 32367 11240
rect 32309 11231 32367 11237
rect 33410 11228 33416 11240
rect 33468 11228 33474 11280
rect 33689 11271 33747 11277
rect 33689 11237 33701 11271
rect 33735 11268 33747 11271
rect 33870 11268 33876 11280
rect 33735 11240 33876 11268
rect 33735 11237 33747 11240
rect 33689 11231 33747 11237
rect 33870 11228 33876 11240
rect 33928 11228 33934 11280
rect 33980 11268 34008 11308
rect 35986 11296 35992 11308
rect 36044 11296 36050 11348
rect 37274 11336 37280 11348
rect 36280 11308 37280 11336
rect 33980 11240 35940 11268
rect 27709 11203 27767 11209
rect 27709 11169 27721 11203
rect 27755 11169 27767 11203
rect 27709 11163 27767 11169
rect 27893 11203 27951 11209
rect 27893 11169 27905 11203
rect 27939 11169 27951 11203
rect 27893 11163 27951 11169
rect 27982 11160 27988 11212
rect 28040 11200 28046 11212
rect 28040 11172 31156 11200
rect 28040 11160 28046 11172
rect 24946 11132 24952 11144
rect 22388 11104 24952 11132
rect 24946 11092 24952 11104
rect 25004 11132 25010 11144
rect 26326 11132 26332 11144
rect 25004 11104 26188 11132
rect 26287 11104 26332 11132
rect 25004 11092 25010 11104
rect 26160 11076 26188 11104
rect 26326 11092 26332 11104
rect 26384 11092 26390 11144
rect 26513 11135 26571 11141
rect 26513 11101 26525 11135
rect 26559 11132 26571 11135
rect 27062 11132 27068 11144
rect 26559 11104 27068 11132
rect 26559 11101 26571 11104
rect 26513 11095 26571 11101
rect 27062 11092 27068 11104
rect 27120 11132 27126 11144
rect 27430 11132 27436 11144
rect 27120 11104 27436 11132
rect 27120 11092 27126 11104
rect 27430 11092 27436 11104
rect 27488 11092 27494 11144
rect 27617 11135 27675 11141
rect 27617 11101 27629 11135
rect 27663 11132 27675 11135
rect 27663 11104 28580 11132
rect 27663 11101 27675 11104
rect 27617 11095 27675 11101
rect 17770 11073 17776 11076
rect 16908 11036 17080 11064
rect 16908 11024 16914 11036
rect 17764 11027 17776 11073
rect 17828 11064 17834 11076
rect 17828 11036 17864 11064
rect 17770 11024 17776 11027
rect 17828 11024 17834 11036
rect 20806 11024 20812 11076
rect 20864 11064 20870 11076
rect 21094 11067 21152 11073
rect 21094 11064 21106 11067
rect 20864 11036 21106 11064
rect 20864 11024 20870 11036
rect 21094 11033 21106 11036
rect 21140 11033 21152 11067
rect 21094 11027 21152 11033
rect 21450 11024 21456 11076
rect 21508 11064 21514 11076
rect 22526 11067 22584 11073
rect 22526 11064 22538 11067
rect 21508 11036 22538 11064
rect 21508 11024 21514 11036
rect 22526 11033 22538 11036
rect 22572 11033 22584 11067
rect 22526 11027 22584 11033
rect 22830 11024 22836 11076
rect 22888 11064 22894 11076
rect 24762 11064 24768 11076
rect 22888 11036 24768 11064
rect 22888 11024 22894 11036
rect 24762 11024 24768 11036
rect 24820 11024 24826 11076
rect 26142 11024 26148 11076
rect 26200 11064 26206 11076
rect 27632 11064 27660 11095
rect 26200 11036 27660 11064
rect 26200 11024 26206 11036
rect 17310 10996 17316 11008
rect 16546 10968 17316 10996
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 18598 10956 18604 11008
rect 18656 10996 18662 11008
rect 18877 10999 18935 11005
rect 18877 10996 18889 10999
rect 18656 10968 18889 10996
rect 18656 10956 18662 10968
rect 18877 10965 18889 10968
rect 18923 10965 18935 10999
rect 18877 10959 18935 10965
rect 19981 10999 20039 11005
rect 19981 10965 19993 10999
rect 20027 10996 20039 10999
rect 20070 10996 20076 11008
rect 20027 10968 20076 10996
rect 20027 10965 20039 10968
rect 19981 10959 20039 10965
rect 20070 10956 20076 10968
rect 20128 10956 20134 11008
rect 23658 10996 23664 11008
rect 23619 10968 23664 10996
rect 23658 10956 23664 10968
rect 23716 10956 23722 11008
rect 27249 10999 27307 11005
rect 27249 10965 27261 10999
rect 27295 10996 27307 10999
rect 27338 10996 27344 11008
rect 27295 10968 27344 10996
rect 27295 10965 27307 10968
rect 27249 10959 27307 10965
rect 27338 10956 27344 10968
rect 27396 10956 27402 11008
rect 28552 10996 28580 11104
rect 28626 11092 28632 11144
rect 28684 11132 28690 11144
rect 28813 11135 28871 11141
rect 28813 11132 28825 11135
rect 28684 11104 28825 11132
rect 28684 11092 28690 11104
rect 28813 11101 28825 11104
rect 28859 11101 28871 11135
rect 28813 11095 28871 11101
rect 29733 11135 29791 11141
rect 29733 11101 29745 11135
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 30009 11135 30067 11141
rect 30009 11101 30021 11135
rect 30055 11132 30067 11135
rect 30558 11132 30564 11144
rect 30055 11104 30420 11132
rect 30519 11104 30564 11132
rect 30055 11101 30067 11104
rect 30009 11095 30067 11101
rect 28718 11064 28724 11076
rect 28679 11036 28724 11064
rect 28718 11024 28724 11036
rect 28776 11024 28782 11076
rect 29638 11064 29644 11076
rect 28828 11036 29644 11064
rect 28828 10996 28856 11036
rect 29638 11024 29644 11036
rect 29696 11024 29702 11076
rect 29748 11064 29776 11095
rect 30190 11064 30196 11076
rect 29748 11036 30196 11064
rect 30190 11024 30196 11036
rect 30248 11024 30254 11076
rect 28552 10968 28856 10996
rect 30392 10996 30420 11104
rect 30558 11092 30564 11104
rect 30616 11092 30622 11144
rect 30742 11141 30748 11144
rect 30740 11132 30748 11141
rect 30703 11104 30748 11132
rect 30740 11095 30748 11104
rect 30742 11092 30748 11095
rect 30800 11092 30806 11144
rect 30834 11092 30840 11144
rect 30892 11132 30898 11144
rect 31018 11141 31024 11144
rect 30975 11135 31024 11141
rect 30892 11104 30937 11132
rect 30892 11092 30898 11104
rect 30975 11101 30987 11135
rect 31021 11101 31024 11135
rect 30975 11095 31024 11101
rect 31018 11092 31024 11095
rect 31076 11092 31082 11144
rect 31128 11132 31156 11172
rect 32858 11160 32864 11212
rect 32916 11200 32922 11212
rect 33137 11203 33195 11209
rect 33137 11200 33149 11203
rect 32916 11172 33149 11200
rect 32916 11160 32922 11172
rect 33137 11169 33149 11172
rect 33183 11169 33195 11203
rect 33137 11163 33195 11169
rect 31478 11132 31484 11144
rect 31128 11104 31484 11132
rect 31478 11092 31484 11104
rect 31536 11092 31542 11144
rect 31662 11132 31668 11144
rect 31623 11104 31668 11132
rect 31662 11092 31668 11104
rect 31720 11092 31726 11144
rect 31846 11132 31852 11144
rect 31807 11104 31852 11132
rect 31846 11092 31852 11104
rect 31904 11092 31910 11144
rect 31941 11135 31999 11141
rect 31941 11101 31953 11135
rect 31987 11101 31999 11135
rect 31941 11095 31999 11101
rect 31956 11064 31984 11095
rect 32030 11092 32036 11144
rect 32088 11132 32094 11144
rect 33321 11135 33379 11141
rect 32088 11104 32133 11132
rect 32088 11092 32094 11104
rect 33321 11101 33333 11135
rect 33367 11132 33379 11135
rect 33502 11132 33508 11144
rect 33367 11104 33508 11132
rect 33367 11101 33379 11104
rect 33321 11095 33379 11101
rect 33502 11092 33508 11104
rect 33560 11092 33566 11144
rect 33594 11092 33600 11144
rect 33652 11132 33658 11144
rect 34149 11135 34207 11141
rect 34149 11132 34161 11135
rect 33652 11104 34161 11132
rect 33652 11092 33658 11104
rect 34149 11101 34161 11104
rect 34195 11101 34207 11135
rect 34330 11132 34336 11144
rect 34291 11104 34336 11132
rect 34149 11095 34207 11101
rect 34330 11092 34336 11104
rect 34388 11092 34394 11144
rect 34790 11092 34796 11144
rect 34848 11132 34854 11144
rect 34977 11135 35035 11141
rect 34977 11132 34989 11135
rect 34848 11104 34989 11132
rect 34848 11092 34854 11104
rect 34977 11101 34989 11104
rect 35023 11132 35035 11135
rect 35802 11132 35808 11144
rect 35023 11104 35808 11132
rect 35023 11101 35035 11104
rect 34977 11095 35035 11101
rect 35802 11092 35808 11104
rect 35860 11092 35866 11144
rect 35912 11132 35940 11240
rect 36078 11228 36084 11280
rect 36136 11268 36142 11280
rect 36280 11277 36308 11308
rect 37274 11296 37280 11308
rect 37332 11296 37338 11348
rect 37366 11296 37372 11348
rect 37424 11336 37430 11348
rect 37826 11336 37832 11348
rect 37424 11308 37832 11336
rect 37424 11296 37430 11308
rect 37826 11296 37832 11308
rect 37884 11296 37890 11348
rect 38378 11296 38384 11348
rect 38436 11336 38442 11348
rect 39117 11339 39175 11345
rect 39117 11336 39129 11339
rect 38436 11308 39129 11336
rect 38436 11296 38442 11308
rect 39117 11305 39129 11308
rect 39163 11305 39175 11339
rect 40034 11336 40040 11348
rect 39995 11308 40040 11336
rect 39117 11299 39175 11305
rect 40034 11296 40040 11308
rect 40092 11296 40098 11348
rect 40954 11336 40960 11348
rect 40915 11308 40960 11336
rect 40954 11296 40960 11308
rect 41012 11296 41018 11348
rect 36265 11271 36323 11277
rect 36265 11268 36277 11271
rect 36136 11240 36277 11268
rect 36136 11228 36142 11240
rect 36265 11237 36277 11240
rect 36311 11237 36323 11271
rect 36265 11231 36323 11237
rect 36446 11228 36452 11280
rect 36504 11268 36510 11280
rect 40405 11271 40463 11277
rect 40405 11268 40417 11271
rect 36504 11240 40417 11268
rect 36504 11228 36510 11240
rect 40405 11237 40417 11240
rect 40451 11237 40463 11271
rect 54202 11268 54208 11280
rect 54163 11240 54208 11268
rect 40405 11231 40463 11237
rect 54202 11228 54208 11240
rect 54260 11228 54266 11280
rect 36357 11203 36415 11209
rect 36357 11169 36369 11203
rect 36403 11200 36415 11203
rect 37366 11200 37372 11212
rect 36403 11172 37372 11200
rect 36403 11169 36415 11172
rect 36357 11163 36415 11169
rect 37366 11160 37372 11172
rect 37424 11160 37430 11212
rect 40310 11200 40316 11212
rect 37476 11172 40316 11200
rect 36173 11135 36231 11141
rect 36173 11132 36185 11135
rect 35912 11104 36185 11132
rect 36173 11101 36185 11104
rect 36219 11101 36231 11135
rect 36449 11135 36507 11141
rect 36449 11134 36461 11135
rect 36372 11132 36461 11134
rect 36173 11095 36231 11101
rect 36280 11106 36461 11132
rect 36280 11104 36400 11106
rect 32582 11064 32588 11076
rect 31956 11036 32588 11064
rect 32582 11024 32588 11036
rect 32640 11024 32646 11076
rect 32950 11024 32956 11076
rect 33008 11064 33014 11076
rect 34241 11067 34299 11073
rect 34241 11064 34253 11067
rect 33008 11036 34253 11064
rect 33008 11024 33014 11036
rect 34241 11033 34253 11036
rect 34287 11033 34299 11067
rect 34241 11027 34299 11033
rect 34698 11024 34704 11076
rect 34756 11064 34762 11076
rect 36280 11064 36308 11104
rect 36449 11101 36461 11106
rect 36495 11101 36507 11135
rect 36630 11132 36636 11144
rect 36591 11104 36636 11132
rect 36449 11095 36507 11101
rect 36630 11092 36636 11104
rect 36688 11092 36694 11144
rect 37182 11092 37188 11144
rect 37240 11141 37246 11144
rect 37476 11141 37504 11172
rect 40310 11160 40316 11172
rect 40368 11160 40374 11212
rect 40494 11200 40500 11212
rect 40455 11172 40500 11200
rect 40494 11160 40500 11172
rect 40552 11160 40558 11212
rect 37240 11135 37289 11141
rect 37240 11101 37243 11135
rect 37277 11101 37289 11135
rect 37240 11095 37289 11101
rect 37461 11135 37519 11141
rect 37461 11101 37473 11135
rect 37507 11101 37519 11135
rect 37589 11135 37647 11141
rect 37589 11132 37601 11135
rect 37461 11095 37519 11101
rect 37568 11101 37601 11132
rect 37635 11101 37647 11135
rect 37568 11095 37647 11101
rect 37737 11135 37795 11141
rect 37737 11101 37749 11135
rect 37783 11132 37795 11135
rect 37826 11132 37832 11144
rect 37783 11104 37832 11132
rect 37783 11101 37795 11104
rect 37737 11095 37795 11101
rect 37240 11092 37246 11095
rect 34756 11036 36308 11064
rect 34756 11024 34762 11036
rect 36998 11024 37004 11076
rect 37056 11064 37062 11076
rect 37366 11064 37372 11076
rect 37056 11036 37228 11064
rect 37327 11036 37372 11064
rect 37056 11024 37062 11036
rect 32674 10996 32680 11008
rect 30392 10968 32680 10996
rect 32674 10956 32680 10968
rect 32732 10956 32738 11008
rect 33226 10996 33232 11008
rect 33187 10968 33232 10996
rect 33226 10956 33232 10968
rect 33284 10956 33290 11008
rect 33686 10956 33692 11008
rect 33744 10996 33750 11008
rect 35529 10999 35587 11005
rect 35529 10996 35541 10999
rect 33744 10968 35541 10996
rect 33744 10956 33750 10968
rect 35529 10965 35541 10968
rect 35575 10996 35587 10999
rect 35618 10996 35624 11008
rect 35575 10968 35624 10996
rect 35575 10965 35587 10968
rect 35529 10959 35587 10965
rect 35618 10956 35624 10968
rect 35676 10956 35682 11008
rect 36446 10956 36452 11008
rect 36504 10996 36510 11008
rect 37093 10999 37151 11005
rect 37093 10996 37105 10999
rect 36504 10968 37105 10996
rect 36504 10956 36510 10968
rect 37093 10965 37105 10968
rect 37139 10965 37151 10999
rect 37200 10996 37228 11036
rect 37366 11024 37372 11036
rect 37424 11024 37430 11076
rect 37568 11064 37596 11095
rect 37826 11092 37832 11104
rect 37884 11132 37890 11144
rect 37884 11104 38312 11132
rect 37884 11092 37890 11104
rect 37476 11036 37596 11064
rect 37476 10996 37504 11036
rect 38102 11024 38108 11076
rect 38160 11064 38166 11076
rect 38197 11067 38255 11073
rect 38197 11064 38209 11067
rect 38160 11036 38209 11064
rect 38160 11024 38166 11036
rect 38197 11033 38209 11036
rect 38243 11033 38255 11067
rect 38284 11064 38312 11104
rect 38378 11092 38384 11144
rect 38436 11132 38442 11144
rect 38562 11132 38568 11144
rect 38436 11104 38481 11132
rect 38523 11104 38568 11132
rect 38436 11092 38442 11104
rect 38562 11092 38568 11104
rect 38620 11092 38626 11144
rect 38654 11092 38660 11144
rect 38712 11132 38718 11144
rect 38712 11104 38757 11132
rect 38712 11092 38718 11104
rect 39206 11092 39212 11144
rect 39264 11132 39270 11144
rect 39301 11135 39359 11141
rect 39301 11132 39313 11135
rect 39264 11104 39313 11132
rect 39264 11092 39270 11104
rect 39301 11101 39313 11104
rect 39347 11101 39359 11135
rect 39301 11095 39359 11101
rect 39758 11092 39764 11144
rect 39816 11132 39822 11144
rect 40221 11135 40279 11141
rect 40221 11132 40233 11135
rect 39816 11104 40233 11132
rect 39816 11092 39822 11104
rect 40221 11101 40233 11104
rect 40267 11101 40279 11135
rect 40221 11095 40279 11101
rect 51074 11092 51080 11144
rect 51132 11132 51138 11144
rect 54021 11135 54079 11141
rect 54021 11132 54033 11135
rect 51132 11104 54033 11132
rect 51132 11092 51138 11104
rect 54021 11101 54033 11104
rect 54067 11101 54079 11135
rect 54021 11095 54079 11101
rect 53561 11067 53619 11073
rect 38284 11036 40264 11064
rect 38197 11027 38255 11033
rect 40236 11008 40264 11036
rect 53561 11033 53573 11067
rect 53607 11033 53619 11067
rect 53561 11027 53619 11033
rect 37200 10968 37504 10996
rect 37093 10959 37151 10965
rect 40218 10956 40224 11008
rect 40276 10956 40282 11008
rect 53576 10996 53604 11027
rect 54202 10996 54208 11008
rect 53576 10968 54208 10996
rect 54202 10956 54208 10968
rect 54260 10956 54266 11008
rect 1104 10906 54832 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 54832 10906
rect 1104 10832 54832 10854
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 14921 10795 14979 10801
rect 14921 10792 14933 10795
rect 11112 10764 14933 10792
rect 11112 10752 11118 10764
rect 14921 10761 14933 10764
rect 14967 10761 14979 10795
rect 14921 10755 14979 10761
rect 16301 10795 16359 10801
rect 16301 10761 16313 10795
rect 16347 10761 16359 10795
rect 16301 10755 16359 10761
rect 13998 10724 14004 10736
rect 13959 10696 14004 10724
rect 13998 10684 14004 10696
rect 14056 10684 14062 10736
rect 16316 10724 16344 10755
rect 16574 10752 16580 10804
rect 16632 10792 16638 10804
rect 16853 10795 16911 10801
rect 16853 10792 16865 10795
rect 16632 10764 16865 10792
rect 16632 10752 16638 10764
rect 16853 10761 16865 10764
rect 16899 10761 16911 10795
rect 16853 10755 16911 10761
rect 20990 10752 20996 10804
rect 21048 10792 21054 10804
rect 24673 10795 24731 10801
rect 21048 10764 24624 10792
rect 21048 10752 21054 10764
rect 17954 10724 17960 10736
rect 16316 10696 17960 10724
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 22830 10724 22836 10736
rect 19996 10696 22836 10724
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10656 1915 10659
rect 15010 10656 15016 10668
rect 1903 10628 15016 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10656 15255 10659
rect 16117 10659 16175 10665
rect 15243 10628 16068 10656
rect 15243 10625 15255 10628
rect 15197 10619 15255 10625
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10588 13599 10591
rect 13814 10588 13820 10600
rect 13587 10560 13820 10588
rect 13587 10557 13599 10560
rect 13541 10551 13599 10557
rect 13814 10548 13820 10560
rect 13872 10588 13878 10600
rect 14918 10588 14924 10600
rect 13872 10560 14924 10588
rect 13872 10548 13878 10560
rect 14918 10548 14924 10560
rect 14976 10588 14982 10600
rect 15105 10591 15163 10597
rect 15105 10588 15117 10591
rect 14976 10560 15117 10588
rect 14976 10548 14982 10560
rect 15105 10557 15117 10560
rect 15151 10557 15163 10591
rect 15286 10588 15292 10600
rect 15247 10560 15292 10588
rect 15105 10551 15163 10557
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 15381 10591 15439 10597
rect 15381 10557 15393 10591
rect 15427 10557 15439 10591
rect 16040 10588 16068 10628
rect 16117 10625 16129 10659
rect 16163 10656 16175 10659
rect 18046 10656 18052 10668
rect 16163 10628 18052 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18230 10616 18236 10668
rect 18288 10656 18294 10668
rect 19996 10665 20024 10696
rect 22830 10684 22836 10696
rect 22888 10684 22894 10736
rect 18397 10659 18455 10665
rect 18397 10656 18409 10659
rect 18288 10628 18409 10656
rect 18288 10616 18294 10628
rect 18397 10625 18409 10628
rect 18443 10625 18455 10659
rect 18397 10619 18455 10625
rect 19981 10659 20039 10665
rect 19981 10625 19993 10659
rect 20027 10625 20039 10659
rect 20990 10656 20996 10668
rect 20951 10628 20996 10656
rect 19981 10619 20039 10625
rect 20990 10616 20996 10628
rect 21048 10616 21054 10668
rect 22738 10656 22744 10668
rect 22699 10628 22744 10656
rect 22738 10616 22744 10628
rect 22796 10616 22802 10668
rect 23382 10656 23388 10668
rect 23295 10628 23388 10656
rect 23382 10616 23388 10628
rect 23440 10656 23446 10668
rect 23440 10628 24256 10656
rect 23440 10616 23446 10628
rect 16040 10560 17264 10588
rect 15381 10551 15439 10557
rect 14274 10520 14280 10532
rect 14235 10492 14280 10520
rect 14274 10480 14280 10492
rect 14332 10480 14338 10532
rect 14366 10480 14372 10532
rect 14424 10520 14430 10532
rect 15396 10520 15424 10551
rect 14424 10492 15424 10520
rect 14424 10480 14430 10492
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 16945 10523 17003 10529
rect 16945 10520 16957 10523
rect 15620 10492 16957 10520
rect 15620 10480 15626 10492
rect 16945 10489 16957 10492
rect 16991 10489 17003 10523
rect 17236 10520 17264 10560
rect 17310 10548 17316 10600
rect 17368 10588 17374 10600
rect 18141 10591 18199 10597
rect 17368 10560 17413 10588
rect 17368 10548 17374 10560
rect 18141 10557 18153 10591
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 18046 10520 18052 10532
rect 17236 10492 18052 10520
rect 16945 10483 17003 10489
rect 18046 10480 18052 10492
rect 18104 10480 18110 10532
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 14461 10455 14519 10461
rect 14461 10421 14473 10455
rect 14507 10452 14519 10455
rect 15194 10452 15200 10464
rect 14507 10424 15200 10452
rect 14507 10421 14519 10424
rect 14461 10415 14519 10421
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 18156 10452 18184 10551
rect 20070 10548 20076 10600
rect 20128 10588 20134 10600
rect 21085 10591 21143 10597
rect 21085 10588 21097 10591
rect 20128 10560 21097 10588
rect 20128 10548 20134 10560
rect 21085 10557 21097 10560
rect 21131 10557 21143 10591
rect 21085 10551 21143 10557
rect 21174 10548 21180 10600
rect 21232 10588 21238 10600
rect 22557 10591 22615 10597
rect 21232 10560 21277 10588
rect 21232 10548 21238 10560
rect 22557 10557 22569 10591
rect 22603 10588 22615 10591
rect 23014 10588 23020 10600
rect 22603 10560 23020 10588
rect 22603 10557 22615 10560
rect 22557 10551 22615 10557
rect 23014 10548 23020 10560
rect 23072 10548 23078 10600
rect 19242 10480 19248 10532
rect 19300 10520 19306 10532
rect 19521 10523 19579 10529
rect 19521 10520 19533 10523
rect 19300 10492 19533 10520
rect 19300 10480 19306 10492
rect 19521 10489 19533 10492
rect 19567 10489 19579 10523
rect 19521 10483 19579 10489
rect 20165 10523 20223 10529
rect 20165 10489 20177 10523
rect 20211 10520 20223 10523
rect 22462 10520 22468 10532
rect 20211 10492 22468 10520
rect 20211 10489 20223 10492
rect 20165 10483 20223 10489
rect 22462 10480 22468 10492
rect 22520 10480 22526 10532
rect 19334 10452 19340 10464
rect 18156 10424 19340 10452
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 20622 10452 20628 10464
rect 20583 10424 20628 10452
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 22097 10455 22155 10461
rect 22097 10421 22109 10455
rect 22143 10452 22155 10455
rect 22554 10452 22560 10464
rect 22143 10424 22560 10452
rect 22143 10421 22155 10424
rect 22097 10415 22155 10421
rect 22554 10412 22560 10424
rect 22612 10412 22618 10464
rect 22925 10455 22983 10461
rect 22925 10421 22937 10455
rect 22971 10452 22983 10455
rect 23842 10452 23848 10464
rect 22971 10424 23848 10452
rect 22971 10421 22983 10424
rect 22925 10415 22983 10421
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 24228 10452 24256 10628
rect 24596 10520 24624 10764
rect 24673 10761 24685 10795
rect 24719 10792 24731 10795
rect 24762 10792 24768 10804
rect 24719 10764 24768 10792
rect 24719 10761 24731 10764
rect 24673 10755 24731 10761
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 26418 10752 26424 10804
rect 26476 10792 26482 10804
rect 26605 10795 26663 10801
rect 26605 10792 26617 10795
rect 26476 10764 26617 10792
rect 26476 10752 26482 10764
rect 26605 10761 26617 10764
rect 26651 10761 26663 10795
rect 29178 10792 29184 10804
rect 29139 10764 29184 10792
rect 26605 10755 26663 10761
rect 29178 10752 29184 10764
rect 29236 10752 29242 10804
rect 30098 10792 30104 10804
rect 29564 10764 30104 10792
rect 26145 10727 26203 10733
rect 26145 10693 26157 10727
rect 26191 10724 26203 10727
rect 27154 10724 27160 10736
rect 26191 10696 27160 10724
rect 26191 10693 26203 10696
rect 26145 10687 26203 10693
rect 27154 10684 27160 10696
rect 27212 10684 27218 10736
rect 26234 10656 26240 10668
rect 26195 10628 26240 10656
rect 26234 10616 26240 10628
rect 26292 10616 26298 10668
rect 27338 10656 27344 10668
rect 27299 10628 27344 10656
rect 27338 10616 27344 10628
rect 27396 10616 27402 10668
rect 28166 10656 28172 10668
rect 28127 10628 28172 10656
rect 28166 10616 28172 10628
rect 28224 10616 28230 10668
rect 28997 10659 29055 10665
rect 28997 10625 29009 10659
rect 29043 10656 29055 10659
rect 29564 10656 29592 10764
rect 30098 10752 30104 10764
rect 30156 10752 30162 10804
rect 30193 10795 30251 10801
rect 30193 10761 30205 10795
rect 30239 10792 30251 10795
rect 31662 10792 31668 10804
rect 30239 10764 31668 10792
rect 30239 10761 30251 10764
rect 30193 10755 30251 10761
rect 31662 10752 31668 10764
rect 31720 10752 31726 10804
rect 32585 10795 32643 10801
rect 32585 10761 32597 10795
rect 32631 10792 32643 10795
rect 32766 10792 32772 10804
rect 32631 10764 32772 10792
rect 32631 10761 32643 10764
rect 32585 10755 32643 10761
rect 32766 10752 32772 10764
rect 32824 10752 32830 10804
rect 33965 10795 34023 10801
rect 33965 10761 33977 10795
rect 34011 10792 34023 10795
rect 34054 10792 34060 10804
rect 34011 10764 34060 10792
rect 34011 10761 34023 10764
rect 33965 10755 34023 10761
rect 34054 10752 34060 10764
rect 34112 10792 34118 10804
rect 35526 10792 35532 10804
rect 34112 10764 35532 10792
rect 34112 10752 34118 10764
rect 35526 10752 35532 10764
rect 35584 10752 35590 10804
rect 37550 10792 37556 10804
rect 37511 10764 37556 10792
rect 37550 10752 37556 10764
rect 37608 10752 37614 10804
rect 37734 10752 37740 10804
rect 37792 10792 37798 10804
rect 38930 10792 38936 10804
rect 37792 10764 38936 10792
rect 37792 10752 37798 10764
rect 38930 10752 38936 10764
rect 38988 10792 38994 10804
rect 40037 10795 40095 10801
rect 40037 10792 40049 10795
rect 38988 10764 40049 10792
rect 38988 10752 38994 10764
rect 40037 10761 40049 10764
rect 40083 10761 40095 10795
rect 40037 10755 40095 10761
rect 40405 10795 40463 10801
rect 40405 10761 40417 10795
rect 40451 10792 40463 10795
rect 40957 10795 41015 10801
rect 40957 10792 40969 10795
rect 40451 10764 40969 10792
rect 40451 10761 40463 10764
rect 40405 10755 40463 10761
rect 40957 10761 40969 10764
rect 41003 10761 41015 10795
rect 40957 10755 41015 10761
rect 41414 10752 41420 10804
rect 41472 10792 41478 10804
rect 41969 10795 42027 10801
rect 41969 10792 41981 10795
rect 41472 10764 41981 10792
rect 41472 10752 41478 10764
rect 41969 10761 41981 10764
rect 42015 10792 42027 10795
rect 42058 10792 42064 10804
rect 42015 10764 42064 10792
rect 42015 10761 42027 10764
rect 41969 10755 42027 10761
rect 42058 10752 42064 10764
rect 42116 10752 42122 10804
rect 29638 10684 29644 10736
rect 29696 10724 29702 10736
rect 29914 10724 29920 10736
rect 29696 10696 29920 10724
rect 29696 10684 29702 10696
rect 29914 10684 29920 10696
rect 29972 10724 29978 10736
rect 31297 10727 31355 10733
rect 29972 10696 30052 10724
rect 29972 10684 29978 10696
rect 29822 10656 29828 10668
rect 29043 10628 29592 10656
rect 29783 10628 29828 10656
rect 29043 10625 29055 10628
rect 28997 10619 29055 10625
rect 29822 10616 29828 10628
rect 29880 10616 29886 10668
rect 30024 10665 30052 10696
rect 31297 10693 31309 10727
rect 31343 10724 31355 10727
rect 31386 10724 31392 10736
rect 31343 10696 31392 10724
rect 31343 10693 31355 10696
rect 31297 10687 31355 10693
rect 31386 10684 31392 10696
rect 31444 10684 31450 10736
rect 31846 10684 31852 10736
rect 31904 10724 31910 10736
rect 37568 10724 37596 10752
rect 48958 10724 48964 10736
rect 31904 10696 37596 10724
rect 40236 10696 48964 10724
rect 31904 10684 31910 10696
rect 30009 10659 30067 10665
rect 30009 10625 30021 10659
rect 30055 10625 30067 10659
rect 30009 10619 30067 10625
rect 30653 10659 30711 10665
rect 30653 10625 30665 10659
rect 30699 10625 30711 10659
rect 30653 10619 30711 10625
rect 26053 10591 26111 10597
rect 26053 10557 26065 10591
rect 26099 10588 26111 10591
rect 26326 10588 26332 10600
rect 26099 10560 26332 10588
rect 26099 10557 26111 10560
rect 26053 10551 26111 10557
rect 26326 10548 26332 10560
rect 26384 10548 26390 10600
rect 27157 10591 27215 10597
rect 27157 10557 27169 10591
rect 27203 10588 27215 10591
rect 28353 10591 28411 10597
rect 28353 10588 28365 10591
rect 27203 10560 28365 10588
rect 27203 10557 27215 10560
rect 27157 10551 27215 10557
rect 28353 10557 28365 10560
rect 28399 10588 28411 10591
rect 29178 10588 29184 10600
rect 28399 10560 29184 10588
rect 28399 10557 28411 10560
rect 28353 10551 28411 10557
rect 29178 10548 29184 10560
rect 29236 10548 29242 10600
rect 29730 10588 29736 10600
rect 29691 10560 29736 10588
rect 29730 10548 29736 10560
rect 29788 10548 29794 10600
rect 29914 10548 29920 10600
rect 29972 10588 29978 10600
rect 30668 10588 30696 10619
rect 30742 10616 30748 10668
rect 30800 10656 30806 10668
rect 30837 10659 30895 10665
rect 30837 10656 30849 10659
rect 30800 10628 30849 10656
rect 30800 10616 30806 10628
rect 30837 10625 30849 10628
rect 30883 10625 30895 10659
rect 30837 10619 30895 10625
rect 30926 10616 30932 10668
rect 30984 10656 30990 10668
rect 31067 10659 31125 10665
rect 30984 10628 31029 10656
rect 30984 10616 30990 10628
rect 31067 10625 31079 10659
rect 31113 10656 31125 10659
rect 31478 10656 31484 10668
rect 31113 10628 31484 10656
rect 31113 10625 31125 10628
rect 31067 10619 31125 10625
rect 31478 10616 31484 10628
rect 31536 10616 31542 10668
rect 32766 10656 32772 10668
rect 32727 10628 32772 10656
rect 32766 10616 32772 10628
rect 32824 10616 32830 10668
rect 32953 10659 33011 10665
rect 32953 10625 32965 10659
rect 32999 10625 33011 10659
rect 32953 10619 33011 10625
rect 33045 10659 33103 10665
rect 33045 10625 33057 10659
rect 33091 10656 33103 10659
rect 33134 10656 33140 10668
rect 33091 10628 33140 10656
rect 33091 10625 33103 10628
rect 33045 10619 33103 10625
rect 32306 10588 32312 10600
rect 29972 10560 30017 10588
rect 30668 10560 32312 10588
rect 29972 10548 29978 10560
rect 32306 10548 32312 10560
rect 32364 10548 32370 10600
rect 32968 10588 32996 10619
rect 33134 10616 33140 10628
rect 33192 10616 33198 10668
rect 34790 10656 34796 10668
rect 33244 10628 34796 10656
rect 33244 10588 33272 10628
rect 34790 10616 34796 10628
rect 34848 10616 34854 10668
rect 35089 10659 35147 10665
rect 35089 10625 35101 10659
rect 35135 10656 35147 10659
rect 35802 10656 35808 10668
rect 35135 10628 35808 10656
rect 35135 10625 35147 10628
rect 35089 10619 35147 10625
rect 35802 10616 35808 10628
rect 35860 10616 35866 10668
rect 36173 10659 36231 10665
rect 36173 10625 36185 10659
rect 36219 10625 36231 10659
rect 36354 10656 36360 10668
rect 36315 10628 36360 10656
rect 36173 10619 36231 10625
rect 35342 10588 35348 10600
rect 32968 10560 33272 10588
rect 35303 10560 35348 10588
rect 35342 10548 35348 10560
rect 35400 10548 35406 10600
rect 32490 10520 32496 10532
rect 24596 10492 32496 10520
rect 32490 10480 32496 10492
rect 32548 10480 32554 10532
rect 36188 10520 36216 10619
rect 36354 10616 36360 10628
rect 36412 10616 36418 10668
rect 36446 10616 36452 10668
rect 36504 10656 36510 10668
rect 36504 10628 36549 10656
rect 36504 10616 36510 10628
rect 36541 10591 36599 10597
rect 36541 10557 36553 10591
rect 36587 10588 36599 10591
rect 36648 10588 36676 10696
rect 36725 10659 36783 10665
rect 36725 10625 36737 10659
rect 36771 10625 36783 10659
rect 37734 10656 37740 10668
rect 37695 10628 37740 10656
rect 36725 10619 36783 10625
rect 36587 10560 36676 10588
rect 36740 10588 36768 10619
rect 37734 10616 37740 10628
rect 37792 10616 37798 10668
rect 38470 10665 38476 10668
rect 38464 10619 38476 10665
rect 38528 10656 38534 10668
rect 40236 10665 40264 10696
rect 48958 10684 48964 10696
rect 49016 10684 49022 10736
rect 54202 10724 54208 10736
rect 54163 10696 54208 10724
rect 54202 10684 54208 10696
rect 54260 10684 54266 10736
rect 40221 10659 40279 10665
rect 38528 10628 38564 10656
rect 38470 10616 38476 10619
rect 38528 10616 38534 10628
rect 40221 10625 40233 10659
rect 40267 10625 40279 10659
rect 40221 10619 40279 10625
rect 40310 10616 40316 10668
rect 40368 10656 40374 10668
rect 40497 10659 40555 10665
rect 40497 10656 40509 10659
rect 40368 10628 40509 10656
rect 40368 10616 40374 10628
rect 40497 10625 40509 10628
rect 40543 10625 40555 10659
rect 40497 10619 40555 10625
rect 41414 10616 41420 10668
rect 41472 10656 41478 10668
rect 53466 10656 53472 10668
rect 41472 10628 41517 10656
rect 53427 10628 53472 10656
rect 41472 10616 41478 10628
rect 53466 10616 53472 10628
rect 53524 10616 53530 10668
rect 37918 10588 37924 10600
rect 36740 10560 37924 10588
rect 36587 10557 36599 10560
rect 36541 10551 36599 10557
rect 37918 10548 37924 10560
rect 37976 10548 37982 10600
rect 38194 10588 38200 10600
rect 38155 10560 38200 10588
rect 38194 10548 38200 10560
rect 38252 10548 38258 10600
rect 36188 10492 38240 10520
rect 25866 10452 25872 10464
rect 24228 10424 25872 10452
rect 25866 10412 25872 10424
rect 25924 10412 25930 10464
rect 27522 10452 27528 10464
rect 27483 10424 27528 10452
rect 27522 10412 27528 10424
rect 27580 10412 27586 10464
rect 27982 10452 27988 10464
rect 27943 10424 27988 10452
rect 27982 10412 27988 10424
rect 28040 10412 28046 10464
rect 30742 10412 30748 10464
rect 30800 10452 30806 10464
rect 36354 10452 36360 10464
rect 30800 10424 36360 10452
rect 30800 10412 30806 10424
rect 36354 10412 36360 10424
rect 36412 10412 36418 10464
rect 36906 10452 36912 10464
rect 36867 10424 36912 10452
rect 36906 10412 36912 10424
rect 36964 10412 36970 10464
rect 38212 10452 38240 10492
rect 53282 10480 53288 10532
rect 53340 10520 53346 10532
rect 54021 10523 54079 10529
rect 54021 10520 54033 10523
rect 53340 10492 54033 10520
rect 53340 10480 53346 10492
rect 54021 10489 54033 10492
rect 54067 10489 54079 10523
rect 54021 10483 54079 10489
rect 38378 10452 38384 10464
rect 38212 10424 38384 10452
rect 38378 10412 38384 10424
rect 38436 10412 38442 10464
rect 39574 10452 39580 10464
rect 39535 10424 39580 10452
rect 39574 10412 39580 10424
rect 39632 10412 39638 10464
rect 41322 10452 41328 10464
rect 41283 10424 41328 10452
rect 41322 10412 41328 10424
rect 41380 10412 41386 10464
rect 53374 10452 53380 10464
rect 53335 10424 53380 10452
rect 53374 10412 53380 10424
rect 53432 10412 53438 10464
rect 1104 10362 54832 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 54832 10362
rect 1104 10288 54832 10310
rect 13725 10251 13783 10257
rect 13725 10217 13737 10251
rect 13771 10248 13783 10251
rect 14366 10248 14372 10260
rect 13771 10220 14372 10248
rect 13771 10217 13783 10220
rect 13725 10211 13783 10217
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 15010 10248 15016 10260
rect 14971 10220 15016 10248
rect 15010 10208 15016 10220
rect 15068 10208 15074 10260
rect 16022 10208 16028 10260
rect 16080 10248 16086 10260
rect 16577 10251 16635 10257
rect 16577 10248 16589 10251
rect 16080 10220 16589 10248
rect 16080 10208 16086 10220
rect 16577 10217 16589 10220
rect 16623 10217 16635 10251
rect 17681 10251 17739 10257
rect 16577 10211 16635 10217
rect 16684 10220 17632 10248
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 13541 10183 13599 10189
rect 13541 10180 13553 10183
rect 13228 10152 13553 10180
rect 13228 10140 13234 10152
rect 13541 10149 13553 10152
rect 13587 10149 13599 10183
rect 13541 10143 13599 10149
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 16684 10180 16712 10220
rect 15344 10152 15516 10180
rect 15344 10140 15350 10152
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10112 13323 10115
rect 13998 10112 14004 10124
rect 13311 10084 14004 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 13998 10072 14004 10084
rect 14056 10072 14062 10124
rect 15381 10115 15439 10121
rect 15381 10081 15393 10115
rect 15427 10112 15439 10115
rect 15488 10112 15516 10152
rect 16040 10152 16712 10180
rect 16761 10183 16819 10189
rect 15654 10112 15660 10124
rect 15427 10084 15660 10112
rect 15427 10081 15439 10084
rect 15381 10075 15439 10081
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 15010 10044 15016 10056
rect 1903 10016 15016 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 15194 10044 15200 10056
rect 15155 10016 15200 10044
rect 15194 10004 15200 10016
rect 15252 10004 15258 10056
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 15304 9976 15332 10007
rect 15470 10004 15476 10056
rect 15528 10044 15534 10056
rect 15528 10016 15573 10044
rect 15528 10004 15534 10016
rect 16040 9976 16068 10152
rect 16761 10149 16773 10183
rect 16807 10180 16819 10183
rect 16850 10180 16856 10192
rect 16807 10152 16856 10180
rect 16807 10149 16819 10152
rect 16761 10143 16819 10149
rect 16850 10140 16856 10152
rect 16908 10140 16914 10192
rect 17604 10180 17632 10220
rect 17681 10217 17693 10251
rect 17727 10248 17739 10251
rect 17770 10248 17776 10260
rect 17727 10220 17776 10248
rect 17727 10217 17739 10220
rect 17681 10211 17739 10217
rect 17770 10208 17776 10220
rect 17828 10208 17834 10260
rect 17862 10208 17868 10260
rect 17920 10248 17926 10260
rect 18141 10251 18199 10257
rect 18141 10248 18153 10251
rect 17920 10220 18153 10248
rect 17920 10208 17926 10220
rect 18141 10217 18153 10220
rect 18187 10217 18199 10251
rect 19426 10248 19432 10260
rect 18141 10211 18199 10217
rect 18616 10220 19432 10248
rect 18616 10180 18644 10220
rect 19426 10208 19432 10220
rect 19484 10208 19490 10260
rect 19978 10208 19984 10260
rect 20036 10248 20042 10260
rect 20625 10251 20683 10257
rect 20625 10248 20637 10251
rect 20036 10220 20637 10248
rect 20036 10208 20042 10220
rect 20625 10217 20637 10220
rect 20671 10217 20683 10251
rect 20625 10211 20683 10217
rect 21634 10208 21640 10260
rect 21692 10248 21698 10260
rect 23566 10248 23572 10260
rect 21692 10220 23428 10248
rect 23527 10220 23572 10248
rect 21692 10208 21698 10220
rect 20990 10180 20996 10192
rect 17604 10152 18644 10180
rect 18708 10152 20996 10180
rect 16117 10115 16175 10121
rect 16117 10081 16129 10115
rect 16163 10112 16175 10115
rect 18708 10112 18736 10152
rect 20990 10140 20996 10152
rect 21048 10140 21054 10192
rect 23400 10180 23428 10220
rect 23566 10208 23572 10220
rect 23624 10208 23630 10260
rect 28350 10248 28356 10260
rect 28311 10220 28356 10248
rect 28350 10208 28356 10220
rect 28408 10208 28414 10260
rect 29181 10251 29239 10257
rect 29181 10217 29193 10251
rect 29227 10248 29239 10251
rect 29270 10248 29276 10260
rect 29227 10220 29276 10248
rect 29227 10217 29239 10220
rect 29181 10211 29239 10217
rect 29270 10208 29276 10220
rect 29328 10208 29334 10260
rect 29730 10208 29736 10260
rect 29788 10248 29794 10260
rect 32677 10251 32735 10257
rect 32677 10248 32689 10251
rect 29788 10220 32689 10248
rect 29788 10208 29794 10220
rect 32677 10217 32689 10220
rect 32723 10217 32735 10251
rect 32677 10211 32735 10217
rect 33686 10208 33692 10260
rect 33744 10248 33750 10260
rect 35805 10251 35863 10257
rect 33744 10220 35572 10248
rect 33744 10208 33750 10220
rect 23400 10152 25084 10180
rect 16163 10084 18736 10112
rect 18785 10115 18843 10121
rect 16163 10081 16175 10084
rect 16117 10075 16175 10081
rect 18785 10081 18797 10115
rect 18831 10112 18843 10115
rect 18874 10112 18880 10124
rect 18831 10084 18880 10112
rect 18831 10081 18843 10084
rect 18785 10075 18843 10081
rect 18874 10072 18880 10084
rect 18932 10112 18938 10124
rect 19981 10115 20039 10121
rect 19981 10112 19993 10115
rect 18932 10084 19993 10112
rect 18932 10072 18938 10084
rect 19981 10081 19993 10084
rect 20027 10112 20039 10115
rect 21174 10112 21180 10124
rect 20027 10084 21180 10112
rect 20027 10081 20039 10084
rect 19981 10075 20039 10081
rect 21174 10072 21180 10084
rect 21232 10072 21238 10124
rect 22094 10112 22100 10124
rect 21652 10084 22100 10112
rect 17037 10047 17095 10053
rect 17037 10013 17049 10047
rect 17083 10044 17095 10047
rect 17126 10044 17132 10056
rect 17083 10016 17132 10044
rect 17083 10013 17095 10016
rect 17037 10007 17095 10013
rect 17126 10004 17132 10016
rect 17184 10004 17190 10056
rect 17497 10047 17555 10053
rect 17497 10013 17509 10047
rect 17543 10044 17555 10047
rect 17862 10044 17868 10056
rect 17543 10016 17868 10044
rect 17543 10013 17555 10016
rect 17497 10007 17555 10013
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 17954 10004 17960 10056
rect 18012 10044 18018 10056
rect 19242 10044 19248 10056
rect 18012 10016 19248 10044
rect 18012 10004 18018 10016
rect 19242 10004 19248 10016
rect 19300 10044 19306 10056
rect 20809 10047 20867 10053
rect 19300 10016 19932 10044
rect 19300 10004 19306 10016
rect 19058 9976 19064 9988
rect 15304 9948 16068 9976
rect 18524 9948 19064 9976
rect 1670 9908 1676 9920
rect 1631 9880 1676 9908
rect 1670 9868 1676 9880
rect 1728 9868 1734 9920
rect 18524 9917 18552 9948
rect 19058 9936 19064 9948
rect 19116 9936 19122 9988
rect 19904 9985 19932 10016
rect 20809 10013 20821 10047
rect 20855 10044 20867 10047
rect 21266 10044 21272 10056
rect 20855 10016 21272 10044
rect 20855 10013 20867 10016
rect 20809 10007 20867 10013
rect 21266 10004 21272 10016
rect 21324 10004 21330 10056
rect 21652 10053 21680 10084
rect 22094 10072 22100 10084
rect 22152 10072 22158 10124
rect 21637 10047 21695 10053
rect 21637 10013 21649 10047
rect 21683 10013 21695 10047
rect 21637 10007 21695 10013
rect 22189 10047 22247 10053
rect 22189 10013 22201 10047
rect 22235 10044 22247 10047
rect 22278 10044 22284 10056
rect 22235 10016 22284 10044
rect 22235 10013 22247 10016
rect 22189 10007 22247 10013
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 22462 10053 22468 10056
rect 22456 10007 22468 10053
rect 22520 10044 22526 10056
rect 22520 10016 22556 10044
rect 22462 10004 22468 10007
rect 22520 10004 22526 10016
rect 23658 10004 23664 10056
rect 23716 10044 23722 10056
rect 24949 10047 25007 10053
rect 24949 10044 24961 10047
rect 23716 10016 24961 10044
rect 23716 10004 23722 10016
rect 24949 10013 24961 10016
rect 24995 10013 25007 10047
rect 24949 10007 25007 10013
rect 19889 9979 19947 9985
rect 19889 9945 19901 9979
rect 19935 9945 19947 9979
rect 19889 9939 19947 9945
rect 22554 9936 22560 9988
rect 22612 9976 22618 9988
rect 23934 9976 23940 9988
rect 22612 9948 23940 9976
rect 22612 9936 22618 9948
rect 23934 9936 23940 9948
rect 23992 9936 23998 9988
rect 25056 9920 25084 10152
rect 29822 10140 29828 10192
rect 29880 10180 29886 10192
rect 30193 10183 30251 10189
rect 30193 10180 30205 10183
rect 29880 10152 30205 10180
rect 29880 10140 29886 10152
rect 30193 10149 30205 10152
rect 30239 10180 30251 10183
rect 30374 10180 30380 10192
rect 30239 10152 30380 10180
rect 30239 10149 30251 10152
rect 30193 10143 30251 10149
rect 30374 10140 30380 10152
rect 30432 10180 30438 10192
rect 30558 10180 30564 10192
rect 30432 10152 30564 10180
rect 30432 10140 30438 10152
rect 30558 10140 30564 10152
rect 30616 10140 30622 10192
rect 30650 10140 30656 10192
rect 30708 10180 30714 10192
rect 31205 10183 31263 10189
rect 31205 10180 31217 10183
rect 30708 10152 31217 10180
rect 30708 10140 30714 10152
rect 31205 10149 31217 10152
rect 31251 10149 31263 10183
rect 33042 10180 33048 10192
rect 31205 10143 31263 10149
rect 31864 10152 33048 10180
rect 31864 10124 31892 10152
rect 33042 10140 33048 10152
rect 33100 10140 33106 10192
rect 33597 10183 33655 10189
rect 33597 10149 33609 10183
rect 33643 10149 33655 10183
rect 33597 10143 33655 10149
rect 25222 10112 25228 10124
rect 25183 10084 25228 10112
rect 25222 10072 25228 10084
rect 25280 10072 25286 10124
rect 27522 10072 27528 10124
rect 27580 10112 27586 10124
rect 31846 10112 31852 10124
rect 27580 10084 31432 10112
rect 31759 10084 31852 10112
rect 27580 10072 27586 10084
rect 25866 10004 25872 10056
rect 25924 10044 25930 10056
rect 26050 10044 26056 10056
rect 25924 10016 26056 10044
rect 25924 10004 25930 10016
rect 26050 10004 26056 10016
rect 26108 10004 26114 10056
rect 28258 10044 28264 10056
rect 28219 10016 28264 10044
rect 28258 10004 28264 10016
rect 28316 10004 28322 10056
rect 28994 10044 29000 10056
rect 28955 10016 29000 10044
rect 28994 10004 29000 10016
rect 29052 10004 29058 10056
rect 30377 10047 30435 10053
rect 30377 10013 30389 10047
rect 30423 10044 30435 10047
rect 30834 10044 30840 10056
rect 30423 10016 30840 10044
rect 30423 10013 30435 10016
rect 30377 10007 30435 10013
rect 30834 10004 30840 10016
rect 30892 10004 30898 10056
rect 31404 10053 31432 10084
rect 31846 10072 31852 10084
rect 31904 10072 31910 10124
rect 33612 10112 33640 10143
rect 34514 10140 34520 10192
rect 34572 10180 34578 10192
rect 35250 10180 35256 10192
rect 34572 10152 35256 10180
rect 34572 10140 34578 10152
rect 35250 10140 35256 10152
rect 35308 10140 35314 10192
rect 35544 10180 35572 10220
rect 35805 10217 35817 10251
rect 35851 10248 35863 10251
rect 36262 10248 36268 10260
rect 35851 10220 36268 10248
rect 35851 10217 35863 10220
rect 35805 10211 35863 10217
rect 36262 10208 36268 10220
rect 36320 10208 36326 10260
rect 38381 10251 38439 10257
rect 36372 10220 37504 10248
rect 36372 10180 36400 10220
rect 35544 10152 36400 10180
rect 37476 10180 37504 10220
rect 38381 10217 38393 10251
rect 38427 10248 38439 10251
rect 38470 10248 38476 10260
rect 38427 10220 38476 10248
rect 38427 10217 38439 10220
rect 38381 10211 38439 10217
rect 38470 10208 38476 10220
rect 38528 10208 38534 10260
rect 41322 10208 41328 10260
rect 41380 10248 41386 10260
rect 48314 10248 48320 10260
rect 41380 10220 48320 10248
rect 41380 10208 41386 10220
rect 48314 10208 48320 10220
rect 48372 10208 48378 10260
rect 54202 10248 54208 10260
rect 54163 10220 54208 10248
rect 54202 10208 54208 10220
rect 54260 10208 54266 10260
rect 38749 10183 38807 10189
rect 38749 10180 38761 10183
rect 37476 10152 38761 10180
rect 38749 10149 38761 10152
rect 38795 10149 38807 10183
rect 53466 10180 53472 10192
rect 53427 10152 53472 10180
rect 38749 10143 38807 10149
rect 53466 10140 53472 10152
rect 53524 10140 53530 10192
rect 34149 10115 34207 10121
rect 34149 10112 34161 10115
rect 32048 10084 33640 10112
rect 33888 10084 34161 10112
rect 32048 10053 32076 10084
rect 31389 10047 31447 10053
rect 31389 10013 31401 10047
rect 31435 10013 31447 10047
rect 31389 10007 31447 10013
rect 32033 10047 32091 10053
rect 32033 10013 32045 10047
rect 32079 10013 32091 10047
rect 32033 10007 32091 10013
rect 32766 10004 32772 10056
rect 32824 10044 32830 10056
rect 32861 10047 32919 10053
rect 32861 10044 32873 10047
rect 32824 10016 32873 10044
rect 32824 10004 32830 10016
rect 32861 10013 32873 10016
rect 32907 10013 32919 10047
rect 33134 10044 33140 10056
rect 33095 10016 33140 10044
rect 32861 10007 32919 10013
rect 33134 10004 33140 10016
rect 33192 10004 33198 10056
rect 33318 10004 33324 10056
rect 33376 10044 33382 10056
rect 33778 10044 33784 10056
rect 33376 10016 33784 10044
rect 33376 10004 33382 10016
rect 33778 10004 33784 10016
rect 33836 10044 33842 10056
rect 33888 10044 33916 10084
rect 34149 10081 34161 10084
rect 34195 10081 34207 10115
rect 34149 10075 34207 10081
rect 39574 10072 39580 10124
rect 39632 10112 39638 10124
rect 40405 10115 40463 10121
rect 40405 10112 40417 10115
rect 39632 10084 40417 10112
rect 39632 10072 39638 10084
rect 40405 10081 40417 10084
rect 40451 10112 40463 10115
rect 53009 10115 53067 10121
rect 40451 10084 41414 10112
rect 40451 10081 40463 10084
rect 40405 10075 40463 10081
rect 33836 10016 33916 10044
rect 33965 10047 34023 10053
rect 33836 10004 33842 10016
rect 33965 10013 33977 10047
rect 34011 10044 34023 10047
rect 34054 10044 34060 10056
rect 34011 10016 34060 10044
rect 34011 10013 34023 10016
rect 33965 10007 34023 10013
rect 26326 9936 26332 9988
rect 26384 9976 26390 9988
rect 27890 9976 27896 9988
rect 26384 9948 27896 9976
rect 26384 9936 26390 9948
rect 27890 9936 27896 9948
rect 27948 9936 27954 9988
rect 29914 9936 29920 9988
rect 29972 9976 29978 9988
rect 30282 9976 30288 9988
rect 29972 9948 30288 9976
rect 29972 9936 29978 9948
rect 30282 9936 30288 9948
rect 30340 9976 30346 9988
rect 30466 9976 30472 9988
rect 30340 9948 30472 9976
rect 30340 9936 30346 9948
rect 30466 9936 30472 9948
rect 30524 9936 30530 9988
rect 30742 9976 30748 9988
rect 30703 9948 30748 9976
rect 30742 9936 30748 9948
rect 30800 9936 30806 9988
rect 33045 9979 33103 9985
rect 33045 9945 33057 9979
rect 33091 9976 33103 9979
rect 33980 9976 34008 10007
rect 34054 10004 34060 10016
rect 34112 10004 34118 10056
rect 34974 10044 34980 10056
rect 34935 10016 34980 10044
rect 34974 10004 34980 10016
rect 35032 10004 35038 10056
rect 35069 10047 35127 10053
rect 35069 10013 35081 10047
rect 35115 10013 35127 10047
rect 35069 10007 35127 10013
rect 33091 9948 34008 9976
rect 33091 9945 33103 9948
rect 33045 9939 33103 9945
rect 34514 9936 34520 9988
rect 34572 9976 34578 9988
rect 35084 9976 35112 10007
rect 35618 10004 35624 10056
rect 35676 10044 35682 10056
rect 35713 10047 35771 10053
rect 35713 10044 35725 10047
rect 35676 10016 35725 10044
rect 35676 10004 35682 10016
rect 35713 10013 35725 10016
rect 35759 10013 35771 10047
rect 35713 10007 35771 10013
rect 35897 10047 35955 10053
rect 35897 10013 35909 10047
rect 35943 10013 35955 10047
rect 35897 10007 35955 10013
rect 36541 10047 36599 10053
rect 36541 10013 36553 10047
rect 36587 10044 36599 10047
rect 38194 10044 38200 10056
rect 36587 10016 38200 10044
rect 36587 10013 36599 10016
rect 36541 10007 36599 10013
rect 35526 9976 35532 9988
rect 34572 9948 35112 9976
rect 35176 9948 35532 9976
rect 34572 9936 34578 9948
rect 14553 9911 14611 9917
rect 14553 9877 14565 9911
rect 14599 9908 14611 9911
rect 18509 9911 18567 9917
rect 18509 9908 18521 9911
rect 14599 9880 18521 9908
rect 14599 9877 14611 9880
rect 14553 9871 14611 9877
rect 18509 9877 18521 9880
rect 18555 9877 18567 9911
rect 18509 9871 18567 9877
rect 18598 9868 18604 9920
rect 18656 9908 18662 9920
rect 19426 9908 19432 9920
rect 18656 9880 18701 9908
rect 19387 9880 19432 9908
rect 18656 9868 18662 9880
rect 19426 9868 19432 9880
rect 19484 9868 19490 9920
rect 19797 9911 19855 9917
rect 19797 9877 19809 9911
rect 19843 9908 19855 9911
rect 19978 9908 19984 9920
rect 19843 9880 19984 9908
rect 19843 9877 19855 9880
rect 19797 9871 19855 9877
rect 19978 9868 19984 9880
rect 20036 9908 20042 9920
rect 20254 9908 20260 9920
rect 20036 9880 20260 9908
rect 20036 9868 20042 9880
rect 20254 9868 20260 9880
rect 20312 9868 20318 9920
rect 21542 9908 21548 9920
rect 21503 9880 21548 9908
rect 21542 9868 21548 9880
rect 21600 9868 21606 9920
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 24581 9911 24639 9917
rect 24581 9908 24593 9911
rect 22152 9880 24593 9908
rect 22152 9868 22158 9880
rect 24581 9877 24593 9880
rect 24627 9877 24639 9911
rect 25038 9908 25044 9920
rect 24999 9880 25044 9908
rect 24581 9871 24639 9877
rect 25038 9868 25044 9880
rect 25096 9868 25102 9920
rect 27525 9911 27583 9917
rect 27525 9877 27537 9911
rect 27571 9908 27583 9911
rect 27614 9908 27620 9920
rect 27571 9880 27620 9908
rect 27571 9877 27583 9880
rect 27525 9871 27583 9877
rect 27614 9868 27620 9880
rect 27672 9868 27678 9920
rect 30374 9868 30380 9920
rect 30432 9908 30438 9920
rect 30561 9911 30619 9917
rect 30561 9908 30573 9911
rect 30432 9880 30573 9908
rect 30432 9868 30438 9880
rect 30561 9877 30573 9880
rect 30607 9877 30619 9911
rect 30561 9871 30619 9877
rect 32217 9911 32275 9917
rect 32217 9877 32229 9911
rect 32263 9908 32275 9911
rect 32950 9908 32956 9920
rect 32263 9880 32956 9908
rect 32263 9877 32275 9880
rect 32217 9871 32275 9877
rect 32950 9868 32956 9880
rect 33008 9868 33014 9920
rect 34054 9868 34060 9920
rect 34112 9908 34118 9920
rect 35176 9908 35204 9948
rect 35526 9936 35532 9948
rect 35584 9936 35590 9988
rect 34112 9880 35204 9908
rect 35253 9911 35311 9917
rect 34112 9868 34118 9880
rect 35253 9877 35265 9911
rect 35299 9908 35311 9911
rect 35434 9908 35440 9920
rect 35299 9880 35440 9908
rect 35299 9877 35311 9880
rect 35253 9871 35311 9877
rect 35434 9868 35440 9880
rect 35492 9868 35498 9920
rect 35912 9908 35940 10007
rect 38194 10004 38200 10016
rect 38252 10004 38258 10056
rect 38378 10004 38384 10056
rect 38436 10044 38442 10056
rect 38565 10047 38623 10053
rect 38565 10044 38577 10047
rect 38436 10016 38577 10044
rect 38436 10004 38442 10016
rect 38565 10013 38577 10016
rect 38611 10013 38623 10047
rect 38565 10007 38623 10013
rect 38841 10047 38899 10053
rect 38841 10013 38853 10047
rect 38887 10044 38899 10047
rect 40037 10047 40095 10053
rect 40037 10044 40049 10047
rect 38887 10016 40049 10044
rect 38887 10013 38899 10016
rect 38841 10007 38899 10013
rect 40037 10013 40049 10016
rect 40083 10013 40095 10047
rect 40218 10044 40224 10056
rect 40179 10016 40224 10044
rect 40037 10007 40095 10013
rect 40218 10004 40224 10016
rect 40276 10004 40282 10056
rect 41386 10044 41414 10084
rect 53009 10081 53021 10115
rect 53055 10112 53067 10115
rect 53558 10112 53564 10124
rect 53055 10084 53564 10112
rect 53055 10081 53067 10084
rect 53009 10075 53067 10081
rect 53558 10072 53564 10084
rect 53616 10072 53622 10124
rect 54021 10047 54079 10053
rect 54021 10044 54033 10047
rect 41386 10016 54033 10044
rect 54021 10013 54033 10016
rect 54067 10013 54079 10047
rect 54021 10007 54079 10013
rect 36808 9979 36866 9985
rect 36808 9945 36820 9979
rect 36854 9976 36866 9979
rect 36906 9976 36912 9988
rect 36854 9948 36912 9976
rect 36854 9945 36866 9948
rect 36808 9939 36866 9945
rect 36906 9936 36912 9948
rect 36964 9936 36970 9988
rect 39298 9976 39304 9988
rect 37752 9948 39304 9976
rect 37752 9908 37780 9948
rect 39298 9936 39304 9948
rect 39356 9936 39362 9988
rect 53374 9976 53380 9988
rect 41386 9948 53380 9976
rect 37918 9908 37924 9920
rect 35912 9880 37780 9908
rect 37879 9880 37924 9908
rect 37918 9868 37924 9880
rect 37976 9868 37982 9920
rect 38010 9868 38016 9920
rect 38068 9908 38074 9920
rect 41386 9908 41414 9948
rect 53374 9936 53380 9948
rect 53432 9936 53438 9988
rect 38068 9880 41414 9908
rect 38068 9868 38074 9880
rect 1104 9818 54832 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 54832 9818
rect 1104 9744 54832 9766
rect 15194 9664 15200 9716
rect 15252 9704 15258 9716
rect 15378 9704 15384 9716
rect 15252 9676 15384 9704
rect 15252 9664 15258 9676
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 17126 9664 17132 9716
rect 17184 9704 17190 9716
rect 17957 9707 18015 9713
rect 17957 9704 17969 9707
rect 17184 9676 17969 9704
rect 17184 9664 17190 9676
rect 17957 9673 17969 9676
rect 18003 9673 18015 9707
rect 17957 9667 18015 9673
rect 19613 9707 19671 9713
rect 19613 9673 19625 9707
rect 19659 9704 19671 9707
rect 20162 9704 20168 9716
rect 19659 9676 20168 9704
rect 19659 9673 19671 9676
rect 19613 9667 19671 9673
rect 20162 9664 20168 9676
rect 20220 9704 20226 9716
rect 20530 9704 20536 9716
rect 20220 9676 20536 9704
rect 20220 9664 20226 9676
rect 20530 9664 20536 9676
rect 20588 9664 20594 9716
rect 22830 9704 22836 9716
rect 22791 9676 22836 9704
rect 22830 9664 22836 9676
rect 22888 9664 22894 9716
rect 23124 9676 23704 9704
rect 13081 9639 13139 9645
rect 13081 9605 13093 9639
rect 13127 9636 13139 9639
rect 13998 9636 14004 9648
rect 13127 9608 14004 9636
rect 13127 9605 13139 9608
rect 13081 9599 13139 9605
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 16206 9636 16212 9648
rect 14292 9608 16212 9636
rect 14292 9577 14320 9608
rect 16206 9596 16212 9608
rect 16264 9596 16270 9648
rect 16301 9639 16359 9645
rect 16301 9605 16313 9639
rect 16347 9636 16359 9639
rect 17310 9636 17316 9648
rect 16347 9608 17172 9636
rect 17271 9608 17316 9636
rect 16347 9605 16359 9608
rect 16301 9599 16359 9605
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9568 1915 9571
rect 14277 9571 14335 9577
rect 1903 9540 14044 9568
rect 1903 9537 1915 9540
rect 1857 9531 1915 9537
rect 14016 9509 14044 9540
rect 14277 9537 14289 9571
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 14550 9568 14556 9580
rect 14507 9540 14556 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 15102 9568 15108 9580
rect 15063 9540 15108 9568
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 15311 9571 15369 9577
rect 15311 9537 15323 9571
rect 15357 9568 15369 9571
rect 15357 9540 17080 9568
rect 15357 9537 15369 9540
rect 15311 9531 15369 9537
rect 14001 9503 14059 9509
rect 14001 9469 14013 9503
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 14090 9460 14096 9512
rect 14148 9500 14154 9512
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 14148 9472 14197 9500
rect 14148 9460 14154 9472
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9500 14427 9503
rect 14642 9500 14648 9512
rect 14415 9472 14648 9500
rect 14415 9469 14427 9472
rect 14369 9463 14427 9469
rect 14642 9460 14648 9472
rect 14700 9500 14706 9512
rect 15197 9503 15255 9509
rect 15197 9500 15209 9503
rect 14700 9472 15209 9500
rect 14700 9460 14706 9472
rect 15197 9469 15209 9472
rect 15243 9469 15255 9503
rect 15197 9463 15255 9469
rect 15389 9503 15447 9509
rect 15389 9469 15401 9503
rect 15435 9500 15447 9503
rect 15746 9500 15752 9512
rect 15435 9472 15752 9500
rect 15435 9469 15447 9472
rect 15389 9463 15447 9469
rect 13354 9432 13360 9444
rect 13315 9404 13360 9432
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 13541 9435 13599 9441
rect 13541 9401 13553 9435
rect 13587 9432 13599 9435
rect 15102 9432 15108 9444
rect 13587 9404 15108 9432
rect 13587 9401 13599 9404
rect 13541 9395 13599 9401
rect 15102 9392 15108 9404
rect 15160 9392 15166 9444
rect 15212 9432 15240 9463
rect 15746 9460 15752 9472
rect 15804 9460 15810 9512
rect 16390 9460 16396 9512
rect 16448 9500 16454 9512
rect 16853 9503 16911 9509
rect 16853 9500 16865 9503
rect 16448 9472 16865 9500
rect 16448 9460 16454 9472
rect 16853 9469 16865 9472
rect 16899 9469 16911 9503
rect 16853 9463 16911 9469
rect 15654 9432 15660 9444
rect 15212 9404 15660 9432
rect 15654 9392 15660 9404
rect 15712 9392 15718 9444
rect 16574 9392 16580 9444
rect 16632 9432 16638 9444
rect 16945 9435 17003 9441
rect 16945 9432 16957 9435
rect 16632 9404 16957 9432
rect 16632 9392 16638 9404
rect 16945 9401 16957 9404
rect 16991 9401 17003 9435
rect 16945 9395 17003 9401
rect 1670 9364 1676 9376
rect 1631 9336 1676 9364
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 15010 9324 15016 9376
rect 15068 9364 15074 9376
rect 15565 9367 15623 9373
rect 15565 9364 15577 9367
rect 15068 9336 15577 9364
rect 15068 9324 15074 9336
rect 15565 9333 15577 9336
rect 15611 9333 15623 9367
rect 17052 9364 17080 9540
rect 17144 9500 17172 9608
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 23124 9636 23152 9676
rect 17788 9608 23152 9636
rect 23201 9639 23259 9645
rect 17788 9580 17816 9608
rect 23201 9605 23213 9639
rect 23247 9636 23259 9639
rect 23566 9636 23572 9648
rect 23247 9608 23572 9636
rect 23247 9605 23259 9608
rect 23201 9599 23259 9605
rect 23566 9596 23572 9608
rect 23624 9596 23630 9648
rect 23676 9636 23704 9676
rect 25038 9664 25044 9716
rect 25096 9704 25102 9716
rect 25096 9676 33088 9704
rect 25096 9664 25102 9676
rect 26326 9636 26332 9648
rect 23676 9608 26332 9636
rect 17770 9568 17776 9580
rect 17683 9540 17776 9568
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 18601 9571 18659 9577
rect 18601 9537 18613 9571
rect 18647 9568 18659 9571
rect 18690 9568 18696 9580
rect 18647 9540 18696 9568
rect 18647 9537 18659 9540
rect 18601 9531 18659 9537
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9568 19763 9571
rect 19978 9568 19984 9580
rect 19751 9540 19984 9568
rect 19751 9537 19763 9540
rect 19705 9531 19763 9537
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 20622 9568 20628 9580
rect 20583 9540 20628 9568
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9568 21327 9571
rect 22094 9568 22100 9580
rect 21315 9540 22100 9568
rect 21315 9537 21327 9540
rect 21269 9531 21327 9537
rect 22094 9528 22100 9540
rect 22152 9528 22158 9580
rect 22186 9528 22192 9580
rect 22244 9568 22250 9580
rect 22244 9540 22289 9568
rect 22244 9528 22250 9540
rect 23474 9528 23480 9580
rect 23532 9568 23538 9580
rect 24596 9577 24624 9608
rect 26326 9596 26332 9608
rect 26384 9596 26390 9648
rect 28350 9636 28356 9648
rect 27632 9608 28356 9636
rect 24121 9571 24179 9577
rect 24121 9568 24133 9571
rect 23532 9540 24133 9568
rect 23532 9528 23538 9540
rect 24121 9537 24133 9540
rect 24167 9537 24179 9571
rect 24121 9531 24179 9537
rect 24581 9571 24639 9577
rect 24581 9537 24593 9571
rect 24627 9537 24639 9571
rect 24581 9531 24639 9537
rect 24762 9528 24768 9580
rect 24820 9568 24826 9580
rect 24820 9540 24865 9568
rect 24820 9528 24826 9540
rect 25866 9528 25872 9580
rect 25924 9568 25930 9580
rect 26053 9571 26111 9577
rect 26053 9568 26065 9571
rect 25924 9540 26065 9568
rect 25924 9528 25930 9540
rect 26053 9537 26065 9540
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 26142 9528 26148 9580
rect 26200 9568 26206 9580
rect 26200 9540 26245 9568
rect 26200 9528 26206 9540
rect 27154 9528 27160 9580
rect 27212 9568 27218 9580
rect 27632 9577 27660 9608
rect 28350 9596 28356 9608
rect 28408 9596 28414 9648
rect 29454 9636 29460 9648
rect 28552 9608 29460 9636
rect 27525 9571 27583 9577
rect 27525 9568 27537 9571
rect 27212 9540 27537 9568
rect 27212 9528 27218 9540
rect 27525 9537 27537 9540
rect 27571 9537 27583 9571
rect 27525 9531 27583 9537
rect 27617 9571 27675 9577
rect 27890 9572 27896 9580
rect 27617 9537 27629 9571
rect 27663 9537 27675 9571
rect 27617 9531 27675 9537
rect 27816 9544 27896 9572
rect 19518 9500 19524 9512
rect 17144 9472 19524 9500
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 19610 9460 19616 9512
rect 19668 9500 19674 9512
rect 19797 9503 19855 9509
rect 19797 9500 19809 9503
rect 19668 9472 19809 9500
rect 19668 9460 19674 9472
rect 19797 9469 19809 9472
rect 19843 9469 19855 9503
rect 19797 9463 19855 9469
rect 23106 9460 23112 9512
rect 23164 9500 23170 9512
rect 23293 9503 23351 9509
rect 23293 9500 23305 9503
rect 23164 9472 23305 9500
rect 23164 9460 23170 9472
rect 23293 9469 23305 9472
rect 23339 9469 23351 9503
rect 23293 9463 23351 9469
rect 23385 9503 23443 9509
rect 23385 9469 23397 9503
rect 23431 9500 23443 9503
rect 23566 9500 23572 9512
rect 23431 9472 23572 9500
rect 23431 9469 23443 9472
rect 23385 9463 23443 9469
rect 23566 9460 23572 9472
rect 23624 9460 23630 9512
rect 24857 9503 24915 9509
rect 24857 9469 24869 9503
rect 24903 9469 24915 9503
rect 26326 9500 26332 9512
rect 26287 9472 26332 9500
rect 24857 9463 24915 9469
rect 18782 9432 18788 9444
rect 18743 9404 18788 9432
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 20070 9432 20076 9444
rect 18892 9404 20076 9432
rect 18892 9364 18920 9404
rect 20070 9392 20076 9404
rect 20128 9392 20134 9444
rect 20806 9432 20812 9444
rect 20767 9404 20812 9432
rect 20806 9392 20812 9404
rect 20864 9392 20870 9444
rect 21450 9432 21456 9444
rect 21411 9404 21456 9432
rect 21450 9392 21456 9404
rect 21508 9392 21514 9444
rect 22373 9435 22431 9441
rect 22373 9401 22385 9435
rect 22419 9432 22431 9435
rect 23750 9432 23756 9444
rect 22419 9404 23756 9432
rect 22419 9401 22431 9404
rect 22373 9395 22431 9401
rect 23750 9392 23756 9404
rect 23808 9392 23814 9444
rect 17052 9336 18920 9364
rect 15565 9327 15623 9333
rect 18966 9324 18972 9376
rect 19024 9364 19030 9376
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 19024 9336 19257 9364
rect 19024 9324 19030 9336
rect 19245 9333 19257 9336
rect 19291 9333 19303 9367
rect 19245 9327 19303 9333
rect 19794 9324 19800 9376
rect 19852 9364 19858 9376
rect 20714 9364 20720 9376
rect 19852 9336 20720 9364
rect 19852 9324 19858 9336
rect 20714 9324 20720 9336
rect 20772 9364 20778 9376
rect 21910 9364 21916 9376
rect 20772 9336 21916 9364
rect 20772 9324 20778 9336
rect 21910 9324 21916 9336
rect 21968 9324 21974 9376
rect 24118 9324 24124 9376
rect 24176 9364 24182 9376
rect 24872 9364 24900 9463
rect 26326 9460 26332 9472
rect 26384 9460 26390 9512
rect 27816 9509 27844 9544
rect 27890 9528 27896 9544
rect 27948 9528 27954 9580
rect 28552 9577 28580 9608
rect 29454 9596 29460 9608
rect 29512 9636 29518 9648
rect 30837 9639 30895 9645
rect 29512 9608 30604 9636
rect 29512 9596 29518 9608
rect 28537 9571 28595 9577
rect 28537 9537 28549 9571
rect 28583 9537 28595 9571
rect 28661 9571 28719 9577
rect 28661 9568 28673 9571
rect 28537 9531 28595 9537
rect 28644 9537 28673 9568
rect 28707 9537 28719 9571
rect 28644 9531 28719 9537
rect 27801 9503 27859 9509
rect 27801 9469 27813 9503
rect 27847 9469 27859 9503
rect 28442 9500 28448 9512
rect 28403 9472 28448 9500
rect 27801 9463 27859 9469
rect 28442 9460 28448 9472
rect 28500 9460 28506 9512
rect 28644 9500 28672 9531
rect 28902 9528 28908 9580
rect 28960 9572 28966 9580
rect 28960 9528 28994 9572
rect 29641 9571 29699 9577
rect 29641 9568 29653 9571
rect 28966 9500 28994 9528
rect 29288 9540 29653 9568
rect 29288 9500 29316 9540
rect 29641 9537 29653 9540
rect 29687 9537 29699 9571
rect 29641 9531 29699 9537
rect 29454 9500 29460 9512
rect 28644 9472 28856 9500
rect 28966 9472 29316 9500
rect 29415 9472 29460 9500
rect 25685 9435 25743 9441
rect 25685 9401 25697 9435
rect 25731 9432 25743 9435
rect 25958 9432 25964 9444
rect 25731 9404 25964 9432
rect 25731 9401 25743 9404
rect 25685 9395 25743 9401
rect 25958 9392 25964 9404
rect 26016 9392 26022 9444
rect 26970 9392 26976 9444
rect 27028 9432 27034 9444
rect 27157 9435 27215 9441
rect 27157 9432 27169 9435
rect 27028 9404 27169 9432
rect 27028 9392 27034 9404
rect 27157 9401 27169 9404
rect 27203 9401 27215 9435
rect 28828 9432 28856 9472
rect 29454 9460 29460 9472
rect 29512 9460 29518 9512
rect 29656 9500 29684 9531
rect 29730 9528 29736 9580
rect 29788 9568 29794 9580
rect 30374 9568 30380 9580
rect 29788 9540 30380 9568
rect 29788 9528 29794 9540
rect 30374 9528 30380 9540
rect 30432 9528 30438 9580
rect 30576 9577 30604 9608
rect 30837 9605 30849 9639
rect 30883 9636 30895 9639
rect 30926 9636 30932 9648
rect 30883 9608 30932 9636
rect 30883 9605 30895 9608
rect 30837 9599 30895 9605
rect 30926 9596 30932 9608
rect 30984 9636 30990 9648
rect 31110 9636 31116 9648
rect 30984 9608 31116 9636
rect 30984 9596 30990 9608
rect 31110 9596 31116 9608
rect 31168 9596 31174 9648
rect 31846 9636 31852 9648
rect 31496 9608 31852 9636
rect 30561 9571 30619 9577
rect 30561 9537 30573 9571
rect 30607 9537 30619 9571
rect 30561 9531 30619 9537
rect 30650 9528 30656 9580
rect 30708 9568 30714 9580
rect 31496 9577 31524 9608
rect 31846 9596 31852 9608
rect 31904 9596 31910 9648
rect 33060 9636 33088 9676
rect 33134 9664 33140 9716
rect 33192 9704 33198 9716
rect 33192 9676 35480 9704
rect 33192 9664 33198 9676
rect 34054 9636 34060 9648
rect 33060 9608 34060 9636
rect 34054 9596 34060 9608
rect 34112 9596 34118 9648
rect 35342 9636 35348 9648
rect 34624 9608 35348 9636
rect 31481 9571 31539 9577
rect 30708 9540 30753 9568
rect 30708 9528 30714 9540
rect 31481 9537 31493 9571
rect 31527 9537 31539 9571
rect 31481 9531 31539 9537
rect 31573 9571 31631 9577
rect 31573 9537 31585 9571
rect 31619 9568 31631 9571
rect 31662 9568 31668 9580
rect 31619 9540 31668 9568
rect 31619 9537 31631 9540
rect 31573 9531 31631 9537
rect 31662 9528 31668 9540
rect 31720 9528 31726 9580
rect 31754 9528 31760 9580
rect 31812 9568 31818 9580
rect 32030 9568 32036 9580
rect 31812 9540 32036 9568
rect 31812 9528 31818 9540
rect 32030 9528 32036 9540
rect 32088 9528 32094 9580
rect 32490 9528 32496 9580
rect 32548 9568 32554 9580
rect 33422 9571 33480 9577
rect 33422 9568 33434 9571
rect 32548 9540 33434 9568
rect 32548 9528 32554 9540
rect 33422 9537 33434 9540
rect 33468 9537 33480 9571
rect 33422 9531 33480 9537
rect 31110 9500 31116 9512
rect 29656 9472 31116 9500
rect 31110 9460 31116 9472
rect 31168 9500 31174 9512
rect 33686 9500 33692 9512
rect 31168 9472 31616 9500
rect 33647 9472 33692 9500
rect 31168 9460 31174 9472
rect 31588 9444 31616 9472
rect 33686 9460 33692 9472
rect 33744 9500 33750 9512
rect 34624 9509 34652 9608
rect 35342 9596 35348 9608
rect 35400 9596 35406 9648
rect 34698 9528 34704 9580
rect 34756 9568 34762 9580
rect 34865 9571 34923 9577
rect 34865 9568 34877 9571
rect 34756 9540 34877 9568
rect 34756 9528 34762 9540
rect 34865 9537 34877 9540
rect 34911 9537 34923 9571
rect 35452 9568 35480 9676
rect 35526 9664 35532 9716
rect 35584 9704 35590 9716
rect 38010 9704 38016 9716
rect 35584 9676 38016 9704
rect 35584 9664 35590 9676
rect 38010 9664 38016 9676
rect 38068 9664 38074 9716
rect 38286 9664 38292 9716
rect 38344 9664 38350 9716
rect 36538 9636 36544 9648
rect 36499 9608 36544 9636
rect 36538 9596 36544 9608
rect 36596 9596 36602 9648
rect 38304 9636 38332 9664
rect 39853 9639 39911 9645
rect 39853 9636 39865 9639
rect 38028 9608 39865 9636
rect 36449 9571 36507 9577
rect 36449 9568 36461 9571
rect 35452 9540 36461 9568
rect 34865 9531 34923 9537
rect 36449 9537 36461 9540
rect 36495 9537 36507 9571
rect 36449 9531 36507 9537
rect 36633 9571 36691 9577
rect 36633 9537 36645 9571
rect 36679 9568 36691 9571
rect 37550 9568 37556 9580
rect 36679 9540 37556 9568
rect 36679 9537 36691 9540
rect 36633 9531 36691 9537
rect 37550 9528 37556 9540
rect 37608 9528 37614 9580
rect 38028 9577 38056 9608
rect 39853 9605 39865 9608
rect 39899 9605 39911 9639
rect 39853 9599 39911 9605
rect 44450 9596 44456 9648
rect 44508 9636 44514 9648
rect 48317 9639 48375 9645
rect 48317 9636 48329 9639
rect 44508 9608 48329 9636
rect 44508 9596 44514 9608
rect 48317 9605 48329 9608
rect 48363 9605 48375 9639
rect 48317 9599 48375 9605
rect 38013 9571 38071 9577
rect 38013 9537 38025 9571
rect 38059 9537 38071 9571
rect 38013 9531 38071 9537
rect 38102 9528 38108 9580
rect 38160 9568 38166 9580
rect 38269 9571 38327 9577
rect 38269 9568 38281 9571
rect 38160 9540 38281 9568
rect 38160 9528 38166 9540
rect 38269 9537 38281 9540
rect 38315 9537 38327 9571
rect 48332 9568 48360 9599
rect 48406 9596 48412 9648
rect 48464 9636 48470 9648
rect 53374 9636 53380 9648
rect 48464 9608 53380 9636
rect 48464 9596 48470 9608
rect 53374 9596 53380 9608
rect 53432 9596 53438 9648
rect 48774 9568 48780 9580
rect 48332 9540 48780 9568
rect 38269 9531 38327 9537
rect 48774 9528 48780 9540
rect 48832 9528 48838 9580
rect 49050 9577 49056 9580
rect 49044 9531 49056 9577
rect 49108 9568 49114 9580
rect 50801 9571 50859 9577
rect 50801 9568 50813 9571
rect 49108 9540 49144 9568
rect 50172 9540 50813 9568
rect 49050 9528 49056 9531
rect 49108 9528 49114 9540
rect 34609 9503 34667 9509
rect 34609 9500 34621 9503
rect 33744 9472 34621 9500
rect 33744 9460 33750 9472
rect 34609 9469 34621 9472
rect 34655 9469 34667 9503
rect 34609 9463 34667 9469
rect 30837 9435 30895 9441
rect 30837 9432 30849 9435
rect 28828 9404 30849 9432
rect 27157 9395 27215 9401
rect 30837 9401 30849 9404
rect 30883 9401 30895 9435
rect 30837 9395 30895 9401
rect 31570 9392 31576 9444
rect 31628 9392 31634 9444
rect 32122 9392 32128 9444
rect 32180 9432 32186 9444
rect 32309 9435 32367 9441
rect 32309 9432 32321 9435
rect 32180 9404 32321 9432
rect 32180 9392 32186 9404
rect 32309 9401 32321 9404
rect 32355 9401 32367 9435
rect 37366 9432 37372 9444
rect 32309 9395 32367 9401
rect 35544 9404 37372 9432
rect 24176 9336 24900 9364
rect 24176 9324 24182 9336
rect 25774 9324 25780 9376
rect 25832 9364 25838 9376
rect 28718 9364 28724 9376
rect 25832 9336 28724 9364
rect 25832 9324 25838 9336
rect 28718 9324 28724 9336
rect 28776 9324 28782 9376
rect 28905 9367 28963 9373
rect 28905 9333 28917 9367
rect 28951 9364 28963 9367
rect 29822 9364 29828 9376
rect 28951 9336 29828 9364
rect 28951 9333 28963 9336
rect 28905 9327 28963 9333
rect 29822 9324 29828 9336
rect 29880 9324 29886 9376
rect 30098 9364 30104 9376
rect 30059 9336 30104 9364
rect 30098 9324 30104 9336
rect 30156 9324 30162 9376
rect 31754 9324 31760 9376
rect 31812 9364 31818 9376
rect 31812 9336 31857 9364
rect 31812 9324 31818 9336
rect 32030 9324 32036 9376
rect 32088 9364 32094 9376
rect 35544 9364 35572 9404
rect 37366 9392 37372 9404
rect 37424 9392 37430 9444
rect 50172 9441 50200 9540
rect 50801 9537 50813 9540
rect 50847 9537 50859 9571
rect 50801 9531 50859 9537
rect 50890 9528 50896 9580
rect 50948 9568 50954 9580
rect 53285 9571 53343 9577
rect 53285 9568 53297 9571
rect 50948 9540 53297 9568
rect 50948 9528 50954 9540
rect 53285 9537 53297 9540
rect 53331 9537 53343 9571
rect 53285 9531 53343 9537
rect 53469 9571 53527 9577
rect 53469 9537 53481 9571
rect 53515 9568 53527 9571
rect 53558 9568 53564 9580
rect 53515 9540 53564 9568
rect 53515 9537 53527 9540
rect 53469 9531 53527 9537
rect 53558 9528 53564 9540
rect 53616 9528 53622 9580
rect 54021 9571 54079 9577
rect 54021 9537 54033 9571
rect 54067 9537 54079 9571
rect 54021 9531 54079 9537
rect 50617 9503 50675 9509
rect 50617 9469 50629 9503
rect 50663 9469 50675 9503
rect 54036 9500 54064 9531
rect 50617 9463 50675 9469
rect 52288 9472 54064 9500
rect 50157 9435 50215 9441
rect 50157 9401 50169 9435
rect 50203 9401 50215 9435
rect 50157 9395 50215 9401
rect 35986 9364 35992 9376
rect 32088 9336 35572 9364
rect 35947 9336 35992 9364
rect 32088 9324 32094 9336
rect 35986 9324 35992 9336
rect 36044 9364 36050 9376
rect 36998 9364 37004 9376
rect 36044 9336 37004 9364
rect 36044 9324 36050 9336
rect 36998 9324 37004 9336
rect 37056 9324 37062 9376
rect 37553 9367 37611 9373
rect 37553 9333 37565 9367
rect 37599 9364 37611 9367
rect 37642 9364 37648 9376
rect 37599 9336 37648 9364
rect 37599 9333 37611 9336
rect 37553 9327 37611 9333
rect 37642 9324 37648 9336
rect 37700 9324 37706 9376
rect 39114 9324 39120 9376
rect 39172 9364 39178 9376
rect 39393 9367 39451 9373
rect 39393 9364 39405 9367
rect 39172 9336 39405 9364
rect 39172 9324 39178 9336
rect 39393 9333 39405 9336
rect 39439 9333 39451 9367
rect 39393 9327 39451 9333
rect 43622 9324 43628 9376
rect 43680 9364 43686 9376
rect 50430 9364 50436 9376
rect 43680 9336 50436 9364
rect 43680 9324 43686 9336
rect 50430 9324 50436 9336
rect 50488 9364 50494 9376
rect 50632 9364 50660 9463
rect 52288 9376 52316 9472
rect 54202 9432 54208 9444
rect 54163 9404 54208 9432
rect 54202 9392 54208 9404
rect 54260 9392 54266 9444
rect 50488 9336 50660 9364
rect 50985 9367 51043 9373
rect 50488 9324 50494 9336
rect 50985 9333 50997 9367
rect 51031 9364 51043 9367
rect 51626 9364 51632 9376
rect 51031 9336 51632 9364
rect 51031 9333 51043 9336
rect 50985 9327 51043 9333
rect 51626 9324 51632 9336
rect 51684 9324 51690 9376
rect 52270 9364 52276 9376
rect 52231 9336 52276 9364
rect 52270 9324 52276 9336
rect 52328 9324 52334 9376
rect 52454 9324 52460 9376
rect 52512 9364 52518 9376
rect 53098 9364 53104 9376
rect 52512 9336 53104 9364
rect 52512 9324 52518 9336
rect 53098 9324 53104 9336
rect 53156 9324 53162 9376
rect 1104 9274 54832 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 54832 9274
rect 1104 9200 54832 9222
rect 13725 9163 13783 9169
rect 13725 9129 13737 9163
rect 13771 9160 13783 9163
rect 14550 9160 14556 9172
rect 13771 9132 14556 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 15473 9163 15531 9169
rect 15473 9129 15485 9163
rect 15519 9160 15531 9163
rect 16393 9163 16451 9169
rect 15519 9132 16344 9160
rect 15519 9129 15531 9132
rect 15473 9123 15531 9129
rect 13262 9052 13268 9104
rect 13320 9092 13326 9104
rect 13541 9095 13599 9101
rect 13541 9092 13553 9095
rect 13320 9064 13553 9092
rect 13320 9052 13326 9064
rect 13541 9061 13553 9064
rect 13587 9061 13599 9095
rect 16206 9092 16212 9104
rect 16167 9064 16212 9092
rect 13541 9055 13599 9061
rect 16206 9052 16212 9064
rect 16264 9052 16270 9104
rect 16316 9092 16344 9132
rect 16393 9129 16405 9163
rect 16439 9160 16451 9163
rect 16482 9160 16488 9172
rect 16439 9132 16488 9160
rect 16439 9129 16451 9132
rect 16393 9123 16451 9129
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 16942 9160 16948 9172
rect 16855 9132 16948 9160
rect 16942 9120 16948 9132
rect 17000 9160 17006 9172
rect 17310 9160 17316 9172
rect 17000 9132 17316 9160
rect 17000 9120 17006 9132
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 18230 9160 18236 9172
rect 18191 9132 18236 9160
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 21358 9120 21364 9172
rect 21416 9160 21422 9172
rect 23017 9163 23075 9169
rect 23017 9160 23029 9163
rect 21416 9132 23029 9160
rect 21416 9120 21422 9132
rect 23017 9129 23029 9132
rect 23063 9129 23075 9163
rect 24026 9160 24032 9172
rect 23987 9132 24032 9160
rect 23017 9123 23075 9129
rect 24026 9120 24032 9132
rect 24084 9120 24090 9172
rect 24762 9120 24768 9172
rect 24820 9160 24826 9172
rect 27985 9163 28043 9169
rect 24820 9132 27752 9160
rect 24820 9120 24826 9132
rect 18322 9092 18328 9104
rect 16316 9064 18328 9092
rect 18322 9052 18328 9064
rect 18380 9052 18386 9104
rect 18414 9052 18420 9104
rect 18472 9092 18478 9104
rect 25774 9092 25780 9104
rect 18472 9064 25780 9092
rect 18472 9052 18478 9064
rect 25774 9052 25780 9064
rect 25832 9052 25838 9104
rect 14277 9027 14335 9033
rect 14277 9024 14289 9027
rect 2746 8996 14289 9024
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8956 1915 8959
rect 2746 8956 2774 8996
rect 14277 8993 14289 8996
rect 14323 8993 14335 9027
rect 14277 8987 14335 8993
rect 14553 9027 14611 9033
rect 14553 8993 14565 9027
rect 14599 9024 14611 9027
rect 17954 9024 17960 9036
rect 14599 8996 17960 9024
rect 14599 8993 14611 8996
rect 14553 8987 14611 8993
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 19426 9024 19432 9036
rect 18064 8996 19432 9024
rect 1903 8928 2774 8956
rect 1903 8925 1915 8928
rect 1857 8919 1915 8925
rect 14090 8916 14096 8968
rect 14148 8956 14154 8968
rect 14461 8959 14519 8965
rect 14461 8956 14473 8959
rect 14148 8928 14473 8956
rect 14148 8916 14154 8928
rect 14461 8925 14473 8928
rect 14507 8925 14519 8959
rect 14642 8956 14648 8968
rect 14603 8928 14648 8956
rect 14461 8919 14519 8925
rect 13265 8891 13323 8897
rect 13265 8857 13277 8891
rect 13311 8857 13323 8891
rect 14476 8888 14504 8919
rect 14642 8916 14648 8928
rect 14700 8916 14706 8968
rect 14734 8916 14740 8968
rect 14792 8956 14798 8968
rect 18064 8965 18092 8996
rect 19426 8984 19432 8996
rect 19484 8984 19490 9036
rect 19518 8984 19524 9036
rect 19576 9024 19582 9036
rect 19981 9027 20039 9033
rect 19981 9024 19993 9027
rect 19576 8996 19993 9024
rect 19576 8984 19582 8996
rect 19981 8993 19993 8996
rect 20027 9024 20039 9027
rect 21542 9024 21548 9036
rect 20027 8996 21548 9024
rect 20027 8993 20039 8996
rect 19981 8987 20039 8993
rect 21542 8984 21548 8996
rect 21600 8984 21606 9036
rect 22830 8984 22836 9036
rect 22888 9024 22894 9036
rect 25041 9027 25099 9033
rect 25041 9024 25053 9027
rect 22888 8996 25053 9024
rect 22888 8984 22894 8996
rect 25041 8993 25053 8996
rect 25087 8993 25099 9027
rect 25041 8987 25099 8993
rect 25130 8984 25136 9036
rect 25188 9024 25194 9036
rect 26418 9024 26424 9036
rect 25188 8996 25233 9024
rect 25332 8996 26424 9024
rect 25188 8984 25194 8996
rect 15289 8959 15347 8965
rect 14792 8928 14837 8956
rect 14792 8916 14798 8928
rect 15289 8925 15301 8959
rect 15335 8956 15347 8959
rect 18049 8959 18107 8965
rect 15335 8928 17540 8956
rect 15335 8925 15347 8928
rect 15289 8919 15347 8925
rect 14550 8888 14556 8900
rect 14476 8860 14556 8888
rect 13265 8851 13323 8857
rect 1670 8820 1676 8832
rect 1631 8792 1676 8820
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 13280 8820 13308 8851
rect 14550 8848 14556 8860
rect 14608 8848 14614 8900
rect 15933 8891 15991 8897
rect 15933 8857 15945 8891
rect 15979 8888 15991 8891
rect 16942 8888 16948 8900
rect 15979 8860 16948 8888
rect 15979 8857 15991 8860
rect 15933 8851 15991 8857
rect 14458 8820 14464 8832
rect 13280 8792 14464 8820
rect 14458 8780 14464 8792
rect 14516 8820 14522 8832
rect 15948 8820 15976 8851
rect 16942 8848 16948 8860
rect 17000 8848 17006 8900
rect 17037 8891 17095 8897
rect 17037 8857 17049 8891
rect 17083 8888 17095 8891
rect 17310 8888 17316 8900
rect 17083 8860 17316 8888
rect 17083 8857 17095 8860
rect 17037 8851 17095 8857
rect 17310 8848 17316 8860
rect 17368 8848 17374 8900
rect 17512 8888 17540 8928
rect 18049 8925 18061 8959
rect 18095 8925 18107 8959
rect 18049 8919 18107 8925
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8956 18751 8959
rect 21361 8959 21419 8965
rect 18739 8928 20208 8956
rect 18739 8925 18751 8928
rect 18693 8919 18751 8925
rect 19794 8888 19800 8900
rect 17512 8860 19472 8888
rect 19755 8860 19800 8888
rect 18874 8820 18880 8832
rect 14516 8792 15976 8820
rect 18835 8792 18880 8820
rect 14516 8780 14522 8792
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 19444 8829 19472 8860
rect 19794 8848 19800 8860
rect 19852 8848 19858 8900
rect 19429 8823 19487 8829
rect 19429 8789 19441 8823
rect 19475 8789 19487 8823
rect 19429 8783 19487 8789
rect 19889 8823 19947 8829
rect 19889 8789 19901 8823
rect 19935 8820 19947 8823
rect 20070 8820 20076 8832
rect 19935 8792 20076 8820
rect 19935 8789 19947 8792
rect 19889 8783 19947 8789
rect 20070 8780 20076 8792
rect 20128 8780 20134 8832
rect 20180 8820 20208 8928
rect 21361 8925 21373 8959
rect 21407 8956 21419 8959
rect 21450 8956 21456 8968
rect 21407 8928 21456 8956
rect 21407 8925 21419 8928
rect 21361 8919 21419 8925
rect 21450 8916 21456 8928
rect 21508 8956 21514 8968
rect 21634 8956 21640 8968
rect 21508 8928 21640 8956
rect 21508 8916 21514 8928
rect 21634 8916 21640 8928
rect 21692 8916 21698 8968
rect 22373 8959 22431 8965
rect 22373 8925 22385 8959
rect 22419 8925 22431 8959
rect 23198 8956 23204 8968
rect 23159 8928 23204 8956
rect 22373 8919 22431 8925
rect 22388 8888 22416 8919
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 23842 8956 23848 8968
rect 23803 8928 23848 8956
rect 23842 8916 23848 8928
rect 23900 8916 23906 8968
rect 25332 8956 25360 8996
rect 26418 8984 26424 8996
rect 26476 8984 26482 9036
rect 27724 9024 27752 9132
rect 27985 9129 27997 9163
rect 28031 9160 28043 9163
rect 28166 9160 28172 9172
rect 28031 9132 28172 9160
rect 28031 9129 28043 9132
rect 27985 9123 28043 9129
rect 28166 9120 28172 9132
rect 28224 9120 28230 9172
rect 28350 9120 28356 9172
rect 28408 9160 28414 9172
rect 28534 9160 28540 9172
rect 28408 9132 28540 9160
rect 28408 9120 28414 9132
rect 28534 9120 28540 9132
rect 28592 9160 28598 9172
rect 31113 9163 31171 9169
rect 31113 9160 31125 9163
rect 28592 9132 31125 9160
rect 28592 9120 28598 9132
rect 31113 9129 31125 9132
rect 31159 9160 31171 9163
rect 31202 9160 31208 9172
rect 31159 9132 31208 9160
rect 31159 9129 31171 9132
rect 31113 9123 31171 9129
rect 31202 9120 31208 9132
rect 31260 9120 31266 9172
rect 31662 9160 31668 9172
rect 31623 9132 31668 9160
rect 31662 9120 31668 9132
rect 31720 9120 31726 9172
rect 34333 9163 34391 9169
rect 34333 9129 34345 9163
rect 34379 9160 34391 9163
rect 34514 9160 34520 9172
rect 34379 9132 34520 9160
rect 34379 9129 34391 9132
rect 34333 9123 34391 9129
rect 34514 9120 34520 9132
rect 34572 9120 34578 9172
rect 35802 9120 35808 9172
rect 35860 9160 35866 9172
rect 36081 9163 36139 9169
rect 36081 9160 36093 9163
rect 35860 9132 36093 9160
rect 35860 9120 35866 9132
rect 36081 9129 36093 9132
rect 36127 9129 36139 9163
rect 36081 9123 36139 9129
rect 38654 9120 38660 9172
rect 38712 9160 38718 9172
rect 38749 9163 38807 9169
rect 38749 9160 38761 9163
rect 38712 9132 38761 9160
rect 38712 9120 38718 9132
rect 38749 9129 38761 9132
rect 38795 9129 38807 9163
rect 38749 9123 38807 9129
rect 48961 9163 49019 9169
rect 48961 9129 48973 9163
rect 49007 9160 49019 9163
rect 49050 9160 49056 9172
rect 49007 9132 49056 9160
rect 49007 9129 49019 9132
rect 48961 9123 49019 9129
rect 49050 9120 49056 9132
rect 49108 9120 49114 9172
rect 49142 9120 49148 9172
rect 49200 9160 49206 9172
rect 49200 9132 52592 9160
rect 49200 9120 49206 9132
rect 35618 9092 35624 9104
rect 35452 9064 35624 9092
rect 28442 9024 28448 9036
rect 27724 8996 28448 9024
rect 28442 8984 28448 8996
rect 28500 8984 28506 9036
rect 28629 9027 28687 9033
rect 28629 8993 28641 9027
rect 28675 9024 28687 9027
rect 29086 9024 29092 9036
rect 28675 8996 29092 9024
rect 28675 8993 28687 8996
rect 28629 8987 28687 8993
rect 29086 8984 29092 8996
rect 29144 9024 29150 9036
rect 29454 9024 29460 9036
rect 29144 8996 29460 9024
rect 29144 8984 29150 8996
rect 29454 8984 29460 8996
rect 29512 8984 29518 9036
rect 31846 8984 31852 9036
rect 31904 9024 31910 9036
rect 32125 9027 32183 9033
rect 32125 9024 32137 9027
rect 31904 8996 32137 9024
rect 31904 8984 31910 8996
rect 32125 8993 32137 8996
rect 32171 8993 32183 9027
rect 32306 9024 32312 9036
rect 32267 8996 32312 9024
rect 32125 8987 32183 8993
rect 32306 8984 32312 8996
rect 32364 8984 32370 9036
rect 32950 8984 32956 9036
rect 33008 9024 33014 9036
rect 33008 8996 33548 9024
rect 33008 8984 33014 8996
rect 27430 8956 27436 8968
rect 23952 8928 25360 8956
rect 25976 8928 27436 8956
rect 23750 8888 23756 8900
rect 22388 8860 23756 8888
rect 23750 8848 23756 8860
rect 23808 8848 23814 8900
rect 20993 8823 21051 8829
rect 20993 8820 21005 8823
rect 20180 8792 21005 8820
rect 20993 8789 21005 8792
rect 21039 8789 21051 8823
rect 20993 8783 21051 8789
rect 21358 8780 21364 8832
rect 21416 8820 21422 8832
rect 21453 8823 21511 8829
rect 21453 8820 21465 8823
rect 21416 8792 21465 8820
rect 21416 8780 21422 8792
rect 21453 8789 21465 8792
rect 21499 8789 21511 8823
rect 22554 8820 22560 8832
rect 22515 8792 22560 8820
rect 21453 8783 21511 8789
rect 22554 8780 22560 8792
rect 22612 8780 22618 8832
rect 23106 8780 23112 8832
rect 23164 8820 23170 8832
rect 23952 8820 23980 8928
rect 25976 8832 26004 8928
rect 27430 8916 27436 8928
rect 27488 8916 27494 8968
rect 27525 8959 27583 8965
rect 27525 8925 27537 8959
rect 27571 8956 27583 8959
rect 27614 8956 27620 8968
rect 27571 8928 27620 8956
rect 27571 8925 27583 8928
rect 27525 8919 27583 8925
rect 27614 8916 27620 8928
rect 27672 8956 27678 8968
rect 29730 8956 29736 8968
rect 27672 8928 29736 8956
rect 27672 8916 27678 8928
rect 29730 8916 29736 8928
rect 29788 8916 29794 8968
rect 29822 8916 29828 8968
rect 29880 8956 29886 8968
rect 29989 8959 30047 8965
rect 29880 8952 29960 8956
rect 29989 8952 30001 8959
rect 29880 8928 30001 8952
rect 29880 8916 29886 8928
rect 29932 8925 30001 8928
rect 30035 8956 30047 8959
rect 32861 8959 32919 8965
rect 30035 8925 30052 8956
rect 29932 8924 30052 8925
rect 32861 8925 32873 8959
rect 32907 8956 32919 8959
rect 33318 8956 33324 8968
rect 32907 8928 33324 8956
rect 32907 8925 32919 8928
rect 29989 8919 30047 8924
rect 32861 8919 32919 8925
rect 33318 8916 33324 8928
rect 33376 8916 33382 8968
rect 33520 8952 33548 8996
rect 33594 8984 33600 9036
rect 33652 9024 33658 9036
rect 33689 9027 33747 9033
rect 33689 9024 33701 9027
rect 33652 8996 33701 9024
rect 33652 8984 33658 8996
rect 33689 8993 33701 8996
rect 33735 9024 33747 9027
rect 33778 9024 33784 9036
rect 33735 8996 33784 9024
rect 33735 8993 33747 8996
rect 33689 8987 33747 8993
rect 33778 8984 33784 8996
rect 33836 8984 33842 9036
rect 35452 9033 35480 9064
rect 35618 9052 35624 9064
rect 35676 9052 35682 9104
rect 35894 9052 35900 9104
rect 35952 9092 35958 9104
rect 42978 9092 42984 9104
rect 35952 9064 42984 9092
rect 35952 9052 35958 9064
rect 42978 9052 42984 9064
rect 43036 9052 43042 9104
rect 46198 9052 46204 9104
rect 46256 9092 46262 9104
rect 52454 9092 52460 9104
rect 46256 9064 52460 9092
rect 46256 9052 46262 9064
rect 52454 9052 52460 9064
rect 52512 9052 52518 9104
rect 52564 9092 52592 9132
rect 52730 9120 52736 9172
rect 52788 9160 52794 9172
rect 53561 9163 53619 9169
rect 53561 9160 53573 9163
rect 52788 9132 53573 9160
rect 52788 9120 52794 9132
rect 53561 9129 53573 9132
rect 53607 9129 53619 9163
rect 53561 9123 53619 9129
rect 53745 9095 53803 9101
rect 53745 9092 53757 9095
rect 52564 9064 53757 9092
rect 53745 9061 53757 9064
rect 53791 9061 53803 9095
rect 53745 9055 53803 9061
rect 35437 9027 35495 9033
rect 35437 8993 35449 9027
rect 35483 8993 35495 9027
rect 37918 9024 37924 9036
rect 37831 8996 37924 9024
rect 35437 8987 35495 8993
rect 37918 8984 37924 8996
rect 37976 9024 37982 9036
rect 52270 9024 52276 9036
rect 37976 8996 52276 9024
rect 37976 8984 37982 8996
rect 52270 8984 52276 8996
rect 52328 8984 52334 9036
rect 36265 8959 36323 8965
rect 36265 8956 36277 8959
rect 33704 8952 36277 8956
rect 33520 8928 36277 8952
rect 33520 8924 33732 8928
rect 36265 8925 36277 8928
rect 36311 8925 36323 8959
rect 36265 8919 36323 8925
rect 36722 8916 36728 8968
rect 36780 8956 36786 8968
rect 38933 8959 38991 8965
rect 36780 8928 36825 8956
rect 36780 8916 36786 8928
rect 38933 8925 38945 8959
rect 38979 8925 38991 8959
rect 39114 8956 39120 8968
rect 39075 8928 39120 8956
rect 38933 8919 38991 8925
rect 27246 8888 27252 8900
rect 27304 8897 27310 8900
rect 27216 8860 27252 8888
rect 27246 8848 27252 8860
rect 27304 8851 27316 8897
rect 31018 8888 31024 8900
rect 27356 8860 31024 8888
rect 27304 8848 27310 8851
rect 24578 8820 24584 8832
rect 23164 8792 23980 8820
rect 24539 8792 24584 8820
rect 23164 8780 23170 8792
rect 24578 8780 24584 8792
rect 24636 8780 24642 8832
rect 24949 8823 25007 8829
rect 24949 8789 24961 8823
rect 24995 8820 25007 8823
rect 25958 8820 25964 8832
rect 24995 8792 25964 8820
rect 24995 8789 25007 8792
rect 24949 8783 25007 8789
rect 25958 8780 25964 8792
rect 26016 8780 26022 8832
rect 26145 8823 26203 8829
rect 26145 8789 26157 8823
rect 26191 8820 26203 8823
rect 26326 8820 26332 8832
rect 26191 8792 26332 8820
rect 26191 8789 26203 8792
rect 26145 8783 26203 8789
rect 26326 8780 26332 8792
rect 26384 8780 26390 8832
rect 26418 8780 26424 8832
rect 26476 8820 26482 8832
rect 27356 8820 27384 8860
rect 31018 8848 31024 8860
rect 31076 8848 31082 8900
rect 37277 8891 37335 8897
rect 37277 8888 37289 8891
rect 33888 8860 37289 8888
rect 33888 8832 33916 8860
rect 37277 8857 37289 8860
rect 37323 8888 37335 8891
rect 38654 8888 38660 8900
rect 37323 8860 38660 8888
rect 37323 8857 37335 8860
rect 37277 8851 37335 8857
rect 38654 8848 38660 8860
rect 38712 8848 38718 8900
rect 38948 8888 38976 8919
rect 39114 8916 39120 8928
rect 39172 8916 39178 8968
rect 42518 8916 42524 8968
rect 42576 8956 42582 8968
rect 48777 8959 48835 8965
rect 48777 8956 48789 8959
rect 42576 8928 48789 8956
rect 42576 8916 42582 8928
rect 48777 8925 48789 8928
rect 48823 8925 48835 8959
rect 48958 8956 48964 8968
rect 48919 8928 48964 8956
rect 48777 8919 48835 8925
rect 40218 8888 40224 8900
rect 38948 8860 40224 8888
rect 40218 8848 40224 8860
rect 40276 8848 40282 8900
rect 48792 8888 48820 8919
rect 48958 8916 48964 8928
rect 49016 8956 49022 8968
rect 51626 8956 51632 8968
rect 49016 8928 51074 8956
rect 51587 8928 51632 8956
rect 49016 8916 49022 8928
rect 50430 8888 50436 8900
rect 48792 8860 49556 8888
rect 50391 8860 50436 8888
rect 26476 8792 27384 8820
rect 28353 8823 28411 8829
rect 26476 8780 26482 8792
rect 28353 8789 28365 8823
rect 28399 8820 28411 8823
rect 28626 8820 28632 8832
rect 28399 8792 28632 8820
rect 28399 8789 28411 8792
rect 28353 8783 28411 8789
rect 28626 8780 28632 8792
rect 28684 8780 28690 8832
rect 28718 8780 28724 8832
rect 28776 8820 28782 8832
rect 31846 8820 31852 8832
rect 28776 8792 31852 8820
rect 28776 8780 28782 8792
rect 31846 8780 31852 8792
rect 31904 8780 31910 8832
rect 32033 8823 32091 8829
rect 32033 8789 32045 8823
rect 32079 8820 32091 8823
rect 32122 8820 32128 8832
rect 32079 8792 32128 8820
rect 32079 8789 32091 8792
rect 32033 8783 32091 8789
rect 32122 8780 32128 8792
rect 32180 8780 32186 8832
rect 33045 8823 33103 8829
rect 33045 8789 33057 8823
rect 33091 8820 33103 8823
rect 33502 8820 33508 8832
rect 33091 8792 33508 8820
rect 33091 8789 33103 8792
rect 33045 8783 33103 8789
rect 33502 8780 33508 8792
rect 33560 8780 33566 8832
rect 33870 8820 33876 8832
rect 33831 8792 33876 8820
rect 33870 8780 33876 8792
rect 33928 8780 33934 8832
rect 33965 8823 34023 8829
rect 33965 8789 33977 8823
rect 34011 8820 34023 8823
rect 34422 8820 34428 8832
rect 34011 8792 34428 8820
rect 34011 8789 34023 8792
rect 33965 8783 34023 8789
rect 34422 8780 34428 8792
rect 34480 8780 34486 8832
rect 34514 8780 34520 8832
rect 34572 8820 34578 8832
rect 34885 8823 34943 8829
rect 34885 8820 34897 8823
rect 34572 8792 34897 8820
rect 34572 8780 34578 8792
rect 34885 8789 34897 8792
rect 34931 8789 34943 8823
rect 34885 8783 34943 8789
rect 34974 8780 34980 8832
rect 35032 8820 35038 8832
rect 35253 8823 35311 8829
rect 35253 8820 35265 8823
rect 35032 8792 35265 8820
rect 35032 8780 35038 8792
rect 35253 8789 35265 8792
rect 35299 8789 35311 8823
rect 35253 8783 35311 8789
rect 35345 8823 35403 8829
rect 35345 8789 35357 8823
rect 35391 8820 35403 8823
rect 36630 8820 36636 8832
rect 35391 8792 36636 8820
rect 35391 8789 35403 8792
rect 35345 8783 35403 8789
rect 36630 8780 36636 8792
rect 36688 8780 36694 8832
rect 36722 8780 36728 8832
rect 36780 8820 36786 8832
rect 48406 8820 48412 8832
rect 36780 8792 48412 8820
rect 36780 8780 36786 8792
rect 48406 8780 48412 8792
rect 48464 8780 48470 8832
rect 49528 8829 49556 8860
rect 50430 8848 50436 8860
rect 50488 8848 50494 8900
rect 51046 8888 51074 8928
rect 51626 8916 51632 8928
rect 51684 8916 51690 8968
rect 52454 8916 52460 8968
rect 52512 8956 52518 8968
rect 52730 8956 52736 8968
rect 52512 8928 52736 8956
rect 52512 8916 52518 8928
rect 52730 8916 52736 8928
rect 52788 8916 52794 8968
rect 52917 8959 52975 8965
rect 52917 8925 52929 8959
rect 52963 8956 52975 8959
rect 52963 8928 53236 8956
rect 52963 8925 52975 8928
rect 52917 8919 52975 8925
rect 53208 8900 53236 8928
rect 52825 8891 52883 8897
rect 52825 8888 52837 8891
rect 51046 8860 52837 8888
rect 52825 8857 52837 8860
rect 52871 8857 52883 8891
rect 52825 8851 52883 8857
rect 53190 8848 53196 8900
rect 53248 8888 53254 8900
rect 53377 8891 53435 8897
rect 53377 8888 53389 8891
rect 53248 8860 53389 8888
rect 53248 8848 53254 8860
rect 53377 8857 53389 8860
rect 53423 8857 53435 8891
rect 53377 8851 53435 8857
rect 49513 8823 49571 8829
rect 49513 8789 49525 8823
rect 49559 8820 49571 8823
rect 49694 8820 49700 8832
rect 49559 8792 49700 8820
rect 49559 8789 49571 8792
rect 49513 8783 49571 8789
rect 49694 8780 49700 8792
rect 49752 8780 49758 8832
rect 51813 8823 51871 8829
rect 51813 8789 51825 8823
rect 51859 8820 51871 8823
rect 52730 8820 52736 8832
rect 51859 8792 52736 8820
rect 51859 8789 51871 8792
rect 51813 8783 51871 8789
rect 52730 8780 52736 8792
rect 52788 8780 52794 8832
rect 53558 8820 53564 8832
rect 53519 8792 53564 8820
rect 53558 8780 53564 8792
rect 53616 8780 53622 8832
rect 1104 8730 54832 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 54832 8730
rect 1104 8656 54832 8678
rect 14829 8619 14887 8625
rect 14829 8585 14841 8619
rect 14875 8616 14887 8619
rect 15470 8616 15476 8628
rect 14875 8588 15476 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 17313 8619 17371 8625
rect 17313 8585 17325 8619
rect 17359 8616 17371 8619
rect 17402 8616 17408 8628
rect 17359 8588 17408 8616
rect 17359 8585 17371 8588
rect 17313 8579 17371 8585
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 22005 8619 22063 8625
rect 18932 8588 20116 8616
rect 18932 8576 18938 8588
rect 14369 8551 14427 8557
rect 14369 8517 14381 8551
rect 14415 8548 14427 8551
rect 14458 8548 14464 8560
rect 14415 8520 14464 8548
rect 14415 8517 14427 8520
rect 14369 8511 14427 8517
rect 14458 8508 14464 8520
rect 14516 8508 14522 8560
rect 16301 8551 16359 8557
rect 16301 8548 16313 8551
rect 15488 8520 16313 8548
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 11054 8480 11060 8492
rect 1903 8452 11060 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 11054 8440 11060 8452
rect 11112 8440 11118 8492
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8480 13967 8483
rect 14642 8480 14648 8492
rect 13955 8452 14648 8480
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 15488 8489 15516 8520
rect 16301 8517 16313 8520
rect 16347 8548 16359 8551
rect 16853 8551 16911 8557
rect 16853 8548 16865 8551
rect 16347 8520 16865 8548
rect 16347 8517 16359 8520
rect 16301 8511 16359 8517
rect 16853 8517 16865 8520
rect 16899 8548 16911 8551
rect 17126 8548 17132 8560
rect 16899 8520 17132 8548
rect 16899 8517 16911 8520
rect 16853 8511 16911 8517
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 19334 8548 19340 8560
rect 18248 8520 19340 8548
rect 18248 8489 18276 8520
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 20088 8548 20116 8588
rect 22005 8585 22017 8619
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 22373 8619 22431 8625
rect 22373 8585 22385 8619
rect 22419 8616 22431 8619
rect 23106 8616 23112 8628
rect 22419 8588 23112 8616
rect 22419 8585 22431 8588
rect 22373 8579 22431 8585
rect 20318 8551 20376 8557
rect 20318 8548 20330 8551
rect 20088 8520 20330 8548
rect 20318 8517 20330 8520
rect 20364 8517 20376 8551
rect 20318 8511 20376 8517
rect 18506 8489 18512 8492
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8449 15531 8483
rect 18233 8483 18291 8489
rect 15473 8443 15531 8449
rect 16776 8452 18184 8480
rect 15102 8372 15108 8424
rect 15160 8412 15166 8424
rect 16776 8412 16804 8452
rect 15160 8384 16804 8412
rect 15160 8372 15166 8384
rect 1670 8344 1676 8356
rect 1631 8316 1676 8344
rect 1670 8304 1676 8316
rect 1728 8304 1734 8356
rect 13630 8304 13636 8356
rect 13688 8344 13694 8356
rect 14645 8347 14703 8353
rect 14645 8344 14657 8347
rect 13688 8316 14657 8344
rect 13688 8304 13694 8316
rect 14645 8313 14657 8316
rect 14691 8313 14703 8347
rect 14645 8307 14703 8313
rect 15286 8304 15292 8356
rect 15344 8344 15350 8356
rect 15657 8347 15715 8353
rect 15657 8344 15669 8347
rect 15344 8316 15669 8344
rect 15344 8304 15350 8316
rect 15657 8313 15669 8316
rect 15703 8344 15715 8347
rect 16666 8344 16672 8356
rect 15703 8316 16672 8344
rect 15703 8313 15715 8316
rect 15657 8307 15715 8313
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 17221 8347 17279 8353
rect 17221 8313 17233 8347
rect 17267 8344 17279 8347
rect 17586 8344 17592 8356
rect 17267 8316 17592 8344
rect 17267 8313 17279 8316
rect 17221 8307 17279 8313
rect 17586 8304 17592 8316
rect 17644 8304 17650 8356
rect 18156 8344 18184 8452
rect 18233 8449 18245 8483
rect 18279 8449 18291 8483
rect 18233 8443 18291 8449
rect 18500 8443 18512 8489
rect 18564 8480 18570 8492
rect 18564 8452 18600 8480
rect 18506 8440 18512 8443
rect 18564 8440 18570 8452
rect 18782 8440 18788 8492
rect 18840 8480 18846 8492
rect 22020 8480 22048 8579
rect 23106 8576 23112 8588
rect 23164 8576 23170 8628
rect 25130 8616 25136 8628
rect 23400 8588 25136 8616
rect 18840 8452 22048 8480
rect 18840 8440 18846 8452
rect 22278 8440 22284 8492
rect 22336 8480 22342 8492
rect 22646 8480 22652 8492
rect 22336 8452 22652 8480
rect 22336 8440 22342 8452
rect 22646 8440 22652 8452
rect 22704 8480 22710 8492
rect 23293 8483 23351 8489
rect 23293 8480 23305 8483
rect 22704 8452 23305 8480
rect 22704 8440 22710 8452
rect 23293 8449 23305 8452
rect 23339 8449 23351 8483
rect 23293 8443 23351 8449
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 19978 8412 19984 8424
rect 19392 8384 19984 8412
rect 19392 8372 19398 8384
rect 19978 8372 19984 8384
rect 20036 8412 20042 8424
rect 20073 8415 20131 8421
rect 20073 8412 20085 8415
rect 20036 8384 20085 8412
rect 20036 8372 20042 8384
rect 20073 8381 20085 8384
rect 20119 8381 20131 8415
rect 20073 8375 20131 8381
rect 21266 8372 21272 8424
rect 21324 8412 21330 8424
rect 22465 8415 22523 8421
rect 22465 8412 22477 8415
rect 21324 8384 22477 8412
rect 21324 8372 21330 8384
rect 22465 8381 22477 8384
rect 22511 8381 22523 8415
rect 22465 8375 22523 8381
rect 22557 8415 22615 8421
rect 22557 8381 22569 8415
rect 22603 8412 22615 8415
rect 23400 8412 23428 8588
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 25682 8576 25688 8628
rect 25740 8616 25746 8628
rect 25777 8619 25835 8625
rect 25777 8616 25789 8619
rect 25740 8588 25789 8616
rect 25740 8576 25746 8588
rect 25777 8585 25789 8588
rect 25823 8585 25835 8619
rect 27982 8616 27988 8628
rect 25777 8579 25835 8585
rect 25976 8588 27988 8616
rect 23566 8489 23572 8492
rect 23560 8443 23572 8489
rect 23624 8480 23630 8492
rect 25133 8483 25191 8489
rect 23624 8452 23660 8480
rect 23566 8440 23572 8443
rect 23624 8440 23630 8452
rect 25133 8449 25145 8483
rect 25179 8480 25191 8483
rect 25976 8480 26004 8588
rect 27982 8576 27988 8588
rect 28040 8576 28046 8628
rect 28442 8576 28448 8628
rect 28500 8616 28506 8628
rect 28537 8619 28595 8625
rect 28537 8616 28549 8619
rect 28500 8588 28549 8616
rect 28500 8576 28506 8588
rect 28537 8585 28549 8588
rect 28583 8616 28595 8619
rect 32030 8616 32036 8628
rect 28583 8588 32036 8616
rect 28583 8585 28595 8588
rect 28537 8579 28595 8585
rect 32030 8576 32036 8588
rect 32088 8576 32094 8628
rect 32490 8616 32496 8628
rect 32451 8588 32496 8616
rect 32490 8576 32496 8588
rect 32548 8576 32554 8628
rect 33686 8616 33692 8628
rect 33428 8588 33692 8616
rect 26237 8551 26295 8557
rect 26237 8517 26249 8551
rect 26283 8548 26295 8551
rect 26418 8548 26424 8560
rect 26283 8520 26424 8548
rect 26283 8517 26295 8520
rect 26237 8511 26295 8517
rect 26418 8508 26424 8520
rect 26476 8508 26482 8560
rect 27614 8548 27620 8560
rect 27172 8520 27620 8548
rect 27172 8489 27200 8520
rect 27614 8508 27620 8520
rect 27672 8508 27678 8560
rect 29730 8548 29736 8560
rect 29380 8520 29736 8548
rect 29380 8489 29408 8520
rect 29730 8508 29736 8520
rect 29788 8548 29794 8560
rect 33428 8548 33456 8588
rect 33686 8576 33692 8588
rect 33744 8576 33750 8628
rect 34698 8576 34704 8628
rect 34756 8616 34762 8628
rect 35253 8619 35311 8625
rect 35253 8616 35265 8619
rect 34756 8588 35265 8616
rect 34756 8576 34762 8588
rect 35253 8585 35265 8588
rect 35299 8585 35311 8619
rect 35253 8579 35311 8585
rect 36541 8619 36599 8625
rect 36541 8585 36553 8619
rect 36587 8616 36599 8619
rect 36814 8616 36820 8628
rect 36587 8588 36820 8616
rect 36587 8585 36599 8588
rect 36541 8579 36599 8585
rect 36814 8576 36820 8588
rect 36872 8576 36878 8628
rect 38105 8619 38163 8625
rect 38105 8585 38117 8619
rect 38151 8616 38163 8619
rect 38286 8616 38292 8628
rect 38151 8588 38292 8616
rect 38151 8585 38163 8588
rect 38105 8579 38163 8585
rect 38286 8576 38292 8588
rect 38344 8616 38350 8628
rect 38565 8619 38623 8625
rect 38565 8616 38577 8619
rect 38344 8588 38577 8616
rect 38344 8576 38350 8588
rect 38565 8585 38577 8588
rect 38611 8585 38623 8619
rect 38565 8579 38623 8585
rect 38654 8576 38660 8628
rect 38712 8616 38718 8628
rect 50890 8616 50896 8628
rect 38712 8588 50896 8616
rect 38712 8576 38718 8588
rect 50890 8576 50896 8588
rect 50948 8576 50954 8628
rect 53377 8619 53435 8625
rect 53377 8616 53389 8619
rect 51046 8588 53389 8616
rect 29788 8520 33456 8548
rect 29788 8508 29794 8520
rect 25179 8452 26004 8480
rect 26145 8483 26203 8489
rect 25179 8449 25191 8452
rect 25133 8443 25191 8449
rect 26145 8449 26157 8483
rect 26191 8449 26203 8483
rect 26145 8443 26203 8449
rect 27157 8483 27215 8489
rect 27157 8449 27169 8483
rect 27203 8449 27215 8483
rect 27413 8483 27471 8489
rect 27413 8480 27425 8483
rect 27157 8443 27215 8449
rect 27264 8452 27425 8480
rect 22603 8384 23428 8412
rect 22603 8381 22615 8384
rect 22557 8375 22615 8381
rect 19610 8344 19616 8356
rect 18156 8316 18276 8344
rect 19571 8316 19616 8344
rect 18248 8276 18276 8316
rect 19610 8304 19616 8316
rect 19668 8344 19674 8356
rect 19886 8344 19892 8356
rect 19668 8316 19892 8344
rect 19668 8304 19674 8316
rect 19886 8304 19892 8316
rect 19944 8304 19950 8356
rect 21358 8344 21364 8356
rect 21008 8316 21364 8344
rect 21008 8276 21036 8316
rect 21358 8304 21364 8316
rect 21416 8344 21422 8356
rect 21453 8347 21511 8353
rect 21453 8344 21465 8347
rect 21416 8316 21465 8344
rect 21416 8304 21422 8316
rect 21453 8313 21465 8316
rect 21499 8313 21511 8347
rect 21453 8307 21511 8313
rect 21542 8304 21548 8356
rect 21600 8344 21606 8356
rect 22002 8344 22008 8356
rect 21600 8316 22008 8344
rect 21600 8304 21606 8316
rect 22002 8304 22008 8316
rect 22060 8344 22066 8356
rect 22572 8344 22600 8375
rect 25406 8372 25412 8424
rect 25464 8412 25470 8424
rect 26160 8412 26188 8443
rect 26418 8412 26424 8424
rect 25464 8384 26188 8412
rect 26379 8384 26424 8412
rect 25464 8372 25470 8384
rect 26418 8372 26424 8384
rect 26476 8372 26482 8424
rect 27264 8412 27292 8452
rect 27413 8449 27425 8452
rect 27459 8449 27471 8483
rect 27413 8443 27471 8449
rect 29365 8483 29423 8489
rect 29365 8449 29377 8483
rect 29411 8449 29423 8483
rect 29365 8443 29423 8449
rect 29454 8440 29460 8492
rect 29512 8480 29518 8492
rect 29621 8483 29679 8489
rect 29621 8480 29633 8483
rect 29512 8452 29633 8480
rect 29512 8440 29518 8452
rect 29621 8449 29633 8452
rect 29667 8449 29679 8483
rect 29621 8443 29679 8449
rect 30098 8440 30104 8492
rect 30156 8480 30162 8492
rect 31389 8483 31447 8489
rect 31389 8480 31401 8483
rect 30156 8452 31401 8480
rect 30156 8440 30162 8452
rect 31389 8449 31401 8452
rect 31435 8449 31447 8483
rect 31389 8443 31447 8449
rect 31754 8440 31760 8492
rect 31812 8480 31818 8492
rect 33428 8489 33456 8520
rect 34422 8508 34428 8560
rect 34480 8548 34486 8560
rect 35986 8548 35992 8560
rect 34480 8520 35992 8548
rect 34480 8508 34486 8520
rect 35986 8508 35992 8520
rect 36044 8508 36050 8560
rect 36630 8508 36636 8560
rect 36688 8548 36694 8560
rect 51046 8548 51074 8588
rect 53377 8585 53389 8588
rect 53423 8585 53435 8619
rect 54202 8616 54208 8628
rect 54163 8588 54208 8616
rect 53377 8579 53435 8585
rect 54202 8576 54208 8588
rect 54260 8576 54266 8628
rect 36688 8520 51074 8548
rect 51184 8520 54064 8548
rect 36688 8508 36694 8520
rect 32309 8483 32367 8489
rect 32309 8480 32321 8483
rect 31812 8452 32321 8480
rect 31812 8440 31818 8452
rect 32309 8449 32321 8452
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 33413 8483 33471 8489
rect 33413 8449 33425 8483
rect 33459 8449 33471 8483
rect 33413 8443 33471 8449
rect 33502 8440 33508 8492
rect 33560 8480 33566 8492
rect 33669 8483 33727 8489
rect 33669 8480 33681 8483
rect 33560 8452 33681 8480
rect 33560 8440 33566 8452
rect 33669 8449 33681 8452
rect 33715 8449 33727 8483
rect 35434 8480 35440 8492
rect 35395 8452 35440 8480
rect 33669 8443 33727 8449
rect 35434 8440 35440 8452
rect 35492 8440 35498 8492
rect 39114 8440 39120 8492
rect 39172 8480 39178 8492
rect 51184 8480 51212 8520
rect 39172 8452 51212 8480
rect 51721 8483 51779 8489
rect 39172 8440 39178 8452
rect 51721 8449 51733 8483
rect 51767 8480 51779 8483
rect 52178 8480 52184 8492
rect 51767 8452 52184 8480
rect 51767 8449 51779 8452
rect 51721 8443 51779 8449
rect 52178 8440 52184 8452
rect 52236 8440 52242 8492
rect 53466 8480 53472 8492
rect 53427 8452 53472 8480
rect 53466 8440 53472 8452
rect 53524 8440 53530 8492
rect 54036 8489 54064 8520
rect 54021 8483 54079 8489
rect 54021 8449 54033 8483
rect 54067 8449 54079 8483
rect 54021 8443 54079 8449
rect 27172 8384 27292 8412
rect 22060 8316 22600 8344
rect 22060 8304 22066 8316
rect 24486 8304 24492 8356
rect 24544 8344 24550 8356
rect 24673 8347 24731 8353
rect 24673 8344 24685 8347
rect 24544 8316 24685 8344
rect 24544 8304 24550 8316
rect 24673 8313 24685 8316
rect 24719 8313 24731 8347
rect 24673 8307 24731 8313
rect 25317 8347 25375 8353
rect 25317 8313 25329 8347
rect 25363 8344 25375 8347
rect 27172 8344 27200 8384
rect 30374 8372 30380 8424
rect 30432 8412 30438 8424
rect 31570 8412 31576 8424
rect 30432 8384 31432 8412
rect 31531 8384 31576 8412
rect 30432 8372 30438 8384
rect 25363 8316 27200 8344
rect 30745 8347 30803 8353
rect 25363 8313 25375 8316
rect 25317 8307 25375 8313
rect 30745 8313 30757 8347
rect 30791 8344 30803 8347
rect 31018 8344 31024 8356
rect 30791 8316 31024 8344
rect 30791 8313 30803 8316
rect 30745 8307 30803 8313
rect 31018 8304 31024 8316
rect 31076 8304 31082 8356
rect 31404 8344 31432 8384
rect 31570 8372 31576 8384
rect 31628 8372 31634 8424
rect 37642 8412 37648 8424
rect 34624 8384 37648 8412
rect 31478 8344 31484 8356
rect 31391 8316 31484 8344
rect 31478 8304 31484 8316
rect 31536 8344 31542 8356
rect 33226 8344 33232 8356
rect 31536 8316 33232 8344
rect 31536 8304 31542 8316
rect 33226 8304 33232 8316
rect 33284 8344 33290 8356
rect 34624 8344 34652 8384
rect 37642 8372 37648 8384
rect 37700 8412 37706 8424
rect 46198 8412 46204 8424
rect 37700 8384 46204 8412
rect 37700 8372 37706 8384
rect 46198 8372 46204 8384
rect 46256 8372 46262 8424
rect 51169 8415 51227 8421
rect 51169 8381 51181 8415
rect 51215 8412 51227 8415
rect 53484 8412 53512 8440
rect 51215 8384 53512 8412
rect 51215 8381 51227 8384
rect 51169 8375 51227 8381
rect 34790 8344 34796 8356
rect 33284 8316 33456 8344
rect 33284 8304 33290 8316
rect 18248 8248 21036 8276
rect 28626 8236 28632 8288
rect 28684 8276 28690 8288
rect 30926 8276 30932 8288
rect 28684 8248 30932 8276
rect 28684 8236 28690 8248
rect 30926 8236 30932 8248
rect 30984 8236 30990 8288
rect 31202 8276 31208 8288
rect 31163 8248 31208 8276
rect 31202 8236 31208 8248
rect 31260 8236 31266 8288
rect 33428 8276 33456 8316
rect 34348 8316 34652 8344
rect 34751 8316 34796 8344
rect 34348 8276 34376 8316
rect 34790 8304 34796 8316
rect 34848 8304 34854 8356
rect 37550 8344 37556 8356
rect 37511 8316 37556 8344
rect 37550 8304 37556 8316
rect 37608 8304 37614 8356
rect 48314 8304 48320 8356
rect 48372 8344 48378 8356
rect 52365 8347 52423 8353
rect 52365 8344 52377 8347
rect 48372 8316 52377 8344
rect 48372 8304 48378 8316
rect 52365 8313 52377 8316
rect 52411 8344 52423 8347
rect 53558 8344 53564 8356
rect 52411 8316 53564 8344
rect 52411 8313 52423 8316
rect 52365 8307 52423 8313
rect 53558 8304 53564 8316
rect 53616 8304 53622 8356
rect 33428 8248 34376 8276
rect 35618 8236 35624 8288
rect 35676 8276 35682 8288
rect 35894 8276 35900 8288
rect 35676 8248 35900 8276
rect 35676 8236 35682 8248
rect 35894 8236 35900 8248
rect 35952 8236 35958 8288
rect 1104 8186 54832 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 54832 8186
rect 1104 8112 54832 8134
rect 14642 8072 14648 8084
rect 12636 8044 13584 8072
rect 14603 8044 14648 8072
rect 12636 7945 12664 8044
rect 12437 7939 12495 7945
rect 12437 7936 12449 7939
rect 2746 7908 12449 7936
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7868 1915 7871
rect 2746 7868 2774 7908
rect 12437 7905 12449 7908
rect 12483 7905 12495 7939
rect 12437 7899 12495 7905
rect 12621 7939 12679 7945
rect 12621 7905 12633 7939
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 12805 7939 12863 7945
rect 12805 7905 12817 7939
rect 12851 7936 12863 7939
rect 12986 7936 12992 7948
rect 12851 7908 12992 7936
rect 12851 7905 12863 7908
rect 12805 7899 12863 7905
rect 12986 7896 12992 7908
rect 13044 7896 13050 7948
rect 13556 7945 13584 8044
rect 14642 8032 14648 8044
rect 14700 8032 14706 8084
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 15657 8075 15715 8081
rect 15657 8072 15669 8075
rect 15252 8044 15669 8072
rect 15252 8032 15258 8044
rect 15657 8041 15669 8044
rect 15703 8041 15715 8075
rect 15657 8035 15715 8041
rect 16761 8075 16819 8081
rect 16761 8041 16773 8075
rect 16807 8072 16819 8075
rect 17126 8072 17132 8084
rect 16807 8044 17132 8072
rect 16807 8041 16819 8044
rect 16761 8035 16819 8041
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 17221 8075 17279 8081
rect 17221 8041 17233 8075
rect 17267 8072 17279 8075
rect 17494 8072 17500 8084
rect 17267 8044 17500 8072
rect 17267 8041 17279 8044
rect 17221 8035 17279 8041
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 22189 8075 22247 8081
rect 18156 8044 20944 8072
rect 17405 8007 17463 8013
rect 17405 7973 17417 8007
rect 17451 8004 17463 8007
rect 18046 8004 18052 8016
rect 17451 7976 18052 8004
rect 17451 7973 17463 7976
rect 17405 7967 17463 7973
rect 18046 7964 18052 7976
rect 18104 7964 18110 8016
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 13722 7936 13728 7948
rect 13587 7908 13728 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 13722 7896 13728 7908
rect 13780 7936 13786 7948
rect 18156 7936 18184 8044
rect 13780 7908 18184 7936
rect 18325 7939 18383 7945
rect 13780 7896 13786 7908
rect 18325 7905 18337 7939
rect 18371 7936 18383 7939
rect 19426 7936 19432 7948
rect 18371 7908 19432 7936
rect 18371 7905 18383 7908
rect 18325 7899 18383 7905
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 1903 7840 2774 7868
rect 12713 7871 12771 7877
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12728 7800 12756 7831
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 19610 7868 19616 7880
rect 12952 7840 12997 7868
rect 17604 7840 19616 7868
rect 12952 7828 12958 7840
rect 17604 7800 17632 7840
rect 19610 7828 19616 7840
rect 19668 7828 19674 7880
rect 19889 7871 19947 7877
rect 19889 7837 19901 7871
rect 19935 7868 19947 7871
rect 19978 7868 19984 7880
rect 19935 7840 19984 7868
rect 19935 7837 19947 7840
rect 19889 7831 19947 7837
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 12728 7772 17632 7800
rect 17681 7803 17739 7809
rect 17681 7769 17693 7803
rect 17727 7769 17739 7803
rect 17681 7763 17739 7769
rect 18417 7803 18475 7809
rect 18417 7769 18429 7803
rect 18463 7800 18475 7803
rect 19242 7800 19248 7812
rect 18463 7772 19248 7800
rect 18463 7769 18475 7772
rect 18417 7763 18475 7769
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 15197 7735 15255 7741
rect 15197 7701 15209 7735
rect 15243 7732 15255 7735
rect 17126 7732 17132 7744
rect 15243 7704 17132 7732
rect 15243 7701 15255 7704
rect 15197 7695 15255 7701
rect 17126 7692 17132 7704
rect 17184 7732 17190 7744
rect 17696 7732 17724 7763
rect 19242 7760 19248 7772
rect 19300 7760 19306 7812
rect 19426 7760 19432 7812
rect 19484 7800 19490 7812
rect 20134 7803 20192 7809
rect 20134 7800 20146 7803
rect 19484 7772 20146 7800
rect 19484 7760 19490 7772
rect 20134 7769 20146 7772
rect 20180 7769 20192 7803
rect 20916 7800 20944 8044
rect 22189 8041 22201 8075
rect 22235 8072 22247 8075
rect 23566 8072 23572 8084
rect 22235 8044 23572 8072
rect 22235 8041 22247 8044
rect 22189 8035 22247 8041
rect 23566 8032 23572 8044
rect 23624 8032 23630 8084
rect 24670 8072 24676 8084
rect 24631 8044 24676 8072
rect 24670 8032 24676 8044
rect 24728 8032 24734 8084
rect 25133 8075 25191 8081
rect 25133 8041 25145 8075
rect 25179 8041 25191 8075
rect 25133 8035 25191 8041
rect 23750 7964 23756 8016
rect 23808 8004 23814 8016
rect 25148 8004 25176 8035
rect 25222 8032 25228 8084
rect 25280 8072 25286 8084
rect 28169 8075 28227 8081
rect 28169 8072 28181 8075
rect 25280 8044 28181 8072
rect 25280 8032 25286 8044
rect 28169 8041 28181 8044
rect 28215 8041 28227 8075
rect 31110 8072 31116 8084
rect 28169 8035 28227 8041
rect 28276 8044 30696 8072
rect 31071 8044 31116 8072
rect 27614 8004 27620 8016
rect 23808 7976 25176 8004
rect 27448 7976 27620 8004
rect 23808 7964 23814 7976
rect 22646 7936 22652 7948
rect 22607 7908 22652 7936
rect 22646 7896 22652 7908
rect 22704 7896 22710 7948
rect 25130 7896 25136 7948
rect 25188 7936 25194 7948
rect 25685 7939 25743 7945
rect 25685 7936 25697 7939
rect 25188 7908 25697 7936
rect 25188 7896 25194 7908
rect 25685 7905 25697 7908
rect 25731 7905 25743 7939
rect 25685 7899 25743 7905
rect 26418 7896 26424 7948
rect 26476 7936 26482 7948
rect 27341 7939 27399 7945
rect 27341 7936 27353 7939
rect 26476 7908 27353 7936
rect 26476 7896 26482 7908
rect 27341 7905 27353 7908
rect 27387 7905 27399 7939
rect 27341 7899 27399 7905
rect 22005 7871 22063 7877
rect 22005 7837 22017 7871
rect 22051 7868 22063 7871
rect 22462 7868 22468 7880
rect 22051 7840 22468 7868
rect 22051 7837 22063 7840
rect 22005 7831 22063 7837
rect 22462 7828 22468 7840
rect 22520 7828 22526 7880
rect 22554 7828 22560 7880
rect 22612 7868 22618 7880
rect 22905 7871 22963 7877
rect 22905 7868 22917 7871
rect 22612 7840 22917 7868
rect 22612 7828 22618 7840
rect 22905 7837 22917 7840
rect 22951 7837 22963 7871
rect 22905 7831 22963 7837
rect 23198 7828 23204 7880
rect 23256 7868 23262 7880
rect 27249 7871 27307 7877
rect 27249 7868 27261 7871
rect 23256 7840 27261 7868
rect 23256 7828 23262 7840
rect 27249 7837 27261 7840
rect 27295 7868 27307 7871
rect 27448 7868 27476 7976
rect 27614 7964 27620 7976
rect 27672 8004 27678 8016
rect 28276 8004 28304 8044
rect 27672 7976 28304 8004
rect 30668 8004 30696 8044
rect 31110 8032 31116 8044
rect 31168 8032 31174 8084
rect 32214 8072 32220 8084
rect 32175 8044 32220 8072
rect 32214 8032 32220 8044
rect 32272 8032 32278 8084
rect 32306 8032 32312 8084
rect 32364 8072 32370 8084
rect 32677 8075 32735 8081
rect 32677 8072 32689 8075
rect 32364 8044 32689 8072
rect 32364 8032 32370 8044
rect 32677 8041 32689 8044
rect 32723 8041 32735 8075
rect 33318 8072 33324 8084
rect 33279 8044 33324 8072
rect 32677 8035 32735 8041
rect 33318 8032 33324 8044
rect 33376 8032 33382 8084
rect 35526 8072 35532 8084
rect 35487 8044 35532 8072
rect 35526 8032 35532 8044
rect 35584 8032 35590 8084
rect 35894 8032 35900 8084
rect 35952 8072 35958 8084
rect 35989 8075 36047 8081
rect 35989 8072 36001 8075
rect 35952 8044 36001 8072
rect 35952 8032 35958 8044
rect 35989 8041 36001 8044
rect 36035 8041 36047 8075
rect 36630 8072 36636 8084
rect 36591 8044 36636 8072
rect 35989 8035 36047 8041
rect 36630 8032 36636 8044
rect 36688 8032 36694 8084
rect 52454 8072 52460 8084
rect 52415 8044 52460 8072
rect 52454 8032 52460 8044
rect 52512 8032 52518 8084
rect 36648 8004 36676 8032
rect 30668 7976 36676 8004
rect 27672 7964 27678 7976
rect 27525 7939 27583 7945
rect 27525 7905 27537 7939
rect 27571 7936 27583 7939
rect 29086 7936 29092 7948
rect 27571 7908 29092 7936
rect 27571 7905 27583 7908
rect 27525 7899 27583 7905
rect 28184 7877 28212 7908
rect 29086 7896 29092 7908
rect 29144 7896 29150 7948
rect 29178 7896 29184 7948
rect 29236 7936 29242 7948
rect 29730 7936 29736 7948
rect 29236 7908 29281 7936
rect 29691 7908 29736 7936
rect 29236 7896 29242 7908
rect 29730 7896 29736 7908
rect 29788 7896 29794 7948
rect 34514 7936 34520 7948
rect 33520 7908 34520 7936
rect 27295 7840 27476 7868
rect 28169 7871 28227 7877
rect 27295 7837 27307 7840
rect 27249 7831 27307 7837
rect 28169 7837 28181 7871
rect 28215 7837 28227 7871
rect 28169 7831 28227 7837
rect 28353 7871 28411 7877
rect 28353 7837 28365 7871
rect 28399 7868 28411 7871
rect 28626 7868 28632 7880
rect 28399 7840 28632 7868
rect 28399 7837 28411 7840
rect 28353 7831 28411 7837
rect 28626 7828 28632 7840
rect 28684 7828 28690 7880
rect 28994 7868 29000 7880
rect 28955 7840 29000 7868
rect 28994 7828 29000 7840
rect 29052 7828 29058 7880
rect 29196 7868 29224 7896
rect 31570 7868 31576 7880
rect 29196 7840 31576 7868
rect 31570 7828 31576 7840
rect 31628 7868 31634 7880
rect 33520 7877 33548 7908
rect 34514 7896 34520 7908
rect 34572 7896 34578 7948
rect 34977 7939 35035 7945
rect 34977 7905 34989 7939
rect 35023 7936 35035 7939
rect 37458 7936 37464 7948
rect 35023 7908 37464 7936
rect 35023 7905 35035 7908
rect 34977 7899 35035 7905
rect 33505 7871 33563 7877
rect 31628 7840 31754 7868
rect 31628 7828 31634 7840
rect 24302 7800 24308 7812
rect 20916 7772 24308 7800
rect 20134 7763 20192 7769
rect 24302 7760 24308 7772
rect 24360 7800 24366 7812
rect 24762 7800 24768 7812
rect 24360 7772 24768 7800
rect 24360 7760 24366 7772
rect 24762 7760 24768 7772
rect 24820 7760 24826 7812
rect 25593 7803 25651 7809
rect 25593 7800 25605 7803
rect 24872 7772 25605 7800
rect 24872 7744 24900 7772
rect 25593 7769 25605 7772
rect 25639 7769 25651 7803
rect 28718 7800 28724 7812
rect 25593 7763 25651 7769
rect 26252 7772 28724 7800
rect 17184 7704 17724 7732
rect 18509 7735 18567 7741
rect 17184 7692 17190 7704
rect 18509 7701 18521 7735
rect 18555 7732 18567 7735
rect 18598 7732 18604 7744
rect 18555 7704 18604 7732
rect 18555 7701 18567 7704
rect 18509 7695 18567 7701
rect 18598 7692 18604 7704
rect 18656 7692 18662 7744
rect 18877 7735 18935 7741
rect 18877 7701 18889 7735
rect 18923 7732 18935 7735
rect 19334 7732 19340 7744
rect 18923 7704 19340 7732
rect 18923 7701 18935 7704
rect 18877 7695 18935 7701
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 21266 7732 21272 7744
rect 21227 7704 21272 7732
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 24029 7735 24087 7741
rect 24029 7701 24041 7735
rect 24075 7732 24087 7735
rect 24854 7732 24860 7744
rect 24075 7704 24860 7732
rect 24075 7701 24087 7704
rect 24029 7695 24087 7701
rect 24854 7692 24860 7704
rect 24912 7692 24918 7744
rect 25501 7735 25559 7741
rect 25501 7701 25513 7735
rect 25547 7732 25559 7735
rect 26252 7732 26280 7772
rect 28718 7760 28724 7772
rect 28776 7760 28782 7812
rect 30000 7803 30058 7809
rect 30000 7769 30012 7803
rect 30046 7800 30058 7803
rect 30374 7800 30380 7812
rect 30046 7772 30380 7800
rect 30046 7769 30058 7772
rect 30000 7763 30058 7769
rect 30374 7760 30380 7772
rect 30432 7760 30438 7812
rect 31726 7800 31754 7840
rect 33505 7837 33517 7871
rect 33551 7837 33563 7871
rect 33505 7831 33563 7837
rect 33689 7871 33747 7877
rect 33689 7837 33701 7871
rect 33735 7868 33747 7871
rect 33870 7868 33876 7880
rect 33735 7840 33876 7868
rect 33735 7837 33747 7840
rect 33689 7831 33747 7837
rect 33704 7800 33732 7831
rect 33870 7828 33876 7840
rect 33928 7868 33934 7880
rect 34992 7868 35020 7899
rect 37458 7896 37464 7908
rect 37516 7896 37522 7948
rect 33928 7840 35020 7868
rect 51813 7871 51871 7877
rect 33928 7828 33934 7840
rect 51813 7837 51825 7871
rect 51859 7868 51871 7871
rect 52270 7868 52276 7880
rect 51859 7840 52276 7868
rect 51859 7837 51871 7840
rect 51813 7831 51871 7837
rect 52270 7828 52276 7840
rect 52328 7828 52334 7880
rect 52914 7868 52920 7880
rect 52875 7840 52920 7868
rect 52914 7828 52920 7840
rect 52972 7828 52978 7880
rect 31726 7772 33732 7800
rect 52730 7760 52736 7812
rect 52788 7800 52794 7812
rect 53162 7803 53220 7809
rect 53162 7800 53174 7803
rect 52788 7772 53174 7800
rect 52788 7760 52794 7772
rect 53162 7769 53174 7772
rect 53208 7769 53220 7803
rect 53162 7763 53220 7769
rect 26418 7732 26424 7744
rect 25547 7704 26280 7732
rect 26379 7704 26424 7732
rect 25547 7701 25559 7704
rect 25501 7695 25559 7701
rect 26418 7692 26424 7704
rect 26476 7692 26482 7744
rect 26878 7732 26884 7744
rect 26839 7704 26884 7732
rect 26878 7692 26884 7704
rect 26936 7692 26942 7744
rect 28350 7692 28356 7744
rect 28408 7732 28414 7744
rect 28813 7735 28871 7741
rect 28813 7732 28825 7735
rect 28408 7704 28825 7732
rect 28408 7692 28414 7704
rect 28813 7701 28825 7704
rect 28859 7701 28871 7735
rect 28813 7695 28871 7701
rect 30190 7692 30196 7744
rect 30248 7732 30254 7744
rect 30558 7732 30564 7744
rect 30248 7704 30564 7732
rect 30248 7692 30254 7704
rect 30558 7692 30564 7704
rect 30616 7732 30622 7744
rect 31573 7735 31631 7741
rect 31573 7732 31585 7735
rect 30616 7704 31585 7732
rect 30616 7692 30622 7704
rect 31573 7701 31585 7704
rect 31619 7701 31631 7735
rect 31573 7695 31631 7701
rect 34054 7692 34060 7744
rect 34112 7732 34118 7744
rect 34149 7735 34207 7741
rect 34149 7732 34161 7735
rect 34112 7704 34161 7732
rect 34112 7692 34118 7704
rect 34149 7701 34161 7704
rect 34195 7732 34207 7735
rect 34238 7732 34244 7744
rect 34195 7704 34244 7732
rect 34195 7701 34207 7704
rect 34149 7695 34207 7701
rect 34238 7692 34244 7704
rect 34296 7692 34302 7744
rect 39666 7692 39672 7744
rect 39724 7732 39730 7744
rect 51074 7732 51080 7744
rect 39724 7704 51080 7732
rect 39724 7692 39730 7704
rect 51074 7692 51080 7704
rect 51132 7692 51138 7744
rect 54294 7732 54300 7744
rect 54255 7704 54300 7732
rect 54294 7692 54300 7704
rect 54352 7692 54358 7744
rect 1104 7642 54832 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 54832 7642
rect 1104 7568 54832 7590
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 12621 7531 12679 7537
rect 12621 7528 12633 7531
rect 11112 7500 12633 7528
rect 11112 7488 11118 7500
rect 12621 7497 12633 7500
rect 12667 7497 12679 7531
rect 13722 7528 13728 7540
rect 13683 7500 13728 7528
rect 12621 7491 12679 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 15746 7528 15752 7540
rect 15707 7500 15752 7528
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 17218 7528 17224 7540
rect 17179 7500 17224 7528
rect 17218 7488 17224 7500
rect 17276 7488 17282 7540
rect 18598 7488 18604 7540
rect 18656 7528 18662 7540
rect 22186 7528 22192 7540
rect 18656 7500 22192 7528
rect 18656 7488 18662 7500
rect 22186 7488 22192 7500
rect 22244 7488 22250 7540
rect 22373 7531 22431 7537
rect 22373 7497 22385 7531
rect 22419 7528 22431 7531
rect 23198 7528 23204 7540
rect 22419 7500 23204 7528
rect 22419 7497 22431 7500
rect 22373 7491 22431 7497
rect 23198 7488 23204 7500
rect 23256 7488 23262 7540
rect 27246 7488 27252 7540
rect 27304 7528 27310 7540
rect 27341 7531 27399 7537
rect 27341 7528 27353 7531
rect 27304 7500 27353 7528
rect 27304 7488 27310 7500
rect 27341 7497 27353 7500
rect 27387 7497 27399 7531
rect 27341 7491 27399 7497
rect 28994 7488 29000 7540
rect 29052 7528 29058 7540
rect 29181 7531 29239 7537
rect 29181 7528 29193 7531
rect 29052 7500 29193 7528
rect 29052 7488 29058 7500
rect 29181 7497 29193 7500
rect 29227 7497 29239 7531
rect 30374 7528 30380 7540
rect 30335 7500 30380 7528
rect 29181 7491 29239 7497
rect 30374 7488 30380 7500
rect 30432 7488 30438 7540
rect 30926 7488 30932 7540
rect 30984 7528 30990 7540
rect 31021 7531 31079 7537
rect 31021 7528 31033 7531
rect 30984 7500 31033 7528
rect 30984 7488 30990 7500
rect 31021 7497 31033 7500
rect 31067 7528 31079 7531
rect 33413 7531 33471 7537
rect 33413 7528 33425 7531
rect 31067 7500 33425 7528
rect 31067 7497 31079 7500
rect 31021 7491 31079 7497
rect 33413 7497 33425 7500
rect 33459 7497 33471 7531
rect 33413 7491 33471 7497
rect 33778 7488 33784 7540
rect 33836 7528 33842 7540
rect 33965 7531 34023 7537
rect 33965 7528 33977 7531
rect 33836 7500 33977 7528
rect 33836 7488 33842 7500
rect 33965 7497 33977 7500
rect 34011 7528 34023 7531
rect 34517 7531 34575 7537
rect 34517 7528 34529 7531
rect 34011 7500 34529 7528
rect 34011 7497 34023 7500
rect 33965 7491 34023 7497
rect 34517 7497 34529 7500
rect 34563 7528 34575 7531
rect 35069 7531 35127 7537
rect 35069 7528 35081 7531
rect 34563 7500 35081 7528
rect 34563 7497 34575 7500
rect 34517 7491 34575 7497
rect 35069 7497 35081 7500
rect 35115 7528 35127 7531
rect 35894 7528 35900 7540
rect 35115 7500 35900 7528
rect 35115 7497 35127 7500
rect 35069 7491 35127 7497
rect 35894 7488 35900 7500
rect 35952 7488 35958 7540
rect 48774 7488 48780 7540
rect 48832 7528 48838 7540
rect 52365 7531 52423 7537
rect 52365 7528 52377 7531
rect 48832 7500 52377 7528
rect 48832 7488 48838 7500
rect 52365 7497 52377 7500
rect 52411 7528 52423 7531
rect 52914 7528 52920 7540
rect 52411 7500 52920 7528
rect 52411 7497 52423 7500
rect 52365 7491 52423 7497
rect 52914 7488 52920 7500
rect 52972 7488 52978 7540
rect 53190 7528 53196 7540
rect 53151 7500 53196 7528
rect 53190 7488 53196 7500
rect 53248 7488 53254 7540
rect 13740 7460 13768 7488
rect 12452 7432 13768 7460
rect 17681 7463 17739 7469
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 11054 7392 11060 7404
rect 1903 7364 11060 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 11054 7352 11060 7364
rect 11112 7352 11118 7404
rect 12452 7324 12480 7432
rect 17681 7429 17693 7463
rect 17727 7429 17739 7463
rect 19978 7460 19984 7472
rect 17681 7423 17739 7429
rect 18248 7432 19984 7460
rect 12526 7352 12532 7404
rect 12584 7392 12590 7404
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 12584 7364 13093 7392
rect 12584 7352 12590 7364
rect 13081 7361 13093 7364
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7392 16359 7395
rect 17126 7392 17132 7404
rect 16347 7364 17132 7392
rect 16347 7361 16359 7364
rect 16301 7355 16359 7361
rect 17126 7352 17132 7364
rect 17184 7392 17190 7404
rect 17494 7392 17500 7404
rect 17184 7364 17500 7392
rect 17184 7352 17190 7364
rect 17494 7352 17500 7364
rect 17552 7392 17558 7404
rect 17696 7392 17724 7423
rect 18248 7401 18276 7432
rect 19978 7420 19984 7432
rect 20036 7460 20042 7472
rect 20036 7432 21496 7460
rect 20036 7420 20042 7432
rect 17552 7364 17724 7392
rect 18233 7395 18291 7401
rect 17552 7352 17558 7364
rect 18233 7361 18245 7395
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 18322 7352 18328 7404
rect 18380 7392 18386 7404
rect 18489 7395 18547 7401
rect 18489 7392 18501 7395
rect 18380 7364 18501 7392
rect 18380 7352 18386 7364
rect 18489 7361 18501 7364
rect 18535 7361 18547 7395
rect 18489 7355 18547 7361
rect 19058 7352 19064 7404
rect 19116 7392 19122 7404
rect 21197 7395 21255 7401
rect 19116 7364 19288 7392
rect 19116 7352 19122 7364
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 12452 7296 12817 7324
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 1670 7188 1676 7200
rect 1631 7160 1676 7188
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 12912 7188 12940 7287
rect 12986 7284 12992 7336
rect 13044 7324 13050 7336
rect 13446 7324 13452 7336
rect 13044 7296 13452 7324
rect 13044 7284 13050 7296
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 17405 7259 17463 7265
rect 15580 7228 17356 7256
rect 15580 7188 15608 7228
rect 12912 7160 15608 7188
rect 17328 7188 17356 7228
rect 17405 7225 17417 7259
rect 17451 7256 17463 7259
rect 17954 7256 17960 7268
rect 17451 7228 17960 7256
rect 17451 7225 17463 7228
rect 17405 7219 17463 7225
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 19260 7256 19288 7364
rect 21197 7361 21209 7395
rect 21243 7392 21255 7395
rect 21358 7392 21364 7404
rect 21243 7364 21364 7392
rect 21243 7361 21255 7364
rect 21197 7355 21255 7361
rect 21358 7352 21364 7364
rect 21416 7352 21422 7404
rect 21468 7333 21496 7432
rect 22278 7420 22284 7472
rect 22336 7460 22342 7472
rect 26878 7460 26884 7472
rect 22336 7432 25084 7460
rect 22336 7420 22342 7432
rect 22002 7352 22008 7404
rect 22060 7392 22066 7404
rect 24785 7395 24843 7401
rect 22060 7364 22600 7392
rect 22060 7352 22066 7364
rect 21453 7327 21511 7333
rect 21453 7293 21465 7327
rect 21499 7324 21511 7327
rect 22278 7324 22284 7336
rect 21499 7296 22284 7324
rect 21499 7293 21511 7296
rect 21453 7287 21511 7293
rect 22278 7284 22284 7296
rect 22336 7284 22342 7336
rect 22572 7333 22600 7364
rect 24785 7361 24797 7395
rect 24831 7392 24843 7395
rect 24946 7392 24952 7404
rect 24831 7364 24952 7392
rect 24831 7361 24843 7364
rect 24785 7355 24843 7361
rect 24946 7352 24952 7364
rect 25004 7352 25010 7404
rect 25056 7401 25084 7432
rect 26252 7432 26884 7460
rect 26252 7401 26280 7432
rect 26878 7420 26884 7432
rect 26936 7420 26942 7472
rect 28629 7463 28687 7469
rect 28629 7429 28641 7463
rect 28675 7460 28687 7463
rect 30650 7460 30656 7472
rect 28675 7432 30656 7460
rect 28675 7429 28687 7432
rect 28629 7423 28687 7429
rect 30650 7420 30656 7432
rect 30708 7420 30714 7472
rect 30742 7420 30748 7472
rect 30800 7460 30806 7472
rect 32309 7463 32367 7469
rect 32309 7460 32321 7463
rect 30800 7432 32321 7460
rect 30800 7420 30806 7432
rect 32309 7429 32321 7432
rect 32355 7429 32367 7463
rect 32309 7423 32367 7429
rect 49694 7420 49700 7472
rect 49752 7460 49758 7472
rect 53837 7463 53895 7469
rect 53837 7460 53849 7463
rect 49752 7432 53849 7460
rect 49752 7420 49758 7432
rect 53837 7429 53849 7432
rect 53883 7429 53895 7463
rect 53837 7423 53895 7429
rect 25041 7395 25099 7401
rect 25041 7361 25053 7395
rect 25087 7361 25099 7395
rect 25041 7355 25099 7361
rect 26237 7395 26295 7401
rect 26237 7361 26249 7395
rect 26283 7361 26295 7395
rect 26237 7355 26295 7361
rect 26421 7395 26479 7401
rect 26421 7361 26433 7395
rect 26467 7392 26479 7395
rect 27157 7395 27215 7401
rect 27157 7392 27169 7395
rect 26467 7364 27169 7392
rect 26467 7361 26479 7364
rect 26421 7355 26479 7361
rect 27157 7361 27169 7364
rect 27203 7361 27215 7395
rect 27157 7355 27215 7361
rect 27893 7395 27951 7401
rect 27893 7361 27905 7395
rect 27939 7392 27951 7395
rect 28350 7392 28356 7404
rect 27939 7364 28356 7392
rect 27939 7361 27951 7364
rect 27893 7355 27951 7361
rect 28350 7352 28356 7364
rect 28408 7352 28414 7404
rect 28534 7392 28540 7404
rect 28495 7364 28540 7392
rect 28534 7352 28540 7364
rect 28592 7352 28598 7404
rect 29178 7392 29184 7404
rect 28644 7364 29184 7392
rect 22465 7327 22523 7333
rect 22465 7293 22477 7327
rect 22511 7293 22523 7327
rect 22465 7287 22523 7293
rect 22557 7327 22615 7333
rect 22557 7293 22569 7327
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 26053 7327 26111 7333
rect 26053 7293 26065 7327
rect 26099 7324 26111 7327
rect 28644 7324 28672 7364
rect 29178 7352 29184 7364
rect 29236 7352 29242 7404
rect 29362 7352 29368 7404
rect 29420 7392 29426 7404
rect 29549 7395 29607 7401
rect 29549 7392 29561 7395
rect 29420 7364 29561 7392
rect 29420 7352 29426 7364
rect 29549 7361 29561 7364
rect 29595 7361 29607 7395
rect 29549 7355 29607 7361
rect 29641 7395 29699 7401
rect 29641 7361 29653 7395
rect 29687 7392 29699 7395
rect 30561 7395 30619 7401
rect 29687 7364 29868 7392
rect 29687 7361 29699 7364
rect 29641 7355 29699 7361
rect 26099 7296 28672 7324
rect 26099 7293 26111 7296
rect 26053 7287 26111 7293
rect 20073 7259 20131 7265
rect 20073 7256 20085 7259
rect 19260 7228 20085 7256
rect 20073 7225 20085 7228
rect 20119 7225 20131 7259
rect 22480 7256 22508 7287
rect 29086 7284 29092 7336
rect 29144 7324 29150 7336
rect 29733 7327 29791 7333
rect 29144 7296 29592 7324
rect 29144 7284 29150 7296
rect 20073 7219 20131 7225
rect 21468 7228 22508 7256
rect 25593 7259 25651 7265
rect 19613 7191 19671 7197
rect 19613 7188 19625 7191
rect 17328 7160 19625 7188
rect 19613 7157 19625 7160
rect 19659 7188 19671 7191
rect 19978 7188 19984 7200
rect 19659 7160 19984 7188
rect 19659 7157 19671 7160
rect 19613 7151 19671 7157
rect 19978 7148 19984 7160
rect 20036 7148 20042 7200
rect 20088 7188 20116 7219
rect 21468 7188 21496 7228
rect 25593 7225 25605 7259
rect 25639 7256 25651 7259
rect 27982 7256 27988 7268
rect 25639 7228 27988 7256
rect 25639 7225 25651 7228
rect 25593 7219 25651 7225
rect 20088 7160 21496 7188
rect 21634 7148 21640 7200
rect 21692 7188 21698 7200
rect 22005 7191 22063 7197
rect 22005 7188 22017 7191
rect 21692 7160 22017 7188
rect 21692 7148 21698 7160
rect 22005 7157 22017 7160
rect 22051 7157 22063 7191
rect 22005 7151 22063 7157
rect 23566 7148 23572 7200
rect 23624 7188 23630 7200
rect 23661 7191 23719 7197
rect 23661 7188 23673 7191
rect 23624 7160 23673 7188
rect 23624 7148 23630 7160
rect 23661 7157 23673 7160
rect 23707 7157 23719 7191
rect 23661 7151 23719 7157
rect 24762 7148 24768 7200
rect 24820 7188 24826 7200
rect 25608 7188 25636 7219
rect 27982 7216 27988 7228
rect 28040 7216 28046 7268
rect 28077 7259 28135 7265
rect 28077 7225 28089 7259
rect 28123 7256 28135 7259
rect 29454 7256 29460 7268
rect 28123 7228 29460 7256
rect 28123 7225 28135 7228
rect 28077 7219 28135 7225
rect 29454 7216 29460 7228
rect 29512 7216 29518 7268
rect 29564 7256 29592 7296
rect 29733 7293 29745 7327
rect 29779 7293 29791 7327
rect 29840 7324 29868 7364
rect 30561 7361 30573 7395
rect 30607 7392 30619 7395
rect 31202 7392 31208 7404
rect 30607 7364 31208 7392
rect 30607 7361 30619 7364
rect 30561 7355 30619 7361
rect 31202 7352 31208 7364
rect 31260 7352 31266 7404
rect 53374 7392 53380 7404
rect 53335 7364 53380 7392
rect 53374 7352 53380 7364
rect 53432 7352 53438 7404
rect 54205 7395 54263 7401
rect 54205 7361 54217 7395
rect 54251 7392 54263 7395
rect 54386 7392 54392 7404
rect 54251 7364 54392 7392
rect 54251 7361 54263 7364
rect 54205 7355 54263 7361
rect 54386 7352 54392 7364
rect 54444 7352 54450 7404
rect 31018 7324 31024 7336
rect 29840 7296 31024 7324
rect 29733 7287 29791 7293
rect 29748 7256 29776 7287
rect 31018 7284 31024 7296
rect 31076 7284 31082 7336
rect 32861 7327 32919 7333
rect 32861 7324 32873 7327
rect 31726 7296 32873 7324
rect 29564 7228 29776 7256
rect 30282 7216 30288 7268
rect 30340 7256 30346 7268
rect 31726 7256 31754 7296
rect 32861 7293 32873 7296
rect 32907 7293 32919 7327
rect 32861 7287 32919 7293
rect 30340 7228 31754 7256
rect 30340 7216 30346 7228
rect 24820 7160 25636 7188
rect 24820 7148 24826 7160
rect 26418 7148 26424 7200
rect 26476 7188 26482 7200
rect 30834 7188 30840 7200
rect 26476 7160 30840 7188
rect 26476 7148 26482 7160
rect 30834 7148 30840 7160
rect 30892 7188 30898 7200
rect 31570 7188 31576 7200
rect 30892 7160 31576 7188
rect 30892 7148 30898 7160
rect 31570 7148 31576 7160
rect 31628 7148 31634 7200
rect 1104 7098 54832 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 54832 7098
rect 1104 7024 54832 7046
rect 18233 6987 18291 6993
rect 18233 6953 18245 6987
rect 18279 6984 18291 6987
rect 18598 6984 18604 6996
rect 18279 6956 18604 6984
rect 18279 6953 18291 6956
rect 18233 6947 18291 6953
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 21358 6944 21364 6996
rect 21416 6984 21422 6996
rect 21453 6987 21511 6993
rect 21453 6984 21465 6987
rect 21416 6956 21465 6984
rect 21416 6944 21422 6956
rect 21453 6953 21465 6956
rect 21499 6953 21511 6987
rect 21453 6947 21511 6953
rect 22186 6944 22192 6996
rect 22244 6984 22250 6996
rect 22244 6956 24900 6984
rect 22244 6944 22250 6956
rect 17221 6919 17279 6925
rect 17221 6885 17233 6919
rect 17267 6885 17279 6919
rect 24872 6916 24900 6956
rect 24946 6944 24952 6996
rect 25004 6984 25010 6996
rect 25777 6987 25835 6993
rect 25777 6984 25789 6987
rect 25004 6956 25789 6984
rect 25004 6944 25010 6956
rect 25777 6953 25789 6956
rect 25823 6953 25835 6987
rect 33870 6984 33876 6996
rect 33831 6956 33876 6984
rect 25777 6947 25835 6953
rect 33870 6944 33876 6956
rect 33928 6944 33934 6996
rect 53374 6944 53380 6996
rect 53432 6984 53438 6996
rect 53469 6987 53527 6993
rect 53469 6984 53481 6987
rect 53432 6956 53481 6984
rect 53432 6944 53438 6956
rect 53469 6953 53481 6956
rect 53515 6953 53527 6987
rect 54110 6984 54116 6996
rect 54071 6956 54116 6984
rect 53469 6947 53527 6953
rect 54110 6944 54116 6956
rect 54168 6944 54174 6996
rect 29362 6916 29368 6928
rect 24872 6888 29368 6916
rect 17221 6879 17279 6885
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 13081 6851 13139 6857
rect 13081 6848 13093 6851
rect 11112 6820 13093 6848
rect 11112 6808 11118 6820
rect 13081 6817 13093 6820
rect 13127 6817 13139 6851
rect 13081 6811 13139 6817
rect 13357 6851 13415 6857
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 17236 6848 17264 6879
rect 29362 6876 29368 6888
rect 29420 6876 29426 6928
rect 17402 6848 17408 6860
rect 13403 6820 14504 6848
rect 17236 6820 17408 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 12986 6780 12992 6792
rect 1903 6752 12992 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 12986 6740 12992 6752
rect 13044 6740 13050 6792
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 13096 6752 13277 6780
rect 13096 6724 13124 6752
rect 13265 6749 13277 6752
rect 13311 6749 13323 6783
rect 13446 6780 13452 6792
rect 13407 6752 13452 6780
rect 13265 6743 13323 6749
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 13538 6740 13544 6792
rect 13596 6780 13602 6792
rect 13596 6752 13641 6780
rect 13596 6740 13602 6752
rect 13078 6672 13084 6724
rect 13136 6672 13142 6724
rect 14369 6715 14427 6721
rect 14369 6712 14381 6715
rect 13280 6684 14381 6712
rect 1670 6644 1676 6656
rect 1631 6616 1676 6644
rect 1670 6604 1676 6616
rect 1728 6604 1734 6656
rect 12066 6604 12072 6656
rect 12124 6644 12130 6656
rect 13280 6644 13308 6684
rect 14369 6681 14381 6684
rect 14415 6681 14427 6715
rect 14476 6712 14504 6820
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 17494 6808 17500 6860
rect 17552 6848 17558 6860
rect 20809 6851 20867 6857
rect 17552 6820 17597 6848
rect 18616 6820 19840 6848
rect 17552 6808 17558 6820
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 15197 6783 15255 6789
rect 15197 6780 15209 6783
rect 14599 6752 15209 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 15197 6749 15209 6752
rect 15243 6780 15255 6783
rect 17512 6780 17540 6808
rect 15243 6752 17540 6780
rect 15243 6749 15255 6752
rect 15197 6743 15255 6749
rect 18616 6712 18644 6820
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6780 18751 6783
rect 18782 6780 18788 6792
rect 18739 6752 18788 6780
rect 18739 6749 18751 6752
rect 18693 6743 18751 6749
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 19426 6740 19432 6792
rect 19484 6740 19490 6792
rect 19812 6780 19840 6820
rect 20809 6817 20821 6851
rect 20855 6848 20867 6851
rect 22278 6848 22284 6860
rect 20855 6820 22284 6848
rect 20855 6817 20867 6820
rect 20809 6811 20867 6817
rect 22278 6808 22284 6820
rect 22336 6808 22342 6860
rect 24765 6851 24823 6857
rect 24765 6817 24777 6851
rect 24811 6848 24823 6851
rect 25130 6848 25136 6860
rect 24811 6820 25136 6848
rect 24811 6817 24823 6820
rect 24765 6811 24823 6817
rect 25130 6808 25136 6820
rect 25188 6808 25194 6860
rect 26510 6848 26516 6860
rect 25424 6820 26096 6848
rect 26471 6820 26516 6848
rect 21634 6780 21640 6792
rect 19812 6752 20668 6780
rect 21595 6752 21640 6780
rect 19444 6712 19472 6740
rect 14476 6684 18644 6712
rect 18892 6684 19472 6712
rect 14369 6675 14427 6681
rect 12124 6616 13308 6644
rect 17037 6647 17095 6653
rect 12124 6604 12130 6616
rect 17037 6613 17049 6647
rect 17083 6644 17095 6647
rect 17678 6644 17684 6656
rect 17083 6616 17684 6644
rect 17083 6613 17095 6616
rect 17037 6607 17095 6613
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 18892 6653 18920 6684
rect 19978 6672 19984 6724
rect 20036 6712 20042 6724
rect 20542 6715 20600 6721
rect 20542 6712 20554 6715
rect 20036 6684 20554 6712
rect 20036 6672 20042 6684
rect 20542 6681 20554 6684
rect 20588 6681 20600 6715
rect 20640 6712 20668 6752
rect 21634 6740 21640 6752
rect 21692 6740 21698 6792
rect 22296 6780 22324 6808
rect 24029 6783 24087 6789
rect 24029 6780 24041 6783
rect 22296 6752 24041 6780
rect 24029 6749 24041 6752
rect 24075 6749 24087 6783
rect 24029 6743 24087 6749
rect 24949 6783 25007 6789
rect 24949 6749 24961 6783
rect 24995 6780 25007 6783
rect 25314 6780 25320 6792
rect 24995 6752 25320 6780
rect 24995 6749 25007 6752
rect 24949 6743 25007 6749
rect 25314 6740 25320 6752
rect 25372 6740 25378 6792
rect 23566 6712 23572 6724
rect 20640 6684 23572 6712
rect 20542 6675 20600 6681
rect 23566 6672 23572 6684
rect 23624 6672 23630 6724
rect 23658 6672 23664 6724
rect 23716 6712 23722 6724
rect 23762 6715 23820 6721
rect 23762 6712 23774 6715
rect 23716 6684 23774 6712
rect 23716 6672 23722 6684
rect 23762 6681 23774 6684
rect 23808 6681 23820 6715
rect 23762 6675 23820 6681
rect 24670 6672 24676 6724
rect 24728 6712 24734 6724
rect 25424 6712 25452 6820
rect 25961 6783 26019 6789
rect 25961 6749 25973 6783
rect 26007 6749 26019 6783
rect 25961 6743 26019 6749
rect 24728 6684 25452 6712
rect 24728 6672 24734 6684
rect 18877 6647 18935 6653
rect 18877 6613 18889 6647
rect 18923 6613 18935 6647
rect 18877 6607 18935 6613
rect 19242 6604 19248 6656
rect 19300 6644 19306 6656
rect 19429 6647 19487 6653
rect 19429 6644 19441 6647
rect 19300 6616 19441 6644
rect 19300 6604 19306 6616
rect 19429 6613 19441 6616
rect 19475 6613 19487 6647
rect 22186 6644 22192 6656
rect 22099 6616 22192 6644
rect 19429 6607 19487 6613
rect 22186 6604 22192 6616
rect 22244 6644 22250 6656
rect 22370 6644 22376 6656
rect 22244 6616 22376 6644
rect 22244 6604 22250 6616
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 22649 6647 22707 6653
rect 22649 6613 22661 6647
rect 22695 6644 22707 6647
rect 22830 6644 22836 6656
rect 22695 6616 22836 6644
rect 22695 6613 22707 6616
rect 22649 6607 22707 6613
rect 22830 6604 22836 6616
rect 22888 6604 22894 6656
rect 23584 6644 23612 6672
rect 24857 6647 24915 6653
rect 24857 6644 24869 6647
rect 23584 6616 24869 6644
rect 24857 6613 24869 6616
rect 24903 6613 24915 6647
rect 24857 6607 24915 6613
rect 25317 6647 25375 6653
rect 25317 6613 25329 6647
rect 25363 6644 25375 6647
rect 25976 6644 26004 6743
rect 26068 6712 26096 6820
rect 26510 6808 26516 6820
rect 26568 6808 26574 6860
rect 27338 6808 27344 6860
rect 27396 6848 27402 6860
rect 27709 6851 27767 6857
rect 27709 6848 27721 6851
rect 27396 6820 27721 6848
rect 27396 6808 27402 6820
rect 27709 6817 27721 6820
rect 27755 6848 27767 6851
rect 27890 6848 27896 6860
rect 27755 6820 27896 6848
rect 27755 6817 27767 6820
rect 27709 6811 27767 6817
rect 27890 6808 27896 6820
rect 27948 6808 27954 6860
rect 29546 6808 29552 6860
rect 29604 6848 29610 6860
rect 29733 6851 29791 6857
rect 29733 6848 29745 6851
rect 29604 6820 29745 6848
rect 29604 6808 29610 6820
rect 29733 6817 29745 6820
rect 29779 6817 29791 6851
rect 29733 6811 29791 6817
rect 30466 6808 30472 6860
rect 30524 6848 30530 6860
rect 30837 6851 30895 6857
rect 30837 6848 30849 6851
rect 30524 6820 30849 6848
rect 30524 6808 30530 6820
rect 30837 6817 30849 6820
rect 30883 6817 30895 6851
rect 30837 6811 30895 6817
rect 31386 6808 31392 6860
rect 31444 6848 31450 6860
rect 31941 6851 31999 6857
rect 31941 6848 31953 6851
rect 31444 6820 31953 6848
rect 31444 6808 31450 6820
rect 31941 6817 31953 6820
rect 31987 6817 31999 6851
rect 33042 6848 33048 6860
rect 33003 6820 33048 6848
rect 31941 6811 31999 6817
rect 33042 6808 33048 6820
rect 33100 6808 33106 6860
rect 43714 6808 43720 6860
rect 43772 6848 43778 6860
rect 51258 6848 51264 6860
rect 43772 6820 51264 6848
rect 43772 6808 43778 6820
rect 51258 6808 51264 6820
rect 51316 6808 51322 6860
rect 30374 6780 30380 6792
rect 30287 6752 30380 6780
rect 30374 6740 30380 6752
rect 30432 6780 30438 6792
rect 31294 6780 31300 6792
rect 30432 6752 31300 6780
rect 30432 6740 30438 6752
rect 31294 6740 31300 6752
rect 31352 6740 31358 6792
rect 44910 6740 44916 6792
rect 44968 6780 44974 6792
rect 49970 6780 49976 6792
rect 44968 6752 49976 6780
rect 44968 6740 44974 6752
rect 49970 6740 49976 6752
rect 50028 6740 50034 6792
rect 54294 6780 54300 6792
rect 54255 6752 54300 6780
rect 54294 6740 54300 6752
rect 54352 6740 54358 6792
rect 26973 6715 27031 6721
rect 26973 6712 26985 6715
rect 26068 6684 26985 6712
rect 26973 6681 26985 6684
rect 27019 6681 27031 6715
rect 26973 6675 27031 6681
rect 27062 6672 27068 6724
rect 27120 6712 27126 6724
rect 29089 6715 29147 6721
rect 29089 6712 29101 6715
rect 27120 6684 29101 6712
rect 27120 6672 27126 6684
rect 29089 6681 29101 6684
rect 29135 6681 29147 6715
rect 29089 6675 29147 6681
rect 29362 6672 29368 6724
rect 29420 6712 29426 6724
rect 30006 6712 30012 6724
rect 29420 6684 30012 6712
rect 29420 6672 29426 6684
rect 30006 6672 30012 6684
rect 30064 6712 30070 6724
rect 31389 6715 31447 6721
rect 31389 6712 31401 6715
rect 30064 6684 31401 6712
rect 30064 6672 30070 6684
rect 31389 6681 31401 6684
rect 31435 6681 31447 6715
rect 31389 6675 31447 6681
rect 31570 6672 31576 6724
rect 31628 6712 31634 6724
rect 32493 6715 32551 6721
rect 32493 6712 32505 6715
rect 31628 6684 32505 6712
rect 31628 6672 31634 6684
rect 32493 6681 32505 6684
rect 32539 6681 32551 6715
rect 32493 6675 32551 6681
rect 25363 6616 26004 6644
rect 28629 6647 28687 6653
rect 25363 6613 25375 6616
rect 25317 6607 25375 6613
rect 28629 6613 28641 6647
rect 28675 6644 28687 6647
rect 28994 6644 29000 6656
rect 28675 6616 29000 6644
rect 28675 6613 28687 6616
rect 28629 6607 28687 6613
rect 28994 6604 29000 6616
rect 29052 6604 29058 6656
rect 1104 6554 54832 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 54832 6554
rect 1104 6480 54832 6502
rect 12526 6440 12532 6452
rect 12487 6412 12532 6440
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 12986 6440 12992 6452
rect 12947 6412 12992 6440
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 14093 6443 14151 6449
rect 14093 6440 14105 6443
rect 13136 6412 14105 6440
rect 13136 6400 13142 6412
rect 8294 6332 8300 6384
rect 8352 6372 8358 6384
rect 12434 6372 12440 6384
rect 8352 6344 12440 6372
rect 8352 6332 8358 6344
rect 12434 6332 12440 6344
rect 12492 6332 12498 6384
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 13078 6304 13084 6316
rect 1903 6276 13084 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13188 6313 13216 6412
rect 14093 6409 14105 6412
rect 14139 6440 14151 6443
rect 14182 6440 14188 6452
rect 14139 6412 14188 6440
rect 14139 6409 14151 6412
rect 14093 6403 14151 6409
rect 14182 6400 14188 6412
rect 14240 6440 14246 6452
rect 14553 6443 14611 6449
rect 14553 6440 14565 6443
rect 14240 6412 14565 6440
rect 14240 6400 14246 6412
rect 14553 6409 14565 6412
rect 14599 6409 14611 6443
rect 14553 6403 14611 6409
rect 17313 6443 17371 6449
rect 17313 6409 17325 6443
rect 17359 6440 17371 6443
rect 17494 6440 17500 6452
rect 17359 6412 17500 6440
rect 17359 6409 17371 6412
rect 17313 6403 17371 6409
rect 17494 6400 17500 6412
rect 17552 6440 17558 6452
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 17552 6412 17785 6440
rect 17552 6400 17558 6412
rect 17773 6409 17785 6412
rect 17819 6409 17831 6443
rect 17773 6403 17831 6409
rect 18506 6400 18512 6452
rect 18564 6440 18570 6452
rect 18693 6443 18751 6449
rect 18693 6440 18705 6443
rect 18564 6412 18705 6440
rect 18564 6400 18570 6412
rect 18693 6409 18705 6412
rect 18739 6409 18751 6443
rect 18693 6403 18751 6409
rect 19521 6443 19579 6449
rect 19521 6409 19533 6443
rect 19567 6440 19579 6443
rect 19978 6440 19984 6452
rect 19567 6412 19984 6440
rect 19567 6409 19579 6412
rect 19521 6403 19579 6409
rect 19978 6400 19984 6412
rect 20036 6400 20042 6452
rect 20162 6440 20168 6452
rect 20123 6412 20168 6440
rect 20162 6400 20168 6412
rect 20220 6400 20226 6452
rect 20714 6440 20720 6452
rect 20675 6412 20720 6440
rect 20714 6400 20720 6412
rect 20772 6400 20778 6452
rect 21450 6440 21456 6452
rect 21411 6412 21456 6440
rect 21450 6400 21456 6412
rect 21508 6400 21514 6452
rect 22465 6443 22523 6449
rect 22465 6409 22477 6443
rect 22511 6440 22523 6443
rect 23106 6440 23112 6452
rect 22511 6412 23112 6440
rect 22511 6409 22523 6412
rect 22465 6403 22523 6409
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 23658 6440 23664 6452
rect 23619 6412 23664 6440
rect 23658 6400 23664 6412
rect 23716 6400 23722 6452
rect 24949 6443 25007 6449
rect 24949 6409 24961 6443
rect 24995 6440 25007 6443
rect 25038 6440 25044 6452
rect 24995 6412 25044 6440
rect 24995 6409 25007 6412
rect 24949 6403 25007 6409
rect 25038 6400 25044 6412
rect 25096 6400 25102 6452
rect 25314 6400 25320 6452
rect 25372 6440 25378 6452
rect 25774 6440 25780 6452
rect 25372 6412 25780 6440
rect 25372 6400 25378 6412
rect 25774 6400 25780 6412
rect 25832 6400 25838 6452
rect 26605 6443 26663 6449
rect 26605 6409 26617 6443
rect 26651 6440 26663 6443
rect 27062 6440 27068 6452
rect 26651 6412 27068 6440
rect 26651 6409 26663 6412
rect 26605 6403 26663 6409
rect 27062 6400 27068 6412
rect 27120 6400 27126 6452
rect 27617 6443 27675 6449
rect 27617 6409 27629 6443
rect 27663 6440 27675 6443
rect 28629 6443 28687 6449
rect 28629 6440 28641 6443
rect 27663 6412 28641 6440
rect 27663 6409 27675 6412
rect 27617 6403 27675 6409
rect 28629 6409 28641 6412
rect 28675 6440 28687 6443
rect 29178 6440 29184 6452
rect 28675 6412 29184 6440
rect 28675 6409 28687 6412
rect 28629 6403 28687 6409
rect 29178 6400 29184 6412
rect 29236 6400 29242 6452
rect 29917 6443 29975 6449
rect 29917 6409 29929 6443
rect 29963 6440 29975 6443
rect 30466 6440 30472 6452
rect 29963 6412 30472 6440
rect 29963 6409 29975 6412
rect 29917 6403 29975 6409
rect 30466 6400 30472 6412
rect 30524 6400 30530 6452
rect 31478 6440 31484 6452
rect 31439 6412 31484 6440
rect 31478 6400 31484 6412
rect 31536 6400 31542 6452
rect 32401 6443 32459 6449
rect 32401 6409 32413 6443
rect 32447 6440 32459 6443
rect 33042 6440 33048 6452
rect 32447 6412 33048 6440
rect 32447 6409 32459 6412
rect 32401 6403 32459 6409
rect 25056 6372 25084 6400
rect 28077 6375 28135 6381
rect 28077 6372 28089 6375
rect 13280 6344 16344 6372
rect 25056 6344 28089 6372
rect 13280 6313 13308 6344
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6273 13231 6307
rect 13173 6267 13231 6273
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6273 13323 6307
rect 13265 6267 13323 6273
rect 12066 6236 12072 6248
rect 12027 6208 12072 6236
rect 12066 6196 12072 6208
rect 12124 6196 12130 6248
rect 12986 6236 12992 6248
rect 12268 6208 12992 6236
rect 10870 6128 10876 6180
rect 10928 6168 10934 6180
rect 12268 6168 12296 6208
rect 12986 6196 12992 6208
rect 13044 6236 13050 6248
rect 13357 6239 13415 6245
rect 13357 6236 13369 6239
rect 13044 6208 13369 6236
rect 13044 6196 13050 6208
rect 13357 6205 13369 6208
rect 13403 6205 13415 6239
rect 13357 6199 13415 6205
rect 13449 6239 13507 6245
rect 13449 6205 13461 6239
rect 13495 6205 13507 6239
rect 16316 6236 16344 6344
rect 28077 6341 28089 6344
rect 28123 6341 28135 6375
rect 28077 6335 28135 6341
rect 31021 6375 31079 6381
rect 31021 6341 31033 6375
rect 31067 6372 31079 6375
rect 31570 6372 31576 6384
rect 31067 6344 31576 6372
rect 31067 6341 31079 6344
rect 31021 6335 31079 6341
rect 31570 6332 31576 6344
rect 31628 6332 31634 6384
rect 18877 6307 18935 6313
rect 18877 6273 18889 6307
rect 18923 6304 18935 6307
rect 18966 6304 18972 6316
rect 18923 6276 18972 6304
rect 18923 6273 18935 6276
rect 18877 6267 18935 6273
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 19334 6304 19340 6316
rect 19295 6276 19340 6304
rect 19334 6264 19340 6276
rect 19392 6264 19398 6316
rect 23477 6307 23535 6313
rect 23477 6273 23489 6307
rect 23523 6304 23535 6307
rect 24578 6304 24584 6316
rect 23523 6276 24584 6304
rect 23523 6273 23535 6276
rect 23477 6267 23535 6273
rect 24578 6264 24584 6276
rect 24636 6264 24642 6316
rect 27430 6264 27436 6316
rect 27488 6304 27494 6316
rect 29730 6304 29736 6316
rect 27488 6276 29736 6304
rect 27488 6264 27494 6276
rect 29730 6264 29736 6276
rect 29788 6304 29794 6316
rect 30282 6304 30288 6316
rect 29788 6276 30288 6304
rect 29788 6264 29794 6276
rect 30282 6264 30288 6276
rect 30340 6264 30346 6316
rect 30469 6307 30527 6313
rect 30469 6273 30481 6307
rect 30515 6304 30527 6307
rect 30558 6304 30564 6316
rect 30515 6276 30564 6304
rect 30515 6273 30527 6276
rect 30469 6267 30527 6273
rect 30558 6264 30564 6276
rect 30616 6264 30622 6316
rect 24486 6236 24492 6248
rect 16316 6208 24492 6236
rect 13449 6199 13507 6205
rect 10928 6140 12296 6168
rect 12345 6171 12403 6177
rect 10928 6128 10934 6140
rect 12345 6137 12357 6171
rect 12391 6168 12403 6171
rect 12710 6168 12716 6180
rect 12391 6140 12716 6168
rect 12391 6137 12403 6140
rect 12345 6131 12403 6137
rect 12710 6128 12716 6140
rect 12768 6128 12774 6180
rect 12802 6128 12808 6180
rect 12860 6168 12866 6180
rect 13464 6168 13492 6199
rect 24486 6196 24492 6208
rect 24544 6236 24550 6248
rect 25041 6239 25099 6245
rect 25041 6236 25053 6239
rect 24544 6208 25053 6236
rect 24544 6196 24550 6208
rect 25041 6205 25053 6208
rect 25087 6205 25099 6239
rect 25041 6199 25099 6205
rect 25130 6196 25136 6248
rect 25188 6236 25194 6248
rect 29365 6239 29423 6245
rect 25188 6208 25233 6236
rect 25188 6196 25194 6208
rect 29365 6205 29377 6239
rect 29411 6236 29423 6239
rect 32416 6236 32444 6403
rect 33042 6400 33048 6412
rect 33100 6400 33106 6452
rect 54297 6443 54355 6449
rect 54297 6409 54309 6443
rect 54343 6440 54355 6443
rect 54386 6440 54392 6452
rect 54343 6412 54392 6440
rect 54343 6409 54355 6412
rect 54297 6403 54355 6409
rect 54386 6400 54392 6412
rect 54444 6400 54450 6452
rect 29411 6208 32444 6236
rect 29411 6205 29423 6208
rect 29365 6199 29423 6205
rect 12860 6140 13492 6168
rect 12860 6128 12866 6140
rect 22462 6128 22468 6180
rect 22520 6168 22526 6180
rect 24581 6171 24639 6177
rect 24581 6168 24593 6171
rect 22520 6140 24593 6168
rect 22520 6128 22526 6140
rect 24581 6137 24593 6140
rect 24627 6137 24639 6171
rect 24581 6131 24639 6137
rect 24670 6128 24676 6180
rect 24728 6168 24734 6180
rect 29380 6168 29408 6199
rect 24728 6140 29408 6168
rect 24728 6128 24734 6140
rect 44818 6128 44824 6180
rect 44876 6168 44882 6180
rect 51534 6168 51540 6180
rect 44876 6140 51540 6168
rect 44876 6128 44882 6140
rect 51534 6128 51540 6140
rect 51592 6128 51598 6180
rect 1670 6100 1676 6112
rect 1631 6072 1676 6100
rect 1670 6060 1676 6072
rect 1728 6060 1734 6112
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 17218 6100 17224 6112
rect 12492 6072 17224 6100
rect 12492 6060 12498 6072
rect 17218 6060 17224 6072
rect 17276 6060 17282 6112
rect 23017 6103 23075 6109
rect 23017 6069 23029 6103
rect 23063 6100 23075 6103
rect 24210 6100 24216 6112
rect 23063 6072 24216 6100
rect 23063 6069 23075 6072
rect 23017 6063 23075 6069
rect 24210 6060 24216 6072
rect 24268 6100 24274 6112
rect 24688 6100 24716 6128
rect 24268 6072 24716 6100
rect 24268 6060 24274 6072
rect 1104 6010 54832 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 54832 6010
rect 1104 5936 54832 5958
rect 12621 5899 12679 5905
rect 12621 5865 12633 5899
rect 12667 5896 12679 5899
rect 12894 5896 12900 5908
rect 12667 5868 12900 5896
rect 12667 5865 12679 5868
rect 12621 5859 12679 5865
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 13078 5896 13084 5908
rect 13039 5868 13084 5896
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 13446 5896 13452 5908
rect 13188 5868 13452 5896
rect 11514 5828 11520 5840
rect 11475 5800 11520 5828
rect 11514 5788 11520 5800
rect 11572 5788 11578 5840
rect 12526 5828 12532 5840
rect 12487 5800 12532 5828
rect 12526 5788 12532 5800
rect 12584 5788 12590 5840
rect 12986 5788 12992 5840
rect 13044 5828 13050 5840
rect 13188 5828 13216 5868
rect 13446 5856 13452 5868
rect 13504 5896 13510 5908
rect 22925 5899 22983 5905
rect 13504 5868 13676 5896
rect 13504 5856 13510 5868
rect 13538 5828 13544 5840
rect 13044 5800 13216 5828
rect 13280 5800 13544 5828
rect 13044 5788 13050 5800
rect 11701 5763 11759 5769
rect 11701 5729 11713 5763
rect 11747 5760 11759 5763
rect 13280 5760 13308 5800
rect 13538 5788 13544 5800
rect 13596 5788 13602 5840
rect 11747 5732 13308 5760
rect 13449 5763 13507 5769
rect 11747 5729 11759 5732
rect 11701 5723 11759 5729
rect 13449 5729 13461 5763
rect 13495 5760 13507 5763
rect 13648 5760 13676 5868
rect 22925 5865 22937 5899
rect 22971 5896 22983 5899
rect 23198 5896 23204 5908
rect 22971 5868 23204 5896
rect 22971 5865 22983 5868
rect 22925 5859 22983 5865
rect 23198 5856 23204 5868
rect 23256 5856 23262 5908
rect 24029 5899 24087 5905
rect 24029 5865 24041 5899
rect 24075 5896 24087 5899
rect 24118 5896 24124 5908
rect 24075 5868 24124 5896
rect 24075 5865 24087 5868
rect 24029 5859 24087 5865
rect 24118 5856 24124 5868
rect 24176 5856 24182 5908
rect 24670 5896 24676 5908
rect 24631 5868 24676 5896
rect 24670 5856 24676 5868
rect 24728 5856 24734 5908
rect 25225 5899 25283 5905
rect 25225 5865 25237 5899
rect 25271 5896 25283 5899
rect 26050 5896 26056 5908
rect 25271 5868 26056 5896
rect 25271 5865 25283 5868
rect 25225 5859 25283 5865
rect 26050 5856 26056 5868
rect 26108 5896 26114 5908
rect 27893 5899 27951 5905
rect 27893 5896 27905 5899
rect 26108 5868 27905 5896
rect 26108 5856 26114 5868
rect 27893 5865 27905 5868
rect 27939 5865 27951 5899
rect 27893 5859 27951 5865
rect 28537 5899 28595 5905
rect 28537 5865 28549 5899
rect 28583 5896 28595 5899
rect 28718 5896 28724 5908
rect 28583 5868 28724 5896
rect 28583 5865 28595 5868
rect 28537 5859 28595 5865
rect 28718 5856 28724 5868
rect 28776 5856 28782 5908
rect 30466 5856 30472 5908
rect 30524 5896 30530 5908
rect 30745 5899 30803 5905
rect 30745 5896 30757 5899
rect 30524 5868 30757 5896
rect 30524 5856 30530 5868
rect 30745 5865 30757 5868
rect 30791 5865 30803 5899
rect 30745 5859 30803 5865
rect 21450 5788 21456 5840
rect 21508 5828 21514 5840
rect 26237 5831 26295 5837
rect 26237 5828 26249 5831
rect 21508 5800 26249 5828
rect 21508 5788 21514 5800
rect 26237 5797 26249 5800
rect 26283 5797 26295 5831
rect 26237 5791 26295 5797
rect 26973 5763 27031 5769
rect 26973 5760 26985 5763
rect 13495 5732 13676 5760
rect 19306 5732 26985 5760
rect 13495 5729 13507 5732
rect 13449 5723 13507 5729
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 12434 5692 12440 5704
rect 1903 5664 12440 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 12434 5652 12440 5664
rect 12492 5652 12498 5704
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 13265 5695 13323 5701
rect 13265 5692 13277 5695
rect 12676 5664 13277 5692
rect 12676 5652 12682 5664
rect 13265 5661 13277 5664
rect 13311 5661 13323 5695
rect 13265 5655 13323 5661
rect 13357 5695 13415 5701
rect 13357 5661 13369 5695
rect 13403 5661 13415 5695
rect 13538 5692 13544 5704
rect 13499 5664 13544 5692
rect 13357 5655 13415 5661
rect 11241 5627 11299 5633
rect 11241 5593 11253 5627
rect 11287 5624 11299 5627
rect 11698 5624 11704 5636
rect 11287 5596 11704 5624
rect 11287 5593 11299 5596
rect 11241 5587 11299 5593
rect 11698 5584 11704 5596
rect 11756 5624 11762 5636
rect 12066 5624 12072 5636
rect 11756 5596 12072 5624
rect 11756 5584 11762 5596
rect 12066 5584 12072 5596
rect 12124 5624 12130 5636
rect 12161 5627 12219 5633
rect 12161 5624 12173 5627
rect 12124 5596 12173 5624
rect 12124 5584 12130 5596
rect 12161 5593 12173 5596
rect 12207 5593 12219 5627
rect 12161 5587 12219 5593
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 10689 5559 10747 5565
rect 10689 5525 10701 5559
rect 10735 5556 10747 5559
rect 11146 5556 11152 5568
rect 10735 5528 11152 5556
rect 10735 5525 10747 5528
rect 10689 5519 10747 5525
rect 11146 5516 11152 5528
rect 11204 5516 11210 5568
rect 13280 5556 13308 5655
rect 13372 5624 13400 5655
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 17218 5652 17224 5704
rect 17276 5692 17282 5704
rect 19306 5692 19334 5732
rect 26973 5729 26985 5732
rect 27019 5760 27031 5763
rect 27154 5760 27160 5772
rect 27019 5732 27160 5760
rect 27019 5729 27031 5732
rect 26973 5723 27031 5729
rect 27154 5720 27160 5732
rect 27212 5720 27218 5772
rect 17276 5664 19334 5692
rect 17276 5652 17282 5664
rect 23106 5652 23112 5704
rect 23164 5692 23170 5704
rect 23385 5695 23443 5701
rect 23385 5692 23397 5695
rect 23164 5664 23397 5692
rect 23164 5652 23170 5664
rect 23385 5661 23397 5664
rect 23431 5661 23443 5695
rect 23385 5655 23443 5661
rect 24302 5652 24308 5704
rect 24360 5692 24366 5704
rect 25777 5695 25835 5701
rect 25777 5692 25789 5695
rect 24360 5664 25789 5692
rect 24360 5652 24366 5664
rect 25777 5661 25789 5664
rect 25823 5692 25835 5695
rect 26142 5692 26148 5704
rect 25823 5664 26148 5692
rect 25823 5661 25835 5664
rect 25777 5655 25835 5661
rect 26142 5652 26148 5664
rect 26200 5652 26206 5704
rect 28994 5692 29000 5704
rect 26252 5664 29000 5692
rect 19242 5624 19248 5636
rect 13372 5596 19248 5624
rect 19242 5584 19248 5596
rect 19300 5584 19306 5636
rect 26252 5624 26280 5664
rect 28994 5652 29000 5664
rect 29052 5652 29058 5704
rect 30285 5695 30343 5701
rect 30285 5661 30297 5695
rect 30331 5692 30343 5695
rect 30466 5692 30472 5704
rect 30331 5664 30472 5692
rect 30331 5661 30343 5664
rect 30285 5655 30343 5661
rect 30466 5652 30472 5664
rect 30524 5652 30530 5704
rect 24136 5596 26280 5624
rect 14369 5559 14427 5565
rect 14369 5556 14381 5559
rect 13280 5528 14381 5556
rect 14369 5525 14381 5528
rect 14415 5556 14427 5559
rect 24136 5556 24164 5596
rect 26326 5584 26332 5636
rect 26384 5624 26390 5636
rect 30009 5627 30067 5633
rect 30009 5624 30021 5627
rect 26384 5596 30021 5624
rect 26384 5584 26390 5596
rect 30009 5593 30021 5596
rect 30055 5624 30067 5627
rect 37458 5624 37464 5636
rect 30055 5596 37464 5624
rect 30055 5593 30067 5596
rect 30009 5587 30067 5593
rect 37458 5584 37464 5596
rect 37516 5584 37522 5636
rect 14415 5528 24164 5556
rect 14415 5525 14427 5528
rect 14369 5519 14427 5525
rect 25774 5516 25780 5568
rect 25832 5556 25838 5568
rect 28997 5559 29055 5565
rect 28997 5556 29009 5559
rect 25832 5528 29009 5556
rect 25832 5516 25838 5528
rect 28997 5525 29009 5528
rect 29043 5525 29055 5559
rect 28997 5519 29055 5525
rect 32766 5516 32772 5568
rect 32824 5556 32830 5568
rect 34606 5556 34612 5568
rect 32824 5528 34612 5556
rect 32824 5516 32830 5528
rect 34606 5516 34612 5528
rect 34664 5516 34670 5568
rect 1104 5466 54832 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 54832 5466
rect 1104 5392 54832 5414
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 12492 5324 12537 5352
rect 12492 5312 12498 5324
rect 16022 5312 16028 5364
rect 16080 5352 16086 5364
rect 22830 5352 22836 5364
rect 16080 5324 22836 5352
rect 16080 5312 16086 5324
rect 22830 5312 22836 5324
rect 22888 5312 22894 5364
rect 24489 5355 24547 5361
rect 24489 5321 24501 5355
rect 24535 5352 24547 5355
rect 25038 5352 25044 5364
rect 24535 5324 25044 5352
rect 24535 5321 24547 5324
rect 24489 5315 24547 5321
rect 25038 5312 25044 5324
rect 25096 5312 25102 5364
rect 25593 5355 25651 5361
rect 25593 5321 25605 5355
rect 25639 5352 25651 5355
rect 25866 5352 25872 5364
rect 25639 5324 25872 5352
rect 25639 5321 25651 5324
rect 25593 5315 25651 5321
rect 25866 5312 25872 5324
rect 25924 5312 25930 5364
rect 25958 5312 25964 5364
rect 26016 5352 26022 5364
rect 26053 5355 26111 5361
rect 26053 5352 26065 5355
rect 26016 5324 26065 5352
rect 26016 5312 26022 5324
rect 26053 5321 26065 5324
rect 26099 5321 26111 5355
rect 26053 5315 26111 5321
rect 27614 5312 27620 5364
rect 27672 5352 27678 5364
rect 27709 5355 27767 5361
rect 27709 5352 27721 5355
rect 27672 5324 27721 5352
rect 27672 5312 27678 5324
rect 27709 5321 27721 5324
rect 27755 5321 27767 5355
rect 27709 5315 27767 5321
rect 28537 5355 28595 5361
rect 28537 5321 28549 5355
rect 28583 5352 28595 5355
rect 28626 5352 28632 5364
rect 28583 5324 28632 5352
rect 28583 5321 28595 5324
rect 28537 5315 28595 5321
rect 28626 5312 28632 5324
rect 28684 5312 28690 5364
rect 30006 5352 30012 5364
rect 29967 5324 30012 5352
rect 30006 5312 30012 5324
rect 30064 5312 30070 5364
rect 30466 5312 30472 5364
rect 30524 5352 30530 5364
rect 30561 5355 30619 5361
rect 30561 5352 30573 5355
rect 30524 5324 30573 5352
rect 30524 5312 30530 5324
rect 30561 5321 30573 5324
rect 30607 5321 30619 5355
rect 30561 5315 30619 5321
rect 14461 5287 14519 5293
rect 14461 5284 14473 5287
rect 12636 5256 13124 5284
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 10502 5216 10508 5228
rect 1903 5188 10508 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 12636 5225 12664 5256
rect 12617 5219 12675 5225
rect 12617 5185 12629 5219
rect 12663 5185 12675 5219
rect 12617 5179 12675 5185
rect 12894 5176 12900 5228
rect 12952 5216 12958 5228
rect 13096 5216 13124 5256
rect 14108 5256 14473 5284
rect 14108 5216 14136 5256
rect 14461 5253 14473 5256
rect 14507 5284 14519 5287
rect 14826 5284 14832 5296
rect 14507 5256 14832 5284
rect 14507 5253 14519 5256
rect 14461 5247 14519 5253
rect 14826 5244 14832 5256
rect 14884 5284 14890 5296
rect 37550 5284 37556 5296
rect 14884 5256 37556 5284
rect 14884 5244 14890 5256
rect 37550 5244 37556 5256
rect 37608 5284 37614 5296
rect 38378 5284 38384 5296
rect 37608 5256 38384 5284
rect 37608 5244 37614 5256
rect 38378 5244 38384 5256
rect 38436 5244 38442 5296
rect 12952 5188 12997 5216
rect 13096 5188 14136 5216
rect 12952 5176 12958 5188
rect 14182 5176 14188 5228
rect 14240 5216 14246 5228
rect 14921 5219 14979 5225
rect 14921 5216 14933 5219
rect 14240 5188 14933 5216
rect 14240 5176 14246 5188
rect 14921 5185 14933 5188
rect 14967 5185 14979 5219
rect 14921 5179 14979 5185
rect 27249 5219 27307 5225
rect 27249 5185 27261 5219
rect 27295 5216 27307 5219
rect 29178 5216 29184 5228
rect 27295 5188 29184 5216
rect 27295 5185 27307 5188
rect 27249 5179 27307 5185
rect 29178 5176 29184 5188
rect 29236 5216 29242 5228
rect 29273 5219 29331 5225
rect 29273 5216 29285 5219
rect 29236 5188 29285 5216
rect 29236 5176 29242 5188
rect 29273 5185 29285 5188
rect 29319 5185 29331 5219
rect 29273 5179 29331 5185
rect 7098 5108 7104 5160
rect 7156 5148 7162 5160
rect 12434 5148 12440 5160
rect 7156 5120 12440 5148
rect 7156 5108 7162 5120
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 12714 5151 12772 5157
rect 12714 5117 12726 5151
rect 12760 5117 12772 5151
rect 12714 5111 12772 5117
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5117 12863 5151
rect 13446 5148 13452 5160
rect 13407 5120 13452 5148
rect 12805 5111 12863 5117
rect 10597 5083 10655 5089
rect 10597 5049 10609 5083
rect 10643 5080 10655 5083
rect 11790 5080 11796 5092
rect 10643 5052 11796 5080
rect 10643 5049 10655 5052
rect 10597 5043 10655 5049
rect 11790 5040 11796 5052
rect 11848 5040 11854 5092
rect 1670 5012 1676 5024
rect 1631 4984 1676 5012
rect 1670 4972 1676 4984
rect 1728 4972 1734 5024
rect 9309 5015 9367 5021
rect 9309 4981 9321 5015
rect 9355 5012 9367 5015
rect 9582 5012 9588 5024
rect 9355 4984 9588 5012
rect 9355 4981 9367 4984
rect 9309 4975 9367 4981
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 9858 5012 9864 5024
rect 9819 4984 9864 5012
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 10744 4984 11161 5012
rect 10744 4972 10750 4984
rect 11149 4981 11161 4984
rect 11195 5012 11207 5015
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11195 4984 11713 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11701 4981 11713 4984
rect 11747 5012 11759 5015
rect 12342 5012 12348 5024
rect 11747 4984 12348 5012
rect 11747 4981 11759 4984
rect 11701 4975 11759 4981
rect 12342 4972 12348 4984
rect 12400 4972 12406 5024
rect 12728 5012 12756 5111
rect 12820 5080 12848 5111
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 25866 5148 25872 5160
rect 13872 5120 25872 5148
rect 13872 5108 13878 5120
rect 25866 5108 25872 5120
rect 25924 5108 25930 5160
rect 12986 5080 12992 5092
rect 12820 5052 12992 5080
rect 12986 5040 12992 5052
rect 13044 5040 13050 5092
rect 13722 5040 13728 5092
rect 13780 5080 13786 5092
rect 13909 5083 13967 5089
rect 13780 5052 13825 5080
rect 13780 5040 13786 5052
rect 13909 5049 13921 5083
rect 13955 5080 13967 5083
rect 14734 5080 14740 5092
rect 13955 5052 14740 5080
rect 13955 5049 13967 5052
rect 13909 5043 13967 5049
rect 14734 5040 14740 5052
rect 14792 5040 14798 5092
rect 18138 5040 18144 5092
rect 18196 5080 18202 5092
rect 26878 5080 26884 5092
rect 18196 5052 26884 5080
rect 18196 5040 18202 5052
rect 26878 5040 26884 5052
rect 26936 5040 26942 5092
rect 16022 5012 16028 5024
rect 12728 4984 16028 5012
rect 16022 4972 16028 4984
rect 16080 4972 16086 5024
rect 24946 5012 24952 5024
rect 24907 4984 24952 5012
rect 24946 4972 24952 4984
rect 25004 4972 25010 5024
rect 1104 4922 54832 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 54832 4922
rect 1104 4848 54832 4870
rect 10502 4808 10508 4820
rect 10463 4780 10508 4808
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 12529 4811 12587 4817
rect 12529 4777 12541 4811
rect 12575 4808 12587 4811
rect 12802 4808 12808 4820
rect 12575 4780 12808 4808
rect 12575 4777 12587 4780
rect 12529 4771 12587 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 12989 4811 13047 4817
rect 12989 4808 13001 4811
rect 12952 4780 13001 4808
rect 12952 4768 12958 4780
rect 12989 4777 13001 4780
rect 13035 4777 13047 4811
rect 12989 4771 13047 4777
rect 25133 4811 25191 4817
rect 25133 4777 25145 4811
rect 25179 4808 25191 4811
rect 25774 4808 25780 4820
rect 25179 4780 25780 4808
rect 25179 4777 25191 4780
rect 25133 4771 25191 4777
rect 25774 4768 25780 4780
rect 25832 4768 25838 4820
rect 26237 4811 26295 4817
rect 26237 4777 26249 4811
rect 26283 4808 26295 4811
rect 28718 4808 28724 4820
rect 26283 4780 28724 4808
rect 26283 4777 26295 4780
rect 26237 4771 26295 4777
rect 28718 4768 28724 4780
rect 28776 4768 28782 4820
rect 38378 4808 38384 4820
rect 38339 4780 38384 4808
rect 38378 4768 38384 4780
rect 38436 4768 38442 4820
rect 41417 4811 41475 4817
rect 41417 4777 41429 4811
rect 41463 4808 41475 4811
rect 41690 4808 41696 4820
rect 41463 4780 41696 4808
rect 41463 4777 41475 4780
rect 41417 4771 41475 4777
rect 41690 4768 41696 4780
rect 41748 4768 41754 4820
rect 42426 4808 42432 4820
rect 42387 4780 42432 4808
rect 42426 4768 42432 4780
rect 42484 4768 42490 4820
rect 42978 4808 42984 4820
rect 42939 4780 42984 4808
rect 42978 4768 42984 4780
rect 43036 4768 43042 4820
rect 11238 4700 11244 4752
rect 11296 4740 11302 4752
rect 12345 4743 12403 4749
rect 12345 4740 12357 4743
rect 11296 4712 12357 4740
rect 11296 4700 11302 4712
rect 12345 4709 12357 4712
rect 12391 4709 12403 4743
rect 13078 4740 13084 4752
rect 13039 4712 13084 4740
rect 12345 4703 12403 4709
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 26878 4700 26884 4752
rect 26936 4740 26942 4752
rect 46934 4740 46940 4752
rect 26936 4712 46940 4740
rect 26936 4700 26942 4712
rect 46934 4700 46940 4712
rect 46992 4700 46998 4752
rect 10781 4675 10839 4681
rect 10781 4641 10793 4675
rect 10827 4672 10839 4675
rect 21266 4672 21272 4684
rect 10827 4644 21272 4672
rect 10827 4641 10839 4644
rect 10781 4635 10839 4641
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 23290 4632 23296 4684
rect 23348 4672 23354 4684
rect 27430 4672 27436 4684
rect 23348 4644 27436 4672
rect 23348 4632 23354 4644
rect 27430 4632 27436 4644
rect 27488 4632 27494 4684
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4604 1915 4607
rect 10502 4604 10508 4616
rect 1903 4576 10508 4604
rect 1903 4573 1915 4576
rect 1857 4567 1915 4573
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 10686 4604 10692 4616
rect 10647 4576 10692 4604
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 10870 4604 10876 4616
rect 10831 4576 10876 4604
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 10962 4564 10968 4616
rect 11020 4604 11026 4616
rect 12802 4604 12808 4616
rect 11020 4576 11065 4604
rect 11164 4576 12808 4604
rect 11020 4564 11026 4576
rect 7377 4539 7435 4545
rect 7377 4505 7389 4539
rect 7423 4536 7435 4539
rect 8662 4536 8668 4548
rect 7423 4508 8668 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 10045 4539 10103 4545
rect 10045 4505 10057 4539
rect 10091 4536 10103 4539
rect 11164 4536 11192 4576
rect 12802 4564 12808 4576
rect 12860 4564 12866 4616
rect 14553 4607 14611 4613
rect 14553 4573 14565 4607
rect 14599 4604 14611 4607
rect 15194 4604 15200 4616
rect 14599 4576 15200 4604
rect 14599 4573 14611 4576
rect 14553 4567 14611 4573
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 45554 4604 45560 4616
rect 45515 4576 45560 4604
rect 45554 4564 45560 4576
rect 45612 4564 45618 4616
rect 10091 4508 11192 4536
rect 10091 4505 10103 4508
rect 10045 4499 10103 4505
rect 11698 4496 11704 4548
rect 11756 4536 11762 4548
rect 12069 4539 12127 4545
rect 12069 4536 12081 4539
rect 11756 4508 12081 4536
rect 11756 4496 11762 4508
rect 12069 4505 12081 4508
rect 12115 4536 12127 4539
rect 13446 4536 13452 4548
rect 12115 4508 13452 4536
rect 12115 4505 12127 4508
rect 12069 4499 12127 4505
rect 13446 4496 13452 4508
rect 13504 4496 13510 4548
rect 13906 4496 13912 4548
rect 13964 4536 13970 4548
rect 15289 4539 15347 4545
rect 15289 4536 15301 4539
rect 13964 4508 15301 4536
rect 13964 4496 13970 4508
rect 15289 4505 15301 4508
rect 15335 4505 15347 4539
rect 15289 4499 15347 4505
rect 22554 4496 22560 4548
rect 22612 4536 22618 4548
rect 22741 4539 22799 4545
rect 22741 4536 22753 4539
rect 22612 4508 22753 4536
rect 22612 4496 22618 4508
rect 22741 4505 22753 4508
rect 22787 4536 22799 4539
rect 32398 4536 32404 4548
rect 22787 4508 32404 4536
rect 22787 4505 22799 4508
rect 22741 4499 22799 4505
rect 32398 4496 32404 4508
rect 32456 4496 32462 4548
rect 1670 4468 1676 4480
rect 1631 4440 1676 4468
rect 1670 4428 1676 4440
rect 1728 4428 1734 4480
rect 7742 4428 7748 4480
rect 7800 4468 7806 4480
rect 8021 4471 8079 4477
rect 8021 4468 8033 4471
rect 7800 4440 8033 4468
rect 7800 4428 7806 4440
rect 8021 4437 8033 4440
rect 8067 4437 8079 4471
rect 8021 4431 8079 4437
rect 9493 4471 9551 4477
rect 9493 4437 9505 4471
rect 9539 4468 9551 4471
rect 10778 4468 10784 4480
rect 9539 4440 10784 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11606 4468 11612 4480
rect 11567 4440 11612 4468
rect 11606 4428 11612 4440
rect 11664 4428 11670 4480
rect 12986 4428 12992 4480
rect 13044 4468 13050 4480
rect 14550 4468 14556 4480
rect 13044 4440 14556 4468
rect 13044 4428 13050 4440
rect 14550 4428 14556 4440
rect 14608 4468 14614 4480
rect 14737 4471 14795 4477
rect 14737 4468 14749 4471
rect 14608 4440 14749 4468
rect 14608 4428 14614 4440
rect 14737 4437 14749 4440
rect 14783 4437 14795 4471
rect 23290 4468 23296 4480
rect 23251 4440 23296 4468
rect 14737 4431 14795 4437
rect 23290 4428 23296 4440
rect 23348 4428 23354 4480
rect 23658 4428 23664 4480
rect 23716 4468 23722 4480
rect 23753 4471 23811 4477
rect 23753 4468 23765 4471
rect 23716 4440 23765 4468
rect 23716 4428 23722 4440
rect 23753 4437 23765 4440
rect 23799 4437 23811 4471
rect 23753 4431 23811 4437
rect 25406 4428 25412 4480
rect 25464 4468 25470 4480
rect 25593 4471 25651 4477
rect 25593 4468 25605 4471
rect 25464 4440 25605 4468
rect 25464 4428 25470 4440
rect 25593 4437 25605 4440
rect 25639 4437 25651 4471
rect 25593 4431 25651 4437
rect 38654 4428 38660 4480
rect 38712 4468 38718 4480
rect 38933 4471 38991 4477
rect 38933 4468 38945 4471
rect 38712 4440 38945 4468
rect 38712 4428 38718 4440
rect 38933 4437 38945 4440
rect 38979 4437 38991 4471
rect 43622 4468 43628 4480
rect 43583 4440 43628 4468
rect 38933 4431 38991 4437
rect 43622 4428 43628 4440
rect 43680 4428 43686 4480
rect 45741 4471 45799 4477
rect 45741 4437 45753 4471
rect 45787 4468 45799 4471
rect 45922 4468 45928 4480
rect 45787 4440 45928 4468
rect 45787 4437 45799 4440
rect 45741 4431 45799 4437
rect 45922 4428 45928 4440
rect 45980 4428 45986 4480
rect 1104 4378 54832 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 54832 4378
rect 1104 4304 54832 4326
rect 10045 4267 10103 4273
rect 10045 4233 10057 4267
rect 10091 4264 10103 4267
rect 10962 4264 10968 4276
rect 10091 4236 10968 4264
rect 10091 4233 10103 4236
rect 10045 4227 10103 4233
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 25314 4224 25320 4276
rect 25372 4264 25378 4276
rect 25409 4267 25467 4273
rect 25409 4264 25421 4267
rect 25372 4236 25421 4264
rect 25372 4224 25378 4236
rect 25409 4233 25421 4236
rect 25455 4264 25467 4267
rect 25455 4236 26832 4264
rect 25455 4233 25467 4236
rect 25409 4227 25467 4233
rect 9125 4199 9183 4205
rect 9125 4165 9137 4199
rect 9171 4196 9183 4199
rect 10318 4196 10324 4208
rect 9171 4168 10324 4196
rect 9171 4165 9183 4168
rect 9125 4159 9183 4165
rect 10318 4156 10324 4168
rect 10376 4196 10382 4208
rect 10376 4168 10640 4196
rect 10376 4156 10382 4168
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 10410 4128 10416 4140
rect 1903 4100 10416 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 9582 4060 9588 4072
rect 9543 4032 9588 4060
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 10502 4060 10508 4072
rect 10463 4032 10508 4060
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 10612 4060 10640 4168
rect 12986 4156 12992 4208
rect 13044 4196 13050 4208
rect 13722 4196 13728 4208
rect 13044 4168 13728 4196
rect 13044 4156 13050 4168
rect 13722 4156 13728 4168
rect 13780 4156 13786 4208
rect 26326 4196 26332 4208
rect 25976 4168 26332 4196
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4128 10839 4131
rect 10827 4100 12296 4128
rect 10827 4097 10839 4100
rect 10781 4091 10839 4097
rect 10686 4060 10692 4072
rect 10612 4032 10692 4060
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 10870 4060 10876 4072
rect 10831 4032 10876 4060
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 10962 4020 10968 4072
rect 11020 4060 11026 4072
rect 11020 4032 11065 4060
rect 11020 4020 11026 4032
rect 11698 4020 11704 4072
rect 11756 4060 11762 4072
rect 11977 4063 12035 4069
rect 11977 4060 11989 4063
rect 11756 4032 11989 4060
rect 11756 4020 11762 4032
rect 11977 4029 11989 4032
rect 12023 4029 12035 4063
rect 12268 4060 12296 4100
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 22094 4128 22100 4140
rect 12400 4100 22100 4128
rect 12400 4088 12406 4100
rect 22094 4088 22100 4100
rect 22152 4128 22158 4140
rect 22649 4131 22707 4137
rect 22649 4128 22661 4131
rect 22152 4100 22661 4128
rect 22152 4088 22158 4100
rect 22649 4097 22661 4100
rect 22695 4128 22707 4131
rect 25976 4128 26004 4168
rect 26326 4156 26332 4168
rect 26384 4156 26390 4208
rect 22695 4100 26004 4128
rect 26053 4131 26111 4137
rect 22695 4097 22707 4100
rect 22649 4091 22707 4097
rect 26053 4097 26065 4131
rect 26099 4128 26111 4131
rect 26234 4128 26240 4140
rect 26099 4100 26240 4128
rect 26099 4097 26111 4100
rect 26053 4091 26111 4097
rect 26234 4088 26240 4100
rect 26292 4128 26298 4140
rect 26694 4128 26700 4140
rect 26292 4100 26700 4128
rect 26292 4088 26298 4100
rect 26694 4088 26700 4100
rect 26752 4088 26758 4140
rect 26804 4128 26832 4236
rect 32398 4224 32404 4276
rect 32456 4264 32462 4276
rect 35710 4264 35716 4276
rect 32456 4236 35716 4264
rect 32456 4224 32462 4236
rect 35710 4224 35716 4236
rect 35768 4224 35774 4276
rect 32766 4196 32772 4208
rect 32727 4168 32772 4196
rect 32766 4156 32772 4168
rect 32824 4156 32830 4208
rect 32858 4156 32864 4208
rect 32916 4196 32922 4208
rect 36170 4196 36176 4208
rect 32916 4168 36176 4196
rect 32916 4156 32922 4168
rect 36170 4156 36176 4168
rect 36228 4156 36234 4208
rect 36630 4156 36636 4208
rect 36688 4196 36694 4208
rect 36725 4199 36783 4205
rect 36725 4196 36737 4199
rect 36688 4168 36737 4196
rect 36688 4156 36694 4168
rect 36725 4165 36737 4168
rect 36771 4165 36783 4199
rect 36725 4159 36783 4165
rect 30374 4128 30380 4140
rect 26804 4100 30380 4128
rect 30374 4088 30380 4100
rect 30432 4088 30438 4140
rect 30926 4088 30932 4140
rect 30984 4128 30990 4140
rect 32490 4128 32496 4140
rect 30984 4100 32496 4128
rect 30984 4088 30990 4100
rect 32490 4088 32496 4100
rect 32548 4088 32554 4140
rect 39853 4131 39911 4137
rect 39853 4128 39865 4131
rect 32600 4100 39865 4128
rect 12437 4063 12495 4069
rect 12268 4032 12388 4060
rect 11977 4023 12035 4029
rect 9766 3952 9772 4004
rect 9824 3992 9830 4004
rect 9861 3995 9919 4001
rect 9861 3992 9873 3995
rect 9824 3964 9873 3992
rect 9824 3952 9830 3964
rect 9861 3961 9873 3964
rect 9907 3961 9919 3995
rect 9861 3955 9919 3961
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 12253 3995 12311 4001
rect 12253 3992 12265 3995
rect 11112 3964 12265 3992
rect 11112 3952 11118 3964
rect 12253 3961 12265 3964
rect 12299 3961 12311 3995
rect 12360 3992 12388 4032
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 13538 4060 13544 4072
rect 12483 4032 13544 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 14642 4020 14648 4072
rect 14700 4060 14706 4072
rect 15197 4063 15255 4069
rect 15197 4060 15209 4063
rect 14700 4032 15209 4060
rect 14700 4020 14706 4032
rect 15197 4029 15209 4032
rect 15243 4060 15255 4063
rect 23106 4060 23112 4072
rect 15243 4032 23112 4060
rect 15243 4029 15255 4032
rect 15197 4023 15255 4029
rect 23106 4020 23112 4032
rect 23164 4020 23170 4072
rect 23934 4020 23940 4072
rect 23992 4060 23998 4072
rect 24305 4063 24363 4069
rect 24305 4060 24317 4063
rect 23992 4032 24317 4060
rect 23992 4020 23998 4032
rect 24305 4029 24317 4032
rect 24351 4060 24363 4063
rect 25130 4060 25136 4072
rect 24351 4032 25136 4060
rect 24351 4029 24363 4032
rect 24305 4023 24363 4029
rect 25130 4020 25136 4032
rect 25188 4020 25194 4072
rect 25498 4020 25504 4072
rect 25556 4060 25562 4072
rect 25866 4060 25872 4072
rect 25556 4032 25872 4060
rect 25556 4020 25562 4032
rect 25866 4020 25872 4032
rect 25924 4060 25930 4072
rect 26513 4063 26571 4069
rect 26513 4060 26525 4063
rect 25924 4032 26525 4060
rect 25924 4020 25930 4032
rect 26513 4029 26525 4032
rect 26559 4029 26571 4063
rect 26513 4023 26571 4029
rect 27982 4020 27988 4072
rect 28040 4060 28046 4072
rect 32600 4060 32628 4100
rect 39853 4097 39865 4100
rect 39899 4128 39911 4131
rect 40034 4128 40040 4140
rect 39899 4100 40040 4128
rect 39899 4097 39911 4100
rect 39853 4091 39911 4097
rect 40034 4088 40040 4100
rect 40092 4128 40098 4140
rect 40957 4131 41015 4137
rect 40957 4128 40969 4131
rect 40092 4100 40969 4128
rect 40092 4088 40098 4100
rect 40957 4097 40969 4100
rect 41003 4097 41015 4131
rect 42702 4128 42708 4140
rect 42663 4100 42708 4128
rect 40957 4091 41015 4097
rect 42702 4088 42708 4100
rect 42760 4128 42766 4140
rect 43901 4131 43959 4137
rect 43901 4128 43913 4131
rect 42760 4100 43913 4128
rect 42760 4088 42766 4100
rect 43901 4097 43913 4100
rect 43947 4128 43959 4131
rect 44545 4131 44603 4137
rect 44545 4128 44557 4131
rect 43947 4100 44557 4128
rect 43947 4097 43959 4100
rect 43901 4091 43959 4097
rect 44545 4097 44557 4100
rect 44591 4128 44603 4131
rect 45189 4131 45247 4137
rect 45189 4128 45201 4131
rect 44591 4100 45201 4128
rect 44591 4097 44603 4100
rect 44545 4091 44603 4097
rect 45189 4097 45201 4100
rect 45235 4128 45247 4131
rect 45554 4128 45560 4140
rect 45235 4100 45560 4128
rect 45235 4097 45247 4100
rect 45189 4091 45247 4097
rect 45554 4088 45560 4100
rect 45612 4128 45618 4140
rect 45833 4131 45891 4137
rect 45833 4128 45845 4131
rect 45612 4100 45845 4128
rect 45612 4088 45618 4100
rect 45833 4097 45845 4100
rect 45879 4128 45891 4131
rect 46477 4131 46535 4137
rect 46477 4128 46489 4131
rect 45879 4100 46489 4128
rect 45879 4097 45891 4100
rect 45833 4091 45891 4097
rect 46477 4097 46489 4100
rect 46523 4097 46535 4131
rect 46477 4091 46535 4097
rect 28040 4032 32628 4060
rect 32692 4032 41414 4060
rect 28040 4020 28046 4032
rect 15102 3992 15108 4004
rect 12360 3964 15108 3992
rect 12253 3955 12311 3961
rect 15102 3952 15108 3964
rect 15160 3952 15166 4004
rect 32692 3992 32720 4032
rect 37458 3992 37464 4004
rect 15212 3964 32720 3992
rect 37419 3964 37464 3992
rect 1670 3924 1676 3936
rect 1631 3896 1676 3924
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 6822 3924 6828 3936
rect 6783 3896 6828 3924
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 7469 3927 7527 3933
rect 7469 3893 7481 3927
rect 7515 3924 7527 3927
rect 7650 3924 7656 3936
rect 7515 3896 7656 3924
rect 7515 3893 7527 3896
rect 7469 3887 7527 3893
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8386 3924 8392 3936
rect 8067 3896 8392 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3924 8539 3927
rect 10042 3924 10048 3936
rect 8527 3896 10048 3924
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 11422 3924 11428 3936
rect 10836 3896 11428 3924
rect 10836 3884 10842 3896
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 12894 3924 12900 3936
rect 12584 3896 12900 3924
rect 12584 3884 12590 3896
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13449 3927 13507 3933
rect 13449 3893 13461 3927
rect 13495 3924 13507 3927
rect 13722 3924 13728 3936
rect 13495 3896 13728 3924
rect 13495 3893 13507 3896
rect 13449 3887 13507 3893
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 14090 3924 14096 3936
rect 14051 3896 14096 3924
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 14645 3927 14703 3933
rect 14645 3893 14657 3927
rect 14691 3924 14703 3927
rect 14826 3924 14832 3936
rect 14691 3896 14832 3924
rect 14691 3893 14703 3896
rect 14645 3887 14703 3893
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 14918 3884 14924 3936
rect 14976 3924 14982 3936
rect 15212 3924 15240 3964
rect 37458 3952 37464 3964
rect 37516 3992 37522 4004
rect 38013 3995 38071 4001
rect 38013 3992 38025 3995
rect 37516 3964 38025 3992
rect 37516 3952 37522 3964
rect 38013 3961 38025 3964
rect 38059 3992 38071 3995
rect 38654 3992 38660 4004
rect 38059 3964 38660 3992
rect 38059 3961 38071 3964
rect 38013 3955 38071 3961
rect 38654 3952 38660 3964
rect 38712 3952 38718 4004
rect 40405 3995 40463 4001
rect 40405 3992 40417 3995
rect 38948 3964 40417 3992
rect 38948 3936 38976 3964
rect 40405 3961 40417 3964
rect 40451 3961 40463 3995
rect 40405 3955 40463 3961
rect 14976 3896 15240 3924
rect 14976 3884 14982 3896
rect 15378 3884 15384 3936
rect 15436 3924 15442 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 15436 3896 15669 3924
rect 15436 3884 15442 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 17773 3927 17831 3933
rect 17773 3893 17785 3927
rect 17819 3924 17831 3927
rect 17862 3924 17868 3936
rect 17819 3896 17868 3924
rect 17819 3893 17831 3896
rect 17773 3887 17831 3893
rect 17862 3884 17868 3896
rect 17920 3884 17926 3936
rect 23201 3927 23259 3933
rect 23201 3893 23213 3927
rect 23247 3924 23259 3927
rect 23474 3924 23480 3936
rect 23247 3896 23480 3924
rect 23247 3893 23259 3896
rect 23201 3887 23259 3893
rect 23474 3884 23480 3896
rect 23532 3884 23538 3936
rect 23750 3924 23756 3936
rect 23711 3896 23756 3924
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 24857 3927 24915 3933
rect 24857 3893 24869 3927
rect 24903 3924 24915 3927
rect 25038 3924 25044 3936
rect 24903 3896 25044 3924
rect 24903 3893 24915 3896
rect 24857 3887 24915 3893
rect 25038 3884 25044 3896
rect 25096 3924 25102 3936
rect 27890 3924 27896 3936
rect 25096 3896 27896 3924
rect 25096 3884 25102 3896
rect 27890 3884 27896 3896
rect 27948 3884 27954 3936
rect 30926 3924 30932 3936
rect 30887 3896 30932 3924
rect 30926 3884 30932 3896
rect 30984 3884 30990 3936
rect 32674 3884 32680 3936
rect 32732 3924 32738 3936
rect 34146 3924 34152 3936
rect 32732 3896 34152 3924
rect 32732 3884 32738 3896
rect 34146 3884 34152 3896
rect 34204 3884 34210 3936
rect 38841 3927 38899 3933
rect 38841 3893 38853 3927
rect 38887 3924 38899 3927
rect 38930 3924 38936 3936
rect 38887 3896 38936 3924
rect 38887 3893 38899 3896
rect 38841 3887 38899 3893
rect 38930 3884 38936 3896
rect 38988 3884 38994 3936
rect 39298 3924 39304 3936
rect 39259 3896 39304 3924
rect 39298 3884 39304 3896
rect 39356 3884 39362 3936
rect 41386 3924 41414 4032
rect 42889 3995 42947 4001
rect 42889 3961 42901 3995
rect 42935 3992 42947 3995
rect 43898 3992 43904 4004
rect 42935 3964 43904 3992
rect 42935 3961 42947 3964
rect 42889 3955 42947 3961
rect 43898 3952 43904 3964
rect 43956 3952 43962 4004
rect 44729 3995 44787 4001
rect 44729 3961 44741 3995
rect 44775 3992 44787 3995
rect 45738 3992 45744 4004
rect 44775 3964 45744 3992
rect 44775 3961 44787 3964
rect 44729 3955 44787 3961
rect 45738 3952 45744 3964
rect 45796 3952 45802 4004
rect 41782 3924 41788 3936
rect 41386 3896 41788 3924
rect 41782 3884 41788 3896
rect 41840 3884 41846 3936
rect 43070 3884 43076 3936
rect 43128 3924 43134 3936
rect 43349 3927 43407 3933
rect 43349 3924 43361 3927
rect 43128 3896 43361 3924
rect 43128 3884 43134 3896
rect 43349 3893 43361 3896
rect 43395 3893 43407 3927
rect 43349 3887 43407 3893
rect 44085 3927 44143 3933
rect 44085 3893 44097 3927
rect 44131 3924 44143 3927
rect 44634 3924 44640 3936
rect 44131 3896 44640 3924
rect 44131 3893 44143 3896
rect 44085 3887 44143 3893
rect 44634 3884 44640 3896
rect 44692 3884 44698 3936
rect 45373 3927 45431 3933
rect 45373 3893 45385 3927
rect 45419 3924 45431 3927
rect 45646 3924 45652 3936
rect 45419 3896 45652 3924
rect 45419 3893 45431 3896
rect 45373 3887 45431 3893
rect 45646 3884 45652 3896
rect 45704 3884 45710 3936
rect 46017 3927 46075 3933
rect 46017 3893 46029 3927
rect 46063 3924 46075 3927
rect 46290 3924 46296 3936
rect 46063 3896 46296 3924
rect 46063 3893 46075 3896
rect 46017 3887 46075 3893
rect 46290 3884 46296 3896
rect 46348 3884 46354 3936
rect 46661 3927 46719 3933
rect 46661 3893 46673 3927
rect 46707 3924 46719 3927
rect 47762 3924 47768 3936
rect 46707 3896 47768 3924
rect 46707 3893 46719 3896
rect 46661 3887 46719 3893
rect 47762 3884 47768 3896
rect 47820 3884 47826 3936
rect 49050 3924 49056 3936
rect 49011 3896 49056 3924
rect 49050 3884 49056 3896
rect 49108 3884 49114 3936
rect 50154 3924 50160 3936
rect 50115 3896 50160 3924
rect 50154 3884 50160 3896
rect 50212 3884 50218 3936
rect 50982 3924 50988 3936
rect 50943 3896 50988 3924
rect 50982 3884 50988 3896
rect 51040 3884 51046 3936
rect 1104 3834 54832 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 54832 3834
rect 1104 3760 54832 3782
rect 7098 3720 7104 3732
rect 7059 3692 7104 3720
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 7929 3723 7987 3729
rect 7929 3689 7941 3723
rect 7975 3720 7987 3723
rect 8294 3720 8300 3732
rect 7975 3692 8300 3720
rect 7975 3689 7987 3692
rect 7929 3683 7987 3689
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 10226 3720 10232 3732
rect 9640 3692 10232 3720
rect 9640 3680 9646 3692
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 10410 3720 10416 3732
rect 10371 3692 10416 3720
rect 10410 3680 10416 3692
rect 10468 3680 10474 3732
rect 12437 3723 12495 3729
rect 12437 3689 12449 3723
rect 12483 3720 12495 3723
rect 12710 3720 12716 3732
rect 12483 3692 12716 3720
rect 12483 3689 12495 3692
rect 12437 3683 12495 3689
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 13354 3680 13360 3732
rect 13412 3720 13418 3732
rect 13541 3723 13599 3729
rect 13541 3720 13553 3723
rect 13412 3692 13553 3720
rect 13412 3680 13418 3692
rect 13541 3689 13553 3692
rect 13587 3689 13599 3723
rect 13541 3683 13599 3689
rect 15838 3680 15844 3732
rect 15896 3720 15902 3732
rect 26786 3720 26792 3732
rect 15896 3692 22094 3720
rect 26747 3692 26792 3720
rect 15896 3680 15902 3692
rect 1872 3624 2774 3652
rect 1872 3525 1900 3624
rect 2746 3584 2774 3624
rect 8478 3612 8484 3664
rect 8536 3652 8542 3664
rect 9769 3655 9827 3661
rect 9769 3652 9781 3655
rect 8536 3624 9781 3652
rect 8536 3612 8542 3624
rect 9769 3621 9781 3624
rect 9815 3621 9827 3655
rect 9769 3615 9827 3621
rect 10318 3612 10324 3664
rect 10376 3652 10382 3664
rect 10870 3652 10876 3664
rect 10376 3624 10456 3652
rect 10376 3612 10382 3624
rect 10134 3584 10140 3596
rect 2746 3556 10140 3584
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10428 3584 10456 3624
rect 10796 3624 10876 3652
rect 10796 3593 10824 3624
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 11609 3655 11667 3661
rect 11609 3621 11621 3655
rect 11655 3652 11667 3655
rect 13078 3652 13084 3664
rect 11655 3624 13084 3652
rect 11655 3621 11667 3624
rect 11609 3615 11667 3621
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 10597 3587 10655 3593
rect 10597 3584 10609 3587
rect 10428 3556 10609 3584
rect 10597 3553 10609 3556
rect 10643 3553 10655 3587
rect 10597 3547 10655 3553
rect 10781 3587 10839 3593
rect 10781 3553 10793 3587
rect 10827 3553 10839 3587
rect 14458 3584 14464 3596
rect 14419 3556 14464 3584
rect 10781 3547 10839 3553
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 14642 3584 14648 3596
rect 14603 3556 14648 3584
rect 14642 3544 14648 3556
rect 14700 3544 14706 3596
rect 14737 3587 14795 3593
rect 14737 3553 14749 3587
rect 14783 3584 14795 3587
rect 19058 3584 19064 3596
rect 14783 3556 19064 3584
rect 14783 3553 14795 3556
rect 14737 3547 14795 3553
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 22066 3584 22094 3692
rect 26786 3680 26792 3692
rect 26844 3680 26850 3732
rect 27433 3723 27491 3729
rect 27433 3689 27445 3723
rect 27479 3720 27491 3723
rect 27798 3720 27804 3732
rect 27479 3692 27804 3720
rect 27479 3689 27491 3692
rect 27433 3683 27491 3689
rect 27798 3680 27804 3692
rect 27856 3680 27862 3732
rect 27890 3680 27896 3732
rect 27948 3720 27954 3732
rect 27985 3723 28043 3729
rect 27985 3720 27997 3723
rect 27948 3692 27997 3720
rect 27948 3680 27954 3692
rect 27985 3689 27997 3692
rect 28031 3720 28043 3723
rect 28074 3720 28080 3732
rect 28031 3692 28080 3720
rect 28031 3689 28043 3692
rect 27985 3683 28043 3689
rect 28074 3680 28080 3692
rect 28132 3680 28138 3732
rect 28626 3720 28632 3732
rect 28587 3692 28632 3720
rect 28626 3680 28632 3692
rect 28684 3680 28690 3732
rect 31297 3723 31355 3729
rect 31297 3689 31309 3723
rect 31343 3720 31355 3723
rect 31754 3720 31760 3732
rect 31343 3692 31760 3720
rect 31343 3689 31355 3692
rect 31297 3683 31355 3689
rect 31754 3680 31760 3692
rect 31812 3720 31818 3732
rect 32398 3720 32404 3732
rect 31812 3692 32404 3720
rect 31812 3680 31818 3692
rect 32398 3680 32404 3692
rect 32456 3680 32462 3732
rect 32769 3723 32827 3729
rect 32769 3689 32781 3723
rect 32815 3720 32827 3723
rect 32858 3720 32864 3732
rect 32815 3692 32864 3720
rect 32815 3689 32827 3692
rect 32769 3683 32827 3689
rect 32858 3680 32864 3692
rect 32916 3680 32922 3732
rect 33318 3720 33324 3732
rect 33279 3692 33324 3720
rect 33318 3680 33324 3692
rect 33376 3680 33382 3732
rect 33778 3680 33784 3732
rect 33836 3720 33842 3732
rect 33873 3723 33931 3729
rect 33873 3720 33885 3723
rect 33836 3692 33885 3720
rect 33836 3680 33842 3692
rect 33873 3689 33885 3692
rect 33919 3720 33931 3723
rect 33962 3720 33968 3732
rect 33919 3692 33968 3720
rect 33919 3689 33931 3692
rect 33873 3683 33931 3689
rect 33962 3680 33968 3692
rect 34020 3680 34026 3732
rect 34514 3680 34520 3732
rect 34572 3720 34578 3732
rect 34885 3723 34943 3729
rect 34885 3720 34897 3723
rect 34572 3692 34897 3720
rect 34572 3680 34578 3692
rect 34885 3689 34897 3692
rect 34931 3689 34943 3723
rect 34885 3683 34943 3689
rect 41417 3723 41475 3729
rect 41417 3689 41429 3723
rect 41463 3720 41475 3723
rect 41690 3720 41696 3732
rect 41463 3692 41696 3720
rect 41463 3689 41475 3692
rect 41417 3683 41475 3689
rect 41690 3680 41696 3692
rect 41748 3680 41754 3732
rect 42702 3680 42708 3732
rect 42760 3720 42766 3732
rect 42981 3723 43039 3729
rect 42981 3720 42993 3723
rect 42760 3692 42993 3720
rect 42760 3680 42766 3692
rect 42981 3689 42993 3692
rect 43027 3689 43039 3723
rect 51166 3720 51172 3732
rect 51127 3692 51172 3720
rect 42981 3683 43039 3689
rect 23106 3652 23112 3664
rect 23065 3624 23112 3652
rect 23106 3612 23112 3624
rect 23164 3661 23170 3664
rect 23164 3655 23213 3661
rect 23164 3621 23167 3655
rect 23201 3652 23213 3655
rect 30282 3652 30288 3664
rect 23201 3624 30288 3652
rect 23201 3621 23213 3624
rect 23164 3615 23213 3621
rect 23164 3612 23170 3615
rect 30282 3612 30288 3624
rect 30340 3612 30346 3664
rect 30374 3612 30380 3664
rect 30432 3652 30438 3664
rect 30561 3655 30619 3661
rect 30561 3652 30573 3655
rect 30432 3624 30573 3652
rect 30432 3612 30438 3624
rect 30561 3621 30573 3624
rect 30607 3652 30619 3655
rect 31662 3652 31668 3664
rect 30607 3624 31668 3652
rect 30607 3621 30619 3624
rect 30561 3615 30619 3621
rect 31662 3612 31668 3624
rect 31720 3612 31726 3664
rect 31846 3612 31852 3664
rect 31904 3652 31910 3664
rect 35342 3652 35348 3664
rect 31904 3624 35348 3652
rect 31904 3612 31910 3624
rect 35342 3612 35348 3624
rect 35400 3612 35406 3664
rect 40865 3655 40923 3661
rect 40865 3621 40877 3655
rect 40911 3652 40923 3655
rect 41506 3652 41512 3664
rect 40911 3624 41512 3652
rect 40911 3621 40923 3624
rect 40865 3615 40923 3621
rect 41506 3612 41512 3624
rect 41564 3612 41570 3664
rect 42996 3652 43024 3683
rect 51166 3680 51172 3692
rect 51224 3680 51230 3732
rect 42996 3624 43668 3652
rect 22066 3556 43116 3584
rect 43088 3528 43116 3556
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3485 1915 3519
rect 1857 3479 1915 3485
rect 6822 3476 6828 3528
rect 6880 3516 6886 3528
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 6880 3488 6929 3516
rect 6880 3476 6886 3488
rect 6917 3485 6929 3488
rect 6963 3485 6975 3519
rect 7742 3516 7748 3528
rect 7703 3488 7748 3516
rect 6917 3479 6975 3485
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 8386 3516 8392 3528
rect 8347 3488 8392 3516
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 10678 3519 10736 3525
rect 8588 3488 10548 3516
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 6457 3383 6515 3389
rect 6457 3349 6469 3383
rect 6503 3380 6515 3383
rect 7006 3380 7012 3392
rect 6503 3352 7012 3380
rect 6503 3349 6515 3352
rect 6457 3343 6515 3349
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 8588 3389 8616 3488
rect 9493 3451 9551 3457
rect 9493 3417 9505 3451
rect 9539 3448 9551 3451
rect 9582 3448 9588 3460
rect 9539 3420 9588 3448
rect 9539 3417 9551 3420
rect 9493 3411 9551 3417
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 8573 3383 8631 3389
rect 8573 3349 8585 3383
rect 8619 3349 8631 3383
rect 8573 3343 8631 3349
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 9674 3380 9680 3392
rect 8996 3352 9680 3380
rect 8996 3340 9002 3352
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 9950 3380 9956 3392
rect 9911 3352 9956 3380
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 10520 3380 10548 3488
rect 10678 3485 10690 3519
rect 10724 3504 10736 3519
rect 10678 3479 10692 3485
rect 10686 3452 10692 3479
rect 10744 3452 10750 3504
rect 10870 3476 10876 3528
rect 10928 3516 10934 3528
rect 11422 3516 11428 3528
rect 10928 3488 10973 3516
rect 11383 3488 11428 3516
rect 10928 3476 10934 3488
rect 11422 3476 11428 3488
rect 11480 3476 11486 3528
rect 11606 3476 11612 3528
rect 11664 3516 11670 3528
rect 12342 3516 12348 3528
rect 11664 3488 12348 3516
rect 11664 3476 11670 3488
rect 12342 3476 12348 3488
rect 12400 3516 12406 3528
rect 12621 3519 12679 3525
rect 12621 3516 12633 3519
rect 12400 3488 12633 3516
rect 12400 3476 12406 3488
rect 12621 3485 12633 3488
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 13446 3476 13452 3528
rect 13504 3516 13510 3528
rect 13722 3516 13728 3528
rect 13504 3488 13728 3516
rect 13504 3476 13510 3488
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 14829 3519 14887 3525
rect 14829 3516 14841 3519
rect 14608 3488 14841 3516
rect 14608 3476 14614 3488
rect 14829 3485 14841 3488
rect 14875 3485 14887 3519
rect 14829 3479 14887 3485
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 19797 3519 19855 3525
rect 14976 3488 15021 3516
rect 14976 3476 14982 3488
rect 19797 3485 19809 3519
rect 19843 3516 19855 3519
rect 19978 3516 19984 3528
rect 19843 3488 19984 3516
rect 19843 3485 19855 3488
rect 19797 3479 19855 3485
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 21637 3519 21695 3525
rect 21637 3485 21649 3519
rect 21683 3516 21695 3519
rect 22465 3519 22523 3525
rect 21683 3488 22324 3516
rect 21683 3485 21695 3488
rect 21637 3479 21695 3485
rect 22094 3408 22100 3460
rect 22152 3448 22158 3460
rect 22296 3457 22324 3488
rect 22465 3485 22477 3519
rect 22511 3516 22523 3519
rect 22925 3519 22983 3525
rect 22925 3516 22937 3519
rect 22511 3488 22937 3516
rect 22511 3485 22523 3488
rect 22465 3479 22523 3485
rect 22925 3485 22937 3488
rect 22971 3485 22983 3519
rect 24946 3516 24952 3528
rect 22925 3479 22983 3485
rect 23400 3488 24952 3516
rect 22281 3451 22339 3457
rect 22152 3420 22197 3448
rect 22152 3408 22158 3420
rect 22281 3417 22293 3451
rect 22327 3448 22339 3451
rect 22738 3448 22744 3460
rect 22327 3420 22744 3448
rect 22327 3417 22339 3420
rect 22281 3411 22339 3417
rect 22738 3408 22744 3420
rect 22796 3408 22802 3460
rect 14642 3380 14648 3392
rect 10520 3352 14648 3380
rect 14642 3340 14648 3352
rect 14700 3340 14706 3392
rect 15933 3383 15991 3389
rect 15933 3349 15945 3383
rect 15979 3380 15991 3383
rect 16114 3380 16120 3392
rect 15979 3352 16120 3380
rect 15979 3349 15991 3352
rect 15933 3343 15991 3349
rect 16114 3340 16120 3352
rect 16172 3340 16178 3392
rect 16390 3380 16396 3392
rect 16351 3352 16396 3380
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 17497 3383 17555 3389
rect 17497 3349 17509 3383
rect 17543 3380 17555 3383
rect 17770 3380 17776 3392
rect 17543 3352 17776 3380
rect 17543 3349 17555 3352
rect 17497 3343 17555 3349
rect 17770 3340 17776 3352
rect 17828 3340 17834 3392
rect 18233 3383 18291 3389
rect 18233 3349 18245 3383
rect 18279 3380 18291 3383
rect 18506 3380 18512 3392
rect 18279 3352 18512 3380
rect 18279 3349 18291 3352
rect 18233 3343 18291 3349
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 18598 3340 18604 3392
rect 18656 3380 18662 3392
rect 23400 3380 23428 3488
rect 24946 3476 24952 3488
rect 25004 3476 25010 3528
rect 25225 3519 25283 3525
rect 25225 3485 25237 3519
rect 25271 3516 25283 3519
rect 25314 3516 25320 3528
rect 25271 3488 25320 3516
rect 25271 3485 25283 3488
rect 25225 3479 25283 3485
rect 25314 3476 25320 3488
rect 25372 3476 25378 3528
rect 34054 3516 34060 3528
rect 25516 3488 34060 3516
rect 23474 3408 23480 3460
rect 23532 3448 23538 3460
rect 25516 3448 25544 3488
rect 34054 3476 34060 3488
rect 34112 3476 34118 3528
rect 37277 3519 37335 3525
rect 37277 3485 37289 3519
rect 37323 3516 37335 3519
rect 37458 3516 37464 3528
rect 37323 3488 37464 3516
rect 37323 3485 37335 3488
rect 37277 3479 37335 3485
rect 37458 3476 37464 3488
rect 37516 3516 37522 3528
rect 37921 3519 37979 3525
rect 37921 3516 37933 3519
rect 37516 3488 37933 3516
rect 37516 3476 37522 3488
rect 37921 3485 37933 3488
rect 37967 3485 37979 3519
rect 38930 3516 38936 3528
rect 38891 3488 38936 3516
rect 37921 3479 37979 3485
rect 38930 3476 38936 3488
rect 38988 3476 38994 3528
rect 40034 3516 40040 3528
rect 39995 3488 40040 3516
rect 40034 3476 40040 3488
rect 40092 3476 40098 3528
rect 40681 3519 40739 3525
rect 40681 3485 40693 3519
rect 40727 3516 40739 3519
rect 41690 3516 41696 3528
rect 40727 3488 41696 3516
rect 40727 3485 40739 3488
rect 40681 3479 40739 3485
rect 41690 3476 41696 3488
rect 41748 3476 41754 3528
rect 41782 3476 41788 3528
rect 41840 3516 41846 3528
rect 41877 3519 41935 3525
rect 41877 3516 41889 3519
rect 41840 3488 41889 3516
rect 41840 3476 41846 3488
rect 41877 3485 41889 3488
rect 41923 3485 41935 3519
rect 43070 3516 43076 3528
rect 43031 3488 43076 3516
rect 41877 3479 41935 3485
rect 23532 3420 25544 3448
rect 26237 3451 26295 3457
rect 23532 3408 23538 3420
rect 26237 3417 26249 3451
rect 26283 3448 26295 3451
rect 26326 3448 26332 3460
rect 26283 3420 26332 3448
rect 26283 3417 26295 3420
rect 26237 3411 26295 3417
rect 26326 3408 26332 3420
rect 26384 3448 26390 3460
rect 27706 3448 27712 3460
rect 26384 3420 27712 3448
rect 26384 3408 26390 3420
rect 27706 3408 27712 3420
rect 27764 3408 27770 3460
rect 28994 3408 29000 3460
rect 29052 3448 29058 3460
rect 39298 3448 39304 3460
rect 29052 3420 39304 3448
rect 29052 3408 29058 3420
rect 39298 3408 39304 3420
rect 39356 3408 39362 3460
rect 41892 3448 41920 3479
rect 43070 3476 43076 3488
rect 43128 3476 43134 3528
rect 43640 3525 43668 3624
rect 43625 3519 43683 3525
rect 43625 3485 43637 3519
rect 43671 3516 43683 3519
rect 44269 3519 44327 3525
rect 44269 3516 44281 3519
rect 43671 3488 44281 3516
rect 43671 3485 43683 3488
rect 43625 3479 43683 3485
rect 44269 3485 44281 3488
rect 44315 3516 44327 3519
rect 45189 3519 45247 3525
rect 45189 3516 45201 3519
rect 44315 3488 45201 3516
rect 44315 3485 44327 3488
rect 44269 3479 44327 3485
rect 45189 3485 45201 3488
rect 45235 3485 45247 3519
rect 45922 3516 45928 3528
rect 45883 3488 45928 3516
rect 45189 3479 45247 3485
rect 45922 3476 45928 3488
rect 45980 3476 45986 3528
rect 46934 3516 46940 3528
rect 46895 3488 46940 3516
rect 46934 3476 46940 3488
rect 46992 3516 46998 3528
rect 47397 3519 47455 3525
rect 47397 3516 47409 3519
rect 46992 3488 47409 3516
rect 46992 3476 46998 3488
rect 47397 3485 47409 3488
rect 47443 3485 47455 3519
rect 47397 3479 47455 3485
rect 41892 3420 43668 3448
rect 43640 3392 43668 3420
rect 50982 3408 50988 3460
rect 51040 3448 51046 3460
rect 51261 3451 51319 3457
rect 51261 3448 51273 3451
rect 51040 3420 51273 3448
rect 51040 3408 51046 3420
rect 51261 3417 51273 3420
rect 51307 3417 51319 3451
rect 51261 3411 51319 3417
rect 18656 3352 23428 3380
rect 18656 3340 18662 3352
rect 24854 3340 24860 3392
rect 24912 3380 24918 3392
rect 25041 3383 25099 3389
rect 25041 3380 25053 3383
rect 24912 3352 25053 3380
rect 24912 3340 24918 3352
rect 25041 3349 25053 3352
rect 25087 3349 25099 3383
rect 25041 3343 25099 3349
rect 35894 3340 35900 3392
rect 35952 3380 35958 3392
rect 35989 3383 36047 3389
rect 35989 3380 36001 3383
rect 35952 3352 36001 3380
rect 35952 3340 35958 3352
rect 35989 3349 36001 3352
rect 36035 3349 36047 3383
rect 35989 3343 36047 3349
rect 36262 3340 36268 3392
rect 36320 3380 36326 3392
rect 36633 3383 36691 3389
rect 36633 3380 36645 3383
rect 36320 3352 36645 3380
rect 36320 3340 36326 3352
rect 36633 3349 36645 3352
rect 36679 3349 36691 3383
rect 36633 3343 36691 3349
rect 37461 3383 37519 3389
rect 37461 3349 37473 3383
rect 37507 3380 37519 3383
rect 37918 3380 37924 3392
rect 37507 3352 37924 3380
rect 37507 3349 37519 3352
rect 37461 3343 37519 3349
rect 37918 3340 37924 3352
rect 37976 3340 37982 3392
rect 38102 3380 38108 3392
rect 38063 3352 38108 3380
rect 38102 3340 38108 3352
rect 38160 3340 38166 3392
rect 39117 3383 39175 3389
rect 39117 3349 39129 3383
rect 39163 3380 39175 3383
rect 40034 3380 40040 3392
rect 39163 3352 40040 3380
rect 39163 3349 39175 3352
rect 39117 3343 39175 3349
rect 40034 3340 40040 3352
rect 40092 3340 40098 3392
rect 40221 3383 40279 3389
rect 40221 3349 40233 3383
rect 40267 3380 40279 3383
rect 40770 3380 40776 3392
rect 40267 3352 40776 3380
rect 40267 3349 40279 3352
rect 40221 3343 40279 3349
rect 40770 3340 40776 3352
rect 40828 3340 40834 3392
rect 42061 3383 42119 3389
rect 42061 3349 42073 3383
rect 42107 3380 42119 3383
rect 42794 3380 42800 3392
rect 42107 3352 42800 3380
rect 42107 3349 42119 3352
rect 42061 3343 42119 3349
rect 42794 3340 42800 3352
rect 42852 3340 42858 3392
rect 43622 3340 43628 3392
rect 43680 3340 43686 3392
rect 43809 3383 43867 3389
rect 43809 3349 43821 3383
rect 43855 3380 43867 3383
rect 44082 3380 44088 3392
rect 43855 3352 44088 3380
rect 43855 3349 43867 3352
rect 43809 3343 43867 3349
rect 44082 3340 44088 3352
rect 44140 3340 44146 3392
rect 44453 3383 44511 3389
rect 44453 3349 44465 3383
rect 44499 3380 44511 3383
rect 45186 3380 45192 3392
rect 44499 3352 45192 3380
rect 44499 3349 44511 3352
rect 44453 3343 44511 3349
rect 45186 3340 45192 3352
rect 45244 3340 45250 3392
rect 45373 3383 45431 3389
rect 45373 3349 45385 3383
rect 45419 3380 45431 3383
rect 45554 3380 45560 3392
rect 45419 3352 45560 3380
rect 45419 3349 45431 3352
rect 45373 3343 45431 3349
rect 45554 3340 45560 3352
rect 45612 3340 45618 3392
rect 45830 3340 45836 3392
rect 45888 3380 45894 3392
rect 46109 3383 46167 3389
rect 46109 3380 46121 3383
rect 45888 3352 46121 3380
rect 45888 3340 45894 3352
rect 46109 3349 46121 3352
rect 46155 3349 46167 3383
rect 46109 3343 46167 3349
rect 46566 3340 46572 3392
rect 46624 3380 46630 3392
rect 46753 3383 46811 3389
rect 46753 3380 46765 3383
rect 46624 3352 46765 3380
rect 46624 3340 46630 3352
rect 46753 3349 46765 3352
rect 46799 3349 46811 3383
rect 46753 3343 46811 3349
rect 47670 3340 47676 3392
rect 47728 3380 47734 3392
rect 48317 3383 48375 3389
rect 48317 3380 48329 3383
rect 47728 3352 48329 3380
rect 47728 3340 47734 3352
rect 48317 3349 48329 3352
rect 48363 3349 48375 3383
rect 48866 3380 48872 3392
rect 48827 3352 48872 3380
rect 48317 3343 48375 3349
rect 48866 3340 48872 3352
rect 48924 3340 48930 3392
rect 49418 3380 49424 3392
rect 49379 3352 49424 3380
rect 49418 3340 49424 3352
rect 49476 3340 49482 3392
rect 49602 3340 49608 3392
rect 49660 3380 49666 3392
rect 50341 3383 50399 3389
rect 50341 3380 50353 3383
rect 49660 3352 50353 3380
rect 49660 3340 49666 3352
rect 50341 3349 50353 3352
rect 50387 3349 50399 3383
rect 51810 3380 51816 3392
rect 51771 3352 51816 3380
rect 50341 3343 50399 3349
rect 51810 3340 51816 3352
rect 51868 3340 51874 3392
rect 51994 3340 52000 3392
rect 52052 3380 52058 3392
rect 52457 3383 52515 3389
rect 52457 3380 52469 3383
rect 52052 3352 52469 3380
rect 52052 3340 52058 3352
rect 52457 3349 52469 3352
rect 52503 3349 52515 3383
rect 52457 3343 52515 3349
rect 1104 3290 54832 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 54832 3290
rect 1104 3216 54832 3238
rect 7650 3136 7656 3188
rect 7708 3176 7714 3188
rect 8294 3176 8300 3188
rect 7708 3148 8300 3176
rect 7708 3136 7714 3148
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 8478 3176 8484 3188
rect 8439 3148 8484 3176
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 9398 3176 9404 3188
rect 8812 3148 9404 3176
rect 8812 3136 8818 3148
rect 9398 3136 9404 3148
rect 9456 3136 9462 3188
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10689 3179 10747 3185
rect 10689 3145 10701 3179
rect 10735 3176 10747 3179
rect 10962 3176 10968 3188
rect 10735 3148 10968 3176
rect 10735 3145 10747 3148
rect 10689 3139 10747 3145
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 11977 3179 12035 3185
rect 11977 3145 11989 3179
rect 12023 3176 12035 3179
rect 12894 3176 12900 3188
rect 12023 3148 12900 3176
rect 12023 3145 12035 3148
rect 11977 3139 12035 3145
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 13265 3179 13323 3185
rect 13265 3145 13277 3179
rect 13311 3176 13323 3179
rect 13630 3176 13636 3188
rect 13311 3148 13636 3176
rect 13311 3145 13323 3148
rect 13265 3139 13323 3145
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 13909 3179 13967 3185
rect 13909 3145 13921 3179
rect 13955 3176 13967 3179
rect 14274 3176 14280 3188
rect 13955 3148 14280 3176
rect 13955 3145 13967 3148
rect 13909 3139 13967 3145
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 14829 3179 14887 3185
rect 14829 3145 14841 3179
rect 14875 3176 14887 3179
rect 14918 3176 14924 3188
rect 14875 3148 14924 3176
rect 14875 3145 14887 3148
rect 14829 3139 14887 3145
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 15562 3176 15568 3188
rect 15523 3148 15568 3176
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 16301 3179 16359 3185
rect 16301 3145 16313 3179
rect 16347 3176 16359 3179
rect 16574 3176 16580 3188
rect 16347 3148 16580 3176
rect 16347 3145 16359 3148
rect 16301 3139 16359 3145
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 16758 3136 16764 3188
rect 16816 3176 16822 3188
rect 16945 3179 17003 3185
rect 16945 3176 16957 3179
rect 16816 3148 16957 3176
rect 16816 3136 16822 3148
rect 16945 3145 16957 3148
rect 16991 3145 17003 3179
rect 17586 3176 17592 3188
rect 17547 3148 17592 3176
rect 16945 3139 17003 3145
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18325 3179 18383 3185
rect 18325 3176 18337 3179
rect 18012 3148 18337 3176
rect 18012 3136 18018 3148
rect 18325 3145 18337 3148
rect 18371 3145 18383 3179
rect 18325 3139 18383 3145
rect 24394 3136 24400 3188
rect 24452 3176 24458 3188
rect 24452 3148 25544 3176
rect 24452 3136 24458 3148
rect 5997 3111 6055 3117
rect 5997 3077 6009 3111
rect 6043 3108 6055 3111
rect 6043 3080 8340 3108
rect 6043 3077 6055 3080
rect 5997 3071 6055 3077
rect 7006 3040 7012 3052
rect 6967 3012 7012 3040
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 7650 3040 7656 3052
rect 7611 3012 7656 3040
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 8312 3049 8340 3080
rect 8386 3068 8392 3120
rect 8444 3108 8450 3120
rect 9030 3108 9036 3120
rect 8444 3080 9036 3108
rect 8444 3068 8450 3080
rect 9030 3068 9036 3080
rect 9088 3068 9094 3120
rect 25406 3108 25412 3120
rect 9508 3080 25412 3108
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 8754 3040 8760 3052
rect 8343 3012 8760 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 8938 3040 8944 3052
rect 8899 3012 8944 3040
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 9508 2972 9536 3080
rect 25406 3068 25412 3080
rect 25464 3068 25470 3120
rect 25516 3108 25544 3148
rect 28810 3136 28816 3188
rect 28868 3176 28874 3188
rect 28997 3179 29055 3185
rect 28997 3176 29009 3179
rect 28868 3148 29009 3176
rect 28868 3136 28874 3148
rect 28997 3145 29009 3148
rect 29043 3145 29055 3179
rect 29638 3176 29644 3188
rect 29599 3148 29644 3176
rect 28997 3139 29055 3145
rect 29638 3136 29644 3148
rect 29696 3136 29702 3188
rect 29914 3136 29920 3188
rect 29972 3176 29978 3188
rect 31573 3179 31631 3185
rect 31573 3176 31585 3179
rect 29972 3148 31585 3176
rect 29972 3136 29978 3148
rect 31573 3145 31585 3148
rect 31619 3145 31631 3179
rect 38930 3176 38936 3188
rect 31573 3139 31631 3145
rect 31726 3148 38936 3176
rect 31726 3108 31754 3148
rect 38930 3136 38936 3148
rect 38988 3136 38994 3188
rect 40126 3136 40132 3188
rect 40184 3176 40190 3188
rect 47854 3176 47860 3188
rect 40184 3148 41092 3176
rect 47815 3148 47860 3176
rect 40184 3136 40190 3148
rect 25516 3080 31754 3108
rect 34422 3068 34428 3120
rect 34480 3108 34486 3120
rect 35069 3111 35127 3117
rect 35069 3108 35081 3111
rect 34480 3080 35081 3108
rect 34480 3068 34486 3080
rect 35069 3077 35081 3080
rect 35115 3077 35127 3111
rect 38948 3108 38976 3136
rect 38948 3080 40356 3108
rect 35069 3071 35127 3077
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3040 9643 3043
rect 9858 3040 9864 3052
rect 9631 3012 9864 3040
rect 9631 3009 9643 3012
rect 9585 3003 9643 3009
rect 9858 3000 9864 3012
rect 9916 3040 9922 3052
rect 10134 3040 10140 3052
rect 9916 3012 10140 3040
rect 9916 3000 9922 3012
rect 10134 3000 10140 3012
rect 10192 3000 10198 3052
rect 10226 3000 10232 3052
rect 10284 3040 10290 3052
rect 11606 3040 11612 3052
rect 10284 3012 11612 3040
rect 10284 3000 10290 3012
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 11790 3040 11796 3052
rect 11751 3012 11796 3040
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3040 12495 3043
rect 12483 3012 12517 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 7208 2944 9536 2972
rect 7208 2913 7236 2944
rect 10318 2932 10324 2984
rect 10376 2972 10382 2984
rect 12452 2972 12480 3003
rect 12894 3000 12900 3052
rect 12952 3040 12958 3052
rect 13081 3043 13139 3049
rect 13081 3040 13093 3043
rect 12952 3012 13093 3040
rect 12952 3000 12958 3012
rect 13081 3009 13093 3012
rect 13127 3040 13139 3043
rect 13630 3040 13636 3052
rect 13127 3012 13636 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3040 13783 3043
rect 14090 3040 14096 3052
rect 13771 3012 14096 3040
rect 13771 3009 13783 3012
rect 13725 3003 13783 3009
rect 14090 3000 14096 3012
rect 14148 3040 14154 3052
rect 14550 3040 14556 3052
rect 14148 3012 14556 3040
rect 14148 3000 14154 3012
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 15378 3040 15384 3052
rect 15339 3012 15384 3040
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3040 16175 3043
rect 16390 3040 16396 3052
rect 16163 3012 16396 3040
rect 16163 3009 16175 3012
rect 16117 3003 16175 3009
rect 16390 3000 16396 3012
rect 16448 3000 16454 3052
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17494 3000 17500 3052
rect 17552 3040 17558 3052
rect 17770 3040 17776 3052
rect 17552 3012 17776 3040
rect 17552 3000 17558 3012
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 18230 3000 18236 3052
rect 18288 3040 18294 3052
rect 18506 3040 18512 3052
rect 18288 3012 18512 3040
rect 18288 3000 18294 3012
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 23658 3040 23664 3052
rect 23619 3012 23664 3040
rect 23658 3000 23664 3012
rect 23716 3000 23722 3052
rect 23750 3000 23756 3052
rect 23808 3040 23814 3052
rect 24397 3043 24455 3049
rect 24397 3040 24409 3043
rect 23808 3012 24409 3040
rect 23808 3000 23814 3012
rect 24397 3009 24409 3012
rect 24443 3009 24455 3043
rect 24397 3003 24455 3009
rect 24857 3043 24915 3049
rect 24857 3009 24869 3043
rect 24903 3040 24915 3043
rect 25038 3040 25044 3052
rect 24903 3012 25044 3040
rect 24903 3009 24915 3012
rect 24857 3003 24915 3009
rect 12710 2972 12716 2984
rect 10376 2944 12716 2972
rect 10376 2932 10382 2944
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 14369 2975 14427 2981
rect 14369 2941 14381 2975
rect 14415 2972 14427 2975
rect 15194 2972 15200 2984
rect 14415 2944 15200 2972
rect 14415 2941 14427 2944
rect 14369 2935 14427 2941
rect 15194 2932 15200 2944
rect 15252 2932 15258 2984
rect 24118 2972 24124 2984
rect 22066 2944 24124 2972
rect 7193 2907 7251 2913
rect 7193 2873 7205 2907
rect 7239 2873 7251 2907
rect 7193 2867 7251 2873
rect 7837 2907 7895 2913
rect 7837 2873 7849 2907
rect 7883 2904 7895 2907
rect 9125 2907 9183 2913
rect 7883 2876 9076 2904
rect 7883 2873 7895 2876
rect 7837 2867 7895 2873
rect 9048 2836 9076 2876
rect 9125 2873 9137 2907
rect 9171 2904 9183 2907
rect 10505 2907 10563 2913
rect 10505 2904 10517 2907
rect 9171 2876 10517 2904
rect 9171 2873 9183 2876
rect 9125 2867 9183 2873
rect 10505 2873 10517 2876
rect 10551 2873 10563 2907
rect 12621 2907 12679 2913
rect 10505 2867 10563 2873
rect 10612 2876 12434 2904
rect 10612 2836 10640 2876
rect 9048 2808 10640 2836
rect 12406 2836 12434 2876
rect 12621 2873 12633 2907
rect 12667 2904 12679 2907
rect 12986 2904 12992 2916
rect 12667 2876 12992 2904
rect 12667 2873 12679 2876
rect 12621 2867 12679 2873
rect 12986 2864 12992 2876
rect 13044 2864 13050 2916
rect 14642 2904 14648 2916
rect 14603 2876 14648 2904
rect 14642 2864 14648 2876
rect 14700 2864 14706 2916
rect 22066 2904 22094 2944
rect 24118 2932 24124 2944
rect 24176 2932 24182 2984
rect 24412 2972 24440 3003
rect 25038 3000 25044 3012
rect 25096 3000 25102 3052
rect 25593 3043 25651 3049
rect 25593 3009 25605 3043
rect 25639 3040 25651 3043
rect 26234 3040 26240 3052
rect 25639 3012 26240 3040
rect 25639 3009 25651 3012
rect 25593 3003 25651 3009
rect 26234 3000 26240 3012
rect 26292 3000 26298 3052
rect 26329 3043 26387 3049
rect 26329 3009 26341 3043
rect 26375 3040 26387 3043
rect 26786 3040 26792 3052
rect 26375 3012 26792 3040
rect 26375 3009 26387 3012
rect 26329 3003 26387 3009
rect 26786 3000 26792 3012
rect 26844 3000 26850 3052
rect 27798 3040 27804 3052
rect 27759 3012 27804 3040
rect 27798 3000 27804 3012
rect 27856 3000 27862 3052
rect 28537 3043 28595 3049
rect 28537 3009 28549 3043
rect 28583 3040 28595 3043
rect 28810 3040 28816 3052
rect 28583 3012 28816 3040
rect 28583 3009 28595 3012
rect 28537 3003 28595 3009
rect 28810 3000 28816 3012
rect 28868 3000 28874 3052
rect 30374 3040 30380 3052
rect 30335 3012 30380 3040
rect 30374 3000 30380 3012
rect 30432 3000 30438 3052
rect 31113 3043 31171 3049
rect 31113 3009 31125 3043
rect 31159 3040 31171 3043
rect 31754 3040 31760 3052
rect 31159 3012 31760 3040
rect 31159 3009 31171 3012
rect 31113 3003 31171 3009
rect 31754 3000 31760 3012
rect 31812 3000 31818 3052
rect 32585 3043 32643 3049
rect 32585 3009 32597 3043
rect 32631 3040 32643 3043
rect 32858 3040 32864 3052
rect 32631 3012 32864 3040
rect 32631 3009 32643 3012
rect 32585 3003 32643 3009
rect 32858 3000 32864 3012
rect 32916 3000 32922 3052
rect 33318 3040 33324 3052
rect 33279 3012 33324 3040
rect 33318 3000 33324 3012
rect 33376 3000 33382 3052
rect 35526 3000 35532 3052
rect 35584 3040 35590 3052
rect 36357 3043 36415 3049
rect 36357 3040 36369 3043
rect 35584 3012 36369 3040
rect 35584 3000 35590 3012
rect 36357 3009 36369 3012
rect 36403 3009 36415 3043
rect 38102 3040 38108 3052
rect 38063 3012 38108 3040
rect 36357 3003 36415 3009
rect 38102 3000 38108 3012
rect 38160 3000 38166 3052
rect 38378 3000 38384 3052
rect 38436 3040 38442 3052
rect 38565 3043 38623 3049
rect 38565 3040 38577 3043
rect 38436 3012 38577 3040
rect 38436 3000 38442 3012
rect 38565 3009 38577 3012
rect 38611 3009 38623 3043
rect 39298 3040 39304 3052
rect 39259 3012 39304 3040
rect 38565 3003 38623 3009
rect 39298 3000 39304 3012
rect 39356 3000 39362 3052
rect 40328 3049 40356 3080
rect 41064 3049 41092 3148
rect 47854 3136 47860 3148
rect 47912 3136 47918 3188
rect 48590 3176 48596 3188
rect 48551 3148 48596 3176
rect 48590 3136 48596 3148
rect 48648 3136 48654 3188
rect 49326 3176 49332 3188
rect 49287 3148 49332 3176
rect 49326 3136 49332 3148
rect 49384 3136 49390 3188
rect 50062 3176 50068 3188
rect 50023 3148 50068 3176
rect 50062 3136 50068 3148
rect 50120 3136 50126 3188
rect 50798 3176 50804 3188
rect 50759 3148 50804 3176
rect 50798 3136 50804 3148
rect 50856 3136 50862 3188
rect 51534 3176 51540 3188
rect 51495 3148 51540 3176
rect 51534 3136 51540 3148
rect 51592 3136 51598 3188
rect 47670 3068 47676 3120
rect 47728 3108 47734 3120
rect 48685 3111 48743 3117
rect 48685 3108 48697 3111
rect 47728 3080 48697 3108
rect 47728 3068 47734 3080
rect 48685 3077 48697 3080
rect 48731 3077 48743 3111
rect 48685 3071 48743 3077
rect 50614 3068 50620 3120
rect 50672 3108 50678 3120
rect 51629 3111 51687 3117
rect 51629 3108 51641 3111
rect 50672 3080 51641 3108
rect 50672 3068 50678 3080
rect 51629 3077 51641 3080
rect 51675 3108 51687 3111
rect 51810 3108 51816 3120
rect 51675 3080 51816 3108
rect 51675 3077 51687 3080
rect 51629 3071 51687 3077
rect 51810 3068 51816 3080
rect 51868 3068 51874 3120
rect 40313 3043 40371 3049
rect 40313 3009 40325 3043
rect 40359 3009 40371 3043
rect 40313 3003 40371 3009
rect 41049 3043 41107 3049
rect 41049 3009 41061 3043
rect 41095 3009 41107 3043
rect 41049 3003 41107 3009
rect 41690 3000 41696 3052
rect 41748 3040 41754 3052
rect 41785 3043 41843 3049
rect 41785 3040 41797 3043
rect 41748 3012 41797 3040
rect 41748 3000 41754 3012
rect 41785 3009 41797 3012
rect 41831 3009 41843 3043
rect 41785 3003 41843 3009
rect 42426 3000 42432 3052
rect 42484 3040 42490 3052
rect 42613 3043 42671 3049
rect 42613 3040 42625 3043
rect 42484 3012 42625 3040
rect 42484 3000 42490 3012
rect 42613 3009 42625 3012
rect 42659 3009 42671 3043
rect 43622 3040 43628 3052
rect 43583 3012 43628 3040
rect 42613 3003 42671 3009
rect 43622 3000 43628 3012
rect 43680 3000 43686 3052
rect 44082 3040 44088 3052
rect 44043 3012 44088 3040
rect 44082 3000 44088 3012
rect 44140 3000 44146 3052
rect 44634 3000 44640 3052
rect 44692 3040 44698 3052
rect 44821 3043 44879 3049
rect 44821 3040 44833 3043
rect 44692 3012 44833 3040
rect 44692 3000 44698 3012
rect 44821 3009 44833 3012
rect 44867 3009 44879 3043
rect 45554 3040 45560 3052
rect 45515 3012 45560 3040
rect 44821 3003 44879 3009
rect 45554 3000 45560 3012
rect 45612 3000 45618 3052
rect 46290 3040 46296 3052
rect 46251 3012 46296 3040
rect 46290 3000 46296 3012
rect 46348 3000 46354 3052
rect 46934 3000 46940 3052
rect 46992 3040 46998 3052
rect 47213 3043 47271 3049
rect 47213 3040 47225 3043
rect 46992 3012 47225 3040
rect 46992 3000 46998 3012
rect 47213 3009 47225 3012
rect 47259 3040 47271 3043
rect 47949 3043 48007 3049
rect 47949 3040 47961 3043
rect 47259 3012 47961 3040
rect 47259 3009 47271 3012
rect 47213 3003 47271 3009
rect 47949 3009 47961 3012
rect 47995 3009 48007 3043
rect 47949 3003 48007 3009
rect 48406 3000 48412 3052
rect 48464 3040 48470 3052
rect 49418 3040 49424 3052
rect 48464 3012 49424 3040
rect 48464 3000 48470 3012
rect 49418 3000 49424 3012
rect 49476 3000 49482 3052
rect 50249 3043 50307 3049
rect 50249 3009 50261 3043
rect 50295 3009 50307 3043
rect 50249 3003 50307 3009
rect 50985 3043 51043 3049
rect 50985 3009 50997 3043
rect 51031 3009 51043 3043
rect 50985 3003 51043 3009
rect 32214 2972 32220 2984
rect 24412 2944 32220 2972
rect 32214 2932 32220 2944
rect 32272 2932 32278 2984
rect 32950 2932 32956 2984
rect 33008 2972 33014 2984
rect 33781 2975 33839 2981
rect 33781 2972 33793 2975
rect 33008 2944 33793 2972
rect 33008 2932 33014 2944
rect 33781 2941 33793 2944
rect 33827 2941 33839 2975
rect 33781 2935 33839 2941
rect 34425 2975 34483 2981
rect 34425 2941 34437 2975
rect 34471 2941 34483 2975
rect 34425 2935 34483 2941
rect 15488 2876 22094 2904
rect 15488 2836 15516 2876
rect 31478 2864 31484 2916
rect 31536 2904 31542 2916
rect 32401 2907 32459 2913
rect 32401 2904 32413 2907
rect 31536 2876 32413 2904
rect 31536 2864 31542 2876
rect 32401 2873 32413 2876
rect 32447 2873 32459 2907
rect 32401 2867 32459 2873
rect 33686 2864 33692 2916
rect 33744 2904 33750 2916
rect 34440 2904 34468 2935
rect 35342 2932 35348 2984
rect 35400 2972 35406 2984
rect 35713 2975 35771 2981
rect 35713 2972 35725 2975
rect 35400 2944 35725 2972
rect 35400 2932 35406 2944
rect 35713 2941 35725 2944
rect 35759 2941 35771 2975
rect 35713 2935 35771 2941
rect 49142 2932 49148 2984
rect 49200 2972 49206 2984
rect 49602 2972 49608 2984
rect 49200 2944 49608 2972
rect 49200 2932 49206 2944
rect 49602 2932 49608 2944
rect 49660 2972 49666 2984
rect 50264 2972 50292 3003
rect 49660 2944 50292 2972
rect 49660 2932 49666 2944
rect 33744 2876 34468 2904
rect 33744 2864 33750 2876
rect 42518 2864 42524 2916
rect 42576 2904 42582 2916
rect 42576 2876 43024 2904
rect 42576 2864 42582 2876
rect 12406 2808 15516 2836
rect 18966 2796 18972 2848
rect 19024 2836 19030 2848
rect 19061 2839 19119 2845
rect 19061 2836 19073 2839
rect 19024 2808 19073 2836
rect 19024 2796 19030 2808
rect 19061 2805 19073 2808
rect 19107 2805 19119 2839
rect 20070 2836 20076 2848
rect 20031 2808 20076 2836
rect 19061 2799 19119 2805
rect 20070 2796 20076 2808
rect 20128 2796 20134 2848
rect 20438 2796 20444 2848
rect 20496 2836 20502 2848
rect 20533 2839 20591 2845
rect 20533 2836 20545 2839
rect 20496 2808 20545 2836
rect 20496 2796 20502 2808
rect 20533 2805 20545 2808
rect 20579 2805 20591 2839
rect 20533 2799 20591 2805
rect 21453 2839 21511 2845
rect 21453 2805 21465 2839
rect 21499 2836 21511 2839
rect 21542 2836 21548 2848
rect 21499 2808 21548 2836
rect 21499 2805 21511 2808
rect 21453 2799 21511 2805
rect 21542 2796 21548 2808
rect 21600 2796 21606 2848
rect 22278 2836 22284 2848
rect 22239 2808 22284 2836
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 22646 2796 22652 2848
rect 22704 2836 22710 2848
rect 22741 2839 22799 2845
rect 22741 2836 22753 2839
rect 22704 2808 22753 2836
rect 22704 2796 22710 2808
rect 22741 2805 22753 2808
rect 22787 2805 22799 2839
rect 22741 2799 22799 2805
rect 23382 2796 23388 2848
rect 23440 2836 23446 2848
rect 23477 2839 23535 2845
rect 23477 2836 23489 2839
rect 23440 2808 23489 2836
rect 23440 2796 23446 2808
rect 23477 2805 23489 2808
rect 23523 2805 23535 2839
rect 23477 2799 23535 2805
rect 24118 2796 24124 2848
rect 24176 2836 24182 2848
rect 24213 2839 24271 2845
rect 24213 2836 24225 2839
rect 24176 2808 24225 2836
rect 24176 2796 24182 2808
rect 24213 2805 24225 2808
rect 24259 2805 24271 2839
rect 24213 2799 24271 2805
rect 25041 2839 25099 2845
rect 25041 2805 25053 2839
rect 25087 2836 25099 2839
rect 25222 2836 25228 2848
rect 25087 2808 25228 2836
rect 25087 2805 25099 2808
rect 25041 2799 25099 2805
rect 25222 2796 25228 2808
rect 25280 2796 25286 2848
rect 25777 2839 25835 2845
rect 25777 2805 25789 2839
rect 25823 2836 25835 2839
rect 25958 2836 25964 2848
rect 25823 2808 25964 2836
rect 25823 2805 25835 2808
rect 25777 2799 25835 2805
rect 25958 2796 25964 2808
rect 26016 2796 26022 2848
rect 26513 2839 26571 2845
rect 26513 2805 26525 2839
rect 26559 2836 26571 2839
rect 26694 2836 26700 2848
rect 26559 2808 26700 2836
rect 26559 2805 26571 2808
rect 26513 2799 26571 2805
rect 26694 2796 26700 2808
rect 26752 2796 26758 2848
rect 27430 2796 27436 2848
rect 27488 2836 27494 2848
rect 27617 2839 27675 2845
rect 27617 2836 27629 2839
rect 27488 2808 27629 2836
rect 27488 2796 27494 2808
rect 27617 2805 27629 2808
rect 27663 2805 27675 2839
rect 27617 2799 27675 2805
rect 28166 2796 28172 2848
rect 28224 2836 28230 2848
rect 28353 2839 28411 2845
rect 28353 2836 28365 2839
rect 28224 2808 28365 2836
rect 28224 2796 28230 2808
rect 28353 2805 28365 2808
rect 28399 2805 28411 2839
rect 28353 2799 28411 2805
rect 30006 2796 30012 2848
rect 30064 2836 30070 2848
rect 30193 2839 30251 2845
rect 30193 2836 30205 2839
rect 30064 2808 30205 2836
rect 30064 2796 30070 2808
rect 30193 2805 30205 2808
rect 30239 2805 30251 2839
rect 30193 2799 30251 2805
rect 30742 2796 30748 2848
rect 30800 2836 30806 2848
rect 30929 2839 30987 2845
rect 30929 2836 30941 2839
rect 30800 2808 30941 2836
rect 30800 2796 30806 2808
rect 30929 2805 30941 2808
rect 30975 2805 30987 2839
rect 30929 2799 30987 2805
rect 32214 2796 32220 2848
rect 32272 2836 32278 2848
rect 33137 2839 33195 2845
rect 33137 2836 33149 2839
rect 32272 2808 33149 2836
rect 32272 2796 32278 2808
rect 33137 2805 33149 2808
rect 33183 2805 33195 2839
rect 33137 2799 33195 2805
rect 37734 2796 37740 2848
rect 37792 2836 37798 2848
rect 37921 2839 37979 2845
rect 37921 2836 37933 2839
rect 37792 2808 37933 2836
rect 37792 2796 37798 2808
rect 37921 2805 37933 2808
rect 37967 2805 37979 2839
rect 37921 2799 37979 2805
rect 38470 2796 38476 2848
rect 38528 2836 38534 2848
rect 38749 2839 38807 2845
rect 38749 2836 38761 2839
rect 38528 2808 38761 2836
rect 38528 2796 38534 2808
rect 38749 2805 38761 2808
rect 38795 2805 38807 2839
rect 38749 2799 38807 2805
rect 38838 2796 38844 2848
rect 38896 2836 38902 2848
rect 39485 2839 39543 2845
rect 39485 2836 39497 2839
rect 38896 2808 39497 2836
rect 38896 2796 38902 2808
rect 39485 2805 39497 2808
rect 39531 2805 39543 2839
rect 39485 2799 39543 2805
rect 39574 2796 39580 2848
rect 39632 2836 39638 2848
rect 40129 2839 40187 2845
rect 40129 2836 40141 2839
rect 39632 2808 40141 2836
rect 39632 2796 39638 2808
rect 40129 2805 40141 2808
rect 40175 2805 40187 2839
rect 40129 2799 40187 2805
rect 40310 2796 40316 2848
rect 40368 2836 40374 2848
rect 40865 2839 40923 2845
rect 40865 2836 40877 2839
rect 40368 2808 40877 2836
rect 40368 2796 40374 2808
rect 40865 2805 40877 2808
rect 40911 2805 40923 2839
rect 40865 2799 40923 2805
rect 41046 2796 41052 2848
rect 41104 2836 41110 2848
rect 41601 2839 41659 2845
rect 41601 2836 41613 2839
rect 41104 2808 41613 2836
rect 41104 2796 41110 2808
rect 41601 2805 41613 2808
rect 41647 2805 41659 2839
rect 41601 2799 41659 2805
rect 41782 2796 41788 2848
rect 41840 2836 41846 2848
rect 42797 2839 42855 2845
rect 42797 2836 42809 2839
rect 41840 2808 42809 2836
rect 41840 2796 41846 2808
rect 42797 2805 42809 2808
rect 42843 2805 42855 2839
rect 42996 2836 43024 2876
rect 43254 2864 43260 2916
rect 43312 2904 43318 2916
rect 43312 2876 43576 2904
rect 43312 2864 43318 2876
rect 43441 2839 43499 2845
rect 43441 2836 43453 2839
rect 42996 2808 43453 2836
rect 42797 2799 42855 2805
rect 43441 2805 43453 2808
rect 43487 2805 43499 2839
rect 43548 2836 43576 2876
rect 43990 2864 43996 2916
rect 44048 2904 44054 2916
rect 45005 2907 45063 2913
rect 45005 2904 45017 2907
rect 44048 2876 45017 2904
rect 44048 2864 44054 2876
rect 45005 2873 45017 2876
rect 45051 2873 45063 2907
rect 45005 2867 45063 2873
rect 45462 2864 45468 2916
rect 45520 2904 45526 2916
rect 46477 2907 46535 2913
rect 46477 2904 46489 2907
rect 45520 2876 46489 2904
rect 45520 2864 45526 2876
rect 46477 2873 46489 2876
rect 46523 2873 46535 2907
rect 46477 2867 46535 2873
rect 49878 2864 49884 2916
rect 49936 2904 49942 2916
rect 51000 2904 51028 3003
rect 52181 2907 52239 2913
rect 52181 2904 52193 2907
rect 49936 2876 52193 2904
rect 49936 2864 49942 2876
rect 52181 2873 52193 2876
rect 52227 2873 52239 2907
rect 52181 2867 52239 2873
rect 44269 2839 44327 2845
rect 44269 2836 44281 2839
rect 43548 2808 44281 2836
rect 43441 2799 43499 2805
rect 44269 2805 44281 2808
rect 44315 2805 44327 2839
rect 44269 2799 44327 2805
rect 44726 2796 44732 2848
rect 44784 2836 44790 2848
rect 45741 2839 45799 2845
rect 45741 2836 45753 2839
rect 44784 2808 45753 2836
rect 44784 2796 44790 2808
rect 45741 2805 45753 2808
rect 45787 2805 45799 2839
rect 45741 2799 45799 2805
rect 1104 2746 54832 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 54832 2746
rect 1104 2672 54832 2694
rect 9861 2635 9919 2641
rect 9861 2601 9873 2635
rect 9907 2632 9919 2635
rect 11054 2632 11060 2644
rect 9907 2604 11060 2632
rect 9907 2601 9919 2604
rect 9861 2595 9919 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 11514 2632 11520 2644
rect 11195 2604 11520 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 11793 2635 11851 2641
rect 11793 2601 11805 2635
rect 11839 2632 11851 2635
rect 12526 2632 12532 2644
rect 11839 2604 12532 2632
rect 11839 2601 11851 2604
rect 11793 2595 11851 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 13078 2632 13084 2644
rect 13039 2604 13084 2632
rect 13078 2592 13084 2604
rect 13136 2592 13142 2644
rect 13725 2635 13783 2641
rect 13725 2601 13737 2635
rect 13771 2632 13783 2635
rect 14274 2632 14280 2644
rect 13771 2604 14280 2632
rect 13771 2601 13783 2604
rect 13725 2595 13783 2601
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 15657 2635 15715 2641
rect 15657 2601 15669 2635
rect 15703 2632 15715 2635
rect 16206 2632 16212 2644
rect 15703 2604 16212 2632
rect 15703 2601 15715 2604
rect 15657 2595 15715 2601
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 16301 2635 16359 2641
rect 16301 2601 16313 2635
rect 16347 2632 16359 2635
rect 17034 2632 17040 2644
rect 16347 2604 17040 2632
rect 16347 2601 16359 2604
rect 16301 2595 16359 2601
rect 17034 2592 17040 2604
rect 17092 2592 17098 2644
rect 17402 2632 17408 2644
rect 17363 2604 17408 2632
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 24302 2632 24308 2644
rect 20088 2604 24308 2632
rect 7193 2567 7251 2573
rect 7193 2533 7205 2567
rect 7239 2564 7251 2567
rect 9217 2567 9275 2573
rect 7239 2536 7880 2564
rect 7239 2533 7251 2536
rect 7193 2527 7251 2533
rect 4893 2499 4951 2505
rect 4893 2465 4905 2499
rect 4939 2496 4951 2499
rect 4939 2468 7604 2496
rect 4939 2465 4951 2468
rect 4893 2459 4951 2465
rect 7576 2440 7604 2468
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 5442 2292 5448 2304
rect 5403 2264 5448 2292
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 5994 2292 6000 2304
rect 5955 2264 6000 2292
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 7024 2292 7052 2391
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7616 2400 7665 2428
rect 7616 2388 7622 2400
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 7852 2360 7880 2536
rect 9217 2533 9229 2567
rect 9263 2564 9275 2567
rect 10318 2564 10324 2576
rect 9263 2536 10324 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 10318 2524 10324 2536
rect 10376 2524 10382 2576
rect 10505 2567 10563 2573
rect 10505 2533 10517 2567
rect 10551 2564 10563 2567
rect 11238 2564 11244 2576
rect 10551 2536 11244 2564
rect 10551 2533 10563 2536
rect 10505 2527 10563 2533
rect 11238 2524 11244 2536
rect 11296 2524 11302 2576
rect 15013 2567 15071 2573
rect 12268 2536 14964 2564
rect 7929 2499 7987 2505
rect 7929 2465 7941 2499
rect 7975 2496 7987 2499
rect 12268 2496 12296 2536
rect 7975 2468 12296 2496
rect 14936 2496 14964 2536
rect 15013 2533 15025 2567
rect 15059 2564 15071 2567
rect 15930 2564 15936 2576
rect 15059 2536 15936 2564
rect 15059 2533 15071 2536
rect 15013 2527 15071 2533
rect 15930 2524 15936 2536
rect 15988 2524 15994 2576
rect 20088 2564 20116 2604
rect 24302 2592 24308 2604
rect 24360 2592 24366 2644
rect 30282 2592 30288 2644
rect 30340 2632 30346 2644
rect 36817 2635 36875 2641
rect 36817 2632 36829 2635
rect 30340 2604 36829 2632
rect 30340 2592 30346 2604
rect 36817 2601 36829 2604
rect 36863 2601 36875 2635
rect 36817 2595 36875 2601
rect 16546 2536 20116 2564
rect 20165 2567 20223 2573
rect 16546 2496 16574 2536
rect 20165 2533 20177 2567
rect 20211 2564 20223 2567
rect 20806 2564 20812 2576
rect 20211 2536 20812 2564
rect 20211 2533 20223 2536
rect 20165 2527 20223 2533
rect 20806 2524 20812 2536
rect 20864 2524 20870 2576
rect 28902 2524 28908 2576
rect 28960 2564 28966 2576
rect 29825 2567 29883 2573
rect 29825 2564 29837 2567
rect 28960 2536 29837 2564
rect 28960 2524 28966 2536
rect 29825 2533 29837 2536
rect 29871 2533 29883 2567
rect 29825 2527 29883 2533
rect 30374 2524 30380 2576
rect 30432 2564 30438 2576
rect 31297 2567 31355 2573
rect 31297 2564 31309 2567
rect 30432 2536 31309 2564
rect 30432 2524 30438 2536
rect 31297 2533 31309 2536
rect 31343 2533 31355 2567
rect 31297 2527 31355 2533
rect 31846 2524 31852 2576
rect 31904 2564 31910 2576
rect 33137 2567 33195 2573
rect 33137 2564 33149 2567
rect 31904 2536 33149 2564
rect 31904 2524 31910 2536
rect 33137 2533 33149 2536
rect 33183 2533 33195 2567
rect 33137 2527 33195 2533
rect 22186 2496 22192 2508
rect 14936 2468 16574 2496
rect 18156 2468 22192 2496
rect 7975 2465 7987 2468
rect 7929 2459 7987 2465
rect 9674 2428 9680 2440
rect 9635 2400 9680 2428
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2428 10379 2431
rect 10870 2428 10876 2440
rect 10367 2400 10876 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2428 11023 2431
rect 11606 2428 11612 2440
rect 11011 2400 11612 2428
rect 11011 2397 11023 2400
rect 10965 2391 11023 2397
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2428 12311 2431
rect 12802 2428 12808 2440
rect 12299 2400 12808 2428
rect 12299 2397 12311 2400
rect 12253 2391 12311 2397
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 12897 2431 12955 2437
rect 12897 2397 12909 2431
rect 12943 2428 12955 2431
rect 13541 2431 13599 2437
rect 12943 2400 13492 2428
rect 12943 2397 12955 2400
rect 12897 2391 12955 2397
rect 13464 2360 13492 2400
rect 13541 2397 13553 2431
rect 13587 2424 13599 2431
rect 13906 2428 13912 2440
rect 13648 2424 13912 2428
rect 13587 2400 13912 2424
rect 13587 2397 13676 2400
rect 13541 2396 13676 2397
rect 13541 2391 13599 2396
rect 13906 2388 13912 2400
rect 13964 2388 13970 2440
rect 14826 2428 14832 2440
rect 14739 2400 14832 2428
rect 14826 2388 14832 2400
rect 14884 2428 14890 2440
rect 15378 2428 15384 2440
rect 14884 2400 15384 2428
rect 14884 2388 14890 2400
rect 15378 2388 15384 2400
rect 15436 2388 15442 2440
rect 15473 2431 15531 2437
rect 15473 2397 15485 2431
rect 15519 2428 15531 2431
rect 16022 2428 16028 2440
rect 15519 2400 16028 2428
rect 15519 2397 15531 2400
rect 15473 2391 15531 2397
rect 14182 2360 14188 2372
rect 7852 2332 13400 2360
rect 13464 2332 14188 2360
rect 8662 2292 8668 2304
rect 7024 2264 8668 2292
rect 8662 2252 8668 2264
rect 8720 2252 8726 2304
rect 12437 2295 12495 2301
rect 12437 2261 12449 2295
rect 12483 2292 12495 2295
rect 13262 2292 13268 2304
rect 12483 2264 13268 2292
rect 12483 2261 12495 2264
rect 12437 2255 12495 2261
rect 13262 2252 13268 2264
rect 13320 2252 13326 2304
rect 13372 2292 13400 2332
rect 14182 2320 14188 2332
rect 14240 2320 14246 2372
rect 14369 2363 14427 2369
rect 14369 2329 14381 2363
rect 14415 2360 14427 2363
rect 15488 2360 15516 2391
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16758 2428 16764 2440
rect 16172 2400 16764 2428
rect 16172 2388 16178 2400
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 17589 2431 17647 2437
rect 17589 2397 17601 2431
rect 17635 2428 17647 2431
rect 17862 2428 17868 2440
rect 17635 2400 17868 2428
rect 17635 2397 17647 2400
rect 17589 2391 17647 2397
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 18156 2360 18184 2468
rect 22186 2456 22192 2468
rect 22244 2456 22250 2508
rect 33410 2456 33416 2508
rect 33468 2496 33474 2508
rect 34885 2499 34943 2505
rect 34885 2496 34897 2499
rect 33468 2468 34897 2496
rect 33468 2456 33474 2468
rect 34885 2465 34897 2468
rect 34931 2465 34943 2499
rect 34885 2459 34943 2465
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 18598 2428 18604 2440
rect 18279 2400 18604 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2428 18935 2431
rect 19334 2428 19340 2440
rect 18923 2400 19340 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19334 2388 19340 2400
rect 19392 2388 19398 2440
rect 20809 2431 20867 2437
rect 20809 2397 20821 2431
rect 20855 2428 20867 2431
rect 21174 2428 21180 2440
rect 20855 2400 21180 2428
rect 20855 2397 20867 2400
rect 20809 2391 20867 2397
rect 21174 2388 21180 2400
rect 21232 2388 21238 2440
rect 21453 2431 21511 2437
rect 21453 2397 21465 2431
rect 21499 2428 21511 2431
rect 21910 2428 21916 2440
rect 21499 2400 21916 2428
rect 21499 2397 21511 2400
rect 21453 2391 21511 2397
rect 21910 2388 21916 2400
rect 21968 2388 21974 2440
rect 22554 2428 22560 2440
rect 22515 2400 22560 2428
rect 22554 2388 22560 2400
rect 22612 2388 22618 2440
rect 23290 2428 23296 2440
rect 23251 2400 23296 2428
rect 23290 2388 23296 2400
rect 23348 2388 23354 2440
rect 23474 2388 23480 2440
rect 23532 2428 23538 2440
rect 23753 2431 23811 2437
rect 23753 2428 23765 2431
rect 23532 2400 23765 2428
rect 23532 2388 23538 2400
rect 23753 2397 23765 2400
rect 23799 2397 23811 2431
rect 23753 2391 23811 2397
rect 24857 2431 24915 2437
rect 24857 2397 24869 2431
rect 24903 2428 24915 2431
rect 25038 2428 25044 2440
rect 24903 2400 25044 2428
rect 24903 2397 24915 2400
rect 24857 2391 24915 2397
rect 25038 2388 25044 2400
rect 25096 2388 25102 2440
rect 25593 2431 25651 2437
rect 25593 2397 25605 2431
rect 25639 2428 25651 2431
rect 25866 2428 25872 2440
rect 25639 2400 25872 2428
rect 25639 2397 25651 2400
rect 25593 2391 25651 2397
rect 25866 2388 25872 2400
rect 25924 2388 25930 2440
rect 26326 2428 26332 2440
rect 26287 2400 26332 2428
rect 26326 2388 26332 2400
rect 26384 2388 26390 2440
rect 27433 2431 27491 2437
rect 27433 2397 27445 2431
rect 27479 2428 27491 2431
rect 27890 2428 27896 2440
rect 27479 2400 27896 2428
rect 27479 2397 27491 2400
rect 27433 2391 27491 2397
rect 27890 2388 27896 2400
rect 27948 2388 27954 2440
rect 28169 2431 28227 2437
rect 28169 2397 28181 2431
rect 28215 2428 28227 2431
rect 28534 2428 28540 2440
rect 28215 2400 28540 2428
rect 28215 2397 28227 2400
rect 28169 2391 28227 2397
rect 28534 2388 28540 2400
rect 28592 2388 28598 2440
rect 29181 2431 29239 2437
rect 29181 2397 29193 2431
rect 29227 2428 29239 2431
rect 29638 2428 29644 2440
rect 29227 2400 29644 2428
rect 29227 2397 29239 2400
rect 29181 2391 29239 2397
rect 29638 2388 29644 2400
rect 29696 2388 29702 2440
rect 29914 2388 29920 2440
rect 29972 2428 29978 2440
rect 30009 2431 30067 2437
rect 30009 2428 30021 2431
rect 29972 2400 30021 2428
rect 29972 2388 29978 2400
rect 30009 2397 30021 2400
rect 30055 2397 30067 2431
rect 30009 2391 30067 2397
rect 30745 2431 30803 2437
rect 30745 2397 30757 2431
rect 30791 2428 30803 2431
rect 30926 2428 30932 2440
rect 30791 2400 30932 2428
rect 30791 2397 30803 2400
rect 30745 2391 30803 2397
rect 30926 2388 30932 2400
rect 30984 2388 30990 2440
rect 31481 2431 31539 2437
rect 31481 2397 31493 2431
rect 31527 2428 31539 2431
rect 31754 2428 31760 2440
rect 31527 2400 31760 2428
rect 31527 2397 31539 2400
rect 31481 2391 31539 2397
rect 31754 2388 31760 2400
rect 31812 2388 31818 2440
rect 32585 2431 32643 2437
rect 32585 2397 32597 2431
rect 32631 2428 32643 2431
rect 32858 2428 32864 2440
rect 32631 2400 32864 2428
rect 32631 2397 32643 2400
rect 32585 2391 32643 2397
rect 32858 2388 32864 2400
rect 32916 2388 32922 2440
rect 33321 2431 33379 2437
rect 33321 2397 33333 2431
rect 33367 2428 33379 2431
rect 33778 2428 33784 2440
rect 33367 2400 33784 2428
rect 33367 2397 33379 2400
rect 33321 2391 33379 2397
rect 33778 2388 33784 2400
rect 33836 2388 33842 2440
rect 34057 2431 34115 2437
rect 34057 2397 34069 2431
rect 34103 2397 34115 2431
rect 34057 2391 34115 2397
rect 14415 2332 15516 2360
rect 16546 2332 18184 2360
rect 18616 2360 18644 2388
rect 19429 2363 19487 2369
rect 19429 2360 19441 2363
rect 18616 2332 19441 2360
rect 14415 2329 14427 2332
rect 14369 2323 14427 2329
rect 16546 2292 16574 2332
rect 19429 2329 19441 2332
rect 19475 2329 19487 2363
rect 34072 2360 34100 2391
rect 34146 2388 34152 2440
rect 34204 2428 34210 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 34204 2400 35541 2428
rect 34204 2388 34210 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 36832 2428 36860 2595
rect 47578 2592 47584 2644
rect 47636 2632 47642 2644
rect 49421 2635 49479 2641
rect 49421 2632 49433 2635
rect 47636 2604 49433 2632
rect 47636 2592 47642 2604
rect 49421 2601 49433 2604
rect 49467 2601 49479 2635
rect 49421 2595 49479 2601
rect 37366 2524 37372 2576
rect 37424 2564 37430 2576
rect 38381 2567 38439 2573
rect 38381 2564 38393 2567
rect 37424 2536 38393 2564
rect 37424 2524 37430 2536
rect 38381 2533 38393 2536
rect 38427 2533 38439 2567
rect 38381 2527 38439 2533
rect 39942 2524 39948 2576
rect 40000 2564 40006 2576
rect 40957 2567 41015 2573
rect 40957 2564 40969 2567
rect 40000 2536 40969 2564
rect 40000 2524 40006 2536
rect 40957 2533 40969 2536
rect 41003 2533 41015 2567
rect 40957 2527 41015 2533
rect 41414 2524 41420 2576
rect 41472 2564 41478 2576
rect 42705 2567 42763 2573
rect 42705 2564 42717 2567
rect 41472 2536 42717 2564
rect 41472 2524 41478 2536
rect 42705 2533 42717 2536
rect 42751 2533 42763 2567
rect 42705 2527 42763 2533
rect 42886 2524 42892 2576
rect 42944 2564 42950 2576
rect 44269 2567 44327 2573
rect 44269 2564 44281 2567
rect 42944 2536 44281 2564
rect 42944 2524 42950 2536
rect 44269 2533 44281 2536
rect 44315 2533 44327 2567
rect 44269 2527 44327 2533
rect 44358 2524 44364 2576
rect 44416 2564 44422 2576
rect 46109 2567 46167 2573
rect 46109 2564 46121 2567
rect 44416 2536 46121 2564
rect 44416 2524 44422 2536
rect 46109 2533 46121 2536
rect 46155 2533 46167 2567
rect 46109 2527 46167 2533
rect 46198 2524 46204 2576
rect 46256 2564 46262 2576
rect 47949 2567 48007 2573
rect 47949 2564 47961 2567
rect 46256 2536 47961 2564
rect 46256 2524 46262 2536
rect 47949 2533 47961 2536
rect 47995 2533 48007 2567
rect 48498 2564 48504 2576
rect 48459 2536 48504 2564
rect 47949 2527 48007 2533
rect 48498 2524 48504 2536
rect 48556 2524 48562 2576
rect 49970 2524 49976 2576
rect 50028 2564 50034 2576
rect 50341 2567 50399 2573
rect 50341 2564 50353 2567
rect 50028 2536 50353 2564
rect 50028 2524 50034 2536
rect 50341 2533 50353 2536
rect 50387 2533 50399 2567
rect 51074 2564 51080 2576
rect 51035 2536 51080 2564
rect 50341 2527 50399 2533
rect 51074 2524 51080 2536
rect 51132 2524 51138 2576
rect 42794 2456 42800 2508
rect 42852 2496 42858 2508
rect 42852 2468 43392 2496
rect 42852 2456 42858 2468
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 36832 2400 37473 2428
rect 35529 2391 35587 2397
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 37918 2388 37924 2440
rect 37976 2428 37982 2440
rect 38197 2431 38255 2437
rect 38197 2428 38209 2431
rect 37976 2400 38209 2428
rect 37976 2388 37982 2400
rect 38197 2397 38209 2400
rect 38243 2397 38255 2431
rect 38197 2391 38255 2397
rect 38746 2388 38752 2440
rect 38804 2428 38810 2440
rect 38933 2431 38991 2437
rect 38933 2428 38945 2431
rect 38804 2400 38945 2428
rect 38804 2388 38810 2400
rect 38933 2397 38945 2400
rect 38979 2397 38991 2431
rect 40034 2428 40040 2440
rect 39995 2400 40040 2428
rect 38933 2391 38991 2397
rect 40034 2388 40040 2400
rect 40092 2388 40098 2440
rect 40770 2428 40776 2440
rect 40731 2400 40776 2428
rect 40770 2388 40776 2400
rect 40828 2388 40834 2440
rect 41506 2428 41512 2440
rect 41467 2400 41512 2428
rect 41506 2388 41512 2400
rect 41564 2388 41570 2440
rect 42889 2431 42947 2437
rect 42889 2397 42901 2431
rect 42935 2428 42947 2431
rect 42978 2428 42984 2440
rect 42935 2400 42984 2428
rect 42935 2397 42947 2400
rect 42889 2391 42947 2397
rect 42978 2388 42984 2400
rect 43036 2388 43042 2440
rect 43364 2437 43392 2468
rect 45646 2456 45652 2508
rect 45704 2496 45710 2508
rect 45704 2468 46704 2496
rect 45704 2456 45710 2468
rect 43349 2431 43407 2437
rect 43349 2397 43361 2431
rect 43395 2397 43407 2431
rect 43349 2391 43407 2397
rect 43898 2388 43904 2440
rect 43956 2428 43962 2440
rect 44085 2431 44143 2437
rect 44085 2428 44097 2431
rect 43956 2400 44097 2428
rect 43956 2388 43962 2400
rect 44085 2397 44097 2400
rect 44131 2397 44143 2431
rect 45186 2428 45192 2440
rect 45147 2400 45192 2428
rect 44085 2391 44143 2397
rect 45186 2388 45192 2400
rect 45244 2388 45250 2440
rect 45738 2388 45744 2440
rect 45796 2428 45802 2440
rect 46676 2437 46704 2468
rect 45925 2431 45983 2437
rect 45925 2428 45937 2431
rect 45796 2400 45937 2428
rect 45796 2388 45802 2400
rect 45925 2397 45937 2400
rect 45971 2397 45983 2431
rect 45925 2391 45983 2397
rect 46661 2431 46719 2437
rect 46661 2397 46673 2431
rect 46707 2397 46719 2431
rect 47762 2428 47768 2440
rect 47723 2400 47768 2428
rect 46661 2391 46719 2397
rect 47762 2388 47768 2400
rect 47820 2388 47826 2440
rect 48038 2388 48044 2440
rect 48096 2428 48102 2440
rect 49050 2428 49056 2440
rect 48096 2400 49056 2428
rect 48096 2388 48102 2400
rect 49050 2388 49056 2400
rect 49108 2428 49114 2440
rect 49237 2431 49295 2437
rect 49237 2428 49249 2431
rect 49108 2400 49249 2428
rect 49108 2388 49114 2400
rect 49237 2397 49249 2400
rect 49283 2397 49295 2431
rect 49237 2391 49295 2397
rect 49694 2388 49700 2440
rect 49752 2428 49758 2440
rect 51261 2431 51319 2437
rect 51261 2428 51273 2431
rect 49752 2400 51273 2428
rect 49752 2388 49758 2400
rect 51261 2397 51273 2400
rect 51307 2428 51319 2431
rect 52917 2431 52975 2437
rect 52917 2428 52929 2431
rect 51307 2400 52929 2428
rect 51307 2397 51319 2400
rect 51261 2391 51319 2397
rect 52917 2397 52929 2400
rect 52963 2397 52975 2431
rect 52917 2391 52975 2397
rect 34514 2360 34520 2372
rect 34072 2332 34520 2360
rect 19429 2323 19487 2329
rect 34514 2320 34520 2332
rect 34572 2320 34578 2372
rect 34790 2320 34796 2372
rect 34848 2360 34854 2372
rect 36173 2363 36231 2369
rect 36173 2360 36185 2363
rect 34848 2332 36185 2360
rect 34848 2320 34854 2332
rect 36173 2329 36185 2332
rect 36219 2329 36231 2363
rect 36173 2323 36231 2329
rect 45094 2320 45100 2372
rect 45152 2360 45158 2372
rect 45152 2332 46888 2360
rect 45152 2320 45158 2332
rect 13372 2264 16574 2292
rect 16945 2295 17003 2301
rect 16945 2261 16957 2295
rect 16991 2292 17003 2295
rect 17126 2292 17132 2304
rect 16991 2264 17132 2292
rect 16991 2261 17003 2264
rect 16945 2255 17003 2261
rect 17126 2252 17132 2264
rect 17184 2252 17190 2304
rect 22373 2295 22431 2301
rect 22373 2261 22385 2295
rect 22419 2292 22431 2295
rect 23014 2292 23020 2304
rect 22419 2264 23020 2292
rect 22419 2261 22431 2264
rect 22373 2255 22431 2261
rect 23014 2252 23020 2264
rect 23072 2252 23078 2304
rect 23109 2295 23167 2301
rect 23109 2261 23121 2295
rect 23155 2292 23167 2295
rect 23750 2292 23756 2304
rect 23155 2264 23756 2292
rect 23155 2261 23167 2264
rect 23109 2255 23167 2261
rect 23750 2252 23756 2264
rect 23808 2252 23814 2304
rect 23937 2295 23995 2301
rect 23937 2261 23949 2295
rect 23983 2292 23995 2295
rect 24486 2292 24492 2304
rect 23983 2264 24492 2292
rect 23983 2261 23995 2264
rect 23937 2255 23995 2261
rect 24486 2252 24492 2264
rect 24544 2252 24550 2304
rect 25041 2295 25099 2301
rect 25041 2261 25053 2295
rect 25087 2292 25099 2295
rect 25590 2292 25596 2304
rect 25087 2264 25596 2292
rect 25087 2261 25099 2264
rect 25041 2255 25099 2261
rect 25590 2252 25596 2264
rect 25648 2252 25654 2304
rect 25777 2295 25835 2301
rect 25777 2261 25789 2295
rect 25823 2292 25835 2295
rect 26326 2292 26332 2304
rect 25823 2264 26332 2292
rect 25823 2261 25835 2264
rect 25777 2255 25835 2261
rect 26326 2252 26332 2264
rect 26384 2252 26390 2304
rect 26513 2295 26571 2301
rect 26513 2261 26525 2295
rect 26559 2292 26571 2295
rect 27062 2292 27068 2304
rect 26559 2264 27068 2292
rect 26559 2261 26571 2264
rect 26513 2255 26571 2261
rect 27062 2252 27068 2264
rect 27120 2252 27126 2304
rect 27617 2295 27675 2301
rect 27617 2261 27629 2295
rect 27663 2292 27675 2295
rect 27798 2292 27804 2304
rect 27663 2264 27804 2292
rect 27663 2261 27675 2264
rect 27617 2255 27675 2261
rect 27798 2252 27804 2264
rect 27856 2252 27862 2304
rect 28353 2295 28411 2301
rect 28353 2261 28365 2295
rect 28399 2292 28411 2295
rect 28534 2292 28540 2304
rect 28399 2264 28540 2292
rect 28399 2261 28411 2264
rect 28353 2255 28411 2261
rect 28534 2252 28540 2264
rect 28592 2252 28598 2304
rect 28997 2295 29055 2301
rect 28997 2261 29009 2295
rect 29043 2292 29055 2295
rect 29270 2292 29276 2304
rect 29043 2264 29276 2292
rect 29043 2261 29055 2264
rect 28997 2255 29055 2261
rect 29270 2252 29276 2264
rect 29328 2252 29334 2304
rect 29638 2252 29644 2304
rect 29696 2292 29702 2304
rect 30561 2295 30619 2301
rect 30561 2292 30573 2295
rect 29696 2264 30573 2292
rect 29696 2252 29702 2264
rect 30561 2261 30573 2264
rect 30607 2261 30619 2295
rect 30561 2255 30619 2261
rect 31110 2252 31116 2304
rect 31168 2292 31174 2304
rect 32401 2295 32459 2301
rect 32401 2292 32413 2295
rect 31168 2264 32413 2292
rect 31168 2252 31174 2264
rect 32401 2261 32413 2264
rect 32447 2261 32459 2295
rect 32401 2255 32459 2261
rect 32582 2252 32588 2304
rect 32640 2292 32646 2304
rect 33873 2295 33931 2301
rect 33873 2292 33885 2295
rect 32640 2264 33885 2292
rect 32640 2252 32646 2264
rect 33873 2261 33885 2264
rect 33919 2261 33931 2295
rect 33873 2255 33931 2261
rect 36998 2252 37004 2304
rect 37056 2292 37062 2304
rect 37645 2295 37703 2301
rect 37645 2292 37657 2295
rect 37056 2264 37657 2292
rect 37056 2252 37062 2264
rect 37645 2261 37657 2264
rect 37691 2261 37703 2295
rect 37645 2255 37703 2261
rect 38102 2252 38108 2304
rect 38160 2292 38166 2304
rect 39117 2295 39175 2301
rect 39117 2292 39129 2295
rect 38160 2264 39129 2292
rect 38160 2252 38166 2264
rect 39117 2261 39129 2264
rect 39163 2261 39175 2295
rect 39117 2255 39175 2261
rect 39206 2252 39212 2304
rect 39264 2292 39270 2304
rect 40221 2295 40279 2301
rect 40221 2292 40233 2295
rect 39264 2264 40233 2292
rect 39264 2252 39270 2264
rect 40221 2261 40233 2264
rect 40267 2261 40279 2295
rect 40221 2255 40279 2261
rect 40678 2252 40684 2304
rect 40736 2292 40742 2304
rect 41693 2295 41751 2301
rect 41693 2292 41705 2295
rect 40736 2264 41705 2292
rect 40736 2252 40742 2264
rect 41693 2261 41705 2264
rect 41739 2261 41751 2295
rect 41693 2255 41751 2261
rect 42150 2252 42156 2304
rect 42208 2292 42214 2304
rect 43533 2295 43591 2301
rect 43533 2292 43545 2295
rect 42208 2264 43545 2292
rect 42208 2252 42214 2264
rect 43533 2261 43545 2264
rect 43579 2261 43591 2295
rect 43533 2255 43591 2261
rect 43622 2252 43628 2304
rect 43680 2292 43686 2304
rect 46860 2301 46888 2332
rect 47302 2320 47308 2372
rect 47360 2360 47366 2372
rect 48685 2363 48743 2369
rect 48685 2360 48697 2363
rect 47360 2332 48697 2360
rect 47360 2320 47366 2332
rect 48685 2329 48697 2332
rect 48731 2360 48743 2363
rect 48866 2360 48872 2372
rect 48731 2332 48872 2360
rect 48731 2329 48743 2332
rect 48685 2323 48743 2329
rect 48866 2320 48872 2332
rect 48924 2320 48930 2372
rect 48958 2320 48964 2372
rect 49016 2360 49022 2372
rect 50154 2360 50160 2372
rect 49016 2332 50160 2360
rect 49016 2320 49022 2332
rect 50154 2320 50160 2332
rect 50212 2360 50218 2372
rect 50525 2363 50583 2369
rect 50525 2360 50537 2363
rect 50212 2332 50537 2360
rect 50212 2320 50218 2332
rect 50525 2329 50537 2332
rect 50571 2329 50583 2363
rect 51810 2360 51816 2372
rect 51771 2332 51816 2360
rect 50525 2323 50583 2329
rect 51810 2320 51816 2332
rect 51868 2320 51874 2372
rect 51994 2360 52000 2372
rect 51955 2332 52000 2360
rect 51994 2320 52000 2332
rect 52052 2320 52058 2372
rect 45373 2295 45431 2301
rect 45373 2292 45385 2295
rect 43680 2264 45385 2292
rect 43680 2252 43686 2264
rect 45373 2261 45385 2264
rect 45419 2261 45431 2295
rect 45373 2255 45431 2261
rect 46845 2295 46903 2301
rect 46845 2261 46857 2295
rect 46891 2261 46903 2295
rect 46845 2255 46903 2261
rect 1104 2202 54832 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 54832 2202
rect 1104 2128 54832 2150
rect 5442 2048 5448 2100
rect 5500 2088 5506 2100
rect 9674 2088 9680 2100
rect 5500 2060 9680 2088
rect 5500 2048 5506 2060
rect 9674 2048 9680 2060
rect 9732 2088 9738 2100
rect 10870 2088 10876 2100
rect 9732 2060 10876 2088
rect 9732 2048 9738 2060
rect 10870 2048 10876 2060
rect 10928 2048 10934 2100
rect 13906 2048 13912 2100
rect 13964 2088 13970 2100
rect 14918 2088 14924 2100
rect 13964 2060 14924 2088
rect 13964 2048 13970 2060
rect 14918 2048 14924 2060
rect 14976 2048 14982 2100
rect 50246 2048 50252 2100
rect 50304 2088 50310 2100
rect 51994 2088 52000 2100
rect 50304 2060 52000 2088
rect 50304 2048 50310 2060
rect 51994 2048 52000 2060
rect 52052 2048 52058 2100
rect 5994 1980 6000 2032
rect 6052 2020 6058 2032
rect 11606 2020 11612 2032
rect 6052 1992 11612 2020
rect 6052 1980 6058 1992
rect 11606 1980 11612 1992
rect 11664 1980 11670 2032
<< via1 >>
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 8576 53227 8628 53236
rect 8576 53193 8585 53227
rect 8585 53193 8619 53227
rect 8619 53193 8628 53227
rect 8576 53184 8628 53193
rect 9312 53227 9364 53236
rect 9312 53193 9321 53227
rect 9321 53193 9355 53227
rect 9355 53193 9364 53227
rect 9312 53184 9364 53193
rect 25596 53184 25648 53236
rect 26608 53227 26660 53236
rect 26608 53193 26617 53227
rect 26617 53193 26651 53227
rect 26651 53193 26660 53227
rect 26608 53184 26660 53193
rect 29184 53227 29236 53236
rect 29184 53193 29193 53227
rect 29193 53193 29227 53227
rect 29227 53193 29236 53227
rect 29184 53184 29236 53193
rect 31760 53227 31812 53236
rect 31760 53193 31769 53227
rect 31769 53193 31803 53227
rect 31803 53193 31812 53227
rect 31760 53184 31812 53193
rect 47124 53227 47176 53236
rect 47124 53193 47133 53227
rect 47133 53193 47167 53227
rect 47167 53193 47176 53227
rect 47124 53184 47176 53193
rect 49700 53227 49752 53236
rect 49700 53193 49709 53227
rect 49709 53193 49743 53227
rect 49743 53193 49752 53227
rect 49700 53184 49752 53193
rect 3148 53159 3200 53168
rect 3148 53125 3157 53159
rect 3157 53125 3191 53159
rect 3191 53125 3200 53159
rect 3148 53116 3200 53125
rect 5448 53159 5500 53168
rect 5448 53125 5457 53159
rect 5457 53125 5491 53159
rect 5491 53125 5500 53159
rect 5448 53116 5500 53125
rect 6644 53159 6696 53168
rect 6644 53125 6653 53159
rect 6653 53125 6687 53159
rect 6687 53125 6696 53159
rect 6644 53116 6696 53125
rect 1676 52980 1728 53032
rect 2596 53023 2648 53032
rect 2596 52989 2605 53023
rect 2605 52989 2639 53023
rect 2639 52989 2648 53023
rect 2596 52980 2648 52989
rect 4068 53048 4120 53100
rect 7748 53091 7800 53100
rect 7748 53057 7757 53091
rect 7757 53057 7791 53091
rect 7791 53057 7800 53091
rect 7748 53048 7800 53057
rect 10140 53091 10192 53100
rect 10140 53057 10149 53091
rect 10149 53057 10183 53091
rect 10183 53057 10192 53091
rect 10140 53048 10192 53057
rect 12532 53091 12584 53100
rect 12532 53057 12541 53091
rect 12541 53057 12575 53091
rect 12575 53057 12584 53091
rect 12532 53048 12584 53057
rect 14832 53091 14884 53100
rect 14832 53057 14841 53091
rect 14841 53057 14875 53091
rect 14875 53057 14884 53091
rect 14832 53048 14884 53057
rect 16304 53091 16356 53100
rect 16304 53057 16313 53091
rect 16313 53057 16347 53091
rect 16347 53057 16356 53091
rect 16304 53048 16356 53057
rect 8208 52980 8260 53032
rect 10416 53023 10468 53032
rect 10416 52989 10425 53023
rect 10425 52989 10459 53023
rect 10459 52989 10468 53023
rect 10416 52980 10468 52989
rect 12808 53023 12860 53032
rect 12808 52989 12817 53023
rect 12817 52989 12851 53023
rect 12851 52989 12860 53023
rect 12808 52980 12860 52989
rect 16028 53023 16080 53032
rect 16028 52989 16037 53023
rect 16037 52989 16071 53023
rect 16071 52989 16080 53023
rect 16028 52980 16080 52989
rect 24492 53116 24544 53168
rect 18420 53048 18472 53100
rect 18788 53048 18840 53100
rect 19432 53048 19484 53100
rect 20904 53091 20956 53100
rect 20904 53057 20913 53091
rect 20913 53057 20947 53091
rect 20947 53057 20956 53091
rect 20904 53048 20956 53057
rect 22008 53048 22060 53100
rect 23296 53091 23348 53100
rect 23296 53057 23305 53091
rect 23305 53057 23339 53091
rect 23339 53057 23348 53091
rect 23296 53048 23348 53057
rect 24584 53091 24636 53100
rect 24584 53057 24593 53091
rect 24593 53057 24627 53091
rect 24627 53057 24636 53091
rect 24584 53048 24636 53057
rect 25688 53091 25740 53100
rect 25688 53057 25697 53091
rect 25697 53057 25731 53091
rect 25731 53057 25740 53091
rect 25688 53048 25740 53057
rect 28264 53091 28316 53100
rect 28264 53057 28273 53091
rect 28273 53057 28307 53091
rect 28307 53057 28316 53091
rect 28264 53048 28316 53057
rect 30656 53091 30708 53100
rect 30656 53057 30665 53091
rect 30665 53057 30699 53091
rect 30699 53057 30708 53091
rect 30656 53048 30708 53057
rect 32220 53116 32272 53168
rect 47032 53116 47084 53168
rect 32772 53048 32824 53100
rect 34244 53091 34296 53100
rect 34244 53057 34253 53091
rect 34253 53057 34287 53091
rect 34287 53057 34296 53091
rect 34244 53048 34296 53057
rect 35440 53091 35492 53100
rect 35440 53057 35449 53091
rect 35449 53057 35483 53091
rect 35483 53057 35492 53091
rect 35440 53048 35492 53057
rect 36636 53091 36688 53100
rect 36636 53057 36645 53091
rect 36645 53057 36679 53091
rect 36679 53057 36688 53091
rect 36636 53048 36688 53057
rect 37832 53091 37884 53100
rect 37832 53057 37841 53091
rect 37841 53057 37875 53091
rect 37875 53057 37884 53091
rect 37832 53048 37884 53057
rect 39028 53091 39080 53100
rect 39028 53057 39037 53091
rect 39037 53057 39071 53091
rect 39071 53057 39080 53091
rect 39028 53048 39080 53057
rect 40040 53048 40092 53100
rect 41420 53091 41472 53100
rect 41420 53057 41429 53091
rect 41429 53057 41463 53091
rect 41463 53057 41472 53091
rect 41420 53048 41472 53057
rect 42340 53048 42392 53100
rect 43628 53091 43680 53100
rect 43628 53057 43637 53091
rect 43637 53057 43671 53091
rect 43671 53057 43680 53091
rect 43628 53048 43680 53057
rect 44732 53048 44784 53100
rect 45192 53091 45244 53100
rect 45192 53057 45201 53091
rect 45201 53057 45235 53091
rect 45235 53057 45244 53091
rect 45192 53048 45244 53057
rect 51080 53116 51132 53168
rect 51448 53116 51500 53168
rect 53196 53091 53248 53100
rect 53196 53057 53205 53091
rect 53205 53057 53239 53091
rect 53239 53057 53248 53091
rect 53196 53048 53248 53057
rect 21456 52980 21508 53032
rect 34796 52980 34848 53032
rect 43904 53023 43956 53032
rect 24032 52912 24084 52964
rect 26700 52912 26752 52964
rect 32128 52912 32180 52964
rect 34704 52912 34756 52964
rect 43904 52989 43913 53023
rect 43913 52989 43947 53023
rect 43947 52989 43956 53023
rect 43904 52980 43956 52989
rect 45468 53023 45520 53032
rect 45468 52989 45477 53023
rect 45477 52989 45511 53023
rect 45511 52989 45520 53023
rect 45468 52980 45520 52989
rect 48044 53023 48096 53032
rect 48044 52989 48053 53023
rect 48053 52989 48087 53023
rect 48087 52989 48096 53023
rect 48044 52980 48096 52989
rect 50160 52980 50212 53032
rect 3240 52887 3292 52896
rect 3240 52853 3249 52887
rect 3249 52853 3283 52887
rect 3283 52853 3292 52887
rect 3240 52844 3292 52853
rect 5540 52887 5592 52896
rect 5540 52853 5549 52887
rect 5549 52853 5583 52887
rect 5583 52853 5592 52887
rect 5540 52844 5592 52853
rect 6736 52887 6788 52896
rect 6736 52853 6745 52887
rect 6745 52853 6779 52887
rect 6779 52853 6788 52887
rect 6736 52844 6788 52853
rect 11704 52844 11756 52896
rect 15016 52887 15068 52896
rect 15016 52853 15025 52887
rect 15025 52853 15059 52887
rect 15059 52853 15068 52887
rect 15016 52844 15068 52853
rect 22284 52887 22336 52896
rect 22284 52853 22293 52887
rect 22293 52853 22327 52887
rect 22327 52853 22336 52887
rect 22284 52844 22336 52853
rect 25412 52844 25464 52896
rect 25964 52844 26016 52896
rect 26976 52844 27028 52896
rect 28080 52887 28132 52896
rect 28080 52853 28089 52887
rect 28089 52853 28123 52887
rect 28123 52853 28132 52887
rect 28080 52844 28132 52853
rect 28724 52844 28776 52896
rect 30104 52844 30156 52896
rect 31208 52844 31260 52896
rect 32588 52844 32640 52896
rect 34336 52844 34388 52896
rect 35348 52844 35400 52896
rect 38844 52887 38896 52896
rect 38844 52853 38853 52887
rect 38853 52853 38887 52887
rect 38887 52853 38896 52887
rect 38844 52844 38896 52853
rect 38936 52844 38988 52896
rect 41236 52887 41288 52896
rect 41236 52853 41245 52887
rect 41245 52853 41279 52887
rect 41279 52853 41288 52887
rect 41236 52844 41288 52853
rect 42616 52887 42668 52896
rect 42616 52853 42625 52887
rect 42625 52853 42659 52887
rect 42659 52853 42668 52887
rect 42616 52844 42668 52853
rect 49516 52844 49568 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 3148 52683 3200 52692
rect 3148 52649 3157 52683
rect 3157 52649 3191 52683
rect 3191 52649 3200 52683
rect 3148 52640 3200 52649
rect 4068 52683 4120 52692
rect 4068 52649 4077 52683
rect 4077 52649 4111 52683
rect 4111 52649 4120 52683
rect 4068 52640 4120 52649
rect 6644 52640 6696 52692
rect 7748 52640 7800 52692
rect 10140 52640 10192 52692
rect 13636 52683 13688 52692
rect 13636 52649 13645 52683
rect 13645 52649 13679 52683
rect 13679 52649 13688 52683
rect 13636 52640 13688 52649
rect 14832 52640 14884 52692
rect 18788 52683 18840 52692
rect 18788 52649 18797 52683
rect 18797 52649 18831 52683
rect 18831 52649 18840 52683
rect 18788 52640 18840 52649
rect 19432 52640 19484 52692
rect 22008 52683 22060 52692
rect 22008 52649 22017 52683
rect 22017 52649 22051 52683
rect 22051 52649 22060 52683
rect 22008 52640 22060 52649
rect 25688 52640 25740 52692
rect 28264 52640 28316 52692
rect 32772 52683 32824 52692
rect 32772 52649 32781 52683
rect 32781 52649 32815 52683
rect 32815 52649 32824 52683
rect 32772 52640 32824 52649
rect 34244 52640 34296 52692
rect 36636 52640 36688 52692
rect 39028 52640 39080 52692
rect 42340 52640 42392 52692
rect 43628 52640 43680 52692
rect 45192 52683 45244 52692
rect 45192 52649 45201 52683
rect 45201 52649 45235 52683
rect 45235 52649 45244 52683
rect 45192 52640 45244 52649
rect 51908 52640 51960 52692
rect 53196 52640 53248 52692
rect 34520 52572 34572 52624
rect 41236 52572 41288 52624
rect 47032 52572 47084 52624
rect 11336 52547 11388 52556
rect 11336 52513 11345 52547
rect 11345 52513 11379 52547
rect 11379 52513 11388 52547
rect 11336 52504 11388 52513
rect 17316 52547 17368 52556
rect 17316 52513 17325 52547
rect 17325 52513 17359 52547
rect 17359 52513 17368 52547
rect 17316 52504 17368 52513
rect 33048 52504 33100 52556
rect 42616 52504 42668 52556
rect 46020 52547 46072 52556
rect 46020 52513 46029 52547
rect 46029 52513 46063 52547
rect 46063 52513 46072 52547
rect 46020 52504 46072 52513
rect 48412 52547 48464 52556
rect 48412 52513 48421 52547
rect 48421 52513 48455 52547
rect 48455 52513 48464 52547
rect 48412 52504 48464 52513
rect 52000 52547 52052 52556
rect 52000 52513 52009 52547
rect 52009 52513 52043 52547
rect 52043 52513 52052 52547
rect 52000 52504 52052 52513
rect 1768 52436 1820 52488
rect 2504 52436 2556 52488
rect 11612 52479 11664 52488
rect 11612 52445 11621 52479
rect 11621 52445 11655 52479
rect 11655 52445 11664 52479
rect 11612 52436 11664 52445
rect 13636 52436 13688 52488
rect 22836 52436 22888 52488
rect 26056 52436 26108 52488
rect 27160 52479 27212 52488
rect 27160 52445 27169 52479
rect 27169 52445 27203 52479
rect 27203 52445 27212 52479
rect 27160 52436 27212 52445
rect 46296 52479 46348 52488
rect 46296 52445 46305 52479
rect 46305 52445 46339 52479
rect 46339 52445 46348 52479
rect 46296 52436 46348 52445
rect 51908 52436 51960 52488
rect 54024 52479 54076 52488
rect 54024 52445 54033 52479
rect 54033 52445 54067 52479
rect 54067 52445 54076 52479
rect 54024 52436 54076 52445
rect 1492 52300 1544 52352
rect 2780 52368 2832 52420
rect 54300 52368 54352 52420
rect 2872 52300 2924 52352
rect 14280 52343 14332 52352
rect 14280 52309 14289 52343
rect 14289 52309 14323 52343
rect 14323 52309 14332 52343
rect 14280 52300 14332 52309
rect 25504 52300 25556 52352
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 2780 52096 2832 52148
rect 24492 52096 24544 52148
rect 2596 52028 2648 52080
rect 1676 52003 1728 52012
rect 1676 51969 1685 52003
rect 1685 51969 1719 52003
rect 1719 51969 1728 52003
rect 1676 51960 1728 51969
rect 26056 52096 26108 52148
rect 46020 52096 46072 52148
rect 51448 52139 51500 52148
rect 51448 52105 51457 52139
rect 51457 52105 51491 52139
rect 51491 52105 51500 52139
rect 51448 52096 51500 52105
rect 54300 52139 54352 52148
rect 54300 52105 54309 52139
rect 54309 52105 54343 52139
rect 54343 52105 54352 52139
rect 54300 52096 54352 52105
rect 25412 52071 25464 52080
rect 25412 52037 25421 52071
rect 25421 52037 25455 52071
rect 25455 52037 25464 52071
rect 25412 52028 25464 52037
rect 27160 52028 27212 52080
rect 28080 52028 28132 52080
rect 25504 52003 25556 52012
rect 25504 51969 25513 52003
rect 25513 51969 25547 52003
rect 25547 51969 25556 52003
rect 25504 51960 25556 51969
rect 9312 51892 9364 51944
rect 27896 52003 27948 52012
rect 27896 51969 27905 52003
rect 27905 51969 27939 52003
rect 27939 51969 27948 52003
rect 27896 51960 27948 51969
rect 1860 51867 1912 51876
rect 1860 51833 1869 51867
rect 1869 51833 1903 51867
rect 1903 51833 1912 51867
rect 1860 51824 1912 51833
rect 32680 51824 32732 51876
rect 49516 51824 49568 51876
rect 27620 51756 27672 51808
rect 29828 51756 29880 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 2872 51595 2924 51604
rect 2872 51561 2881 51595
rect 2881 51561 2915 51595
rect 2915 51561 2924 51595
rect 2872 51552 2924 51561
rect 25504 51552 25556 51604
rect 27896 51552 27948 51604
rect 29644 51552 29696 51604
rect 1676 51323 1728 51332
rect 1676 51289 1685 51323
rect 1685 51289 1719 51323
rect 1719 51289 1728 51323
rect 1676 51280 1728 51289
rect 54392 51280 54444 51332
rect 2688 51212 2740 51264
rect 26056 51255 26108 51264
rect 26056 51221 26065 51255
rect 26065 51221 26099 51255
rect 26099 51221 26108 51255
rect 26056 51212 26108 51221
rect 54300 51255 54352 51264
rect 54300 51221 54309 51255
rect 54309 51221 54343 51255
rect 54343 51221 54352 51255
rect 54300 51212 54352 51221
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 54392 50872 54444 50924
rect 2320 50804 2372 50856
rect 2780 50804 2832 50856
rect 53564 50711 53616 50720
rect 53564 50677 53573 50711
rect 53573 50677 53607 50711
rect 53607 50677 53616 50711
rect 53564 50668 53616 50677
rect 53932 50668 53984 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 16028 50396 16080 50448
rect 25136 50396 25188 50448
rect 52276 50396 52328 50448
rect 8208 50328 8260 50380
rect 25412 50328 25464 50380
rect 29920 50328 29972 50380
rect 45468 50328 45520 50380
rect 2136 50303 2188 50312
rect 2136 50269 2145 50303
rect 2145 50269 2179 50303
rect 2179 50269 2188 50303
rect 2136 50260 2188 50269
rect 2780 50260 2832 50312
rect 54300 50303 54352 50312
rect 54300 50269 54309 50303
rect 54309 50269 54343 50303
rect 54343 50269 54352 50303
rect 54300 50260 54352 50269
rect 54484 50192 54536 50244
rect 53104 50167 53156 50176
rect 53104 50133 53113 50167
rect 53113 50133 53147 50167
rect 53147 50133 53156 50167
rect 53104 50124 53156 50133
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 48136 49852 48188 49904
rect 1676 49827 1728 49836
rect 1676 49793 1685 49827
rect 1685 49793 1719 49827
rect 1719 49793 1728 49827
rect 1676 49784 1728 49793
rect 53656 49827 53708 49836
rect 53656 49793 53665 49827
rect 53665 49793 53699 49827
rect 53699 49793 53708 49827
rect 53656 49784 53708 49793
rect 54484 49784 54536 49836
rect 2044 49716 2096 49768
rect 51172 49716 51224 49768
rect 52920 49623 52972 49632
rect 52920 49589 52929 49623
rect 52929 49589 52963 49623
rect 52963 49589 52972 49623
rect 52920 49580 52972 49589
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 2320 49172 2372 49224
rect 2780 49172 2832 49224
rect 38660 49172 38712 49224
rect 52644 49172 52696 49224
rect 53104 49172 53156 49224
rect 53564 49172 53616 49224
rect 52368 49104 52420 49156
rect 32864 49036 32916 49088
rect 33508 49036 33560 49088
rect 52460 49036 52512 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 52184 48832 52236 48884
rect 53472 48764 53524 48816
rect 52368 48739 52420 48748
rect 52368 48705 52377 48739
rect 52377 48705 52411 48739
rect 52411 48705 52420 48739
rect 52368 48696 52420 48705
rect 2228 48628 2280 48680
rect 2780 48628 2832 48680
rect 38752 48628 38804 48680
rect 53472 48671 53524 48680
rect 53472 48637 53481 48671
rect 53481 48637 53515 48671
rect 53515 48637 53524 48671
rect 53472 48628 53524 48637
rect 32864 48560 32916 48612
rect 2136 48492 2188 48544
rect 33140 48492 33192 48544
rect 33232 48535 33284 48544
rect 33232 48501 33241 48535
rect 33241 48501 33275 48535
rect 33275 48501 33284 48535
rect 33232 48492 33284 48501
rect 34060 48492 34112 48544
rect 34428 48535 34480 48544
rect 34428 48501 34437 48535
rect 34437 48501 34471 48535
rect 34471 48501 34480 48535
rect 34428 48492 34480 48501
rect 35624 48492 35676 48544
rect 51264 48492 51316 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 31116 48220 31168 48272
rect 33416 48220 33468 48272
rect 38844 48220 38896 48272
rect 51264 48220 51316 48272
rect 2780 48084 2832 48136
rect 30472 48016 30524 48068
rect 2688 47948 2740 48000
rect 52828 48152 52880 48204
rect 33416 48127 33468 48136
rect 31852 47991 31904 48000
rect 31852 47957 31861 47991
rect 31861 47957 31895 47991
rect 31895 47957 31904 47991
rect 31852 47948 31904 47957
rect 33416 48093 33425 48127
rect 33425 48093 33459 48127
rect 33459 48093 33468 48127
rect 33416 48084 33468 48093
rect 33508 48084 33560 48136
rect 33968 48084 34020 48136
rect 33232 48016 33284 48068
rect 51816 48084 51868 48136
rect 52184 48127 52236 48136
rect 52184 48093 52193 48127
rect 52193 48093 52227 48127
rect 52227 48093 52236 48127
rect 52184 48084 52236 48093
rect 52644 48127 52696 48136
rect 52644 48093 52653 48127
rect 52653 48093 52687 48127
rect 52687 48093 52696 48127
rect 52644 48084 52696 48093
rect 51356 48016 51408 48068
rect 34152 47948 34204 48000
rect 34888 47991 34940 48000
rect 34888 47957 34897 47991
rect 34897 47957 34931 47991
rect 34931 47957 34940 47991
rect 34888 47948 34940 47957
rect 51264 47948 51316 48000
rect 51632 47948 51684 48000
rect 52000 47991 52052 48000
rect 52000 47957 52009 47991
rect 52009 47957 52043 47991
rect 52043 47957 52052 47991
rect 52000 47948 52052 47957
rect 53012 47948 53064 48000
rect 53196 47948 53248 48000
rect 53840 47991 53892 48000
rect 53840 47957 53849 47991
rect 53849 47957 53883 47991
rect 53883 47957 53892 47991
rect 53840 47948 53892 47957
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 29644 47787 29696 47796
rect 29644 47753 29653 47787
rect 29653 47753 29687 47787
rect 29687 47753 29696 47787
rect 29644 47744 29696 47753
rect 33324 47744 33376 47796
rect 32772 47676 32824 47728
rect 33232 47676 33284 47728
rect 35348 47744 35400 47796
rect 35440 47744 35492 47796
rect 52000 47744 52052 47796
rect 52092 47744 52144 47796
rect 29092 47608 29144 47660
rect 2780 47540 2832 47592
rect 33140 47651 33192 47660
rect 33140 47617 33150 47651
rect 33150 47617 33184 47651
rect 33184 47617 33192 47651
rect 38936 47676 38988 47728
rect 51724 47676 51776 47728
rect 52828 47676 52880 47728
rect 33140 47608 33192 47617
rect 33508 47608 33560 47660
rect 34060 47608 34112 47660
rect 34520 47651 34572 47660
rect 34520 47617 34529 47651
rect 34529 47617 34563 47651
rect 34563 47617 34572 47651
rect 34520 47608 34572 47617
rect 2320 47472 2372 47524
rect 32036 47472 32088 47524
rect 33876 47472 33928 47524
rect 34244 47472 34296 47524
rect 35440 47472 35492 47524
rect 51448 47608 51500 47660
rect 51264 47540 51316 47592
rect 52276 47608 52328 47660
rect 53288 47540 53340 47592
rect 53564 47540 53616 47592
rect 51172 47472 51224 47524
rect 51356 47515 51408 47524
rect 51356 47481 51365 47515
rect 51365 47481 51399 47515
rect 51399 47481 51408 47515
rect 51356 47472 51408 47481
rect 51816 47515 51868 47524
rect 51816 47481 51825 47515
rect 51825 47481 51859 47515
rect 51859 47481 51868 47515
rect 51816 47472 51868 47481
rect 52736 47472 52788 47524
rect 28264 47404 28316 47456
rect 31116 47404 31168 47456
rect 31668 47447 31720 47456
rect 31668 47413 31677 47447
rect 31677 47413 31711 47447
rect 31711 47413 31720 47447
rect 31668 47404 31720 47413
rect 32404 47404 32456 47456
rect 33692 47447 33744 47456
rect 33692 47413 33701 47447
rect 33701 47413 33735 47447
rect 33735 47413 33744 47447
rect 33692 47404 33744 47413
rect 34060 47404 34112 47456
rect 34888 47404 34940 47456
rect 35808 47447 35860 47456
rect 35808 47413 35817 47447
rect 35817 47413 35851 47447
rect 35851 47413 35860 47447
rect 35808 47404 35860 47413
rect 51724 47404 51776 47456
rect 53564 47404 53616 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 29092 47243 29144 47252
rect 29092 47209 29101 47243
rect 29101 47209 29135 47243
rect 29135 47209 29144 47243
rect 29092 47200 29144 47209
rect 31852 47200 31904 47252
rect 2688 47064 2740 47116
rect 2780 46996 2832 47048
rect 31300 47132 31352 47184
rect 29644 47064 29696 47116
rect 30104 47039 30156 47048
rect 30104 47005 30113 47039
rect 30113 47005 30147 47039
rect 30147 47005 30156 47039
rect 30104 46996 30156 47005
rect 31208 47039 31260 47048
rect 30012 46971 30064 46980
rect 30012 46937 30021 46971
rect 30021 46937 30055 46971
rect 30055 46937 30064 46971
rect 30012 46928 30064 46937
rect 30472 46928 30524 46980
rect 31208 47005 31217 47039
rect 31217 47005 31251 47039
rect 31251 47005 31260 47039
rect 31208 46996 31260 47005
rect 31668 46996 31720 47048
rect 32036 47039 32088 47048
rect 32036 47005 32046 47039
rect 32046 47005 32080 47039
rect 32080 47005 32088 47039
rect 32588 47064 32640 47116
rect 32036 46996 32088 47005
rect 32404 46996 32456 47048
rect 33508 47064 33560 47116
rect 33784 47175 33836 47184
rect 33784 47141 33793 47175
rect 33793 47141 33827 47175
rect 33827 47141 33836 47175
rect 33784 47132 33836 47141
rect 35808 47132 35860 47184
rect 51540 47132 51592 47184
rect 53656 47132 53708 47184
rect 53840 47064 53892 47116
rect 33140 47039 33192 47048
rect 33140 47005 33149 47039
rect 33149 47005 33183 47039
rect 33183 47005 33192 47039
rect 33140 46996 33192 47005
rect 33324 47039 33376 47048
rect 33324 47005 33331 47039
rect 33331 47005 33376 47039
rect 33324 46996 33376 47005
rect 34060 46996 34112 47048
rect 34428 46996 34480 47048
rect 48228 46996 48280 47048
rect 50896 47039 50948 47048
rect 50896 47005 50905 47039
rect 50905 47005 50939 47039
rect 50939 47005 50948 47039
rect 50896 46996 50948 47005
rect 31116 46971 31168 46980
rect 31116 46937 31125 46971
rect 31125 46937 31159 46971
rect 31159 46937 31168 46971
rect 31116 46928 31168 46937
rect 30932 46860 30984 46912
rect 33232 46860 33284 46912
rect 34704 46928 34756 46980
rect 51448 46928 51500 46980
rect 33600 46860 33652 46912
rect 34520 46860 34572 46912
rect 51264 46860 51316 46912
rect 51908 46996 51960 47048
rect 52460 46996 52512 47048
rect 52828 47039 52880 47048
rect 51816 46971 51868 46980
rect 51816 46937 51825 46971
rect 51825 46937 51859 46971
rect 51859 46937 51868 46971
rect 51816 46928 51868 46937
rect 52092 46928 52144 46980
rect 52828 47005 52837 47039
rect 52837 47005 52871 47039
rect 52871 47005 52880 47039
rect 52828 46996 52880 47005
rect 53012 47039 53064 47048
rect 53012 47005 53021 47039
rect 53021 47005 53055 47039
rect 53055 47005 53064 47039
rect 53012 46996 53064 47005
rect 53656 46996 53708 47048
rect 52920 46928 52972 46980
rect 54116 46928 54168 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 30472 46699 30524 46708
rect 30472 46665 30481 46699
rect 30481 46665 30515 46699
rect 30515 46665 30524 46699
rect 30472 46656 30524 46665
rect 30012 46588 30064 46640
rect 2596 46520 2648 46572
rect 32772 46588 32824 46640
rect 2780 46452 2832 46504
rect 33324 46520 33376 46572
rect 34244 46656 34296 46708
rect 34336 46656 34388 46708
rect 47032 46588 47084 46640
rect 33968 46563 34020 46572
rect 33968 46529 33977 46563
rect 33977 46529 34011 46563
rect 34011 46529 34020 46563
rect 33968 46520 34020 46529
rect 34244 46520 34296 46572
rect 2228 46384 2280 46436
rect 31208 46359 31260 46368
rect 31208 46325 31217 46359
rect 31217 46325 31251 46359
rect 31251 46325 31260 46359
rect 33968 46384 34020 46436
rect 31208 46316 31260 46325
rect 33048 46316 33100 46368
rect 33416 46316 33468 46368
rect 51080 46452 51132 46504
rect 53472 46495 53524 46504
rect 53472 46461 53481 46495
rect 53481 46461 53515 46495
rect 53515 46461 53524 46495
rect 53472 46452 53524 46461
rect 48136 46316 48188 46368
rect 51264 46316 51316 46368
rect 53012 46359 53064 46368
rect 53012 46325 53021 46359
rect 53021 46325 53055 46359
rect 53055 46325 53064 46359
rect 53012 46316 53064 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 33140 46112 33192 46164
rect 35624 46112 35676 46164
rect 2412 46044 2464 46096
rect 31392 46087 31444 46096
rect 31392 46053 31401 46087
rect 31401 46053 31435 46087
rect 31435 46053 31444 46087
rect 31392 46044 31444 46053
rect 34244 46044 34296 46096
rect 2320 45908 2372 45960
rect 2780 45908 2832 45960
rect 26792 45840 26844 45892
rect 31392 45840 31444 45892
rect 32404 45951 32456 45960
rect 32404 45917 32413 45951
rect 32413 45917 32447 45951
rect 32447 45917 32456 45951
rect 32404 45908 32456 45917
rect 32772 45951 32824 45960
rect 32772 45917 32781 45951
rect 32781 45917 32815 45951
rect 32815 45917 32824 45951
rect 32772 45908 32824 45917
rect 52644 45976 52696 46028
rect 48228 45908 48280 45960
rect 52184 45951 52236 45960
rect 52184 45917 52193 45951
rect 52193 45917 52227 45951
rect 52227 45917 52236 45951
rect 52184 45908 52236 45917
rect 52552 45908 52604 45960
rect 53380 45908 53432 45960
rect 32404 45772 32456 45824
rect 33508 45815 33560 45824
rect 33508 45781 33517 45815
rect 33517 45781 33551 45815
rect 33551 45781 33560 45815
rect 33508 45772 33560 45781
rect 51264 45772 51316 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 33508 45568 33560 45620
rect 51172 45568 51224 45620
rect 26424 45500 26476 45552
rect 29644 45500 29696 45552
rect 33324 45500 33376 45552
rect 53748 45475 53800 45484
rect 2780 45364 2832 45416
rect 28540 45364 28592 45416
rect 53748 45441 53757 45475
rect 53757 45441 53791 45475
rect 53791 45441 53800 45475
rect 53748 45432 53800 45441
rect 22192 45296 22244 45348
rect 53564 45364 53616 45416
rect 31852 45228 31904 45280
rect 32772 45228 32824 45280
rect 53012 45271 53064 45280
rect 53012 45237 53021 45271
rect 53021 45237 53055 45271
rect 53055 45237 53064 45271
rect 53012 45228 53064 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 27436 45067 27488 45076
rect 27436 45033 27445 45067
rect 27445 45033 27479 45067
rect 27479 45033 27488 45067
rect 27436 45024 27488 45033
rect 31208 45024 31260 45076
rect 28632 44956 28684 45008
rect 52920 44956 52972 45008
rect 52460 44931 52512 44940
rect 52460 44897 52469 44931
rect 52469 44897 52503 44931
rect 52503 44897 52512 44931
rect 52460 44888 52512 44897
rect 2780 44820 2832 44872
rect 28356 44820 28408 44872
rect 47032 44820 47084 44872
rect 52184 44863 52236 44872
rect 52184 44829 52193 44863
rect 52193 44829 52227 44863
rect 52227 44829 52236 44863
rect 52184 44820 52236 44829
rect 22928 44752 22980 44804
rect 53656 44820 53708 44872
rect 53748 44863 53800 44872
rect 53748 44829 53757 44863
rect 53757 44829 53791 44863
rect 53791 44829 53800 44863
rect 53748 44820 53800 44829
rect 26884 44727 26936 44736
rect 26884 44693 26893 44727
rect 26893 44693 26927 44727
rect 26927 44693 26936 44727
rect 26884 44684 26936 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 28632 44523 28684 44532
rect 28632 44489 28641 44523
rect 28641 44489 28675 44523
rect 28675 44489 28684 44523
rect 28632 44480 28684 44489
rect 53472 44480 53524 44532
rect 22284 44412 22336 44464
rect 27068 44412 27120 44464
rect 27436 44412 27488 44464
rect 26424 44344 26476 44396
rect 26884 44344 26936 44396
rect 52644 44412 52696 44464
rect 53104 44344 53156 44396
rect 2228 44276 2280 44328
rect 2780 44276 2832 44328
rect 10416 44276 10468 44328
rect 27804 44276 27856 44328
rect 52092 44319 52144 44328
rect 52092 44285 52101 44319
rect 52101 44285 52135 44319
rect 52135 44285 52144 44319
rect 52092 44276 52144 44285
rect 53472 44319 53524 44328
rect 24768 44208 24820 44260
rect 32312 44251 32364 44260
rect 32312 44217 32321 44251
rect 32321 44217 32355 44251
rect 32355 44217 32364 44251
rect 32312 44208 32364 44217
rect 53472 44285 53481 44319
rect 53481 44285 53515 44319
rect 53515 44285 53524 44319
rect 53472 44276 53524 44285
rect 27988 44183 28040 44192
rect 27988 44149 27997 44183
rect 27997 44149 28031 44183
rect 28031 44149 28040 44183
rect 27988 44140 28040 44149
rect 30840 44140 30892 44192
rect 31024 44183 31076 44192
rect 31024 44149 31033 44183
rect 31033 44149 31067 44183
rect 31067 44149 31076 44183
rect 31024 44140 31076 44149
rect 32772 44140 32824 44192
rect 53012 44183 53064 44192
rect 53012 44149 53021 44183
rect 53021 44149 53055 44183
rect 53055 44149 53064 44183
rect 53012 44140 53064 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 32956 43936 33008 43988
rect 12808 43868 12860 43920
rect 30012 43868 30064 43920
rect 51356 43868 51408 43920
rect 53748 43868 53800 43920
rect 2320 43800 2372 43852
rect 2136 43775 2188 43784
rect 2136 43741 2145 43775
rect 2145 43741 2179 43775
rect 2179 43741 2188 43775
rect 2136 43732 2188 43741
rect 2780 43732 2832 43784
rect 25320 43596 25372 43648
rect 27436 43775 27488 43784
rect 27436 43741 27445 43775
rect 27445 43741 27479 43775
rect 27479 43741 27488 43775
rect 28632 43800 28684 43852
rect 27436 43732 27488 43741
rect 28080 43732 28132 43784
rect 52736 43800 52788 43852
rect 28908 43664 28960 43716
rect 30472 43664 30524 43716
rect 26608 43596 26660 43648
rect 29000 43639 29052 43648
rect 29000 43605 29009 43639
rect 29009 43605 29043 43639
rect 29043 43605 29052 43639
rect 29000 43596 29052 43605
rect 30564 43596 30616 43648
rect 31944 43639 31996 43648
rect 31944 43605 31953 43639
rect 31953 43605 31987 43639
rect 31987 43605 31996 43639
rect 31944 43596 31996 43605
rect 32680 43596 32732 43648
rect 32772 43596 32824 43648
rect 33600 43596 33652 43648
rect 33968 43596 34020 43648
rect 52920 43707 52972 43716
rect 52920 43673 52929 43707
rect 52929 43673 52963 43707
rect 52963 43673 52972 43707
rect 52920 43664 52972 43673
rect 52552 43596 52604 43648
rect 52828 43639 52880 43648
rect 52828 43605 52837 43639
rect 52837 43605 52871 43639
rect 52871 43605 52880 43639
rect 52828 43596 52880 43605
rect 53564 43732 53616 43784
rect 53748 43596 53800 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 1860 43324 1912 43376
rect 32680 43392 32732 43444
rect 34612 43435 34664 43444
rect 34612 43401 34621 43435
rect 34621 43401 34655 43435
rect 34655 43401 34664 43435
rect 34612 43392 34664 43401
rect 25412 43367 25464 43376
rect 25412 43333 25421 43367
rect 25421 43333 25455 43367
rect 25455 43333 25464 43367
rect 25412 43324 25464 43333
rect 26056 43367 26108 43376
rect 26056 43333 26065 43367
rect 26065 43333 26099 43367
rect 26099 43333 26108 43367
rect 26056 43324 26108 43333
rect 26792 43324 26844 43376
rect 27252 43324 27304 43376
rect 28264 43367 28316 43376
rect 28264 43333 28273 43367
rect 28273 43333 28307 43367
rect 28307 43333 28316 43367
rect 28264 43324 28316 43333
rect 29184 43324 29236 43376
rect 52092 43392 52144 43444
rect 2504 43256 2556 43308
rect 2688 43256 2740 43308
rect 29000 43256 29052 43308
rect 32036 43256 32088 43308
rect 32588 43256 32640 43308
rect 2780 43188 2832 43240
rect 29644 43231 29696 43240
rect 29644 43197 29653 43231
rect 29653 43197 29687 43231
rect 29687 43197 29696 43231
rect 29644 43188 29696 43197
rect 32404 43231 32456 43240
rect 32404 43197 32413 43231
rect 32413 43197 32447 43231
rect 32447 43197 32456 43231
rect 53564 43256 53616 43308
rect 32404 43188 32456 43197
rect 53656 43188 53708 43240
rect 1768 43120 1820 43172
rect 32588 43120 32640 43172
rect 52644 43120 52696 43172
rect 27712 43052 27764 43104
rect 28448 43052 28500 43104
rect 29092 43095 29144 43104
rect 29092 43061 29101 43095
rect 29101 43061 29135 43095
rect 29135 43061 29144 43095
rect 29092 43052 29144 43061
rect 30196 43095 30248 43104
rect 30196 43061 30205 43095
rect 30205 43061 30239 43095
rect 30239 43061 30248 43095
rect 30196 43052 30248 43061
rect 30748 43095 30800 43104
rect 30748 43061 30757 43095
rect 30757 43061 30791 43095
rect 30791 43061 30800 43095
rect 30748 43052 30800 43061
rect 31484 43052 31536 43104
rect 34336 43052 34388 43104
rect 35440 43052 35492 43104
rect 53380 43052 53432 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 26056 42848 26108 42900
rect 30748 42848 30800 42900
rect 52552 42848 52604 42900
rect 25780 42780 25832 42832
rect 27896 42780 27948 42832
rect 30564 42780 30616 42832
rect 2596 42712 2648 42764
rect 25872 42712 25924 42764
rect 26424 42712 26476 42764
rect 28356 42755 28408 42764
rect 28356 42721 28365 42755
rect 28365 42721 28399 42755
rect 28399 42721 28408 42755
rect 28356 42712 28408 42721
rect 29644 42712 29696 42764
rect 2780 42644 2832 42696
rect 23848 42644 23900 42696
rect 26240 42644 26292 42696
rect 28448 42644 28500 42696
rect 30840 42712 30892 42764
rect 32312 42712 32364 42764
rect 23388 42576 23440 42628
rect 26332 42576 26384 42628
rect 28264 42576 28316 42628
rect 29460 42576 29512 42628
rect 30012 42687 30064 42696
rect 30012 42653 30021 42687
rect 30021 42653 30055 42687
rect 30055 42653 30064 42687
rect 30288 42687 30340 42696
rect 30012 42644 30064 42653
rect 30288 42653 30297 42687
rect 30297 42653 30331 42687
rect 30331 42653 30340 42687
rect 30288 42644 30340 42653
rect 32496 42687 32548 42696
rect 32496 42653 32505 42687
rect 32505 42653 32539 42687
rect 32539 42653 32548 42687
rect 32496 42644 32548 42653
rect 32864 42687 32916 42696
rect 32864 42653 32873 42687
rect 32873 42653 32907 42687
rect 32907 42653 32916 42687
rect 32864 42644 32916 42653
rect 35532 42712 35584 42764
rect 53748 42755 53800 42764
rect 53748 42721 53757 42755
rect 53757 42721 53791 42755
rect 53791 42721 53800 42755
rect 53748 42712 53800 42721
rect 32772 42619 32824 42628
rect 32772 42585 32781 42619
rect 32781 42585 32815 42619
rect 32815 42585 32824 42619
rect 32772 42576 32824 42585
rect 26792 42508 26844 42560
rect 27896 42508 27948 42560
rect 29552 42508 29604 42560
rect 30288 42508 30340 42560
rect 30840 42551 30892 42560
rect 30840 42517 30849 42551
rect 30849 42517 30883 42551
rect 30883 42517 30892 42551
rect 30840 42508 30892 42517
rect 31576 42508 31628 42560
rect 33140 42644 33192 42696
rect 52368 42644 52420 42696
rect 53472 42687 53524 42696
rect 53472 42653 53481 42687
rect 53481 42653 53515 42687
rect 53515 42653 53524 42687
rect 53472 42644 53524 42653
rect 33600 42619 33652 42628
rect 33600 42585 33609 42619
rect 33609 42585 33643 42619
rect 33643 42585 33652 42619
rect 33600 42576 33652 42585
rect 34060 42576 34112 42628
rect 34244 42576 34296 42628
rect 34796 42576 34848 42628
rect 33508 42508 33560 42560
rect 33968 42508 34020 42560
rect 35532 42551 35584 42560
rect 35532 42517 35541 42551
rect 35541 42517 35575 42551
rect 35575 42517 35584 42551
rect 35532 42508 35584 42517
rect 52368 42551 52420 42560
rect 52368 42517 52377 42551
rect 52377 42517 52411 42551
rect 52411 42517 52420 42551
rect 52368 42508 52420 42517
rect 52460 42508 52512 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 25412 42304 25464 42356
rect 24860 42211 24912 42220
rect 24860 42177 24869 42211
rect 24869 42177 24903 42211
rect 24903 42177 24912 42211
rect 24860 42168 24912 42177
rect 25596 42236 25648 42288
rect 26056 42236 26108 42288
rect 29184 42304 29236 42356
rect 29460 42304 29512 42356
rect 30288 42304 30340 42356
rect 2320 42100 2372 42152
rect 2780 42100 2832 42152
rect 24216 42100 24268 42152
rect 23848 42007 23900 42016
rect 23848 41973 23857 42007
rect 23857 41973 23891 42007
rect 23891 41973 23900 42007
rect 23848 41964 23900 41973
rect 26332 42168 26384 42220
rect 27712 42168 27764 42220
rect 27988 42168 28040 42220
rect 28172 42168 28224 42220
rect 29000 42236 29052 42288
rect 30380 42279 30432 42288
rect 30380 42245 30389 42279
rect 30389 42245 30423 42279
rect 30423 42245 30432 42279
rect 30380 42236 30432 42245
rect 31392 42304 31444 42356
rect 31944 42304 31996 42356
rect 28632 42168 28684 42220
rect 28816 42211 28868 42220
rect 28816 42177 28825 42211
rect 28825 42177 28859 42211
rect 28859 42177 28868 42211
rect 28816 42168 28868 42177
rect 30564 42168 30616 42220
rect 32404 42236 32456 42288
rect 32864 42279 32916 42288
rect 32864 42245 32873 42279
rect 32873 42245 32907 42279
rect 32907 42245 32916 42279
rect 32864 42236 32916 42245
rect 33600 42304 33652 42356
rect 28908 42100 28960 42152
rect 32588 42211 32640 42220
rect 32588 42177 32598 42211
rect 32598 42177 32632 42211
rect 32632 42177 32640 42211
rect 32772 42211 32824 42220
rect 32588 42168 32640 42177
rect 32772 42177 32781 42211
rect 32781 42177 32815 42211
rect 32815 42177 32824 42211
rect 32772 42168 32824 42177
rect 31208 42100 31260 42152
rect 31576 42100 31628 42152
rect 33508 42236 33560 42288
rect 34796 42304 34848 42356
rect 35532 42304 35584 42356
rect 35440 42236 35492 42288
rect 33232 42168 33284 42220
rect 33968 42211 34020 42220
rect 33968 42177 33977 42211
rect 33977 42177 34011 42211
rect 34011 42177 34020 42211
rect 33968 42168 34020 42177
rect 38660 42304 38712 42356
rect 52552 42168 52604 42220
rect 53472 42143 53524 42152
rect 27436 42032 27488 42084
rect 29644 42032 29696 42084
rect 30196 42032 30248 42084
rect 33324 42032 33376 42084
rect 33508 42032 33560 42084
rect 53472 42109 53481 42143
rect 53481 42109 53515 42143
rect 53515 42109 53524 42143
rect 53472 42100 53524 42109
rect 34704 42075 34756 42084
rect 34704 42041 34713 42075
rect 34713 42041 34747 42075
rect 34747 42041 34756 42075
rect 34704 42032 34756 42041
rect 48044 42032 48096 42084
rect 54300 42032 54352 42084
rect 26516 42007 26568 42016
rect 26516 41973 26525 42007
rect 26525 41973 26559 42007
rect 26559 41973 26568 42007
rect 26516 41964 26568 41973
rect 27528 41964 27580 42016
rect 27988 41964 28040 42016
rect 28264 42007 28316 42016
rect 28264 41973 28273 42007
rect 28273 41973 28307 42007
rect 28307 41973 28316 42007
rect 28264 41964 28316 41973
rect 30012 41964 30064 42016
rect 31944 41964 31996 42016
rect 32588 41964 32640 42016
rect 32772 41964 32824 42016
rect 32864 41964 32916 42016
rect 34612 41964 34664 42016
rect 35348 41964 35400 42016
rect 52276 42007 52328 42016
rect 52276 41973 52285 42007
rect 52285 41973 52319 42007
rect 52319 41973 52328 42007
rect 52276 41964 52328 41973
rect 53012 42007 53064 42016
rect 53012 41973 53021 42007
rect 53021 41973 53055 42007
rect 53055 41973 53064 42007
rect 53012 41964 53064 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 24860 41760 24912 41812
rect 25044 41692 25096 41744
rect 26792 41692 26844 41744
rect 27988 41760 28040 41812
rect 28540 41760 28592 41812
rect 29828 41692 29880 41744
rect 24492 41624 24544 41676
rect 25872 41624 25924 41676
rect 26148 41624 26200 41676
rect 28816 41624 28868 41676
rect 29460 41624 29512 41676
rect 30104 41624 30156 41676
rect 2780 41556 2832 41608
rect 26884 41556 26936 41608
rect 27252 41599 27304 41608
rect 27252 41565 27261 41599
rect 27261 41565 27295 41599
rect 27295 41565 27304 41599
rect 27252 41556 27304 41565
rect 24676 41531 24728 41540
rect 24676 41497 24685 41531
rect 24685 41497 24719 41531
rect 24719 41497 24728 41531
rect 24676 41488 24728 41497
rect 25412 41488 25464 41540
rect 27804 41599 27856 41608
rect 27804 41565 27814 41599
rect 27814 41565 27848 41599
rect 27848 41565 27856 41599
rect 28080 41599 28132 41608
rect 27804 41556 27856 41565
rect 28080 41565 28089 41599
rect 28089 41565 28123 41599
rect 28123 41565 28132 41599
rect 28080 41556 28132 41565
rect 28448 41556 28500 41608
rect 29276 41556 29328 41608
rect 27988 41531 28040 41540
rect 27988 41497 27997 41531
rect 27997 41497 28031 41531
rect 28031 41497 28040 41531
rect 27988 41488 28040 41497
rect 24400 41420 24452 41472
rect 24952 41463 25004 41472
rect 24952 41429 24961 41463
rect 24961 41429 24995 41463
rect 24995 41429 25004 41463
rect 24952 41420 25004 41429
rect 27252 41420 27304 41472
rect 29736 41463 29788 41472
rect 29736 41429 29745 41463
rect 29745 41429 29779 41463
rect 29779 41429 29788 41463
rect 29736 41420 29788 41429
rect 30104 41531 30156 41540
rect 30104 41497 30113 41531
rect 30113 41497 30147 41531
rect 30147 41497 30156 41531
rect 30104 41488 30156 41497
rect 30564 41556 30616 41608
rect 32036 41760 32088 41812
rect 32496 41760 32548 41812
rect 35348 41760 35400 41812
rect 31208 41624 31260 41676
rect 31392 41599 31444 41608
rect 31392 41565 31400 41599
rect 31400 41565 31434 41599
rect 31434 41565 31444 41599
rect 31392 41556 31444 41565
rect 32588 41599 32640 41608
rect 32588 41565 32592 41599
rect 32592 41565 32626 41599
rect 32626 41565 32640 41599
rect 32588 41556 32640 41565
rect 32680 41599 32732 41608
rect 32680 41565 32689 41599
rect 32689 41565 32723 41599
rect 32723 41565 32732 41599
rect 33324 41624 33376 41676
rect 32680 41556 32732 41565
rect 33876 41692 33928 41744
rect 34336 41692 34388 41744
rect 53288 41692 53340 41744
rect 33600 41556 33652 41608
rect 30472 41488 30524 41540
rect 33232 41488 33284 41540
rect 33876 41531 33928 41540
rect 33876 41497 33885 41531
rect 33885 41497 33919 41531
rect 33919 41497 33928 41531
rect 33876 41488 33928 41497
rect 34796 41556 34848 41608
rect 36268 41556 36320 41608
rect 36820 41624 36872 41676
rect 38752 41624 38804 41676
rect 52460 41624 52512 41676
rect 52368 41599 52420 41608
rect 52368 41565 52377 41599
rect 52377 41565 52411 41599
rect 52411 41565 52420 41599
rect 52368 41556 52420 41565
rect 53012 41599 53064 41608
rect 53012 41565 53021 41599
rect 53021 41565 53055 41599
rect 53055 41565 53064 41599
rect 53012 41556 53064 41565
rect 33324 41420 33376 41472
rect 34060 41420 34112 41472
rect 35440 41488 35492 41540
rect 35348 41420 35400 41472
rect 35624 41420 35676 41472
rect 36268 41420 36320 41472
rect 36820 41463 36872 41472
rect 36820 41429 36829 41463
rect 36829 41429 36863 41463
rect 36863 41429 36872 41463
rect 36820 41420 36872 41429
rect 52276 41420 52328 41472
rect 54300 41599 54352 41608
rect 54300 41565 54309 41599
rect 54309 41565 54343 41599
rect 54343 41565 54352 41599
rect 54300 41556 54352 41565
rect 53656 41420 53708 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 24492 41259 24544 41268
rect 24492 41225 24501 41259
rect 24501 41225 24535 41259
rect 24535 41225 24544 41259
rect 24492 41216 24544 41225
rect 26332 41259 26384 41268
rect 26332 41225 26341 41259
rect 26341 41225 26375 41259
rect 26375 41225 26384 41259
rect 26332 41216 26384 41225
rect 26516 41216 26568 41268
rect 24400 41148 24452 41200
rect 28632 41216 28684 41268
rect 29368 41216 29420 41268
rect 30564 41216 30616 41268
rect 32220 41216 32272 41268
rect 32680 41216 32732 41268
rect 24032 41123 24084 41132
rect 2780 41012 2832 41064
rect 24032 41089 24041 41123
rect 24041 41089 24075 41123
rect 24075 41089 24084 41123
rect 28724 41148 28776 41200
rect 32772 41148 32824 41200
rect 33232 41216 33284 41268
rect 35256 41216 35308 41268
rect 36544 41216 36596 41268
rect 50160 41216 50212 41268
rect 33692 41148 33744 41200
rect 51172 41148 51224 41200
rect 24032 41080 24084 41089
rect 26424 41080 26476 41132
rect 27068 41080 27120 41132
rect 27712 41123 27764 41132
rect 27712 41089 27721 41123
rect 27721 41089 27755 41123
rect 27755 41089 27764 41123
rect 27712 41080 27764 41089
rect 28632 41123 28684 41132
rect 25780 40944 25832 40996
rect 27436 40944 27488 40996
rect 28632 41089 28641 41123
rect 28641 41089 28675 41123
rect 28675 41089 28684 41123
rect 28632 41080 28684 41089
rect 29092 41080 29144 41132
rect 29184 41080 29236 41132
rect 28632 40944 28684 40996
rect 29276 40944 29328 40996
rect 30196 41080 30248 41132
rect 31852 41080 31904 41132
rect 30104 41012 30156 41064
rect 30748 40944 30800 40996
rect 33232 41080 33284 41132
rect 33968 41080 34020 41132
rect 35256 41123 35308 41132
rect 35256 41089 35265 41123
rect 35265 41089 35299 41123
rect 35299 41089 35308 41123
rect 35256 41080 35308 41089
rect 33876 41012 33928 41064
rect 25872 40876 25924 40928
rect 26516 40876 26568 40928
rect 27252 40876 27304 40928
rect 27712 40876 27764 40928
rect 29460 40876 29512 40928
rect 29920 40919 29972 40928
rect 29920 40885 29929 40919
rect 29929 40885 29963 40919
rect 29963 40885 29972 40919
rect 29920 40876 29972 40885
rect 30196 40876 30248 40928
rect 31760 40876 31812 40928
rect 31944 40876 31996 40928
rect 32772 40919 32824 40928
rect 32772 40885 32781 40919
rect 32781 40885 32815 40919
rect 32815 40885 32824 40919
rect 32772 40876 32824 40885
rect 33416 40944 33468 40996
rect 35900 40944 35952 40996
rect 53104 41080 53156 41132
rect 53472 41055 53524 41064
rect 53472 41021 53481 41055
rect 53481 41021 53515 41055
rect 53515 41021 53524 41055
rect 53472 41012 53524 41021
rect 54300 40944 54352 40996
rect 34244 40919 34296 40928
rect 34244 40885 34253 40919
rect 34253 40885 34287 40919
rect 34287 40885 34296 40919
rect 34244 40876 34296 40885
rect 52920 40919 52972 40928
rect 52920 40885 52929 40919
rect 52929 40885 52963 40919
rect 52963 40885 52972 40919
rect 52920 40876 52972 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 23388 40715 23440 40724
rect 23388 40681 23397 40715
rect 23397 40681 23431 40715
rect 23431 40681 23440 40715
rect 23388 40672 23440 40681
rect 2136 40511 2188 40520
rect 2136 40477 2145 40511
rect 2145 40477 2179 40511
rect 2179 40477 2188 40511
rect 2136 40468 2188 40477
rect 2780 40468 2832 40520
rect 24676 40468 24728 40520
rect 26148 40511 26200 40520
rect 26148 40477 26157 40511
rect 26157 40477 26191 40511
rect 26191 40477 26200 40511
rect 26148 40468 26200 40477
rect 26424 40511 26476 40520
rect 26424 40477 26433 40511
rect 26433 40477 26467 40511
rect 26467 40477 26476 40511
rect 26424 40468 26476 40477
rect 26516 40511 26568 40520
rect 26516 40477 26525 40511
rect 26525 40477 26559 40511
rect 26559 40477 26568 40511
rect 26516 40468 26568 40477
rect 26884 40468 26936 40520
rect 36544 40672 36596 40724
rect 27896 40647 27948 40656
rect 27896 40613 27905 40647
rect 27905 40613 27939 40647
rect 27939 40613 27948 40647
rect 27896 40604 27948 40613
rect 28816 40604 28868 40656
rect 30288 40604 30340 40656
rect 30564 40604 30616 40656
rect 24492 40400 24544 40452
rect 27528 40443 27580 40452
rect 27528 40409 27537 40443
rect 27537 40409 27571 40443
rect 27571 40409 27580 40443
rect 27528 40400 27580 40409
rect 23572 40332 23624 40384
rect 25504 40375 25556 40384
rect 25504 40341 25513 40375
rect 25513 40341 25547 40375
rect 25547 40341 25556 40375
rect 25504 40332 25556 40341
rect 25596 40332 25648 40384
rect 26148 40332 26200 40384
rect 26884 40332 26936 40384
rect 28264 40468 28316 40520
rect 28724 40536 28776 40588
rect 30104 40536 30156 40588
rect 28080 40400 28132 40452
rect 29092 40468 29144 40520
rect 33140 40604 33192 40656
rect 33232 40604 33284 40656
rect 33876 40604 33928 40656
rect 35808 40604 35860 40656
rect 51908 40672 51960 40724
rect 53196 40672 53248 40724
rect 54116 40715 54168 40724
rect 54116 40681 54125 40715
rect 54125 40681 54159 40715
rect 54159 40681 54168 40715
rect 54116 40672 54168 40681
rect 52644 40604 52696 40656
rect 32680 40536 32732 40588
rect 32220 40468 32272 40520
rect 32588 40511 32640 40520
rect 32588 40477 32592 40511
rect 32592 40477 32626 40511
rect 32626 40477 32640 40511
rect 32588 40468 32640 40477
rect 33048 40511 33100 40520
rect 33048 40477 33057 40511
rect 33057 40477 33091 40511
rect 33091 40477 33100 40511
rect 33048 40468 33100 40477
rect 33324 40468 33376 40520
rect 35348 40468 35400 40520
rect 32128 40400 32180 40452
rect 33692 40443 33744 40452
rect 33692 40409 33701 40443
rect 33701 40409 33735 40443
rect 33735 40409 33744 40443
rect 33692 40400 33744 40409
rect 34796 40400 34848 40452
rect 52368 40511 52420 40520
rect 52368 40477 52377 40511
rect 52377 40477 52411 40511
rect 52411 40477 52420 40511
rect 52368 40468 52420 40477
rect 52920 40468 52972 40520
rect 53656 40511 53708 40520
rect 53656 40477 53665 40511
rect 53665 40477 53699 40511
rect 53699 40477 53708 40511
rect 53656 40468 53708 40477
rect 54300 40511 54352 40520
rect 54300 40477 54309 40511
rect 54309 40477 54343 40511
rect 54343 40477 54352 40511
rect 54300 40468 54352 40477
rect 29092 40332 29144 40384
rect 29644 40332 29696 40384
rect 29828 40332 29880 40384
rect 32220 40332 32272 40384
rect 32404 40375 32456 40384
rect 32404 40341 32413 40375
rect 32413 40341 32447 40375
rect 32447 40341 32456 40375
rect 32404 40332 32456 40341
rect 32496 40332 32548 40384
rect 33600 40332 33652 40384
rect 33876 40375 33928 40384
rect 33876 40341 33885 40375
rect 33885 40341 33919 40375
rect 33919 40341 33928 40375
rect 33876 40332 33928 40341
rect 34612 40332 34664 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 24400 40171 24452 40180
rect 24400 40137 24409 40171
rect 24409 40137 24443 40171
rect 24443 40137 24452 40171
rect 24400 40128 24452 40137
rect 25044 40171 25096 40180
rect 25044 40137 25053 40171
rect 25053 40137 25087 40171
rect 25087 40137 25096 40171
rect 25044 40128 25096 40137
rect 25504 40128 25556 40180
rect 26240 40128 26292 40180
rect 26700 40128 26752 40180
rect 23388 39992 23440 40044
rect 23848 40035 23900 40044
rect 23848 40001 23857 40035
rect 23857 40001 23891 40035
rect 23891 40001 23900 40035
rect 23848 39992 23900 40001
rect 2780 39924 2832 39976
rect 19340 39924 19392 39976
rect 25688 40060 25740 40112
rect 28448 40128 28500 40180
rect 28908 40128 28960 40180
rect 25044 39992 25096 40044
rect 26148 39992 26200 40044
rect 26332 39992 26384 40044
rect 26516 39992 26568 40044
rect 27804 40060 27856 40112
rect 27344 40035 27396 40044
rect 27344 40001 27351 40035
rect 27351 40001 27396 40035
rect 25780 39924 25832 39976
rect 27344 39992 27396 40001
rect 27436 40035 27488 40044
rect 27436 40001 27445 40035
rect 27445 40001 27479 40035
rect 27479 40001 27488 40035
rect 27436 39992 27488 40001
rect 28080 39992 28132 40044
rect 28172 39992 28224 40044
rect 29736 40060 29788 40112
rect 30104 40128 30156 40180
rect 32496 40128 32548 40180
rect 31300 40103 31352 40112
rect 31300 40069 31309 40103
rect 31309 40069 31343 40103
rect 31343 40069 31352 40103
rect 31300 40060 31352 40069
rect 28448 39924 28500 39976
rect 22744 39856 22796 39908
rect 17224 39788 17276 39840
rect 25228 39788 25280 39840
rect 25412 39788 25464 39840
rect 28356 39856 28408 39908
rect 29460 39924 29512 39976
rect 30564 39992 30616 40044
rect 31484 40035 31536 40044
rect 31484 40001 31493 40035
rect 31493 40001 31527 40035
rect 31527 40001 31536 40035
rect 31484 39992 31536 40001
rect 32496 40035 32548 40044
rect 32496 40001 32500 40035
rect 32500 40001 32534 40035
rect 32534 40001 32548 40035
rect 32496 39992 32548 40001
rect 33232 40060 33284 40112
rect 33508 40060 33560 40112
rect 33968 40060 34020 40112
rect 28908 39856 28960 39908
rect 30196 39924 30248 39976
rect 31852 39924 31904 39976
rect 32864 39992 32916 40044
rect 34152 40060 34204 40112
rect 30932 39856 30984 39908
rect 46112 39992 46164 40044
rect 35532 39924 35584 39976
rect 53564 39924 53616 39976
rect 36084 39856 36136 39908
rect 53656 39856 53708 39908
rect 27528 39788 27580 39840
rect 27804 39831 27856 39840
rect 27804 39797 27813 39831
rect 27813 39797 27847 39831
rect 27847 39797 27856 39831
rect 27804 39788 27856 39797
rect 29000 39788 29052 39840
rect 30472 39831 30524 39840
rect 30472 39797 30481 39831
rect 30481 39797 30515 39831
rect 30515 39797 30524 39831
rect 30472 39788 30524 39797
rect 31668 39831 31720 39840
rect 31668 39797 31677 39831
rect 31677 39797 31711 39831
rect 31711 39797 31720 39831
rect 31668 39788 31720 39797
rect 32312 39831 32364 39840
rect 32312 39797 32321 39831
rect 32321 39797 32355 39831
rect 32355 39797 32364 39831
rect 32312 39788 32364 39797
rect 32680 39788 32732 39840
rect 53380 39788 53432 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 22192 39584 22244 39636
rect 25688 39627 25740 39636
rect 24584 39516 24636 39568
rect 25320 39448 25372 39500
rect 25688 39593 25697 39627
rect 25697 39593 25731 39627
rect 25731 39593 25740 39627
rect 25688 39584 25740 39593
rect 27620 39584 27672 39636
rect 28172 39584 28224 39636
rect 31392 39584 31444 39636
rect 26240 39516 26292 39568
rect 2780 39380 2832 39432
rect 25044 39423 25096 39432
rect 25044 39389 25053 39423
rect 25053 39389 25087 39423
rect 25087 39389 25096 39423
rect 25044 39380 25096 39389
rect 22928 39312 22980 39364
rect 25228 39380 25280 39432
rect 25320 39355 25372 39364
rect 25320 39321 25329 39355
rect 25329 39321 25363 39355
rect 25363 39321 25372 39355
rect 25320 39312 25372 39321
rect 23480 39287 23532 39296
rect 23480 39253 23489 39287
rect 23489 39253 23523 39287
rect 23523 39253 23532 39287
rect 23480 39244 23532 39253
rect 23940 39287 23992 39296
rect 23940 39253 23949 39287
rect 23949 39253 23983 39287
rect 23983 39253 23992 39287
rect 23940 39244 23992 39253
rect 24308 39244 24360 39296
rect 25228 39244 25280 39296
rect 25964 39448 26016 39500
rect 26148 39423 26200 39432
rect 26148 39389 26157 39423
rect 26157 39389 26191 39423
rect 26191 39389 26200 39423
rect 26148 39380 26200 39389
rect 27252 39448 27304 39500
rect 27068 39380 27120 39432
rect 27344 39380 27396 39432
rect 27712 39423 27764 39432
rect 27712 39389 27721 39423
rect 27721 39389 27755 39423
rect 27755 39389 27764 39423
rect 27712 39380 27764 39389
rect 34428 39516 34480 39568
rect 46112 39584 46164 39636
rect 53748 39516 53800 39568
rect 28264 39380 28316 39432
rect 29092 39380 29144 39432
rect 29276 39380 29328 39432
rect 30564 39380 30616 39432
rect 32680 39448 32732 39500
rect 33600 39448 33652 39500
rect 46296 39448 46348 39500
rect 32312 39380 32364 39432
rect 32404 39380 32456 39432
rect 32864 39380 32916 39432
rect 26056 39244 26108 39296
rect 26976 39312 27028 39364
rect 26792 39287 26844 39296
rect 26792 39253 26801 39287
rect 26801 39253 26835 39287
rect 26835 39253 26844 39287
rect 26792 39244 26844 39253
rect 26884 39244 26936 39296
rect 27528 39244 27580 39296
rect 29460 39244 29512 39296
rect 29736 39287 29788 39296
rect 29736 39253 29745 39287
rect 29745 39253 29779 39287
rect 29779 39253 29788 39287
rect 29736 39244 29788 39253
rect 30748 39244 30800 39296
rect 31208 39287 31260 39296
rect 31208 39253 31217 39287
rect 31217 39253 31251 39287
rect 31251 39253 31260 39287
rect 31208 39244 31260 39253
rect 32864 39287 32916 39296
rect 32864 39253 32873 39287
rect 32873 39253 32907 39287
rect 32907 39253 32916 39287
rect 32864 39244 32916 39253
rect 33324 39287 33376 39296
rect 33324 39253 33333 39287
rect 33333 39253 33367 39287
rect 33367 39253 33376 39287
rect 33324 39244 33376 39253
rect 33784 39380 33836 39432
rect 34244 39380 34296 39432
rect 53012 39423 53064 39432
rect 53012 39389 53021 39423
rect 53021 39389 53055 39423
rect 53055 39389 53064 39423
rect 53012 39380 53064 39389
rect 53472 39423 53524 39432
rect 53472 39389 53481 39423
rect 53481 39389 53515 39423
rect 53515 39389 53524 39423
rect 53472 39380 53524 39389
rect 53656 39380 53708 39432
rect 36544 39312 36596 39364
rect 51080 39244 51132 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 11704 39040 11756 39092
rect 22928 39083 22980 39092
rect 2780 38836 2832 38888
rect 14832 38836 14884 38888
rect 17316 38904 17368 38956
rect 22928 39049 22937 39083
rect 22937 39049 22971 39083
rect 22971 39049 22980 39083
rect 22928 39040 22980 39049
rect 23572 39083 23624 39092
rect 23572 39049 23581 39083
rect 23581 39049 23615 39083
rect 23615 39049 23624 39083
rect 23572 39040 23624 39049
rect 24308 39040 24360 39092
rect 22744 38972 22796 39024
rect 24952 39040 25004 39092
rect 26056 39040 26108 39092
rect 26148 39040 26200 39092
rect 27988 39040 28040 39092
rect 28908 39040 28960 39092
rect 24584 39015 24636 39024
rect 24584 38981 24593 39015
rect 24593 38981 24627 39015
rect 24627 38981 24636 39015
rect 30656 39040 30708 39092
rect 24584 38972 24636 38981
rect 26608 38947 26660 38956
rect 26608 38913 26617 38947
rect 26617 38913 26651 38947
rect 26651 38913 26660 38947
rect 26608 38904 26660 38913
rect 27528 38947 27580 38956
rect 27528 38913 27537 38947
rect 27537 38913 27571 38947
rect 27571 38913 27580 38947
rect 27528 38904 27580 38913
rect 27620 38904 27672 38956
rect 28264 38904 28316 38956
rect 28356 38904 28408 38956
rect 28816 38947 28868 38956
rect 28816 38913 28825 38947
rect 28825 38913 28859 38947
rect 28859 38913 28868 38947
rect 28816 38904 28868 38913
rect 29644 38972 29696 39024
rect 29736 38972 29788 39024
rect 30564 38972 30616 39024
rect 31668 39015 31720 39024
rect 31668 38981 31677 39015
rect 31677 38981 31711 39015
rect 31711 38981 31720 39015
rect 31668 38972 31720 38981
rect 32772 38972 32824 39024
rect 29276 38947 29328 38956
rect 29276 38913 29290 38947
rect 29290 38913 29324 38947
rect 29324 38913 29328 38947
rect 29276 38904 29328 38913
rect 29460 38904 29512 38956
rect 33692 38972 33744 39024
rect 33876 39015 33928 39024
rect 33876 38981 33885 39015
rect 33885 38981 33919 39015
rect 33919 38981 33928 39015
rect 33876 38972 33928 38981
rect 52092 38947 52144 38956
rect 52092 38913 52101 38947
rect 52101 38913 52135 38947
rect 52135 38913 52144 38947
rect 52092 38904 52144 38913
rect 23020 38836 23072 38888
rect 29736 38836 29788 38888
rect 23940 38768 23992 38820
rect 26976 38768 27028 38820
rect 28724 38768 28776 38820
rect 24400 38700 24452 38752
rect 24860 38700 24912 38752
rect 25320 38700 25372 38752
rect 25504 38700 25556 38752
rect 25872 38700 25924 38752
rect 26056 38700 26108 38752
rect 26240 38743 26292 38752
rect 26240 38709 26249 38743
rect 26249 38709 26283 38743
rect 26283 38709 26292 38743
rect 26240 38700 26292 38709
rect 26884 38700 26936 38752
rect 27252 38700 27304 38752
rect 27988 38700 28040 38752
rect 29368 38700 29420 38752
rect 29736 38700 29788 38752
rect 29828 38700 29880 38752
rect 35992 38768 36044 38820
rect 53380 38836 53432 38888
rect 32036 38700 32088 38752
rect 32128 38700 32180 38752
rect 34520 38700 34572 38752
rect 53012 38743 53064 38752
rect 53012 38709 53021 38743
rect 53021 38709 53055 38743
rect 53055 38709 53064 38743
rect 53012 38700 53064 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 24860 38539 24912 38548
rect 24860 38505 24869 38539
rect 24869 38505 24903 38539
rect 24903 38505 24912 38539
rect 24860 38496 24912 38505
rect 27252 38496 27304 38548
rect 29460 38496 29512 38548
rect 29828 38496 29880 38548
rect 31852 38496 31904 38548
rect 26240 38428 26292 38480
rect 21916 38360 21968 38412
rect 26424 38335 26476 38344
rect 26424 38301 26433 38335
rect 26433 38301 26467 38335
rect 26467 38301 26476 38335
rect 26424 38292 26476 38301
rect 26608 38335 26660 38344
rect 26608 38301 26617 38335
rect 26617 38301 26651 38335
rect 26651 38301 26660 38335
rect 26608 38292 26660 38301
rect 26792 38335 26844 38344
rect 26792 38301 26801 38335
rect 26801 38301 26835 38335
rect 26835 38301 26844 38335
rect 26792 38292 26844 38301
rect 1676 38267 1728 38276
rect 1676 38233 1685 38267
rect 1685 38233 1719 38267
rect 1719 38233 1728 38267
rect 1676 38224 1728 38233
rect 5540 38224 5592 38276
rect 26056 38224 26108 38276
rect 26976 38224 27028 38276
rect 27436 38267 27488 38276
rect 27436 38233 27445 38267
rect 27445 38233 27479 38267
rect 27479 38233 27488 38267
rect 27436 38224 27488 38233
rect 28172 38360 28224 38412
rect 27712 38335 27764 38344
rect 27712 38301 27721 38335
rect 27721 38301 27755 38335
rect 27755 38301 27764 38335
rect 27712 38292 27764 38301
rect 28540 38428 28592 38480
rect 28954 38428 29006 38480
rect 29736 38428 29788 38480
rect 28816 38360 28868 38412
rect 29000 38292 29052 38344
rect 30932 38360 30984 38412
rect 31484 38360 31536 38412
rect 31576 38360 31628 38412
rect 32680 38360 32732 38412
rect 34428 38360 34480 38412
rect 53748 38403 53800 38412
rect 53748 38369 53757 38403
rect 53757 38369 53791 38403
rect 53791 38369 53800 38403
rect 53748 38360 53800 38369
rect 29920 38292 29972 38344
rect 31208 38292 31260 38344
rect 32864 38292 32916 38344
rect 33324 38292 33376 38344
rect 52184 38335 52236 38344
rect 52184 38301 52193 38335
rect 52193 38301 52227 38335
rect 52227 38301 52236 38335
rect 52184 38292 52236 38301
rect 28816 38224 28868 38276
rect 30104 38224 30156 38276
rect 31484 38224 31536 38276
rect 53748 38224 53800 38276
rect 4344 38156 4396 38208
rect 17316 38156 17368 38208
rect 21456 38156 21508 38208
rect 24032 38199 24084 38208
rect 24032 38165 24041 38199
rect 24041 38165 24075 38199
rect 24075 38165 24084 38199
rect 24032 38156 24084 38165
rect 25228 38156 25280 38208
rect 25872 38156 25924 38208
rect 26792 38156 26844 38208
rect 28356 38156 28408 38208
rect 28540 38156 28592 38208
rect 28724 38156 28776 38208
rect 29000 38156 29052 38208
rect 29920 38156 29972 38208
rect 30196 38199 30248 38208
rect 30196 38165 30205 38199
rect 30205 38165 30239 38199
rect 30239 38165 30248 38199
rect 30196 38156 30248 38165
rect 31668 38156 31720 38208
rect 32864 38156 32916 38208
rect 33416 38199 33468 38208
rect 33416 38165 33425 38199
rect 33425 38165 33459 38199
rect 33459 38165 33468 38199
rect 33416 38156 33468 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 25688 37952 25740 38004
rect 2136 37884 2188 37936
rect 1584 37859 1636 37868
rect 1584 37825 1593 37859
rect 1593 37825 1627 37859
rect 1627 37825 1636 37859
rect 1584 37816 1636 37825
rect 23112 37884 23164 37936
rect 26608 37995 26660 38004
rect 26608 37961 26617 37995
rect 26617 37961 26651 37995
rect 26651 37961 26660 37995
rect 26608 37952 26660 37961
rect 22008 37816 22060 37868
rect 28172 37952 28224 38004
rect 28908 37884 28960 37936
rect 4344 37748 4396 37800
rect 24308 37748 24360 37800
rect 24768 37859 24820 37868
rect 24768 37825 24777 37859
rect 24777 37825 24811 37859
rect 24811 37825 24820 37859
rect 25412 37859 25464 37868
rect 24768 37816 24820 37825
rect 25412 37825 25421 37859
rect 25421 37825 25455 37859
rect 25455 37825 25464 37859
rect 25412 37816 25464 37825
rect 25596 37859 25648 37868
rect 25596 37825 25605 37859
rect 25605 37825 25639 37859
rect 25639 37825 25648 37859
rect 25596 37816 25648 37825
rect 26056 37859 26108 37868
rect 26056 37825 26065 37859
rect 26065 37825 26099 37859
rect 26099 37825 26108 37859
rect 26056 37816 26108 37825
rect 27344 37859 27396 37868
rect 25964 37748 26016 37800
rect 14832 37680 14884 37732
rect 23112 37723 23164 37732
rect 23112 37689 23121 37723
rect 23121 37689 23155 37723
rect 23155 37689 23164 37723
rect 23112 37680 23164 37689
rect 26240 37680 26292 37732
rect 27344 37825 27353 37859
rect 27353 37825 27387 37859
rect 27387 37825 27396 37859
rect 27344 37816 27396 37825
rect 26700 37748 26752 37800
rect 27160 37748 27212 37800
rect 28080 37816 28132 37868
rect 28724 37816 28776 37868
rect 29828 37952 29880 38004
rect 30104 37995 30156 38004
rect 30104 37961 30113 37995
rect 30113 37961 30147 37995
rect 30147 37961 30156 37995
rect 30104 37952 30156 37961
rect 29276 37927 29328 37936
rect 29276 37893 29285 37927
rect 29285 37893 29319 37927
rect 29319 37893 29328 37927
rect 29276 37884 29328 37893
rect 29460 37884 29512 37936
rect 29092 37816 29144 37868
rect 29736 37884 29788 37936
rect 32588 37952 32640 38004
rect 32680 37995 32732 38004
rect 32680 37961 32689 37995
rect 32689 37961 32723 37995
rect 32723 37961 32732 37995
rect 34336 37995 34388 38004
rect 32680 37952 32732 37961
rect 34336 37961 34345 37995
rect 34345 37961 34379 37995
rect 34379 37961 34388 37995
rect 34336 37952 34388 37961
rect 30840 37884 30892 37936
rect 31024 37884 31076 37936
rect 29644 37859 29696 37868
rect 29644 37825 29653 37859
rect 29653 37825 29687 37859
rect 29687 37825 29696 37859
rect 29644 37816 29696 37825
rect 29828 37816 29880 37868
rect 30564 37859 30616 37868
rect 30564 37825 30609 37859
rect 30609 37825 30616 37859
rect 30564 37816 30616 37825
rect 30932 37816 30984 37868
rect 31208 37859 31260 37868
rect 31208 37825 31217 37859
rect 31217 37825 31251 37859
rect 31251 37825 31260 37859
rect 31208 37816 31260 37825
rect 33048 37816 33100 37868
rect 33232 37859 33284 37868
rect 33232 37825 33241 37859
rect 33241 37825 33275 37859
rect 33275 37825 33284 37859
rect 33232 37816 33284 37825
rect 51356 37952 51408 38004
rect 53656 37884 53708 37936
rect 2780 37612 2832 37664
rect 23572 37612 23624 37664
rect 25228 37655 25280 37664
rect 25228 37621 25237 37655
rect 25237 37621 25271 37655
rect 25271 37621 25280 37655
rect 25228 37612 25280 37621
rect 25596 37655 25648 37664
rect 25596 37621 25605 37655
rect 25605 37621 25639 37655
rect 25639 37621 25648 37655
rect 25596 37612 25648 37621
rect 26148 37612 26200 37664
rect 26700 37612 26752 37664
rect 28264 37612 28316 37664
rect 53656 37748 53708 37800
rect 29828 37612 29880 37664
rect 32128 37612 32180 37664
rect 33048 37612 33100 37664
rect 34612 37612 34664 37664
rect 53012 37655 53064 37664
rect 53012 37621 53021 37655
rect 53021 37621 53055 37655
rect 53055 37621 53064 37655
rect 53012 37612 53064 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2320 37408 2372 37460
rect 24032 37451 24084 37460
rect 24032 37417 24041 37451
rect 24041 37417 24075 37451
rect 24075 37417 24084 37451
rect 24032 37408 24084 37417
rect 24676 37451 24728 37460
rect 24676 37417 24685 37451
rect 24685 37417 24719 37451
rect 24719 37417 24728 37451
rect 24676 37408 24728 37417
rect 24768 37408 24820 37460
rect 27344 37408 27396 37460
rect 27436 37408 27488 37460
rect 28172 37408 28224 37460
rect 30104 37408 30156 37460
rect 30380 37408 30432 37460
rect 32128 37451 32180 37460
rect 32128 37417 32137 37451
rect 32137 37417 32171 37451
rect 32171 37417 32180 37451
rect 32128 37408 32180 37417
rect 32312 37408 32364 37460
rect 2780 37272 2832 37324
rect 22376 37315 22428 37324
rect 22376 37281 22385 37315
rect 22385 37281 22419 37315
rect 22419 37281 22428 37315
rect 22376 37272 22428 37281
rect 26424 37340 26476 37392
rect 53564 37408 53616 37460
rect 27436 37272 27488 37324
rect 23940 37204 23992 37256
rect 25228 37204 25280 37256
rect 26884 37247 26936 37256
rect 26884 37213 26893 37247
rect 26893 37213 26927 37247
rect 26927 37213 26936 37247
rect 26884 37204 26936 37213
rect 27068 37247 27120 37256
rect 27068 37213 27076 37247
rect 27076 37213 27110 37247
rect 27110 37213 27120 37247
rect 27068 37204 27120 37213
rect 27160 37247 27212 37256
rect 27160 37213 27169 37247
rect 27169 37213 27203 37247
rect 27203 37213 27212 37247
rect 27160 37204 27212 37213
rect 27344 37204 27396 37256
rect 27620 37204 27672 37256
rect 28448 37272 28500 37324
rect 28816 37315 28868 37324
rect 28816 37281 28825 37315
rect 28825 37281 28859 37315
rect 28859 37281 28868 37315
rect 28816 37272 28868 37281
rect 28908 37272 28960 37324
rect 29828 37272 29880 37324
rect 30196 37272 30248 37324
rect 28172 37247 28224 37256
rect 28172 37213 28180 37247
rect 28180 37213 28214 37247
rect 28214 37213 28224 37247
rect 28172 37204 28224 37213
rect 28724 37247 28776 37256
rect 26056 37179 26108 37188
rect 26056 37145 26065 37179
rect 26065 37145 26099 37179
rect 26099 37145 26108 37179
rect 26792 37179 26844 37188
rect 26056 37136 26108 37145
rect 26792 37145 26801 37179
rect 26801 37145 26835 37179
rect 26835 37145 26844 37179
rect 26792 37136 26844 37145
rect 27896 37179 27948 37188
rect 27896 37145 27908 37179
rect 27908 37145 27942 37179
rect 27942 37145 27948 37179
rect 27896 37136 27948 37145
rect 23020 37068 23072 37120
rect 25504 37068 25556 37120
rect 25596 37068 25648 37120
rect 26700 37068 26752 37120
rect 28724 37213 28733 37247
rect 28733 37213 28767 37247
rect 28767 37213 28776 37247
rect 28724 37204 28776 37213
rect 29092 37111 29144 37120
rect 29092 37077 29101 37111
rect 29101 37077 29135 37111
rect 29135 37077 29144 37111
rect 29092 37068 29144 37077
rect 29828 37068 29880 37120
rect 30104 37179 30156 37188
rect 30104 37145 30113 37179
rect 30113 37145 30147 37179
rect 30147 37145 30156 37179
rect 30380 37247 30432 37256
rect 30380 37213 30389 37247
rect 30389 37213 30423 37247
rect 30423 37213 30432 37247
rect 31576 37272 31628 37324
rect 33784 37315 33836 37324
rect 33784 37281 33793 37315
rect 33793 37281 33827 37315
rect 33827 37281 33836 37315
rect 33784 37272 33836 37281
rect 53472 37315 53524 37324
rect 53472 37281 53481 37315
rect 53481 37281 53515 37315
rect 53515 37281 53524 37315
rect 53472 37272 53524 37281
rect 30380 37204 30432 37213
rect 44180 37204 44232 37256
rect 53012 37247 53064 37256
rect 53012 37213 53021 37247
rect 53021 37213 53055 37247
rect 53055 37213 53064 37247
rect 53012 37204 53064 37213
rect 53564 37204 53616 37256
rect 30104 37136 30156 37145
rect 30840 37136 30892 37188
rect 33232 37136 33284 37188
rect 30288 37068 30340 37120
rect 33048 37111 33100 37120
rect 33048 37077 33057 37111
rect 33057 37077 33091 37111
rect 33091 37077 33100 37111
rect 33048 37068 33100 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 23664 36864 23716 36916
rect 17224 36728 17276 36780
rect 2780 36660 2832 36712
rect 13452 36524 13504 36576
rect 26700 36864 26752 36916
rect 28724 36907 28776 36916
rect 28724 36873 28733 36907
rect 28733 36873 28767 36907
rect 28767 36873 28776 36907
rect 28724 36864 28776 36873
rect 31852 36864 31904 36916
rect 28356 36796 28408 36848
rect 30840 36796 30892 36848
rect 35900 36864 35952 36916
rect 53012 36907 53064 36916
rect 53012 36873 53021 36907
rect 53021 36873 53055 36907
rect 53055 36873 53064 36907
rect 53012 36864 53064 36873
rect 25412 36771 25464 36780
rect 25412 36737 25421 36771
rect 25421 36737 25455 36771
rect 25455 36737 25464 36771
rect 25872 36771 25924 36780
rect 25412 36728 25464 36737
rect 25872 36737 25881 36771
rect 25881 36737 25915 36771
rect 25915 36737 25924 36771
rect 25872 36728 25924 36737
rect 26056 36771 26108 36780
rect 26056 36737 26065 36771
rect 26065 36737 26099 36771
rect 26099 36737 26108 36771
rect 26056 36728 26108 36737
rect 26240 36771 26292 36780
rect 26240 36737 26249 36771
rect 26249 36737 26283 36771
rect 26283 36737 26292 36771
rect 26240 36728 26292 36737
rect 27344 36771 27396 36780
rect 27344 36737 27353 36771
rect 27353 36737 27387 36771
rect 27387 36737 27396 36771
rect 27344 36728 27396 36737
rect 27620 36728 27672 36780
rect 28264 36771 28316 36780
rect 28264 36737 28273 36771
rect 28273 36737 28307 36771
rect 28307 36737 28316 36771
rect 28264 36728 28316 36737
rect 27896 36660 27948 36712
rect 22560 36635 22612 36644
rect 22560 36601 22569 36635
rect 22569 36601 22603 36635
rect 22603 36601 22612 36635
rect 22560 36592 22612 36601
rect 26148 36592 26200 36644
rect 27436 36592 27488 36644
rect 28540 36771 28592 36780
rect 28540 36737 28549 36771
rect 28549 36737 28583 36771
rect 28583 36737 28592 36771
rect 28540 36728 28592 36737
rect 29736 36728 29788 36780
rect 31944 36728 31996 36780
rect 28724 36660 28776 36712
rect 53564 36728 53616 36780
rect 53748 36703 53800 36712
rect 53748 36669 53757 36703
rect 53757 36669 53791 36703
rect 53791 36669 53800 36703
rect 53748 36660 53800 36669
rect 28908 36592 28960 36644
rect 31208 36635 31260 36644
rect 31208 36601 31217 36635
rect 31217 36601 31251 36635
rect 31251 36601 31260 36635
rect 31208 36592 31260 36601
rect 49608 36592 49660 36644
rect 53564 36592 53616 36644
rect 22652 36524 22704 36576
rect 23664 36524 23716 36576
rect 24676 36524 24728 36576
rect 26700 36524 26752 36576
rect 29276 36567 29328 36576
rect 29276 36533 29285 36567
rect 29285 36533 29319 36567
rect 29319 36533 29328 36567
rect 29276 36524 29328 36533
rect 33232 36524 33284 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 23480 36363 23532 36372
rect 23480 36329 23489 36363
rect 23489 36329 23523 36363
rect 23523 36329 23532 36363
rect 23480 36320 23532 36329
rect 25136 36320 25188 36372
rect 25228 36320 25280 36372
rect 26424 36320 26476 36372
rect 27620 36320 27672 36372
rect 28908 36320 28960 36372
rect 31944 36363 31996 36372
rect 13452 36252 13504 36304
rect 17316 36252 17368 36304
rect 22284 36295 22336 36304
rect 22284 36261 22293 36295
rect 22293 36261 22327 36295
rect 22327 36261 22336 36295
rect 22284 36252 22336 36261
rect 31944 36329 31953 36363
rect 31953 36329 31987 36363
rect 31987 36329 31996 36363
rect 31944 36320 31996 36329
rect 33048 36320 33100 36372
rect 2780 36116 2832 36168
rect 2044 36048 2096 36100
rect 26700 36227 26752 36236
rect 25228 36159 25280 36168
rect 25228 36125 25237 36159
rect 25237 36125 25271 36159
rect 25271 36125 25280 36159
rect 25228 36116 25280 36125
rect 26700 36193 26709 36227
rect 26709 36193 26743 36227
rect 26743 36193 26752 36227
rect 26700 36184 26752 36193
rect 25596 36159 25648 36168
rect 25596 36125 25605 36159
rect 25605 36125 25639 36159
rect 25639 36125 25648 36159
rect 25596 36116 25648 36125
rect 25964 36116 26016 36168
rect 26424 36116 26476 36168
rect 27896 36184 27948 36236
rect 21272 36091 21324 36100
rect 21272 36057 21281 36091
rect 21281 36057 21315 36091
rect 21315 36057 21324 36091
rect 21272 36048 21324 36057
rect 25412 36048 25464 36100
rect 27344 36159 27396 36168
rect 27344 36125 27353 36159
rect 27353 36125 27387 36159
rect 27387 36125 27396 36159
rect 27344 36116 27396 36125
rect 27528 36159 27580 36168
rect 27528 36125 27537 36159
rect 27537 36125 27571 36159
rect 27571 36125 27580 36159
rect 27528 36116 27580 36125
rect 28080 36116 28132 36168
rect 28816 36184 28868 36236
rect 29000 36184 29052 36236
rect 31760 36252 31812 36304
rect 32312 36252 32364 36304
rect 53748 36320 53800 36372
rect 49608 36184 49660 36236
rect 26884 36048 26936 36100
rect 27436 36091 27488 36100
rect 27436 36057 27445 36091
rect 27445 36057 27479 36091
rect 27479 36057 27488 36091
rect 27436 36048 27488 36057
rect 28632 36116 28684 36168
rect 29460 36116 29512 36168
rect 52368 36159 52420 36168
rect 52368 36125 52377 36159
rect 52377 36125 52411 36159
rect 52411 36125 52420 36159
rect 52368 36116 52420 36125
rect 53472 36159 53524 36168
rect 53472 36125 53481 36159
rect 53481 36125 53515 36159
rect 53515 36125 53524 36159
rect 53472 36116 53524 36125
rect 29000 36048 29052 36100
rect 32312 36048 32364 36100
rect 15108 35980 15160 36032
rect 22928 36023 22980 36032
rect 22928 35989 22937 36023
rect 22937 35989 22971 36023
rect 22971 35989 22980 36023
rect 22928 35980 22980 35989
rect 23572 35980 23624 36032
rect 25596 35980 25648 36032
rect 25964 35980 26016 36032
rect 27896 35980 27948 36032
rect 28172 36023 28224 36032
rect 28172 35989 28181 36023
rect 28181 35989 28215 36023
rect 28215 35989 28224 36023
rect 28172 35980 28224 35989
rect 28724 35980 28776 36032
rect 29644 35980 29696 36032
rect 29736 35980 29788 36032
rect 31208 35980 31260 36032
rect 32588 36023 32640 36032
rect 32588 35989 32597 36023
rect 32597 35989 32631 36023
rect 32631 35989 32640 36023
rect 32588 35980 32640 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 20812 35776 20864 35828
rect 22284 35776 22336 35828
rect 23296 35776 23348 35828
rect 23664 35776 23716 35828
rect 23480 35708 23532 35760
rect 24032 35776 24084 35828
rect 24216 35819 24268 35828
rect 24216 35785 24225 35819
rect 24225 35785 24259 35819
rect 24259 35785 24268 35819
rect 24216 35776 24268 35785
rect 25320 35776 25372 35828
rect 24400 35708 24452 35760
rect 25044 35751 25096 35760
rect 15108 35640 15160 35692
rect 23572 35683 23624 35692
rect 23572 35649 23581 35683
rect 23581 35649 23615 35683
rect 23615 35649 23624 35683
rect 23572 35640 23624 35649
rect 2780 35572 2832 35624
rect 23756 35640 23808 35692
rect 24584 35640 24636 35692
rect 25044 35717 25053 35751
rect 25053 35717 25087 35751
rect 25087 35717 25096 35751
rect 25044 35708 25096 35717
rect 24860 35640 24912 35692
rect 2504 35436 2556 35488
rect 22560 35547 22612 35556
rect 22560 35513 22569 35547
rect 22569 35513 22603 35547
rect 22603 35513 22612 35547
rect 26148 35640 26200 35692
rect 26424 35683 26476 35692
rect 25596 35572 25648 35624
rect 26424 35649 26433 35683
rect 26433 35649 26467 35683
rect 26467 35649 26476 35683
rect 26424 35640 26476 35649
rect 27160 35776 27212 35828
rect 27528 35751 27580 35760
rect 27528 35717 27537 35751
rect 27537 35717 27571 35751
rect 27571 35717 27580 35751
rect 27528 35708 27580 35717
rect 27436 35683 27488 35692
rect 27436 35649 27445 35683
rect 27445 35649 27479 35683
rect 27479 35649 27488 35683
rect 27436 35640 27488 35649
rect 28724 35751 28776 35760
rect 28724 35717 28733 35751
rect 28733 35717 28767 35751
rect 28767 35717 28776 35751
rect 28724 35708 28776 35717
rect 29092 35708 29144 35760
rect 28356 35683 28408 35692
rect 28356 35649 28365 35683
rect 28365 35649 28399 35683
rect 28399 35649 28408 35683
rect 28356 35640 28408 35649
rect 28540 35640 28592 35692
rect 29644 35640 29696 35692
rect 30012 35683 30064 35692
rect 30012 35649 30021 35683
rect 30021 35649 30055 35683
rect 30055 35649 30064 35683
rect 30012 35640 30064 35649
rect 22560 35504 22612 35513
rect 26148 35504 26200 35556
rect 20812 35479 20864 35488
rect 20812 35445 20821 35479
rect 20821 35445 20855 35479
rect 20855 35445 20864 35479
rect 20812 35436 20864 35445
rect 23020 35436 23072 35488
rect 23296 35436 23348 35488
rect 24216 35436 24268 35488
rect 25872 35436 25924 35488
rect 25964 35436 26016 35488
rect 28632 35572 28684 35624
rect 29460 35572 29512 35624
rect 30288 35683 30340 35692
rect 30288 35649 30297 35683
rect 30297 35649 30331 35683
rect 30331 35649 30340 35683
rect 30288 35640 30340 35649
rect 26516 35504 26568 35556
rect 27160 35479 27212 35488
rect 27160 35445 27169 35479
rect 27169 35445 27203 35479
rect 27203 35445 27212 35479
rect 27160 35436 27212 35445
rect 28632 35436 28684 35488
rect 28908 35436 28960 35488
rect 29092 35436 29144 35488
rect 30288 35504 30340 35556
rect 31392 35572 31444 35624
rect 33692 35776 33744 35828
rect 54024 35776 54076 35828
rect 44180 35640 44232 35692
rect 33692 35572 33744 35624
rect 53472 35615 53524 35624
rect 53472 35581 53481 35615
rect 53481 35581 53515 35615
rect 53515 35581 53524 35615
rect 53472 35572 53524 35581
rect 29644 35436 29696 35488
rect 30840 35436 30892 35488
rect 31024 35479 31076 35488
rect 31024 35445 31033 35479
rect 31033 35445 31067 35479
rect 31067 35445 31076 35479
rect 31024 35436 31076 35445
rect 31484 35436 31536 35488
rect 53564 35436 53616 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 15108 35232 15160 35284
rect 16672 35232 16724 35284
rect 27620 35232 27672 35284
rect 28448 35232 28500 35284
rect 29184 35275 29236 35284
rect 15016 35164 15068 35216
rect 26516 35164 26568 35216
rect 27068 35207 27120 35216
rect 27068 35173 27077 35207
rect 27077 35173 27111 35207
rect 27111 35173 27120 35207
rect 27068 35164 27120 35173
rect 14556 35096 14608 35148
rect 1584 35071 1636 35080
rect 1584 35037 1593 35071
rect 1593 35037 1627 35071
rect 1627 35037 1636 35071
rect 21180 35139 21232 35148
rect 21180 35105 21189 35139
rect 21189 35105 21223 35139
rect 21223 35105 21232 35139
rect 21180 35096 21232 35105
rect 1584 35028 1636 35037
rect 1768 34935 1820 34944
rect 1768 34901 1777 34935
rect 1777 34901 1811 34935
rect 1811 34901 1820 34935
rect 1768 34892 1820 34901
rect 2780 34892 2832 34944
rect 14556 34892 14608 34944
rect 15660 35028 15712 35080
rect 19340 35028 19392 35080
rect 21732 35071 21784 35080
rect 21732 35037 21741 35071
rect 21741 35037 21775 35071
rect 21775 35037 21784 35071
rect 21732 35028 21784 35037
rect 23112 35028 23164 35080
rect 23296 35028 23348 35080
rect 23480 35071 23532 35080
rect 23480 35037 23499 35071
rect 23499 35037 23532 35071
rect 25596 35096 25648 35148
rect 23480 35028 23532 35037
rect 23848 35071 23900 35080
rect 23848 35037 23857 35071
rect 23857 35037 23891 35071
rect 23891 35037 23900 35071
rect 23848 35028 23900 35037
rect 25872 35071 25924 35080
rect 25872 35037 25881 35071
rect 25881 35037 25915 35071
rect 25915 35037 25924 35071
rect 25872 35028 25924 35037
rect 27160 35096 27212 35148
rect 26516 35071 26568 35080
rect 26516 35037 26525 35071
rect 26525 35037 26559 35071
rect 26559 35037 26568 35071
rect 26516 35028 26568 35037
rect 26700 35071 26752 35080
rect 26700 35037 26709 35071
rect 26709 35037 26743 35071
rect 26743 35037 26752 35071
rect 26700 35028 26752 35037
rect 26792 35071 26844 35080
rect 26792 35037 26801 35071
rect 26801 35037 26835 35071
rect 26835 35037 26844 35071
rect 26792 35028 26844 35037
rect 29184 35241 29193 35275
rect 29193 35241 29227 35275
rect 29227 35241 29236 35275
rect 29184 35232 29236 35241
rect 29092 35164 29144 35216
rect 29644 35164 29696 35216
rect 31024 35232 31076 35284
rect 30380 35164 30432 35216
rect 35808 35164 35860 35216
rect 15016 34960 15068 35012
rect 23664 35003 23716 35012
rect 23664 34969 23673 35003
rect 23673 34969 23707 35003
rect 23707 34969 23716 35003
rect 23664 34960 23716 34969
rect 25964 34960 26016 35012
rect 26332 34960 26384 35012
rect 27068 34960 27120 35012
rect 27160 34960 27212 35012
rect 28264 34960 28316 35012
rect 28724 34960 28776 35012
rect 29644 35028 29696 35080
rect 30656 35028 30708 35080
rect 25044 34935 25096 34944
rect 25044 34901 25053 34935
rect 25053 34901 25087 34935
rect 25087 34901 25096 34935
rect 25044 34892 25096 34901
rect 29736 34960 29788 35012
rect 30380 35003 30432 35012
rect 30380 34969 30389 35003
rect 30389 34969 30423 35003
rect 30423 34969 30432 35003
rect 30380 34960 30432 34969
rect 29000 34892 29052 34944
rect 30104 34892 30156 34944
rect 30564 34892 30616 34944
rect 30932 35028 30984 35080
rect 31116 35028 31168 35080
rect 53288 35028 53340 35080
rect 53564 35028 53616 35080
rect 30840 34892 30892 34944
rect 33508 34892 33560 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 1768 34688 1820 34740
rect 23480 34688 23532 34740
rect 23572 34688 23624 34740
rect 25688 34688 25740 34740
rect 25780 34688 25832 34740
rect 22560 34620 22612 34672
rect 2780 34484 2832 34536
rect 13452 34527 13504 34536
rect 13452 34493 13461 34527
rect 13461 34493 13495 34527
rect 13495 34493 13504 34527
rect 14280 34595 14332 34604
rect 14280 34561 14289 34595
rect 14289 34561 14323 34595
rect 14323 34561 14332 34595
rect 14280 34552 14332 34561
rect 14740 34552 14792 34604
rect 15660 34595 15712 34604
rect 15660 34561 15669 34595
rect 15669 34561 15703 34595
rect 15703 34561 15712 34595
rect 15660 34552 15712 34561
rect 15016 34527 15068 34536
rect 13452 34484 13504 34493
rect 15016 34493 15025 34527
rect 15025 34493 15059 34527
rect 15059 34493 15068 34527
rect 15016 34484 15068 34493
rect 16672 34484 16724 34536
rect 17868 34484 17920 34536
rect 23940 34620 23992 34672
rect 24216 34663 24268 34672
rect 24216 34629 24225 34663
rect 24225 34629 24259 34663
rect 24259 34629 24268 34663
rect 24216 34620 24268 34629
rect 25320 34663 25372 34672
rect 25320 34629 25329 34663
rect 25329 34629 25363 34663
rect 25363 34629 25372 34663
rect 25320 34620 25372 34629
rect 25964 34620 26016 34672
rect 26240 34663 26292 34672
rect 26240 34629 26249 34663
rect 26249 34629 26283 34663
rect 26283 34629 26292 34663
rect 26240 34620 26292 34629
rect 23480 34552 23532 34604
rect 24308 34595 24360 34604
rect 24308 34561 24317 34595
rect 24317 34561 24351 34595
rect 24351 34561 24360 34595
rect 24308 34552 24360 34561
rect 25504 34552 25556 34604
rect 27620 34620 27672 34672
rect 28540 34688 28592 34740
rect 29736 34688 29788 34740
rect 29920 34688 29972 34740
rect 31484 34688 31536 34740
rect 24584 34484 24636 34536
rect 27068 34552 27120 34604
rect 28080 34552 28132 34604
rect 28540 34595 28592 34604
rect 28540 34561 28549 34595
rect 28549 34561 28583 34595
rect 28583 34561 28592 34595
rect 28540 34552 28592 34561
rect 28632 34595 28684 34604
rect 28632 34561 28641 34595
rect 28641 34561 28675 34595
rect 28675 34561 28684 34595
rect 29276 34595 29328 34604
rect 28632 34552 28684 34561
rect 29276 34561 29285 34595
rect 29285 34561 29319 34595
rect 29319 34561 29328 34595
rect 29276 34552 29328 34561
rect 23020 34459 23072 34468
rect 23020 34425 23029 34459
rect 23029 34425 23063 34459
rect 23063 34425 23072 34459
rect 23020 34416 23072 34425
rect 29460 34552 29512 34604
rect 29644 34595 29696 34604
rect 29644 34561 29653 34595
rect 29653 34561 29687 34595
rect 29687 34561 29696 34595
rect 29644 34552 29696 34561
rect 29920 34552 29972 34604
rect 30380 34595 30432 34604
rect 30380 34561 30389 34595
rect 30389 34561 30423 34595
rect 30423 34561 30432 34595
rect 30380 34552 30432 34561
rect 30472 34595 30524 34604
rect 30472 34561 30481 34595
rect 30481 34561 30515 34595
rect 30515 34561 30524 34595
rect 32312 34620 32364 34672
rect 30472 34552 30524 34561
rect 30380 34416 30432 34468
rect 30932 34484 30984 34536
rect 31484 34484 31536 34536
rect 43904 34552 43956 34604
rect 53472 34595 53524 34604
rect 53472 34561 53481 34595
rect 53481 34561 53515 34595
rect 53515 34561 53524 34595
rect 53472 34552 53524 34561
rect 53012 34527 53064 34536
rect 53012 34493 53021 34527
rect 53021 34493 53055 34527
rect 53055 34493 53064 34527
rect 53012 34484 53064 34493
rect 31116 34416 31168 34468
rect 53656 34416 53708 34468
rect 22836 34348 22888 34400
rect 23664 34348 23716 34400
rect 24216 34348 24268 34400
rect 26424 34348 26476 34400
rect 29092 34348 29144 34400
rect 30932 34391 30984 34400
rect 30932 34357 30941 34391
rect 30941 34357 30975 34391
rect 30975 34357 30984 34391
rect 30932 34348 30984 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 14740 34187 14792 34196
rect 14740 34153 14749 34187
rect 14749 34153 14783 34187
rect 14783 34153 14792 34187
rect 14740 34144 14792 34153
rect 22008 34144 22060 34196
rect 22836 34187 22888 34196
rect 22836 34153 22845 34187
rect 22845 34153 22879 34187
rect 22879 34153 22888 34187
rect 22836 34144 22888 34153
rect 23480 34187 23532 34196
rect 23480 34153 23489 34187
rect 23489 34153 23523 34187
rect 23523 34153 23532 34187
rect 23480 34144 23532 34153
rect 24216 34144 24268 34196
rect 24676 34144 24728 34196
rect 26700 34144 26752 34196
rect 28264 34144 28316 34196
rect 31208 34144 31260 34196
rect 31300 34144 31352 34196
rect 32312 34144 32364 34196
rect 23848 34076 23900 34128
rect 26056 34076 26108 34128
rect 28080 34076 28132 34128
rect 28356 34076 28408 34128
rect 29552 34076 29604 34128
rect 30288 34076 30340 34128
rect 22652 34008 22704 34060
rect 26332 34008 26384 34060
rect 26976 34008 27028 34060
rect 29460 34008 29512 34060
rect 2780 33940 2832 33992
rect 25320 33983 25372 33992
rect 25320 33949 25329 33983
rect 25329 33949 25363 33983
rect 25363 33949 25372 33983
rect 25320 33940 25372 33949
rect 26516 33940 26568 33992
rect 27068 33940 27120 33992
rect 27344 33983 27396 33992
rect 27344 33949 27353 33983
rect 27353 33949 27387 33983
rect 27387 33949 27396 33983
rect 27344 33940 27396 33949
rect 27988 33983 28040 33992
rect 26700 33872 26752 33924
rect 27252 33872 27304 33924
rect 27988 33949 27997 33983
rect 27997 33949 28031 33983
rect 28031 33949 28040 33983
rect 27988 33940 28040 33949
rect 30656 34008 30708 34060
rect 31760 34076 31812 34128
rect 53380 34119 53432 34128
rect 53380 34085 53389 34119
rect 53389 34085 53423 34119
rect 53423 34085 53432 34119
rect 53380 34076 53432 34085
rect 30288 33983 30340 33992
rect 30288 33949 30297 33983
rect 30297 33949 30331 33983
rect 30331 33949 30340 33983
rect 30288 33940 30340 33949
rect 30380 33983 30432 33992
rect 30380 33949 30389 33983
rect 30389 33949 30423 33983
rect 30423 33949 30432 33983
rect 30380 33940 30432 33949
rect 31208 33940 31260 33992
rect 31760 33872 31812 33924
rect 53104 33940 53156 33992
rect 53656 33983 53708 33992
rect 53656 33949 53665 33983
rect 53665 33949 53699 33983
rect 53699 33949 53708 33983
rect 53932 33983 53984 33992
rect 53656 33940 53708 33949
rect 53932 33949 53941 33983
rect 53941 33949 53975 33983
rect 53975 33949 53984 33983
rect 53932 33940 53984 33949
rect 24952 33804 25004 33856
rect 25872 33804 25924 33856
rect 26884 33804 26936 33856
rect 28448 33804 28500 33856
rect 30564 33804 30616 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 23112 33600 23164 33652
rect 24032 33600 24084 33652
rect 24216 33643 24268 33652
rect 24216 33609 24225 33643
rect 24225 33609 24259 33643
rect 24259 33609 24268 33643
rect 24216 33600 24268 33609
rect 24768 33600 24820 33652
rect 26976 33600 27028 33652
rect 27068 33600 27120 33652
rect 28264 33600 28316 33652
rect 51264 33600 51316 33652
rect 53104 33643 53156 33652
rect 53104 33609 53113 33643
rect 53113 33609 53147 33643
rect 53147 33609 53156 33643
rect 53104 33600 53156 33609
rect 6736 33464 6788 33516
rect 23480 33464 23532 33516
rect 26516 33532 26568 33584
rect 26700 33532 26752 33584
rect 24952 33507 25004 33516
rect 2780 33396 2832 33448
rect 13544 33328 13596 33380
rect 15108 33260 15160 33312
rect 24952 33473 24961 33507
rect 24961 33473 24995 33507
rect 24995 33473 25004 33507
rect 24952 33464 25004 33473
rect 25412 33464 25464 33516
rect 26240 33464 26292 33516
rect 25136 33396 25188 33448
rect 25872 33396 25924 33448
rect 26424 33464 26476 33516
rect 29092 33507 29144 33516
rect 29092 33473 29101 33507
rect 29101 33473 29135 33507
rect 29135 33473 29144 33507
rect 29092 33464 29144 33473
rect 29736 33507 29788 33516
rect 29736 33473 29745 33507
rect 29745 33473 29779 33507
rect 29779 33473 29788 33507
rect 29736 33464 29788 33473
rect 27344 33396 27396 33448
rect 24584 33328 24636 33380
rect 25320 33328 25372 33380
rect 26884 33328 26936 33380
rect 29000 33328 29052 33380
rect 29460 33396 29512 33448
rect 30656 33328 30708 33380
rect 53380 33328 53432 33380
rect 31760 33260 31812 33312
rect 54300 33303 54352 33312
rect 54300 33269 54309 33303
rect 54309 33269 54343 33303
rect 54343 33269 54352 33303
rect 54300 33260 54352 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 23480 33056 23532 33108
rect 25780 33056 25832 33108
rect 26148 33056 26200 33108
rect 27988 33056 28040 33108
rect 29000 33099 29052 33108
rect 29000 33065 29009 33099
rect 29009 33065 29043 33099
rect 29043 33065 29052 33099
rect 29000 33056 29052 33065
rect 26700 32988 26752 33040
rect 25320 32963 25372 32972
rect 25320 32929 25329 32963
rect 25329 32929 25363 32963
rect 25363 32929 25372 32963
rect 25320 32920 25372 32929
rect 26424 32920 26476 32972
rect 27620 32920 27672 32972
rect 1584 32895 1636 32904
rect 1584 32861 1593 32895
rect 1593 32861 1627 32895
rect 1627 32861 1636 32895
rect 1584 32852 1636 32861
rect 15108 32784 15160 32836
rect 26240 32852 26292 32904
rect 26884 32852 26936 32904
rect 27344 32852 27396 32904
rect 28080 32895 28132 32904
rect 28080 32861 28089 32895
rect 28089 32861 28123 32895
rect 28123 32861 28132 32895
rect 28080 32852 28132 32861
rect 28448 32895 28500 32904
rect 28448 32861 28457 32895
rect 28457 32861 28491 32895
rect 28491 32861 28500 32895
rect 54300 32895 54352 32904
rect 28448 32852 28500 32861
rect 54300 32861 54309 32895
rect 54309 32861 54343 32895
rect 54343 32861 54352 32895
rect 54300 32852 54352 32861
rect 2780 32716 2832 32768
rect 24032 32716 24084 32768
rect 27068 32784 27120 32836
rect 26332 32759 26384 32768
rect 26332 32725 26341 32759
rect 26341 32725 26375 32759
rect 26375 32725 26384 32759
rect 26332 32716 26384 32725
rect 29920 32716 29972 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 24032 32512 24084 32564
rect 24860 32512 24912 32564
rect 29736 32512 29788 32564
rect 24584 32487 24636 32496
rect 24584 32453 24593 32487
rect 24593 32453 24627 32487
rect 24627 32453 24636 32487
rect 24584 32444 24636 32453
rect 26516 32444 26568 32496
rect 26884 32444 26936 32496
rect 25872 32376 25924 32428
rect 26240 32376 26292 32428
rect 26976 32376 27028 32428
rect 27620 32444 27672 32496
rect 2780 32308 2832 32360
rect 26424 32351 26476 32360
rect 26424 32317 26433 32351
rect 26433 32317 26467 32351
rect 26467 32317 26476 32351
rect 32588 32376 32640 32428
rect 47860 32376 47912 32428
rect 26424 32308 26476 32317
rect 24952 32240 25004 32292
rect 27436 32240 27488 32292
rect 23020 32172 23072 32224
rect 24860 32215 24912 32224
rect 24860 32181 24869 32215
rect 24869 32181 24903 32215
rect 24903 32181 24912 32215
rect 24860 32172 24912 32181
rect 26976 32172 27028 32224
rect 27252 32172 27304 32224
rect 51172 32172 51224 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 24952 32011 25004 32020
rect 24952 31977 24961 32011
rect 24961 31977 24995 32011
rect 24995 31977 25004 32011
rect 24952 31968 25004 31977
rect 25964 31968 26016 32020
rect 2136 31807 2188 31816
rect 2136 31773 2145 31807
rect 2145 31773 2179 31807
rect 2179 31773 2188 31807
rect 2136 31764 2188 31773
rect 2780 31764 2832 31816
rect 26608 31807 26660 31816
rect 26608 31773 26617 31807
rect 26617 31773 26651 31807
rect 26651 31773 26660 31807
rect 26608 31764 26660 31773
rect 27436 31968 27488 32020
rect 26976 31807 27028 31816
rect 26976 31773 26985 31807
rect 26985 31773 27019 31807
rect 27019 31773 27028 31807
rect 26976 31764 27028 31773
rect 54300 31807 54352 31816
rect 25688 31696 25740 31748
rect 25964 31696 26016 31748
rect 24860 31628 24912 31680
rect 26148 31628 26200 31680
rect 54300 31773 54309 31807
rect 54309 31773 54343 31807
rect 54343 31773 54352 31807
rect 54300 31764 54352 31773
rect 27804 31696 27856 31748
rect 28356 31628 28408 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 26424 31467 26476 31476
rect 26424 31433 26433 31467
rect 26433 31433 26467 31467
rect 26467 31433 26476 31467
rect 26424 31424 26476 31433
rect 25872 31356 25924 31408
rect 26332 31399 26384 31408
rect 26332 31365 26341 31399
rect 26341 31365 26375 31399
rect 26375 31365 26384 31399
rect 26332 31356 26384 31365
rect 26608 31356 26660 31408
rect 27068 31356 27120 31408
rect 20812 31288 20864 31340
rect 25504 31288 25556 31340
rect 28356 31331 28408 31340
rect 2780 31220 2832 31272
rect 25780 31263 25832 31272
rect 25780 31229 25789 31263
rect 25789 31229 25823 31263
rect 25823 31229 25832 31263
rect 25780 31220 25832 31229
rect 28356 31297 28365 31331
rect 28365 31297 28399 31331
rect 28399 31297 28408 31331
rect 28356 31288 28408 31297
rect 26056 31220 26108 31272
rect 27988 31220 28040 31272
rect 33784 31152 33836 31204
rect 49332 31152 49384 31204
rect 30380 31084 30432 31136
rect 52828 31084 52880 31136
rect 54300 31127 54352 31136
rect 54300 31093 54309 31127
rect 54309 31093 54343 31127
rect 54343 31093 54352 31127
rect 54300 31084 54352 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 27712 30880 27764 30932
rect 30748 30880 30800 30932
rect 32404 30880 32456 30932
rect 26148 30812 26200 30864
rect 17868 30744 17920 30796
rect 26056 30744 26108 30796
rect 2780 30676 2832 30728
rect 26148 30583 26200 30592
rect 26148 30549 26157 30583
rect 26157 30549 26191 30583
rect 26191 30549 26200 30583
rect 26148 30540 26200 30549
rect 26976 30651 27028 30660
rect 26976 30617 26985 30651
rect 26985 30617 27019 30651
rect 27019 30617 27028 30651
rect 26976 30608 27028 30617
rect 44824 30540 44876 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 2136 30336 2188 30388
rect 26976 30336 27028 30388
rect 22376 30200 22428 30252
rect 2228 30132 2280 30184
rect 37648 29996 37700 30048
rect 54208 30039 54260 30048
rect 54208 30005 54217 30039
rect 54217 30005 54251 30039
rect 54251 30005 54260 30039
rect 54208 29996 54260 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2228 29835 2280 29844
rect 2228 29801 2237 29835
rect 2237 29801 2271 29835
rect 2271 29801 2280 29835
rect 2228 29792 2280 29801
rect 27344 29792 27396 29844
rect 27804 29792 27856 29844
rect 23296 29656 23348 29708
rect 47584 29656 47636 29708
rect 1584 29631 1636 29640
rect 1584 29597 1593 29631
rect 1593 29597 1627 29631
rect 1627 29597 1636 29631
rect 1584 29588 1636 29597
rect 4528 29588 4580 29640
rect 13820 29520 13872 29572
rect 24308 29588 24360 29640
rect 50804 29588 50856 29640
rect 54208 29631 54260 29640
rect 54208 29597 54217 29631
rect 54217 29597 54251 29631
rect 54251 29597 54260 29631
rect 54208 29588 54260 29597
rect 25964 29520 26016 29572
rect 27804 29520 27856 29572
rect 28356 29520 28408 29572
rect 30104 29520 30156 29572
rect 22744 29452 22796 29504
rect 30472 29452 30524 29504
rect 53564 29452 53616 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 25964 29291 26016 29300
rect 25964 29257 25973 29291
rect 25973 29257 26007 29291
rect 26007 29257 26016 29291
rect 25964 29248 26016 29257
rect 11060 29180 11112 29232
rect 4528 29112 4580 29164
rect 13820 29155 13872 29164
rect 13820 29121 13829 29155
rect 13829 29121 13863 29155
rect 13863 29121 13872 29155
rect 13820 29112 13872 29121
rect 14188 29155 14240 29164
rect 2780 29044 2832 29096
rect 13360 29044 13412 29096
rect 14188 29121 14197 29155
rect 14197 29121 14231 29155
rect 14231 29121 14240 29155
rect 14188 29112 14240 29121
rect 24400 29112 24452 29164
rect 26148 29112 26200 29164
rect 27344 29155 27396 29164
rect 21916 29044 21968 29096
rect 27344 29121 27353 29155
rect 27353 29121 27387 29155
rect 27387 29121 27396 29155
rect 27344 29112 27396 29121
rect 27528 29155 27580 29164
rect 27528 29121 27537 29155
rect 27537 29121 27571 29155
rect 27571 29121 27580 29155
rect 27528 29112 27580 29121
rect 30380 29248 30432 29300
rect 30472 29248 30524 29300
rect 53564 29248 53616 29300
rect 54208 29291 54260 29300
rect 54208 29257 54217 29291
rect 54217 29257 54251 29291
rect 54251 29257 54260 29291
rect 54208 29248 54260 29257
rect 27344 28976 27396 29028
rect 27528 28976 27580 29028
rect 35900 28976 35952 29028
rect 28080 28908 28132 28960
rect 54208 28908 54260 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 25412 28704 25464 28756
rect 26700 28568 26752 28620
rect 29920 28704 29972 28756
rect 29552 28636 29604 28688
rect 2780 28500 2832 28552
rect 24584 28500 24636 28552
rect 24676 28432 24728 28484
rect 26516 28475 26568 28484
rect 26516 28441 26525 28475
rect 26525 28441 26559 28475
rect 26559 28441 26568 28475
rect 26516 28432 26568 28441
rect 27528 28432 27580 28484
rect 28356 28543 28408 28552
rect 28356 28509 28365 28543
rect 28365 28509 28399 28543
rect 28399 28509 28408 28543
rect 28356 28500 28408 28509
rect 29828 28500 29880 28552
rect 54208 28543 54260 28552
rect 54208 28509 54217 28543
rect 54217 28509 54251 28543
rect 54251 28509 54260 28543
rect 54208 28500 54260 28509
rect 27804 28432 27856 28484
rect 33508 28432 33560 28484
rect 48596 28432 48648 28484
rect 53472 28475 53524 28484
rect 53472 28441 53481 28475
rect 53481 28441 53515 28475
rect 53515 28441 53524 28475
rect 53472 28432 53524 28441
rect 14188 28364 14240 28416
rect 15108 28364 15160 28416
rect 25228 28364 25280 28416
rect 27068 28364 27120 28416
rect 27620 28364 27672 28416
rect 30104 28407 30156 28416
rect 30104 28373 30113 28407
rect 30113 28373 30147 28407
rect 30147 28373 30156 28407
rect 30104 28364 30156 28373
rect 53196 28364 53248 28416
rect 53564 28364 53616 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 24676 28203 24728 28212
rect 24676 28169 24685 28203
rect 24685 28169 24719 28203
rect 24719 28169 24728 28203
rect 24676 28160 24728 28169
rect 25228 28135 25280 28144
rect 25228 28101 25237 28135
rect 25237 28101 25271 28135
rect 25271 28101 25280 28135
rect 25228 28092 25280 28101
rect 25872 28135 25924 28144
rect 25872 28101 25881 28135
rect 25881 28101 25915 28135
rect 25915 28101 25924 28135
rect 25872 28092 25924 28101
rect 26516 28160 26568 28212
rect 27804 28203 27856 28212
rect 27804 28169 27813 28203
rect 27813 28169 27847 28203
rect 27847 28169 27856 28203
rect 27804 28160 27856 28169
rect 33048 28160 33100 28212
rect 53564 28160 53616 28212
rect 54208 28203 54260 28212
rect 54208 28169 54217 28203
rect 54217 28169 54251 28203
rect 54251 28169 54260 28203
rect 54208 28160 54260 28169
rect 27528 28135 27580 28144
rect 2688 28024 2740 28076
rect 26424 28067 26476 28076
rect 26424 28033 26433 28067
rect 26433 28033 26467 28067
rect 26467 28033 26476 28067
rect 26424 28024 26476 28033
rect 27528 28101 27537 28135
rect 27537 28101 27571 28135
rect 27571 28101 27580 28135
rect 27528 28092 27580 28101
rect 2228 27956 2280 28008
rect 15108 27956 15160 28008
rect 25228 27956 25280 28008
rect 25780 27956 25832 28008
rect 27344 28024 27396 28076
rect 27620 28067 27672 28076
rect 27620 28033 27634 28067
rect 27634 28033 27668 28067
rect 27668 28033 27672 28067
rect 28264 28067 28316 28076
rect 27620 28024 27672 28033
rect 28264 28033 28273 28067
rect 28273 28033 28307 28067
rect 28307 28033 28316 28067
rect 28264 28024 28316 28033
rect 28172 27956 28224 28008
rect 28356 27999 28408 28008
rect 28356 27965 28365 27999
rect 28365 27965 28399 27999
rect 28399 27965 28408 27999
rect 28356 27956 28408 27965
rect 26608 27888 26660 27940
rect 27344 27888 27396 27940
rect 28080 27820 28132 27872
rect 28632 27863 28684 27872
rect 28632 27829 28641 27863
rect 28641 27829 28675 27863
rect 28675 27829 28684 27863
rect 28632 27820 28684 27829
rect 37464 27820 37516 27872
rect 52828 27956 52880 28008
rect 53472 27863 53524 27872
rect 53472 27829 53481 27863
rect 53481 27829 53515 27863
rect 53515 27829 53524 27863
rect 53472 27820 53524 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2228 27659 2280 27668
rect 2228 27625 2237 27659
rect 2237 27625 2271 27659
rect 2271 27625 2280 27659
rect 2228 27616 2280 27625
rect 24400 27548 24452 27600
rect 26424 27591 26476 27600
rect 26424 27557 26433 27591
rect 26433 27557 26467 27591
rect 26467 27557 26476 27591
rect 26424 27548 26476 27557
rect 28356 27548 28408 27600
rect 23940 27480 23992 27532
rect 1584 27455 1636 27464
rect 1584 27421 1593 27455
rect 1593 27421 1627 27455
rect 1627 27421 1636 27455
rect 1584 27412 1636 27421
rect 25228 27455 25280 27464
rect 11060 27344 11112 27396
rect 25228 27421 25237 27455
rect 25237 27421 25271 27455
rect 25271 27421 25280 27455
rect 25228 27412 25280 27421
rect 25872 27455 25924 27464
rect 25872 27421 25881 27455
rect 25881 27421 25915 27455
rect 25915 27421 25924 27455
rect 25872 27412 25924 27421
rect 26516 27412 26568 27464
rect 27068 27412 27120 27464
rect 28632 27480 28684 27532
rect 27712 27455 27764 27464
rect 27712 27421 27720 27455
rect 27720 27421 27754 27455
rect 27754 27421 27764 27455
rect 27712 27412 27764 27421
rect 27896 27412 27948 27464
rect 29828 27412 29880 27464
rect 30104 27412 30156 27464
rect 53472 27455 53524 27464
rect 53472 27421 53481 27455
rect 53481 27421 53515 27455
rect 53515 27421 53524 27455
rect 53472 27412 53524 27421
rect 53656 27412 53708 27464
rect 26056 27387 26108 27396
rect 26056 27353 26065 27387
rect 26065 27353 26099 27387
rect 26099 27353 26108 27387
rect 26056 27344 26108 27353
rect 26148 27387 26200 27396
rect 26148 27353 26157 27387
rect 26157 27353 26191 27387
rect 26191 27353 26200 27387
rect 26148 27344 26200 27353
rect 25412 27319 25464 27328
rect 25412 27285 25421 27319
rect 25421 27285 25455 27319
rect 25455 27285 25464 27319
rect 25412 27276 25464 27285
rect 27068 27276 27120 27328
rect 33784 27276 33836 27328
rect 52828 27276 52880 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 24400 27115 24452 27124
rect 24400 27081 24409 27115
rect 24409 27081 24443 27115
rect 24443 27081 24452 27115
rect 24400 27072 24452 27081
rect 25228 27072 25280 27124
rect 25872 27072 25924 27124
rect 34520 27115 34572 27124
rect 25412 27004 25464 27056
rect 25964 26936 26016 26988
rect 2780 26868 2832 26920
rect 25688 26868 25740 26920
rect 27068 26936 27120 26988
rect 27436 26936 27488 26988
rect 26516 26911 26568 26920
rect 26516 26877 26525 26911
rect 26525 26877 26559 26911
rect 26559 26877 26568 26911
rect 26516 26868 26568 26877
rect 26884 26868 26936 26920
rect 23940 26800 23992 26852
rect 25780 26800 25832 26852
rect 34520 27081 34529 27115
rect 34529 27081 34563 27115
rect 34563 27081 34572 27115
rect 34520 27072 34572 27081
rect 36084 27072 36136 27124
rect 54208 27047 54260 27056
rect 54208 27013 54217 27047
rect 54217 27013 54251 27047
rect 54251 27013 54260 27047
rect 54208 27004 54260 27013
rect 53564 26936 53616 26988
rect 31760 26868 31812 26920
rect 48504 26868 48556 26920
rect 39580 26800 39632 26852
rect 52552 26800 52604 26852
rect 26424 26732 26476 26784
rect 26608 26732 26660 26784
rect 28264 26775 28316 26784
rect 28264 26741 28273 26775
rect 28273 26741 28307 26775
rect 28307 26741 28316 26775
rect 28264 26732 28316 26741
rect 34336 26732 34388 26784
rect 35716 26732 35768 26784
rect 52368 26732 52420 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 23664 26528 23716 26580
rect 27160 26528 27212 26580
rect 34336 26571 34388 26580
rect 34336 26537 34345 26571
rect 34345 26537 34379 26571
rect 34379 26537 34388 26571
rect 34336 26528 34388 26537
rect 35992 26571 36044 26580
rect 35992 26537 36001 26571
rect 36001 26537 36035 26571
rect 36035 26537 36044 26571
rect 35992 26528 36044 26537
rect 36176 26528 36228 26580
rect 36544 26571 36596 26580
rect 36544 26537 36553 26571
rect 36553 26537 36587 26571
rect 36587 26537 36596 26571
rect 36544 26528 36596 26537
rect 37464 26528 37516 26580
rect 42616 26528 42668 26580
rect 52368 26528 52420 26580
rect 54208 26571 54260 26580
rect 54208 26537 54217 26571
rect 54217 26537 54251 26571
rect 54251 26537 54260 26571
rect 54208 26528 54260 26537
rect 2688 26460 2740 26512
rect 26700 26460 26752 26512
rect 28264 26460 28316 26512
rect 2228 26324 2280 26376
rect 26148 26392 26200 26444
rect 26608 26392 26660 26444
rect 27436 26392 27488 26444
rect 24584 26324 24636 26376
rect 26424 26324 26476 26376
rect 27712 26324 27764 26376
rect 35900 26460 35952 26512
rect 43352 26460 43404 26512
rect 52552 26460 52604 26512
rect 44088 26392 44140 26444
rect 25964 26256 26016 26308
rect 26240 26256 26292 26308
rect 27528 26299 27580 26308
rect 27528 26265 27537 26299
rect 27537 26265 27571 26299
rect 27571 26265 27580 26299
rect 27528 26256 27580 26265
rect 42432 26324 42484 26376
rect 53564 26367 53616 26376
rect 53564 26333 53573 26367
rect 53573 26333 53607 26367
rect 53607 26333 53616 26367
rect 53564 26324 53616 26333
rect 44916 26256 44968 26308
rect 52920 26256 52972 26308
rect 31944 26188 31996 26240
rect 34428 26188 34480 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 2228 26027 2280 26036
rect 2228 25993 2237 26027
rect 2237 25993 2271 26027
rect 2271 25993 2280 26027
rect 2228 25984 2280 25993
rect 26332 25984 26384 26036
rect 27252 26027 27304 26036
rect 27252 25993 27261 26027
rect 27261 25993 27295 26027
rect 27295 25993 27304 26027
rect 27252 25984 27304 25993
rect 32864 25984 32916 26036
rect 33416 25984 33468 26036
rect 33600 26027 33652 26036
rect 33600 25993 33609 26027
rect 33609 25993 33643 26027
rect 33643 25993 33652 26027
rect 33600 25984 33652 25993
rect 35716 25984 35768 26036
rect 38200 26027 38252 26036
rect 38200 25993 38209 26027
rect 38209 25993 38243 26027
rect 38243 25993 38252 26027
rect 38200 25984 38252 25993
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 25412 25891 25464 25900
rect 25412 25857 25421 25891
rect 25421 25857 25455 25891
rect 25455 25857 25464 25891
rect 25412 25848 25464 25857
rect 26700 25848 26752 25900
rect 29000 25848 29052 25900
rect 34520 25891 34572 25900
rect 34520 25857 34529 25891
rect 34529 25857 34563 25891
rect 34563 25857 34572 25891
rect 34520 25848 34572 25857
rect 35440 25848 35492 25900
rect 21640 25780 21692 25832
rect 33048 25780 33100 25832
rect 14556 25712 14608 25764
rect 14924 25712 14976 25764
rect 28264 25712 28316 25764
rect 32864 25712 32916 25764
rect 34428 25780 34480 25832
rect 53472 25823 53524 25832
rect 53472 25789 53481 25823
rect 53481 25789 53515 25823
rect 53515 25789 53524 25823
rect 53472 25780 53524 25789
rect 53748 25823 53800 25832
rect 53748 25789 53757 25823
rect 53757 25789 53791 25823
rect 53791 25789 53800 25823
rect 53748 25780 53800 25789
rect 35532 25712 35584 25764
rect 52828 25712 52880 25764
rect 25228 25687 25280 25696
rect 25228 25653 25237 25687
rect 25237 25653 25271 25687
rect 25271 25653 25280 25687
rect 25228 25644 25280 25653
rect 34704 25687 34756 25696
rect 34704 25653 34713 25687
rect 34713 25653 34747 25687
rect 34747 25653 34756 25687
rect 34704 25644 34756 25653
rect 35348 25644 35400 25696
rect 39028 25644 39080 25696
rect 52920 25687 52972 25696
rect 52920 25653 52929 25687
rect 52929 25653 52963 25687
rect 52963 25653 52972 25687
rect 52920 25644 52972 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1584 25440 1636 25492
rect 26240 25440 26292 25492
rect 29000 25483 29052 25492
rect 29000 25449 29009 25483
rect 29009 25449 29043 25483
rect 29043 25449 29052 25483
rect 29000 25440 29052 25449
rect 31944 25483 31996 25492
rect 31944 25449 31953 25483
rect 31953 25449 31987 25483
rect 31987 25449 31996 25483
rect 31944 25440 31996 25449
rect 32404 25483 32456 25492
rect 32404 25449 32413 25483
rect 32413 25449 32447 25483
rect 32447 25449 32456 25483
rect 32404 25440 32456 25449
rect 35440 25440 35492 25492
rect 37648 25483 37700 25492
rect 37648 25449 37657 25483
rect 37657 25449 37691 25483
rect 37691 25449 37700 25483
rect 37648 25440 37700 25449
rect 39028 25440 39080 25492
rect 54208 25483 54260 25492
rect 25780 25304 25832 25356
rect 26424 25304 26476 25356
rect 29000 25304 29052 25356
rect 30012 25304 30064 25356
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 24860 25279 24912 25288
rect 24860 25245 24869 25279
rect 24869 25245 24903 25279
rect 24903 25245 24912 25279
rect 24860 25236 24912 25245
rect 26608 25279 26660 25288
rect 26608 25245 26617 25279
rect 26617 25245 26651 25279
rect 26651 25245 26660 25279
rect 26608 25236 26660 25245
rect 26700 25236 26752 25288
rect 27528 25279 27580 25288
rect 27528 25245 27537 25279
rect 27537 25245 27571 25279
rect 27571 25245 27580 25279
rect 27528 25236 27580 25245
rect 28172 25279 28224 25288
rect 28172 25245 28181 25279
rect 28181 25245 28215 25279
rect 28215 25245 28224 25279
rect 28172 25236 28224 25245
rect 33140 25279 33192 25288
rect 33140 25245 33149 25279
rect 33149 25245 33183 25279
rect 33183 25245 33192 25279
rect 33140 25236 33192 25245
rect 33600 25236 33652 25288
rect 35808 25372 35860 25424
rect 40132 25372 40184 25424
rect 34704 25304 34756 25356
rect 54208 25449 54217 25483
rect 54217 25449 54251 25483
rect 54251 25449 54260 25483
rect 54208 25440 54260 25449
rect 13452 25168 13504 25220
rect 28540 25168 28592 25220
rect 32588 25168 32640 25220
rect 33968 25211 34020 25220
rect 33968 25177 33977 25211
rect 33977 25177 34011 25211
rect 34011 25177 34020 25211
rect 33968 25168 34020 25177
rect 25044 25143 25096 25152
rect 25044 25109 25053 25143
rect 25053 25109 25087 25143
rect 25087 25109 25096 25143
rect 25044 25100 25096 25109
rect 25872 25143 25924 25152
rect 25872 25109 25881 25143
rect 25881 25109 25915 25143
rect 25915 25109 25924 25143
rect 25872 25100 25924 25109
rect 26792 25100 26844 25152
rect 33324 25143 33376 25152
rect 33324 25109 33333 25143
rect 33333 25109 33367 25143
rect 33367 25109 33376 25143
rect 33324 25100 33376 25109
rect 33876 25100 33928 25152
rect 34336 25236 34388 25288
rect 34428 25236 34480 25288
rect 34980 25279 35032 25288
rect 34980 25245 34989 25279
rect 34989 25245 35023 25279
rect 35023 25245 35032 25279
rect 34980 25236 35032 25245
rect 38384 25279 38436 25288
rect 38384 25245 38393 25279
rect 38393 25245 38427 25279
rect 38427 25245 38436 25279
rect 38384 25236 38436 25245
rect 39764 25236 39816 25288
rect 41420 25236 41472 25288
rect 38200 25168 38252 25220
rect 35716 25143 35768 25152
rect 35716 25109 35725 25143
rect 35725 25109 35759 25143
rect 35759 25109 35768 25143
rect 35716 25100 35768 25109
rect 35808 25100 35860 25152
rect 36820 25100 36872 25152
rect 37832 25100 37884 25152
rect 38660 25100 38712 25152
rect 53472 25143 53524 25152
rect 53472 25109 53481 25143
rect 53481 25109 53515 25143
rect 53515 25109 53524 25143
rect 53472 25100 53524 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 26608 24896 26660 24948
rect 28540 24939 28592 24948
rect 28540 24905 28549 24939
rect 28549 24905 28583 24939
rect 28583 24905 28592 24939
rect 28540 24896 28592 24905
rect 31944 24896 31996 24948
rect 33140 24939 33192 24948
rect 33140 24905 33149 24939
rect 33149 24905 33183 24939
rect 33183 24905 33192 24939
rect 33140 24896 33192 24905
rect 25044 24828 25096 24880
rect 33324 24828 33376 24880
rect 1676 24803 1728 24812
rect 1676 24769 1685 24803
rect 1685 24769 1719 24803
rect 1719 24769 1728 24803
rect 1676 24760 1728 24769
rect 4068 24556 4120 24608
rect 24308 24556 24360 24608
rect 28172 24760 28224 24812
rect 30932 24760 30984 24812
rect 32864 24803 32916 24812
rect 32864 24769 32873 24803
rect 32873 24769 32907 24803
rect 32907 24769 32916 24803
rect 32864 24760 32916 24769
rect 33692 24760 33744 24812
rect 34152 24760 34204 24812
rect 35532 24896 35584 24948
rect 35716 24871 35768 24880
rect 35716 24837 35750 24871
rect 35750 24837 35768 24871
rect 35716 24828 35768 24837
rect 36268 24828 36320 24880
rect 37740 24803 37792 24812
rect 37740 24769 37749 24803
rect 37749 24769 37783 24803
rect 37783 24769 37792 24803
rect 37740 24760 37792 24769
rect 38660 24803 38712 24812
rect 38660 24769 38694 24803
rect 38694 24769 38712 24803
rect 38660 24760 38712 24769
rect 40408 24803 40460 24812
rect 25044 24735 25096 24744
rect 25044 24701 25053 24735
rect 25053 24701 25087 24735
rect 25087 24701 25096 24735
rect 25044 24692 25096 24701
rect 26884 24692 26936 24744
rect 33600 24735 33652 24744
rect 33600 24701 33609 24735
rect 33609 24701 33643 24735
rect 33643 24701 33652 24735
rect 33600 24692 33652 24701
rect 25780 24556 25832 24608
rect 26424 24556 26476 24608
rect 31300 24556 31352 24608
rect 33600 24556 33652 24608
rect 38292 24692 38344 24744
rect 40408 24769 40417 24803
rect 40417 24769 40451 24803
rect 40451 24769 40460 24803
rect 40408 24760 40460 24769
rect 42064 24760 42116 24812
rect 53564 24760 53616 24812
rect 42892 24692 42944 24744
rect 44088 24692 44140 24744
rect 37280 24624 37332 24676
rect 37648 24624 37700 24676
rect 34980 24556 35032 24608
rect 35624 24556 35676 24608
rect 35716 24556 35768 24608
rect 37924 24599 37976 24608
rect 37924 24565 37933 24599
rect 37933 24565 37967 24599
rect 37967 24565 37976 24599
rect 37924 24556 37976 24565
rect 49884 24624 49936 24676
rect 38568 24556 38620 24608
rect 39028 24556 39080 24608
rect 40592 24599 40644 24608
rect 40592 24565 40601 24599
rect 40601 24565 40635 24599
rect 40635 24565 40644 24599
rect 40592 24556 40644 24565
rect 53472 24599 53524 24608
rect 53472 24565 53481 24599
rect 53481 24565 53515 24599
rect 53515 24565 53524 24599
rect 53472 24556 53524 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 14648 24395 14700 24404
rect 14648 24361 14657 24395
rect 14657 24361 14691 24395
rect 14691 24361 14700 24395
rect 14648 24352 14700 24361
rect 15108 24352 15160 24404
rect 24584 24352 24636 24404
rect 23388 24216 23440 24268
rect 15108 24148 15160 24200
rect 25688 24352 25740 24404
rect 26700 24352 26752 24404
rect 28172 24352 28224 24404
rect 30932 24395 30984 24404
rect 30932 24361 30941 24395
rect 30941 24361 30975 24395
rect 30975 24361 30984 24395
rect 30932 24352 30984 24361
rect 33692 24395 33744 24404
rect 33692 24361 33701 24395
rect 33701 24361 33735 24395
rect 33735 24361 33744 24395
rect 33692 24352 33744 24361
rect 33876 24352 33928 24404
rect 34244 24352 34296 24404
rect 35900 24352 35952 24404
rect 37464 24352 37516 24404
rect 25044 24148 25096 24200
rect 26884 24191 26936 24200
rect 26884 24157 26893 24191
rect 26893 24157 26927 24191
rect 26927 24157 26936 24191
rect 26884 24148 26936 24157
rect 31208 24284 31260 24336
rect 29644 24216 29696 24268
rect 31944 24216 31996 24268
rect 1676 24123 1728 24132
rect 1676 24089 1685 24123
rect 1685 24089 1719 24123
rect 1719 24089 1728 24123
rect 1676 24080 1728 24089
rect 25228 24123 25280 24132
rect 25228 24089 25262 24123
rect 25262 24089 25280 24123
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 14464 24012 14516 24064
rect 23572 24055 23624 24064
rect 23572 24021 23581 24055
rect 23581 24021 23615 24055
rect 23615 24021 23624 24055
rect 23572 24012 23624 24021
rect 25228 24080 25280 24089
rect 25320 24080 25372 24132
rect 31576 24191 31628 24200
rect 27160 24123 27212 24132
rect 27160 24089 27194 24123
rect 27194 24089 27212 24123
rect 31576 24157 31585 24191
rect 31585 24157 31619 24191
rect 31619 24157 31628 24191
rect 31576 24148 31628 24157
rect 34704 24284 34756 24336
rect 37740 24352 37792 24404
rect 38752 24352 38804 24404
rect 40316 24352 40368 24404
rect 41420 24395 41472 24404
rect 41420 24361 41429 24395
rect 41429 24361 41463 24395
rect 41463 24361 41472 24395
rect 53564 24395 53616 24404
rect 41420 24352 41472 24361
rect 53564 24361 53573 24395
rect 53573 24361 53607 24395
rect 53607 24361 53616 24395
rect 53564 24352 53616 24361
rect 33600 24216 33652 24268
rect 33876 24191 33928 24200
rect 33876 24157 33885 24191
rect 33885 24157 33919 24191
rect 33919 24157 33928 24191
rect 33876 24148 33928 24157
rect 34152 24148 34204 24200
rect 27160 24080 27212 24089
rect 32312 24080 32364 24132
rect 34060 24123 34112 24132
rect 34060 24089 34069 24123
rect 34069 24089 34103 24123
rect 34103 24089 34112 24123
rect 34060 24080 34112 24089
rect 26516 24012 26568 24064
rect 31392 24012 31444 24064
rect 32220 24055 32272 24064
rect 32220 24021 32229 24055
rect 32229 24021 32263 24055
rect 32263 24021 32272 24055
rect 32220 24012 32272 24021
rect 33232 24055 33284 24064
rect 33232 24021 33241 24055
rect 33241 24021 33275 24055
rect 33275 24021 33284 24055
rect 33232 24012 33284 24021
rect 33876 24012 33928 24064
rect 34612 24148 34664 24200
rect 37832 24216 37884 24268
rect 38292 24216 38344 24268
rect 40040 24259 40092 24268
rect 40040 24225 40049 24259
rect 40049 24225 40083 24259
rect 40083 24225 40092 24259
rect 40040 24216 40092 24225
rect 36360 24148 36412 24200
rect 36820 24148 36872 24200
rect 38752 24191 38804 24200
rect 38752 24157 38761 24191
rect 38761 24157 38795 24191
rect 38795 24157 38804 24191
rect 38752 24148 38804 24157
rect 35348 24080 35400 24132
rect 40132 24148 40184 24200
rect 54208 24191 54260 24200
rect 54208 24157 54217 24191
rect 54217 24157 54251 24191
rect 54251 24157 54260 24191
rect 54208 24148 54260 24157
rect 44088 24080 44140 24132
rect 52920 24080 52972 24132
rect 34336 24012 34388 24064
rect 34796 24012 34848 24064
rect 39304 24012 39356 24064
rect 40132 24012 40184 24064
rect 54116 24055 54168 24064
rect 54116 24021 54125 24055
rect 54125 24021 54159 24055
rect 54159 24021 54168 24055
rect 54116 24012 54168 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 4068 23808 4120 23860
rect 1768 23740 1820 23792
rect 23664 23715 23716 23724
rect 23664 23681 23673 23715
rect 23673 23681 23707 23715
rect 23707 23681 23716 23715
rect 23664 23672 23716 23681
rect 1676 23511 1728 23520
rect 1676 23477 1685 23511
rect 1685 23477 1719 23511
rect 1719 23477 1728 23511
rect 1676 23468 1728 23477
rect 14648 23468 14700 23520
rect 23388 23511 23440 23520
rect 23388 23477 23397 23511
rect 23397 23477 23431 23511
rect 23431 23477 23440 23511
rect 23388 23468 23440 23477
rect 25412 23808 25464 23860
rect 26424 23808 26476 23860
rect 31208 23808 31260 23860
rect 31760 23851 31812 23860
rect 31760 23817 31769 23851
rect 31769 23817 31803 23851
rect 31803 23817 31812 23851
rect 31760 23808 31812 23817
rect 31944 23808 31996 23860
rect 32404 23808 32456 23860
rect 34520 23808 34572 23860
rect 35808 23808 35860 23860
rect 24584 23783 24636 23792
rect 24584 23749 24593 23783
rect 24593 23749 24627 23783
rect 24627 23749 24636 23783
rect 24584 23740 24636 23749
rect 26332 23740 26384 23792
rect 37464 23808 37516 23860
rect 38384 23808 38436 23860
rect 39304 23808 39356 23860
rect 40316 23808 40368 23860
rect 54024 23808 54076 23860
rect 25320 23672 25372 23724
rect 25872 23672 25924 23724
rect 27252 23672 27304 23724
rect 24308 23647 24360 23656
rect 24308 23613 24317 23647
rect 24317 23613 24351 23647
rect 24351 23613 24360 23647
rect 24308 23604 24360 23613
rect 25412 23604 25464 23656
rect 25504 23604 25556 23656
rect 26976 23604 27028 23656
rect 27712 23647 27764 23656
rect 27712 23613 27721 23647
rect 27721 23613 27755 23647
rect 27755 23613 27764 23647
rect 27712 23604 27764 23613
rect 24400 23536 24452 23588
rect 27252 23468 27304 23520
rect 27436 23536 27488 23588
rect 30012 23715 30064 23724
rect 30012 23681 30021 23715
rect 30021 23681 30055 23715
rect 30055 23681 30064 23715
rect 30012 23672 30064 23681
rect 31208 23672 31260 23724
rect 31760 23672 31812 23724
rect 34060 23715 34112 23724
rect 32128 23604 32180 23656
rect 32404 23647 32456 23656
rect 32404 23613 32413 23647
rect 32413 23613 32447 23647
rect 32447 23613 32456 23647
rect 32404 23604 32456 23613
rect 34060 23681 34069 23715
rect 34069 23681 34103 23715
rect 34103 23681 34112 23715
rect 34060 23672 34112 23681
rect 34244 23715 34296 23724
rect 34244 23681 34253 23715
rect 34253 23681 34287 23715
rect 34287 23681 34296 23715
rect 34244 23672 34296 23681
rect 35532 23715 35584 23724
rect 35532 23681 35541 23715
rect 35541 23681 35575 23715
rect 35575 23681 35584 23715
rect 37740 23740 37792 23792
rect 37924 23740 37976 23792
rect 35532 23672 35584 23681
rect 36728 23715 36780 23724
rect 36728 23681 36737 23715
rect 36737 23681 36771 23715
rect 36771 23681 36780 23715
rect 36728 23672 36780 23681
rect 37648 23715 37700 23724
rect 37648 23681 37657 23715
rect 37657 23681 37691 23715
rect 37691 23681 37700 23715
rect 37648 23672 37700 23681
rect 38292 23715 38344 23724
rect 38292 23681 38301 23715
rect 38301 23681 38335 23715
rect 38335 23681 38344 23715
rect 38292 23672 38344 23681
rect 40132 23740 40184 23792
rect 40592 23740 40644 23792
rect 43996 23740 44048 23792
rect 54116 23740 54168 23792
rect 54208 23783 54260 23792
rect 54208 23749 54217 23783
rect 54217 23749 54251 23783
rect 54251 23749 54260 23783
rect 54208 23740 54260 23749
rect 34336 23536 34388 23588
rect 28908 23468 28960 23520
rect 29184 23468 29236 23520
rect 30196 23511 30248 23520
rect 30196 23477 30205 23511
rect 30205 23477 30239 23511
rect 30239 23477 30248 23511
rect 30196 23468 30248 23477
rect 30840 23511 30892 23520
rect 30840 23477 30849 23511
rect 30849 23477 30883 23511
rect 30883 23477 30892 23511
rect 30840 23468 30892 23477
rect 34428 23468 34480 23520
rect 35624 23604 35676 23656
rect 35532 23536 35584 23588
rect 40040 23672 40092 23724
rect 40684 23715 40736 23724
rect 40684 23681 40693 23715
rect 40693 23681 40727 23715
rect 40727 23681 40736 23715
rect 40684 23672 40736 23681
rect 42800 23672 42852 23724
rect 44088 23672 44140 23724
rect 53564 23672 53616 23724
rect 37832 23536 37884 23588
rect 37280 23468 37332 23520
rect 38936 23468 38988 23520
rect 42064 23579 42116 23588
rect 42064 23545 42073 23579
rect 42073 23545 42107 23579
rect 42107 23545 42116 23579
rect 42064 23536 42116 23545
rect 53288 23579 53340 23588
rect 53288 23545 53297 23579
rect 53297 23545 53331 23579
rect 53331 23545 53340 23579
rect 53288 23536 53340 23545
rect 53472 23536 53524 23588
rect 54024 23647 54076 23656
rect 54024 23613 54033 23647
rect 54033 23613 54067 23647
rect 54067 23613 54076 23647
rect 54024 23604 54076 23613
rect 40316 23468 40368 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 22928 23264 22980 23316
rect 23388 23264 23440 23316
rect 25780 23264 25832 23316
rect 27160 23264 27212 23316
rect 28908 23264 28960 23316
rect 29092 23307 29144 23316
rect 29092 23273 29101 23307
rect 29101 23273 29135 23307
rect 29135 23273 29144 23307
rect 29092 23264 29144 23273
rect 30840 23264 30892 23316
rect 32404 23264 32456 23316
rect 33784 23264 33836 23316
rect 34060 23264 34112 23316
rect 34428 23264 34480 23316
rect 37648 23264 37700 23316
rect 38200 23264 38252 23316
rect 40408 23307 40460 23316
rect 24584 23128 24636 23180
rect 25504 23128 25556 23180
rect 26332 23128 26384 23180
rect 27712 23128 27764 23180
rect 28724 23128 28776 23180
rect 33784 23171 33836 23180
rect 33784 23137 33793 23171
rect 33793 23137 33827 23171
rect 33827 23137 33836 23171
rect 33784 23128 33836 23137
rect 34980 23171 35032 23180
rect 2320 23060 2372 23112
rect 23572 23060 23624 23112
rect 25872 23060 25924 23112
rect 26240 23103 26292 23112
rect 26240 23069 26249 23103
rect 26249 23069 26283 23103
rect 26283 23069 26292 23103
rect 26240 23060 26292 23069
rect 27252 23103 27304 23112
rect 27252 23069 27261 23103
rect 27261 23069 27295 23103
rect 27295 23069 27304 23103
rect 27252 23060 27304 23069
rect 30380 23060 30432 23112
rect 33600 23060 33652 23112
rect 30196 22992 30248 23044
rect 31300 22992 31352 23044
rect 34980 23137 34989 23171
rect 34989 23137 35023 23171
rect 35023 23137 35032 23171
rect 34980 23128 35032 23137
rect 38660 23196 38712 23248
rect 40408 23273 40417 23307
rect 40417 23273 40451 23307
rect 40451 23273 40460 23307
rect 40408 23264 40460 23273
rect 43260 23264 43312 23316
rect 54208 23307 54260 23316
rect 54208 23273 54217 23307
rect 54217 23273 54251 23307
rect 54251 23273 54260 23307
rect 54208 23264 54260 23273
rect 42340 23239 42392 23248
rect 37464 23060 37516 23112
rect 37740 23103 37792 23112
rect 37740 23069 37749 23103
rect 37749 23069 37783 23103
rect 37783 23069 37792 23103
rect 37740 23060 37792 23069
rect 38016 23060 38068 23112
rect 38568 23103 38620 23112
rect 38568 23069 38577 23103
rect 38577 23069 38611 23103
rect 38611 23069 38620 23103
rect 38568 23060 38620 23069
rect 42340 23205 42349 23239
rect 42349 23205 42383 23239
rect 42383 23205 42392 23239
rect 53564 23239 53616 23248
rect 42340 23196 42392 23205
rect 40132 23128 40184 23180
rect 40684 23128 40736 23180
rect 40224 23103 40276 23112
rect 40224 23069 40233 23103
rect 40233 23069 40267 23103
rect 40267 23069 40276 23103
rect 40224 23060 40276 23069
rect 41512 23060 41564 23112
rect 53564 23205 53573 23239
rect 53573 23205 53607 23239
rect 53607 23205 53616 23239
rect 53564 23196 53616 23205
rect 35992 22992 36044 23044
rect 1676 22967 1728 22976
rect 1676 22933 1685 22967
rect 1685 22933 1719 22967
rect 1719 22933 1728 22967
rect 1676 22924 1728 22933
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 23020 22967 23072 22976
rect 23020 22933 23029 22967
rect 23029 22933 23063 22967
rect 23063 22933 23072 22967
rect 23020 22924 23072 22933
rect 23480 22924 23532 22976
rect 23756 22924 23808 22976
rect 26424 22924 26476 22976
rect 27344 22924 27396 22976
rect 31208 22967 31260 22976
rect 31208 22933 31217 22967
rect 31217 22933 31251 22967
rect 31251 22933 31260 22967
rect 31208 22924 31260 22933
rect 33140 22924 33192 22976
rect 35164 22967 35216 22976
rect 35164 22933 35173 22967
rect 35173 22933 35207 22967
rect 35207 22933 35216 22967
rect 35164 22924 35216 22933
rect 35808 22924 35860 22976
rect 39028 22924 39080 22976
rect 39948 22924 40000 22976
rect 41420 22924 41472 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 2320 22763 2372 22772
rect 2320 22729 2329 22763
rect 2329 22729 2363 22763
rect 2363 22729 2372 22763
rect 2320 22720 2372 22729
rect 1860 22627 1912 22636
rect 1860 22593 1869 22627
rect 1869 22593 1903 22627
rect 1903 22593 1912 22627
rect 1860 22584 1912 22593
rect 14556 22652 14608 22704
rect 14740 22584 14792 22636
rect 17224 22720 17276 22772
rect 22928 22763 22980 22772
rect 22928 22729 22937 22763
rect 22937 22729 22971 22763
rect 22971 22729 22980 22763
rect 22928 22720 22980 22729
rect 24308 22720 24360 22772
rect 18788 22652 18840 22704
rect 24860 22720 24912 22772
rect 25688 22763 25740 22772
rect 25688 22729 25697 22763
rect 25697 22729 25731 22763
rect 25731 22729 25740 22763
rect 25688 22720 25740 22729
rect 30012 22720 30064 22772
rect 31760 22763 31812 22772
rect 31760 22729 31769 22763
rect 31769 22729 31803 22763
rect 31803 22729 31812 22763
rect 32312 22763 32364 22772
rect 31760 22720 31812 22729
rect 32312 22729 32321 22763
rect 32321 22729 32355 22763
rect 32355 22729 32364 22763
rect 32312 22720 32364 22729
rect 33140 22720 33192 22772
rect 33324 22720 33376 22772
rect 35532 22763 35584 22772
rect 35532 22729 35541 22763
rect 35541 22729 35575 22763
rect 35575 22729 35584 22763
rect 35532 22720 35584 22729
rect 36728 22720 36780 22772
rect 37464 22720 37516 22772
rect 23480 22627 23532 22636
rect 23480 22593 23489 22627
rect 23489 22593 23523 22627
rect 23523 22593 23532 22627
rect 23480 22584 23532 22593
rect 2596 22516 2648 22568
rect 1676 22423 1728 22432
rect 1676 22389 1685 22423
rect 1685 22389 1719 22423
rect 1719 22389 1728 22423
rect 1676 22380 1728 22389
rect 14096 22380 14148 22432
rect 14648 22380 14700 22432
rect 15292 22423 15344 22432
rect 15292 22389 15301 22423
rect 15301 22389 15335 22423
rect 15335 22389 15344 22423
rect 15292 22380 15344 22389
rect 23480 22380 23532 22432
rect 26332 22652 26384 22704
rect 27528 22627 27580 22636
rect 27528 22593 27537 22627
rect 27537 22593 27571 22627
rect 27571 22593 27580 22627
rect 27528 22584 27580 22593
rect 27344 22559 27396 22568
rect 27344 22525 27353 22559
rect 27353 22525 27387 22559
rect 27387 22525 27396 22559
rect 29644 22627 29696 22636
rect 29644 22593 29653 22627
rect 29653 22593 29687 22627
rect 29687 22593 29696 22627
rect 29644 22584 29696 22593
rect 30932 22652 30984 22704
rect 33416 22652 33468 22704
rect 34244 22652 34296 22704
rect 34520 22652 34572 22704
rect 35716 22652 35768 22704
rect 30380 22627 30432 22636
rect 30380 22593 30389 22627
rect 30389 22593 30423 22627
rect 30423 22593 30432 22627
rect 30380 22584 30432 22593
rect 32220 22584 32272 22636
rect 32404 22584 32456 22636
rect 27344 22516 27396 22525
rect 32128 22516 32180 22568
rect 32772 22559 32824 22568
rect 32772 22525 32781 22559
rect 32781 22525 32815 22559
rect 32815 22525 32824 22559
rect 32772 22516 32824 22525
rect 32864 22559 32916 22568
rect 32864 22525 32873 22559
rect 32873 22525 32907 22559
rect 32907 22525 32916 22559
rect 34704 22584 34756 22636
rect 35256 22584 35308 22636
rect 35532 22584 35584 22636
rect 36176 22652 36228 22704
rect 37740 22720 37792 22772
rect 38752 22720 38804 22772
rect 40224 22720 40276 22772
rect 40408 22720 40460 22772
rect 53288 22720 53340 22772
rect 53472 22763 53524 22772
rect 53472 22729 53481 22763
rect 53481 22729 53515 22763
rect 53515 22729 53524 22763
rect 53472 22720 53524 22729
rect 54208 22763 54260 22772
rect 54208 22729 54217 22763
rect 54217 22729 54251 22763
rect 54251 22729 54260 22763
rect 54208 22720 54260 22729
rect 38384 22652 38436 22704
rect 39764 22695 39816 22704
rect 39764 22661 39773 22695
rect 39773 22661 39807 22695
rect 39807 22661 39816 22695
rect 39764 22652 39816 22661
rect 43260 22695 43312 22704
rect 43260 22661 43269 22695
rect 43269 22661 43303 22695
rect 43303 22661 43312 22695
rect 43260 22652 43312 22661
rect 36084 22584 36136 22636
rect 36452 22627 36504 22636
rect 36452 22593 36461 22627
rect 36461 22593 36495 22627
rect 36495 22593 36504 22627
rect 36452 22584 36504 22593
rect 32864 22516 32916 22525
rect 34796 22516 34848 22568
rect 34980 22516 35032 22568
rect 25688 22448 25740 22500
rect 27436 22448 27488 22500
rect 32588 22448 32640 22500
rect 35624 22448 35676 22500
rect 36084 22448 36136 22500
rect 38016 22584 38068 22636
rect 38660 22584 38712 22636
rect 38936 22516 38988 22568
rect 39212 22584 39264 22636
rect 39948 22627 40000 22636
rect 39948 22593 39957 22627
rect 39957 22593 39991 22627
rect 39991 22593 40000 22627
rect 39948 22584 40000 22593
rect 40316 22584 40368 22636
rect 40684 22627 40736 22636
rect 40684 22593 40693 22627
rect 40693 22593 40727 22627
rect 40727 22593 40736 22627
rect 40684 22584 40736 22593
rect 40132 22559 40184 22568
rect 40132 22525 40141 22559
rect 40141 22525 40175 22559
rect 40175 22525 40184 22559
rect 40132 22516 40184 22525
rect 40592 22516 40644 22568
rect 26516 22423 26568 22432
rect 26516 22389 26525 22423
rect 26525 22389 26559 22423
rect 26559 22389 26568 22423
rect 26516 22380 26568 22389
rect 28172 22423 28224 22432
rect 28172 22389 28181 22423
rect 28181 22389 28215 22423
rect 28215 22389 28224 22423
rect 28172 22380 28224 22389
rect 29644 22380 29696 22432
rect 31300 22380 31352 22432
rect 40040 22448 40092 22500
rect 42708 22584 42760 22636
rect 39764 22380 39816 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 14740 22219 14792 22228
rect 14740 22185 14749 22219
rect 14749 22185 14783 22219
rect 14783 22185 14792 22219
rect 14740 22176 14792 22185
rect 22928 22176 22980 22228
rect 24308 22176 24360 22228
rect 24768 22176 24820 22228
rect 25044 22176 25096 22228
rect 26884 22176 26936 22228
rect 27436 22176 27488 22228
rect 30932 22219 30984 22228
rect 30932 22185 30941 22219
rect 30941 22185 30975 22219
rect 30975 22185 30984 22219
rect 30932 22176 30984 22185
rect 32772 22176 32824 22228
rect 40408 22176 40460 22228
rect 43352 22219 43404 22228
rect 1860 22108 1912 22160
rect 23020 22108 23072 22160
rect 23480 22108 23532 22160
rect 15292 22040 15344 22092
rect 2412 21972 2464 22024
rect 21180 21972 21232 22024
rect 1676 21879 1728 21888
rect 1676 21845 1685 21879
rect 1685 21845 1719 21879
rect 1719 21845 1728 21879
rect 1676 21836 1728 21845
rect 22560 21972 22612 22024
rect 23756 22015 23808 22024
rect 23756 21981 23765 22015
rect 23765 21981 23799 22015
rect 23799 21981 23808 22015
rect 23756 21972 23808 21981
rect 24768 22015 24820 22024
rect 24768 21981 24777 22015
rect 24777 21981 24811 22015
rect 24811 21981 24820 22015
rect 24768 21972 24820 21981
rect 27344 22108 27396 22160
rect 30288 22108 30340 22160
rect 27436 22083 27488 22092
rect 27436 22049 27445 22083
rect 27445 22049 27479 22083
rect 27479 22049 27488 22083
rect 27436 22040 27488 22049
rect 28540 22040 28592 22092
rect 30840 22040 30892 22092
rect 32864 22108 32916 22160
rect 36360 22108 36412 22160
rect 36636 22108 36688 22160
rect 36820 22108 36872 22160
rect 37556 22083 37608 22092
rect 22284 21904 22336 21956
rect 25504 21904 25556 21956
rect 27160 21972 27212 22024
rect 28172 21972 28224 22024
rect 26608 21947 26660 21956
rect 26608 21913 26617 21947
rect 26617 21913 26651 21947
rect 26651 21913 26660 21947
rect 26608 21904 26660 21913
rect 26792 21947 26844 21956
rect 26792 21913 26801 21947
rect 26801 21913 26835 21947
rect 26835 21913 26844 21947
rect 26792 21904 26844 21913
rect 22100 21836 22152 21888
rect 22192 21836 22244 21888
rect 23572 21879 23624 21888
rect 23572 21845 23581 21879
rect 23581 21845 23615 21879
rect 23615 21845 23624 21879
rect 23572 21836 23624 21845
rect 23664 21836 23716 21888
rect 24676 21836 24728 21888
rect 26332 21836 26384 21888
rect 31208 21972 31260 22024
rect 31760 21972 31812 22024
rect 32312 21972 32364 22024
rect 33140 21972 33192 22024
rect 33324 21972 33376 22024
rect 37556 22049 37565 22083
rect 37565 22049 37599 22083
rect 37599 22049 37608 22083
rect 37556 22040 37608 22049
rect 38660 22108 38712 22160
rect 38752 22108 38804 22160
rect 41052 22108 41104 22160
rect 36912 22015 36964 22024
rect 36912 21981 36921 22015
rect 36921 21981 36955 22015
rect 36955 21981 36964 22015
rect 36912 21972 36964 21981
rect 37096 21972 37148 22024
rect 38614 21972 38666 22024
rect 39028 21972 39080 22024
rect 40040 22015 40092 22024
rect 40040 21981 40049 22015
rect 40049 21981 40083 22015
rect 40083 21981 40092 22015
rect 40040 21972 40092 21981
rect 40408 22015 40460 22024
rect 40408 21981 40417 22015
rect 40417 21981 40451 22015
rect 40451 21981 40460 22015
rect 40408 21972 40460 21981
rect 40592 21972 40644 22024
rect 40960 21972 41012 22024
rect 41144 21972 41196 22024
rect 43352 22185 43361 22219
rect 43361 22185 43395 22219
rect 43395 22185 43404 22219
rect 43352 22176 43404 22185
rect 41512 22040 41564 22092
rect 42800 22083 42852 22092
rect 42800 22049 42809 22083
rect 42809 22049 42843 22083
rect 42843 22049 42852 22083
rect 42800 22040 42852 22049
rect 41328 21972 41380 22024
rect 42064 22015 42116 22024
rect 42064 21981 42073 22015
rect 42073 21981 42107 22015
rect 42107 21981 42116 22015
rect 42064 21972 42116 21981
rect 42248 22015 42300 22024
rect 42248 21981 42257 22015
rect 42257 21981 42291 22015
rect 42291 21981 42300 22015
rect 42248 21972 42300 21981
rect 53564 21972 53616 22024
rect 54208 22015 54260 22024
rect 54208 21981 54217 22015
rect 54217 21981 54251 22015
rect 54251 21981 54260 22015
rect 54208 21972 54260 21981
rect 27804 21836 27856 21888
rect 28816 21879 28868 21888
rect 28816 21845 28825 21879
rect 28825 21845 28859 21879
rect 28859 21845 28868 21879
rect 28816 21836 28868 21845
rect 29828 21836 29880 21888
rect 30472 21879 30524 21888
rect 30472 21845 30481 21879
rect 30481 21845 30515 21879
rect 30515 21845 30524 21879
rect 30472 21836 30524 21845
rect 31392 21879 31444 21888
rect 31392 21845 31401 21879
rect 31401 21845 31435 21879
rect 31435 21845 31444 21879
rect 31392 21836 31444 21845
rect 31576 21836 31628 21888
rect 32588 21879 32640 21888
rect 32588 21845 32597 21879
rect 32597 21845 32631 21879
rect 32631 21845 32640 21879
rect 32588 21836 32640 21845
rect 33692 21836 33744 21888
rect 34704 21836 34756 21888
rect 35440 21836 35492 21888
rect 39948 21904 40000 21956
rect 40224 21947 40276 21956
rect 40224 21913 40233 21947
rect 40233 21913 40267 21947
rect 40267 21913 40276 21947
rect 40224 21904 40276 21913
rect 42340 21904 42392 21956
rect 53288 21947 53340 21956
rect 53288 21913 53297 21947
rect 53297 21913 53331 21947
rect 53331 21913 53340 21947
rect 53288 21904 53340 21913
rect 53472 21947 53524 21956
rect 53472 21913 53481 21947
rect 53481 21913 53515 21947
rect 53515 21913 53524 21947
rect 53472 21904 53524 21913
rect 54024 21947 54076 21956
rect 54024 21913 54033 21947
rect 54033 21913 54067 21947
rect 54067 21913 54076 21947
rect 54024 21904 54076 21913
rect 37464 21836 37516 21888
rect 38660 21836 38712 21888
rect 40132 21836 40184 21888
rect 41052 21836 41104 21888
rect 43720 21836 43772 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 2412 21675 2464 21684
rect 2412 21641 2421 21675
rect 2421 21641 2455 21675
rect 2455 21641 2464 21675
rect 2412 21632 2464 21641
rect 2504 21632 2556 21684
rect 23572 21632 23624 21684
rect 22284 21564 22336 21616
rect 2412 21496 2464 21548
rect 14096 21539 14148 21548
rect 14096 21505 14105 21539
rect 14105 21505 14139 21539
rect 14139 21505 14148 21539
rect 14096 21496 14148 21505
rect 21364 21428 21416 21480
rect 23664 21496 23716 21548
rect 24584 21564 24636 21616
rect 25044 21564 25096 21616
rect 27528 21632 27580 21684
rect 29828 21632 29880 21684
rect 31668 21632 31720 21684
rect 35440 21675 35492 21684
rect 35440 21641 35449 21675
rect 35449 21641 35483 21675
rect 35483 21641 35492 21675
rect 35440 21632 35492 21641
rect 36084 21632 36136 21684
rect 26148 21564 26200 21616
rect 27804 21496 27856 21548
rect 21180 21360 21232 21412
rect 26516 21428 26568 21480
rect 27436 21428 27488 21480
rect 29368 21496 29420 21548
rect 30288 21496 30340 21548
rect 31208 21496 31260 21548
rect 32496 21496 32548 21548
rect 28540 21471 28592 21480
rect 28540 21437 28549 21471
rect 28549 21437 28583 21471
rect 28583 21437 28592 21471
rect 28540 21428 28592 21437
rect 28632 21471 28684 21480
rect 28632 21437 28641 21471
rect 28641 21437 28675 21471
rect 28675 21437 28684 21471
rect 28632 21428 28684 21437
rect 28816 21428 28868 21480
rect 32404 21471 32456 21480
rect 32404 21437 32413 21471
rect 32413 21437 32447 21471
rect 32447 21437 32456 21471
rect 32404 21428 32456 21437
rect 1676 21335 1728 21344
rect 1676 21301 1685 21335
rect 1685 21301 1719 21335
rect 1719 21301 1728 21335
rect 1676 21292 1728 21301
rect 13912 21335 13964 21344
rect 13912 21301 13921 21335
rect 13921 21301 13955 21335
rect 13955 21301 13964 21335
rect 13912 21292 13964 21301
rect 18144 21292 18196 21344
rect 22100 21292 22152 21344
rect 22376 21335 22428 21344
rect 22376 21301 22385 21335
rect 22385 21301 22419 21335
rect 22419 21301 22428 21335
rect 22376 21292 22428 21301
rect 22836 21292 22888 21344
rect 23296 21292 23348 21344
rect 26884 21360 26936 21412
rect 28724 21360 28776 21412
rect 25136 21292 25188 21344
rect 25504 21292 25556 21344
rect 27620 21292 27672 21344
rect 29092 21335 29144 21344
rect 29092 21301 29101 21335
rect 29101 21301 29135 21335
rect 29135 21301 29144 21335
rect 29092 21292 29144 21301
rect 30104 21292 30156 21344
rect 30932 21292 30984 21344
rect 31852 21360 31904 21412
rect 32036 21360 32088 21412
rect 36360 21564 36412 21616
rect 35532 21539 35584 21548
rect 35532 21505 35541 21539
rect 35541 21505 35575 21539
rect 35575 21505 35584 21539
rect 35532 21496 35584 21505
rect 36176 21496 36228 21548
rect 34704 21471 34756 21480
rect 34704 21437 34713 21471
rect 34713 21437 34747 21471
rect 34747 21437 34756 21471
rect 34704 21428 34756 21437
rect 34796 21428 34848 21480
rect 36728 21539 36780 21548
rect 36728 21505 36737 21539
rect 36737 21505 36771 21539
rect 36771 21505 36780 21539
rect 38568 21539 38620 21548
rect 36728 21496 36780 21505
rect 38568 21505 38586 21539
rect 38586 21505 38620 21539
rect 38568 21496 38620 21505
rect 38844 21539 38896 21548
rect 38844 21505 38853 21539
rect 38853 21505 38887 21539
rect 38887 21505 38896 21539
rect 38844 21496 38896 21505
rect 39212 21632 39264 21684
rect 39764 21607 39816 21616
rect 39764 21573 39773 21607
rect 39773 21573 39807 21607
rect 39807 21573 39816 21607
rect 39764 21564 39816 21573
rect 42064 21632 42116 21684
rect 42248 21632 42300 21684
rect 42708 21632 42760 21684
rect 53564 21675 53616 21684
rect 53564 21641 53573 21675
rect 53573 21641 53607 21675
rect 53607 21641 53616 21675
rect 53564 21632 53616 21641
rect 54208 21675 54260 21684
rect 54208 21641 54217 21675
rect 54217 21641 54251 21675
rect 54251 21641 54260 21675
rect 54208 21632 54260 21641
rect 39948 21564 40000 21616
rect 37372 21428 37424 21480
rect 39120 21428 39172 21480
rect 40408 21496 40460 21548
rect 42708 21496 42760 21548
rect 40224 21428 40276 21480
rect 40684 21471 40736 21480
rect 40684 21437 40693 21471
rect 40693 21437 40727 21471
rect 40727 21437 40736 21471
rect 40684 21428 40736 21437
rect 36912 21403 36964 21412
rect 36912 21369 36921 21403
rect 36921 21369 36955 21403
rect 36955 21369 36964 21403
rect 36912 21360 36964 21369
rect 41696 21360 41748 21412
rect 32864 21292 32916 21344
rect 35900 21292 35952 21344
rect 36544 21292 36596 21344
rect 37464 21335 37516 21344
rect 37464 21301 37473 21335
rect 37473 21301 37507 21335
rect 37507 21301 37516 21335
rect 37464 21292 37516 21301
rect 37648 21292 37700 21344
rect 41788 21292 41840 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2412 21131 2464 21140
rect 2412 21097 2421 21131
rect 2421 21097 2455 21131
rect 2455 21097 2464 21131
rect 2412 21088 2464 21097
rect 21364 21088 21416 21140
rect 23296 21088 23348 21140
rect 19984 21020 20036 21072
rect 26332 21088 26384 21140
rect 26608 21131 26660 21140
rect 26608 21097 26617 21131
rect 26617 21097 26651 21131
rect 26651 21097 26660 21131
rect 26608 21088 26660 21097
rect 26884 21088 26936 21140
rect 32588 21088 32640 21140
rect 34612 21088 34664 21140
rect 28632 21020 28684 21072
rect 29092 21020 29144 21072
rect 35900 21088 35952 21140
rect 37556 21088 37608 21140
rect 38568 21088 38620 21140
rect 43996 21131 44048 21140
rect 22376 20952 22428 21004
rect 13912 20884 13964 20936
rect 23848 20927 23900 20936
rect 23848 20893 23857 20927
rect 23857 20893 23891 20927
rect 23891 20893 23900 20927
rect 23848 20884 23900 20893
rect 1676 20791 1728 20800
rect 1676 20757 1685 20791
rect 1685 20757 1719 20791
rect 1719 20757 1728 20791
rect 1676 20748 1728 20757
rect 21456 20791 21508 20800
rect 21456 20757 21465 20791
rect 21465 20757 21499 20791
rect 21499 20757 21508 20791
rect 24400 20884 24452 20936
rect 24584 20927 24636 20936
rect 24584 20893 24593 20927
rect 24593 20893 24627 20927
rect 24627 20893 24636 20927
rect 24584 20884 24636 20893
rect 27068 20952 27120 21004
rect 28540 20995 28592 21004
rect 21456 20748 21508 20757
rect 28540 20961 28549 20995
rect 28549 20961 28583 20995
rect 28583 20961 28592 20995
rect 28540 20952 28592 20961
rect 31300 20952 31352 21004
rect 32312 20995 32364 21004
rect 32312 20961 32321 20995
rect 32321 20961 32355 20995
rect 32355 20961 32364 20995
rect 32312 20952 32364 20961
rect 33784 20995 33836 21004
rect 33784 20961 33793 20995
rect 33793 20961 33827 20995
rect 33827 20961 33836 20995
rect 33784 20952 33836 20961
rect 25136 20748 25188 20800
rect 26516 20748 26568 20800
rect 28632 20859 28684 20868
rect 28632 20825 28641 20859
rect 28641 20825 28675 20859
rect 28675 20825 28684 20859
rect 28632 20816 28684 20825
rect 30012 20884 30064 20936
rect 30288 20927 30340 20936
rect 30288 20893 30297 20927
rect 30297 20893 30331 20927
rect 30331 20893 30340 20927
rect 30288 20884 30340 20893
rect 32036 20884 32088 20936
rect 32864 20884 32916 20936
rect 35348 20952 35400 21004
rect 35900 20952 35952 21004
rect 36360 20952 36412 21004
rect 37004 20884 37056 20936
rect 43996 21097 44005 21131
rect 44005 21097 44039 21131
rect 44039 21097 44048 21131
rect 43996 21088 44048 21097
rect 54208 21063 54260 21072
rect 34704 20816 34756 20868
rect 35716 20816 35768 20868
rect 38200 20859 38252 20868
rect 29736 20791 29788 20800
rect 29736 20757 29745 20791
rect 29745 20757 29779 20791
rect 29779 20757 29788 20791
rect 29736 20748 29788 20757
rect 30196 20748 30248 20800
rect 32864 20748 32916 20800
rect 34612 20748 34664 20800
rect 34796 20748 34848 20800
rect 38200 20825 38209 20859
rect 38209 20825 38243 20859
rect 38243 20825 38252 20859
rect 38200 20816 38252 20825
rect 38752 20816 38804 20868
rect 39120 20859 39172 20868
rect 39120 20825 39129 20859
rect 39129 20825 39163 20859
rect 39163 20825 39172 20859
rect 39120 20816 39172 20825
rect 39304 20893 39313 20912
rect 39313 20893 39347 20912
rect 39347 20893 39356 20912
rect 39304 20860 39356 20893
rect 40132 20884 40184 20936
rect 40684 20884 40736 20936
rect 42340 20884 42392 20936
rect 43444 20927 43496 20936
rect 43444 20893 43453 20927
rect 43453 20893 43487 20927
rect 43487 20893 43496 20927
rect 43444 20884 43496 20893
rect 54208 21029 54217 21063
rect 54217 21029 54251 21063
rect 54251 21029 54260 21063
rect 54208 21020 54260 21029
rect 36544 20748 36596 20800
rect 39304 20748 39356 20800
rect 42248 20748 42300 20800
rect 42708 20748 42760 20800
rect 53564 20791 53616 20800
rect 53564 20757 53573 20791
rect 53573 20757 53607 20791
rect 53607 20757 53616 20791
rect 53564 20748 53616 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 23848 20544 23900 20596
rect 19616 20408 19668 20460
rect 18972 20340 19024 20392
rect 21456 20340 21508 20392
rect 22192 20451 22244 20460
rect 22192 20417 22201 20451
rect 22201 20417 22235 20451
rect 22235 20417 22244 20451
rect 22192 20408 22244 20417
rect 24400 20544 24452 20596
rect 26516 20544 26568 20596
rect 27160 20587 27212 20596
rect 27160 20553 27169 20587
rect 27169 20553 27203 20587
rect 27203 20553 27212 20587
rect 27160 20544 27212 20553
rect 27804 20587 27856 20596
rect 27804 20553 27813 20587
rect 27813 20553 27847 20587
rect 27847 20553 27856 20587
rect 27804 20544 27856 20553
rect 28816 20544 28868 20596
rect 29644 20544 29696 20596
rect 30288 20544 30340 20596
rect 37464 20544 37516 20596
rect 40684 20544 40736 20596
rect 24860 20476 24912 20528
rect 25136 20408 25188 20460
rect 25780 20476 25832 20528
rect 25320 20408 25372 20460
rect 26608 20408 26660 20460
rect 29828 20476 29880 20528
rect 30104 20476 30156 20528
rect 42800 20544 42852 20596
rect 23480 20340 23532 20392
rect 24216 20340 24268 20392
rect 25044 20340 25096 20392
rect 26792 20340 26844 20392
rect 29092 20408 29144 20460
rect 29184 20451 29236 20460
rect 29184 20417 29193 20451
rect 29193 20417 29227 20451
rect 29227 20417 29236 20451
rect 29184 20408 29236 20417
rect 29644 20408 29696 20460
rect 30012 20451 30064 20460
rect 30012 20417 30021 20451
rect 30021 20417 30055 20451
rect 30055 20417 30064 20451
rect 30012 20408 30064 20417
rect 34152 20408 34204 20460
rect 34428 20408 34480 20460
rect 34612 20408 34664 20460
rect 35348 20408 35400 20460
rect 36728 20451 36780 20460
rect 27528 20340 27580 20392
rect 32220 20340 32272 20392
rect 33600 20383 33652 20392
rect 20536 20272 20588 20324
rect 22836 20272 22888 20324
rect 30012 20272 30064 20324
rect 30472 20272 30524 20324
rect 33600 20349 33609 20383
rect 33609 20349 33643 20383
rect 33643 20349 33652 20383
rect 33600 20340 33652 20349
rect 34336 20340 34388 20392
rect 36728 20417 36737 20451
rect 36737 20417 36771 20451
rect 36771 20417 36780 20451
rect 36728 20408 36780 20417
rect 37188 20408 37240 20460
rect 54208 20519 54260 20528
rect 54208 20485 54217 20519
rect 54217 20485 54251 20519
rect 54251 20485 54260 20519
rect 54208 20476 54260 20485
rect 41512 20451 41564 20460
rect 37096 20340 37148 20392
rect 38752 20340 38804 20392
rect 38936 20340 38988 20392
rect 1676 20247 1728 20256
rect 1676 20213 1685 20247
rect 1685 20213 1719 20247
rect 1719 20213 1728 20247
rect 1676 20204 1728 20213
rect 19248 20247 19300 20256
rect 19248 20213 19257 20247
rect 19257 20213 19291 20247
rect 19291 20213 19300 20247
rect 19248 20204 19300 20213
rect 20628 20204 20680 20256
rect 29460 20204 29512 20256
rect 29644 20204 29696 20256
rect 34244 20247 34296 20256
rect 34244 20213 34253 20247
rect 34253 20213 34287 20247
rect 34287 20213 34296 20247
rect 34244 20204 34296 20213
rect 36820 20272 36872 20324
rect 39396 20272 39448 20324
rect 39488 20204 39540 20256
rect 40500 20340 40552 20392
rect 41512 20417 41521 20451
rect 41521 20417 41555 20451
rect 41555 20417 41564 20451
rect 41512 20408 41564 20417
rect 41788 20451 41840 20460
rect 41328 20272 41380 20324
rect 41788 20417 41797 20451
rect 41797 20417 41831 20451
rect 41831 20417 41840 20451
rect 41788 20408 41840 20417
rect 43720 20451 43772 20460
rect 43720 20417 43729 20451
rect 43729 20417 43763 20451
rect 43763 20417 43772 20451
rect 43720 20408 43772 20417
rect 53288 20451 53340 20460
rect 53288 20417 53297 20451
rect 53297 20417 53331 20451
rect 53331 20417 53340 20451
rect 53288 20408 53340 20417
rect 53564 20408 53616 20460
rect 42616 20247 42668 20256
rect 42616 20213 42625 20247
rect 42625 20213 42659 20247
rect 42659 20213 42668 20247
rect 42616 20204 42668 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2504 20000 2556 20052
rect 19616 20043 19668 20052
rect 19616 20009 19625 20043
rect 19625 20009 19659 20043
rect 19659 20009 19668 20043
rect 19616 20000 19668 20009
rect 21272 20000 21324 20052
rect 20812 19932 20864 19984
rect 21916 19932 21968 19984
rect 15844 19864 15896 19916
rect 20168 19864 20220 19916
rect 21272 19864 21324 19916
rect 14464 19839 14516 19848
rect 14464 19805 14473 19839
rect 14473 19805 14507 19839
rect 14507 19805 14516 19839
rect 14464 19796 14516 19805
rect 19984 19839 20036 19848
rect 19984 19805 19993 19839
rect 19993 19805 20027 19839
rect 20027 19805 20036 19839
rect 19984 19796 20036 19805
rect 24768 20000 24820 20052
rect 26148 20000 26200 20052
rect 27620 20000 27672 20052
rect 30012 20000 30064 20052
rect 29736 19932 29788 19984
rect 22836 19864 22888 19916
rect 24860 19864 24912 19916
rect 25136 19907 25188 19916
rect 25136 19873 25145 19907
rect 25145 19873 25179 19907
rect 25179 19873 25188 19907
rect 25136 19864 25188 19873
rect 25780 19907 25832 19916
rect 25780 19873 25789 19907
rect 25789 19873 25823 19907
rect 25823 19873 25832 19907
rect 25780 19864 25832 19873
rect 29184 19864 29236 19916
rect 30288 19864 30340 19916
rect 30840 19907 30892 19916
rect 30840 19873 30849 19907
rect 30849 19873 30883 19907
rect 30883 19873 30892 19907
rect 30840 19864 30892 19873
rect 22284 19728 22336 19780
rect 1676 19703 1728 19712
rect 1676 19669 1685 19703
rect 1685 19669 1719 19703
rect 1719 19669 1728 19703
rect 1676 19660 1728 19669
rect 14280 19703 14332 19712
rect 14280 19669 14289 19703
rect 14289 19669 14323 19703
rect 14323 19669 14332 19703
rect 14280 19660 14332 19669
rect 20076 19703 20128 19712
rect 20076 19669 20085 19703
rect 20085 19669 20119 19703
rect 20119 19669 20128 19703
rect 20076 19660 20128 19669
rect 20812 19703 20864 19712
rect 20812 19669 20821 19703
rect 20821 19669 20855 19703
rect 20855 19669 20864 19703
rect 20812 19660 20864 19669
rect 21548 19703 21600 19712
rect 21548 19669 21557 19703
rect 21557 19669 21591 19703
rect 21591 19669 21600 19703
rect 21548 19660 21600 19669
rect 22100 19660 22152 19712
rect 25044 19703 25096 19712
rect 25044 19669 25053 19703
rect 25053 19669 25087 19703
rect 25087 19669 25096 19703
rect 25044 19660 25096 19669
rect 26056 19771 26108 19780
rect 26056 19737 26090 19771
rect 26090 19737 26108 19771
rect 27804 19796 27856 19848
rect 28448 19796 28500 19848
rect 29828 19796 29880 19848
rect 30748 19796 30800 19848
rect 31116 19839 31168 19848
rect 31116 19805 31150 19839
rect 31150 19805 31168 19839
rect 32312 20000 32364 20052
rect 35532 20000 35584 20052
rect 32496 19932 32548 19984
rect 39396 20000 39448 20052
rect 42064 20000 42116 20052
rect 43444 20000 43496 20052
rect 54208 20043 54260 20052
rect 54208 20009 54217 20043
rect 54217 20009 54251 20043
rect 54251 20009 54260 20043
rect 54208 20000 54260 20009
rect 37464 19975 37516 19984
rect 37464 19941 37473 19975
rect 37473 19941 37507 19975
rect 37507 19941 37516 19975
rect 37464 19932 37516 19941
rect 37832 19932 37884 19984
rect 53564 19975 53616 19984
rect 53564 19941 53573 19975
rect 53573 19941 53607 19975
rect 53607 19941 53616 19975
rect 53564 19932 53616 19941
rect 38844 19907 38896 19916
rect 31116 19796 31168 19805
rect 34336 19796 34388 19848
rect 36268 19839 36320 19848
rect 36268 19805 36277 19839
rect 36277 19805 36311 19839
rect 36311 19805 36320 19839
rect 36268 19796 36320 19805
rect 26056 19728 26108 19737
rect 26148 19660 26200 19712
rect 29552 19660 29604 19712
rect 30288 19660 30340 19712
rect 34796 19660 34848 19712
rect 38844 19873 38853 19907
rect 38853 19873 38887 19907
rect 38887 19873 38896 19907
rect 38844 19864 38896 19873
rect 36820 19796 36872 19848
rect 37004 19796 37056 19848
rect 39488 19839 39540 19848
rect 39488 19805 39497 19839
rect 39497 19805 39531 19839
rect 39531 19805 39540 19839
rect 39488 19796 39540 19805
rect 40316 19728 40368 19780
rect 41144 19728 41196 19780
rect 41420 19728 41472 19780
rect 38108 19660 38160 19712
rect 40132 19660 40184 19712
rect 40776 19660 40828 19712
rect 40960 19660 41012 19712
rect 42248 19839 42300 19848
rect 42248 19805 42257 19839
rect 42257 19805 42291 19839
rect 42291 19805 42300 19839
rect 42248 19796 42300 19805
rect 44732 19796 44784 19848
rect 42708 19728 42760 19780
rect 42616 19660 42668 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 17040 19456 17092 19508
rect 20076 19499 20128 19508
rect 20076 19465 20085 19499
rect 20085 19465 20119 19499
rect 20119 19465 20128 19499
rect 20076 19456 20128 19465
rect 20168 19456 20220 19508
rect 22284 19456 22336 19508
rect 22560 19456 22612 19508
rect 26056 19456 26108 19508
rect 26516 19456 26568 19508
rect 28080 19456 28132 19508
rect 14280 19320 14332 19372
rect 19340 19388 19392 19440
rect 22468 19388 22520 19440
rect 19248 19320 19300 19372
rect 1676 19159 1728 19168
rect 1676 19125 1685 19159
rect 1685 19125 1719 19159
rect 1719 19125 1728 19159
rect 1676 19116 1728 19125
rect 20628 19320 20680 19372
rect 21548 19320 21600 19372
rect 23480 19388 23532 19440
rect 24584 19388 24636 19440
rect 25044 19388 25096 19440
rect 28356 19388 28408 19440
rect 24124 19363 24176 19372
rect 24124 19329 24133 19363
rect 24133 19329 24167 19363
rect 24167 19329 24176 19363
rect 24124 19320 24176 19329
rect 24216 19363 24268 19372
rect 24216 19329 24225 19363
rect 24225 19329 24259 19363
rect 24259 19329 24268 19363
rect 27528 19363 27580 19372
rect 24216 19320 24268 19329
rect 27528 19329 27537 19363
rect 27537 19329 27571 19363
rect 27571 19329 27580 19363
rect 27528 19320 27580 19329
rect 27620 19320 27672 19372
rect 28448 19320 28500 19372
rect 29092 19456 29144 19508
rect 30472 19499 30524 19508
rect 30472 19465 30481 19499
rect 30481 19465 30515 19499
rect 30515 19465 30524 19499
rect 30472 19456 30524 19465
rect 29920 19388 29972 19440
rect 31208 19456 31260 19508
rect 32220 19456 32272 19508
rect 35716 19499 35768 19508
rect 35716 19465 35725 19499
rect 35725 19465 35759 19499
rect 35759 19465 35768 19499
rect 35716 19456 35768 19465
rect 36728 19456 36780 19508
rect 37832 19456 37884 19508
rect 38108 19499 38160 19508
rect 38108 19465 38117 19499
rect 38117 19465 38151 19499
rect 38151 19465 38160 19499
rect 38108 19456 38160 19465
rect 38752 19456 38804 19508
rect 30748 19388 30800 19440
rect 29092 19320 29144 19372
rect 29552 19363 29604 19372
rect 29552 19329 29561 19363
rect 29561 19329 29595 19363
rect 29595 19329 29604 19363
rect 29552 19320 29604 19329
rect 21180 19295 21232 19304
rect 21180 19261 21189 19295
rect 21189 19261 21223 19295
rect 21223 19261 21232 19295
rect 21180 19252 21232 19261
rect 21272 19295 21324 19304
rect 21272 19261 21281 19295
rect 21281 19261 21315 19295
rect 21315 19261 21324 19295
rect 21272 19252 21324 19261
rect 24952 19252 25004 19304
rect 26516 19295 26568 19304
rect 26516 19261 26525 19295
rect 26525 19261 26559 19295
rect 26559 19261 26568 19295
rect 26516 19252 26568 19261
rect 27804 19252 27856 19304
rect 21456 19184 21508 19236
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 28264 19184 28316 19236
rect 29184 19252 29236 19304
rect 30196 19184 30248 19236
rect 23572 19116 23624 19168
rect 23664 19116 23716 19168
rect 28448 19116 28500 19168
rect 31116 19320 31168 19372
rect 31392 19320 31444 19372
rect 31024 19295 31076 19304
rect 31024 19261 31033 19295
rect 31033 19261 31067 19295
rect 31067 19261 31076 19295
rect 31024 19252 31076 19261
rect 31668 19320 31720 19372
rect 32128 19252 32180 19304
rect 34244 19388 34296 19440
rect 37280 19388 37332 19440
rect 39856 19456 39908 19508
rect 41420 19456 41472 19508
rect 54208 19499 54260 19508
rect 54208 19465 54217 19499
rect 54217 19465 54251 19499
rect 54251 19465 54260 19499
rect 54208 19456 54260 19465
rect 40776 19431 40828 19440
rect 33140 19320 33192 19372
rect 39304 19363 39356 19372
rect 34336 19295 34388 19304
rect 34336 19261 34345 19295
rect 34345 19261 34379 19295
rect 34379 19261 34388 19295
rect 34336 19252 34388 19261
rect 35992 19252 36044 19304
rect 36268 19252 36320 19304
rect 37372 19252 37424 19304
rect 38292 19295 38344 19304
rect 38292 19261 38301 19295
rect 38301 19261 38335 19295
rect 38335 19261 38344 19295
rect 39304 19329 39313 19363
rect 39313 19329 39347 19363
rect 39347 19329 39356 19363
rect 39304 19320 39356 19329
rect 38292 19252 38344 19261
rect 33692 19184 33744 19236
rect 32312 19116 32364 19168
rect 33416 19116 33468 19168
rect 37096 19184 37148 19236
rect 39212 19184 39264 19236
rect 40776 19397 40785 19431
rect 40785 19397 40819 19431
rect 40819 19397 40828 19431
rect 40776 19388 40828 19397
rect 38660 19116 38712 19168
rect 40408 19252 40460 19304
rect 41144 19320 41196 19372
rect 41236 19252 41288 19304
rect 44732 19388 44784 19440
rect 41604 19320 41656 19372
rect 40040 19184 40092 19236
rect 40132 19116 40184 19168
rect 42340 19116 42392 19168
rect 42616 19159 42668 19168
rect 42616 19125 42625 19159
rect 42625 19125 42659 19159
rect 42659 19125 42668 19159
rect 42616 19116 42668 19125
rect 54208 19116 54260 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2596 18912 2648 18964
rect 25320 18912 25372 18964
rect 26516 18955 26568 18964
rect 26516 18921 26525 18955
rect 26525 18921 26559 18955
rect 26559 18921 26568 18955
rect 26516 18912 26568 18921
rect 28632 18912 28684 18964
rect 29184 18912 29236 18964
rect 32036 18912 32088 18964
rect 34336 18955 34388 18964
rect 34336 18921 34345 18955
rect 34345 18921 34379 18955
rect 34379 18921 34388 18955
rect 34336 18912 34388 18921
rect 35992 18955 36044 18964
rect 35992 18921 36001 18955
rect 36001 18921 36035 18955
rect 36035 18921 36044 18955
rect 35992 18912 36044 18921
rect 36912 18912 36964 18964
rect 37096 18912 37148 18964
rect 40040 18955 40092 18964
rect 15476 18844 15528 18896
rect 21180 18844 21232 18896
rect 28448 18844 28500 18896
rect 33048 18844 33100 18896
rect 34888 18887 34940 18896
rect 22468 18819 22520 18828
rect 22468 18785 22477 18819
rect 22477 18785 22511 18819
rect 22511 18785 22520 18819
rect 22468 18776 22520 18785
rect 23940 18776 23992 18828
rect 27160 18776 27212 18828
rect 20352 18708 20404 18760
rect 20720 18708 20772 18760
rect 23664 18751 23716 18760
rect 23664 18717 23673 18751
rect 23673 18717 23707 18751
rect 23707 18717 23716 18751
rect 23664 18708 23716 18717
rect 24676 18751 24728 18760
rect 24676 18717 24685 18751
rect 24685 18717 24719 18751
rect 24719 18717 24728 18751
rect 24676 18708 24728 18717
rect 27620 18776 27672 18828
rect 27804 18776 27856 18828
rect 28172 18708 28224 18760
rect 28356 18776 28408 18828
rect 30840 18776 30892 18828
rect 32864 18776 32916 18828
rect 33508 18819 33560 18828
rect 33508 18785 33517 18819
rect 33517 18785 33551 18819
rect 33551 18785 33560 18819
rect 34888 18853 34897 18887
rect 34897 18853 34931 18887
rect 34931 18853 34940 18887
rect 34888 18844 34940 18853
rect 35348 18844 35400 18896
rect 39304 18844 39356 18896
rect 40040 18921 40049 18955
rect 40049 18921 40083 18955
rect 40083 18921 40092 18955
rect 40040 18912 40092 18921
rect 41512 18844 41564 18896
rect 42524 18887 42576 18896
rect 42524 18853 42533 18887
rect 42533 18853 42567 18887
rect 42567 18853 42576 18887
rect 42524 18844 42576 18853
rect 33508 18776 33560 18785
rect 33876 18776 33928 18828
rect 36268 18819 36320 18828
rect 36268 18785 36277 18819
rect 36277 18785 36311 18819
rect 36311 18785 36320 18819
rect 36268 18776 36320 18785
rect 36912 18776 36964 18828
rect 37832 18776 37884 18828
rect 38660 18776 38712 18828
rect 30104 18708 30156 18760
rect 30288 18751 30340 18760
rect 30288 18717 30297 18751
rect 30297 18717 30331 18751
rect 30331 18717 30340 18751
rect 30288 18708 30340 18717
rect 31668 18751 31720 18760
rect 31668 18717 31702 18751
rect 31702 18717 31720 18751
rect 31668 18708 31720 18717
rect 32496 18708 32548 18760
rect 33784 18708 33836 18760
rect 34520 18708 34572 18760
rect 36176 18751 36228 18760
rect 36176 18717 36185 18751
rect 36185 18717 36219 18751
rect 36219 18717 36228 18751
rect 36176 18708 36228 18717
rect 36360 18751 36412 18760
rect 36360 18717 36369 18751
rect 36369 18717 36403 18751
rect 36403 18717 36412 18751
rect 36360 18708 36412 18717
rect 36636 18708 36688 18760
rect 38292 18751 38344 18760
rect 38292 18717 38301 18751
rect 38301 18717 38335 18751
rect 38335 18717 38344 18751
rect 38292 18708 38344 18717
rect 17224 18640 17276 18692
rect 20536 18640 20588 18692
rect 1676 18615 1728 18624
rect 1676 18581 1685 18615
rect 1685 18581 1719 18615
rect 1719 18581 1728 18615
rect 1676 18572 1728 18581
rect 18328 18615 18380 18624
rect 18328 18581 18337 18615
rect 18337 18581 18371 18615
rect 18371 18581 18380 18615
rect 18328 18572 18380 18581
rect 19432 18572 19484 18624
rect 27620 18640 27672 18692
rect 28356 18640 28408 18692
rect 28540 18640 28592 18692
rect 38844 18708 38896 18760
rect 40040 18776 40092 18828
rect 42708 18776 42760 18828
rect 39212 18708 39264 18760
rect 39304 18708 39356 18760
rect 41880 18708 41932 18760
rect 42064 18751 42116 18760
rect 42064 18717 42073 18751
rect 42073 18717 42107 18751
rect 42107 18717 42116 18751
rect 42064 18708 42116 18717
rect 54208 18751 54260 18760
rect 54208 18717 54217 18751
rect 54217 18717 54251 18751
rect 54251 18717 54260 18751
rect 54208 18708 54260 18717
rect 38660 18640 38712 18692
rect 25320 18615 25372 18624
rect 25320 18581 25329 18615
rect 25329 18581 25363 18615
rect 25363 18581 25372 18615
rect 25320 18572 25372 18581
rect 28264 18572 28316 18624
rect 30840 18615 30892 18624
rect 30840 18581 30849 18615
rect 30849 18581 30883 18615
rect 30883 18581 30892 18615
rect 30840 18572 30892 18581
rect 31852 18572 31904 18624
rect 32680 18572 32732 18624
rect 33692 18572 33744 18624
rect 38108 18615 38160 18624
rect 38108 18581 38117 18615
rect 38117 18581 38151 18615
rect 38151 18581 38160 18615
rect 38108 18572 38160 18581
rect 38292 18572 38344 18624
rect 40224 18640 40276 18692
rect 40500 18640 40552 18692
rect 40960 18640 41012 18692
rect 41420 18640 41472 18692
rect 49700 18640 49752 18692
rect 53472 18683 53524 18692
rect 53472 18649 53481 18683
rect 53481 18649 53515 18683
rect 53515 18649 53524 18683
rect 53472 18640 53524 18649
rect 39948 18572 40000 18624
rect 40316 18572 40368 18624
rect 42708 18572 42760 18624
rect 44088 18572 44140 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 18328 18368 18380 18420
rect 19340 18300 19392 18352
rect 20352 18368 20404 18420
rect 31392 18368 31444 18420
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 17960 18164 18012 18216
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22468 18232 22520 18241
rect 23480 18300 23532 18352
rect 23204 18232 23256 18284
rect 24860 18232 24912 18284
rect 26516 18300 26568 18352
rect 27436 18300 27488 18352
rect 28080 18343 28132 18352
rect 28080 18309 28089 18343
rect 28089 18309 28123 18343
rect 28123 18309 28132 18343
rect 28080 18300 28132 18309
rect 28356 18300 28408 18352
rect 28632 18300 28684 18352
rect 30104 18300 30156 18352
rect 30748 18343 30800 18352
rect 30748 18309 30757 18343
rect 30757 18309 30791 18343
rect 30791 18309 30800 18343
rect 30748 18300 30800 18309
rect 30932 18343 30984 18352
rect 30932 18309 30941 18343
rect 30941 18309 30975 18343
rect 30975 18309 30984 18343
rect 30932 18300 30984 18309
rect 31024 18300 31076 18352
rect 37832 18368 37884 18420
rect 38292 18368 38344 18420
rect 40132 18368 40184 18420
rect 40224 18368 40276 18420
rect 41512 18368 41564 18420
rect 41696 18368 41748 18420
rect 42616 18368 42668 18420
rect 43260 18411 43312 18420
rect 43260 18377 43269 18411
rect 43269 18377 43303 18411
rect 43303 18377 43312 18411
rect 43260 18368 43312 18377
rect 54208 18411 54260 18420
rect 54208 18377 54217 18411
rect 54217 18377 54251 18411
rect 54251 18377 54260 18411
rect 54208 18368 54260 18377
rect 25228 18275 25280 18284
rect 25228 18241 25262 18275
rect 25262 18241 25280 18275
rect 25228 18232 25280 18241
rect 27988 18232 28040 18284
rect 28540 18232 28592 18284
rect 20720 18164 20772 18216
rect 21272 18207 21324 18216
rect 21272 18173 21281 18207
rect 21281 18173 21315 18207
rect 21315 18173 21324 18207
rect 21272 18164 21324 18173
rect 22008 18164 22060 18216
rect 33508 18300 33560 18352
rect 34888 18300 34940 18352
rect 34980 18300 35032 18352
rect 53196 18300 53248 18352
rect 31760 18275 31812 18284
rect 31760 18241 31769 18275
rect 31769 18241 31803 18275
rect 31803 18241 31812 18275
rect 32496 18275 32548 18284
rect 31760 18232 31812 18241
rect 32496 18241 32505 18275
rect 32505 18241 32539 18275
rect 32539 18241 32548 18275
rect 32496 18232 32548 18241
rect 32680 18275 32732 18284
rect 32680 18241 32689 18275
rect 32689 18241 32723 18275
rect 32723 18241 32732 18275
rect 32680 18232 32732 18241
rect 32864 18275 32916 18284
rect 32864 18241 32873 18275
rect 32873 18241 32907 18275
rect 32907 18241 32916 18275
rect 32864 18232 32916 18241
rect 33876 18232 33928 18284
rect 34336 18232 34388 18284
rect 17224 18028 17276 18080
rect 18420 18028 18472 18080
rect 21640 18096 21692 18148
rect 33232 18164 33284 18216
rect 33600 18164 33652 18216
rect 36176 18232 36228 18284
rect 37648 18275 37700 18284
rect 37648 18241 37657 18275
rect 37657 18241 37691 18275
rect 37691 18241 37700 18275
rect 37648 18232 37700 18241
rect 27528 18096 27580 18148
rect 28632 18096 28684 18148
rect 20628 18028 20680 18080
rect 22652 18071 22704 18080
rect 22652 18037 22661 18071
rect 22661 18037 22695 18071
rect 22695 18037 22704 18071
rect 22652 18028 22704 18037
rect 24952 18028 25004 18080
rect 29276 18096 29328 18148
rect 33140 18096 33192 18148
rect 36544 18164 36596 18216
rect 38108 18164 38160 18216
rect 38936 18232 38988 18284
rect 39856 18275 39908 18284
rect 39856 18241 39865 18275
rect 39865 18241 39899 18275
rect 39899 18241 39908 18275
rect 39856 18232 39908 18241
rect 39948 18232 40000 18284
rect 41328 18232 41380 18284
rect 41604 18232 41656 18284
rect 41880 18232 41932 18284
rect 49884 18232 49936 18284
rect 39304 18164 39356 18216
rect 39764 18164 39816 18216
rect 40408 18164 40460 18216
rect 40500 18207 40552 18216
rect 40500 18173 40509 18207
rect 40509 18173 40543 18207
rect 40543 18173 40552 18207
rect 40500 18164 40552 18173
rect 35808 18139 35860 18148
rect 28816 18028 28868 18080
rect 30288 18028 30340 18080
rect 32312 18071 32364 18080
rect 32312 18037 32321 18071
rect 32321 18037 32355 18071
rect 32355 18037 32364 18071
rect 35808 18105 35817 18139
rect 35817 18105 35851 18139
rect 35851 18105 35860 18139
rect 35808 18096 35860 18105
rect 36820 18096 36872 18148
rect 32312 18028 32364 18037
rect 34428 18028 34480 18080
rect 36360 18028 36412 18080
rect 37832 18028 37884 18080
rect 38108 18028 38160 18080
rect 38292 18028 38344 18080
rect 38476 18096 38528 18148
rect 41696 18096 41748 18148
rect 41512 18028 41564 18080
rect 43260 18028 43312 18080
rect 53472 18071 53524 18080
rect 53472 18037 53481 18071
rect 53481 18037 53515 18071
rect 53515 18037 53524 18071
rect 53472 18028 53524 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 22468 17824 22520 17876
rect 24124 17824 24176 17876
rect 25044 17824 25096 17876
rect 18236 17731 18288 17740
rect 18236 17697 18245 17731
rect 18245 17697 18279 17731
rect 18279 17697 18288 17731
rect 18236 17688 18288 17697
rect 19340 17688 19392 17740
rect 15384 17620 15436 17672
rect 23204 17756 23256 17808
rect 23848 17756 23900 17808
rect 26884 17756 26936 17808
rect 27988 17824 28040 17876
rect 54116 17824 54168 17876
rect 34520 17756 34572 17808
rect 22008 17688 22060 17740
rect 21640 17663 21692 17672
rect 21640 17629 21649 17663
rect 21649 17629 21683 17663
rect 21683 17629 21692 17663
rect 21640 17620 21692 17629
rect 22560 17620 22612 17672
rect 18236 17552 18288 17604
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 17132 17527 17184 17536
rect 17132 17493 17141 17527
rect 17141 17493 17175 17527
rect 17175 17493 17184 17527
rect 17132 17484 17184 17493
rect 17684 17527 17736 17536
rect 17684 17493 17693 17527
rect 17693 17493 17727 17527
rect 17727 17493 17736 17527
rect 17684 17484 17736 17493
rect 19248 17484 19300 17536
rect 19432 17552 19484 17604
rect 24032 17688 24084 17740
rect 25136 17731 25188 17740
rect 25136 17697 25145 17731
rect 25145 17697 25179 17731
rect 25179 17697 25188 17731
rect 25136 17688 25188 17697
rect 27528 17731 27580 17740
rect 27528 17697 27537 17731
rect 27537 17697 27571 17731
rect 27571 17697 27580 17731
rect 27528 17688 27580 17697
rect 27712 17731 27764 17740
rect 27712 17697 27721 17731
rect 27721 17697 27755 17731
rect 27755 17697 27764 17731
rect 27712 17688 27764 17697
rect 28356 17688 28408 17740
rect 28908 17688 28960 17740
rect 29368 17688 29420 17740
rect 30104 17688 30156 17740
rect 30288 17688 30340 17740
rect 30380 17688 30432 17740
rect 33140 17688 33192 17740
rect 37004 17756 37056 17808
rect 38016 17756 38068 17808
rect 41328 17756 41380 17808
rect 41420 17756 41472 17808
rect 41604 17756 41656 17808
rect 35532 17731 35584 17740
rect 35532 17697 35541 17731
rect 35541 17697 35575 17731
rect 35575 17697 35584 17731
rect 35532 17688 35584 17697
rect 23388 17663 23440 17672
rect 23388 17629 23397 17663
rect 23397 17629 23431 17663
rect 23431 17629 23440 17663
rect 23388 17620 23440 17629
rect 24676 17620 24728 17672
rect 28816 17663 28868 17672
rect 24584 17552 24636 17604
rect 28816 17629 28825 17663
rect 28825 17629 28859 17663
rect 28859 17629 28868 17663
rect 28816 17620 28868 17629
rect 29460 17620 29512 17672
rect 20720 17484 20772 17536
rect 21732 17527 21784 17536
rect 21732 17493 21741 17527
rect 21741 17493 21775 17527
rect 21775 17493 21784 17527
rect 21732 17484 21784 17493
rect 21824 17484 21876 17536
rect 23848 17484 23900 17536
rect 24032 17527 24084 17536
rect 24032 17493 24041 17527
rect 24041 17493 24075 17527
rect 24075 17493 24084 17527
rect 24032 17484 24084 17493
rect 24124 17484 24176 17536
rect 24952 17527 25004 17536
rect 24952 17493 24961 17527
rect 24961 17493 24995 17527
rect 24995 17493 25004 17527
rect 24952 17484 25004 17493
rect 25044 17527 25096 17536
rect 25044 17493 25053 17527
rect 25053 17493 25087 17527
rect 25087 17493 25096 17527
rect 25044 17484 25096 17493
rect 26148 17484 26200 17536
rect 27896 17527 27948 17536
rect 27896 17493 27905 17527
rect 27905 17493 27939 17527
rect 27939 17493 27948 17527
rect 27896 17484 27948 17493
rect 27988 17484 28040 17536
rect 29092 17484 29144 17536
rect 29828 17484 29880 17536
rect 30380 17484 30432 17536
rect 31392 17620 31444 17672
rect 32312 17620 32364 17672
rect 34428 17620 34480 17672
rect 34520 17620 34572 17672
rect 35808 17620 35860 17672
rect 38108 17688 38160 17740
rect 40132 17688 40184 17740
rect 40224 17688 40276 17740
rect 49700 17756 49752 17808
rect 54208 17799 54260 17808
rect 54208 17765 54217 17799
rect 54217 17765 54251 17799
rect 54251 17765 54260 17799
rect 54208 17756 54260 17765
rect 37464 17620 37516 17672
rect 37924 17620 37976 17672
rect 38660 17663 38712 17672
rect 38660 17629 38669 17663
rect 38669 17629 38703 17663
rect 38703 17629 38712 17663
rect 38660 17620 38712 17629
rect 38844 17663 38896 17672
rect 38844 17629 38853 17663
rect 38853 17629 38887 17663
rect 38887 17629 38896 17663
rect 38844 17620 38896 17629
rect 39304 17620 39356 17672
rect 30748 17552 30800 17604
rect 31852 17527 31904 17536
rect 31852 17493 31861 17527
rect 31861 17493 31895 17527
rect 31895 17493 31904 17527
rect 31852 17484 31904 17493
rect 32404 17484 32456 17536
rect 34796 17484 34848 17536
rect 35164 17484 35216 17536
rect 35348 17527 35400 17536
rect 35348 17493 35357 17527
rect 35357 17493 35391 17527
rect 35391 17493 35400 17527
rect 35348 17484 35400 17493
rect 36084 17527 36136 17536
rect 36084 17493 36093 17527
rect 36093 17493 36127 17527
rect 36127 17493 36136 17527
rect 36084 17484 36136 17493
rect 36636 17527 36688 17536
rect 36636 17493 36645 17527
rect 36645 17493 36679 17527
rect 36679 17493 36688 17527
rect 36636 17484 36688 17493
rect 38476 17552 38528 17604
rect 38936 17595 38988 17604
rect 38936 17561 38945 17595
rect 38945 17561 38979 17595
rect 38979 17561 38988 17595
rect 40132 17595 40184 17604
rect 38936 17552 38988 17561
rect 40132 17561 40141 17595
rect 40141 17561 40175 17595
rect 40175 17561 40184 17595
rect 40132 17552 40184 17561
rect 40316 17663 40368 17672
rect 40316 17629 40325 17663
rect 40325 17629 40359 17663
rect 40359 17629 40368 17663
rect 40316 17620 40368 17629
rect 41144 17620 41196 17672
rect 41328 17620 41380 17672
rect 41696 17663 41748 17672
rect 41696 17629 41705 17663
rect 41705 17629 41739 17663
rect 41739 17629 41748 17663
rect 41696 17620 41748 17629
rect 39028 17484 39080 17536
rect 39120 17484 39172 17536
rect 39304 17484 39356 17536
rect 43260 17527 43312 17536
rect 43260 17493 43269 17527
rect 43269 17493 43303 17527
rect 43303 17493 43312 17527
rect 43260 17484 43312 17493
rect 54208 17484 54260 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 17224 17323 17276 17332
rect 17224 17289 17233 17323
rect 17233 17289 17267 17323
rect 17267 17289 17276 17323
rect 17224 17280 17276 17289
rect 19340 17280 19392 17332
rect 18144 17212 18196 17264
rect 21364 17212 21416 17264
rect 16488 17144 16540 17196
rect 17132 17144 17184 17196
rect 21824 17144 21876 17196
rect 24400 17280 24452 17332
rect 24676 17323 24728 17332
rect 24676 17289 24685 17323
rect 24685 17289 24719 17323
rect 24719 17289 24728 17323
rect 24676 17280 24728 17289
rect 22652 17212 22704 17264
rect 22376 17144 22428 17196
rect 18328 17119 18380 17128
rect 18328 17085 18337 17119
rect 18337 17085 18371 17119
rect 18371 17085 18380 17119
rect 18328 17076 18380 17085
rect 20904 17119 20956 17128
rect 20904 17085 20913 17119
rect 20913 17085 20947 17119
rect 20947 17085 20956 17119
rect 20904 17076 20956 17085
rect 20076 17008 20128 17060
rect 22192 17076 22244 17128
rect 23940 17144 23992 17196
rect 24676 17144 24728 17196
rect 27896 17280 27948 17332
rect 25412 17212 25464 17264
rect 25964 17212 26016 17264
rect 26148 17212 26200 17264
rect 26516 17212 26568 17264
rect 28448 17144 28500 17196
rect 28908 17144 28960 17196
rect 1676 16983 1728 16992
rect 1676 16949 1685 16983
rect 1685 16949 1719 16983
rect 1719 16949 1728 16983
rect 1676 16940 1728 16949
rect 16672 16940 16724 16992
rect 17684 16940 17736 16992
rect 22652 17008 22704 17060
rect 23756 17008 23808 17060
rect 24676 17008 24728 17060
rect 21824 16940 21876 16992
rect 24032 16940 24084 16992
rect 25228 16983 25280 16992
rect 25228 16949 25237 16983
rect 25237 16949 25271 16983
rect 25271 16949 25280 16983
rect 25228 16940 25280 16949
rect 27712 17119 27764 17128
rect 27712 17085 27721 17119
rect 27721 17085 27755 17119
rect 27755 17085 27764 17119
rect 27712 17076 27764 17085
rect 26884 17008 26936 17060
rect 29828 17076 29880 17128
rect 30748 17212 30800 17264
rect 33232 17212 33284 17264
rect 31024 17144 31076 17196
rect 36084 17212 36136 17264
rect 36912 17280 36964 17332
rect 37556 17323 37608 17332
rect 37556 17289 37565 17323
rect 37565 17289 37599 17323
rect 37599 17289 37608 17323
rect 37556 17280 37608 17289
rect 38568 17280 38620 17332
rect 38936 17280 38988 17332
rect 38660 17212 38712 17264
rect 39028 17212 39080 17264
rect 39764 17212 39816 17264
rect 54116 17323 54168 17332
rect 54116 17289 54125 17323
rect 54125 17289 54159 17323
rect 54159 17289 54168 17323
rect 54116 17280 54168 17289
rect 54208 17255 54260 17264
rect 54208 17221 54217 17255
rect 54217 17221 54251 17255
rect 54251 17221 54260 17255
rect 54208 17212 54260 17221
rect 34704 17076 34756 17128
rect 35992 17144 36044 17196
rect 39120 17144 39172 17196
rect 36820 17076 36872 17128
rect 37280 17076 37332 17128
rect 39212 17076 39264 17128
rect 40316 17076 40368 17128
rect 40868 17187 40920 17196
rect 40868 17153 40877 17187
rect 40877 17153 40911 17187
rect 40911 17153 40920 17187
rect 40868 17144 40920 17153
rect 41420 17076 41472 17128
rect 27712 16940 27764 16992
rect 32312 16983 32364 16992
rect 32312 16949 32321 16983
rect 32321 16949 32355 16983
rect 32355 16949 32364 16983
rect 32312 16940 32364 16949
rect 34520 17008 34572 17060
rect 53564 17144 53616 17196
rect 53288 17051 53340 17060
rect 35164 16940 35216 16992
rect 35900 16940 35952 16992
rect 36912 16940 36964 16992
rect 53288 17017 53297 17051
rect 53297 17017 53331 17051
rect 53331 17017 53340 17051
rect 53288 17008 53340 17017
rect 42064 16940 42116 16992
rect 42708 16983 42760 16992
rect 42708 16949 42717 16983
rect 42717 16949 42751 16983
rect 42751 16949 42760 16983
rect 42708 16940 42760 16949
rect 43260 16940 43312 16992
rect 44180 16940 44232 16992
rect 44456 16940 44508 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 18236 16736 18288 16788
rect 16120 16643 16172 16652
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 16764 16643 16816 16652
rect 16764 16609 16773 16643
rect 16773 16609 16807 16643
rect 16807 16609 16816 16643
rect 16764 16600 16816 16609
rect 16948 16600 17000 16652
rect 22192 16736 22244 16788
rect 22376 16779 22428 16788
rect 22376 16745 22385 16779
rect 22385 16745 22419 16779
rect 22419 16745 22428 16779
rect 22376 16736 22428 16745
rect 23112 16736 23164 16788
rect 23756 16736 23808 16788
rect 24124 16736 24176 16788
rect 24584 16779 24636 16788
rect 24584 16745 24593 16779
rect 24593 16745 24627 16779
rect 24627 16745 24636 16779
rect 24584 16736 24636 16745
rect 24676 16736 24728 16788
rect 29552 16736 29604 16788
rect 30380 16736 30432 16788
rect 31024 16779 31076 16788
rect 31024 16745 31033 16779
rect 31033 16745 31067 16779
rect 31067 16745 31076 16779
rect 31024 16736 31076 16745
rect 33140 16779 33192 16788
rect 33140 16745 33149 16779
rect 33149 16745 33183 16779
rect 33183 16745 33192 16779
rect 33140 16736 33192 16745
rect 16580 16532 16632 16584
rect 17224 16575 17276 16584
rect 17224 16541 17233 16575
rect 17233 16541 17267 16575
rect 17267 16541 17276 16575
rect 17224 16532 17276 16541
rect 14832 16464 14884 16516
rect 18236 16575 18288 16584
rect 18236 16541 18245 16575
rect 18245 16541 18279 16575
rect 18279 16541 18288 16575
rect 18236 16532 18288 16541
rect 22100 16532 22152 16584
rect 27436 16711 27488 16720
rect 27436 16677 27445 16711
rect 27445 16677 27479 16711
rect 27479 16677 27488 16711
rect 27436 16668 27488 16677
rect 29092 16668 29144 16720
rect 31576 16668 31628 16720
rect 25044 16643 25096 16652
rect 23756 16532 23808 16584
rect 24216 16532 24268 16584
rect 25044 16609 25053 16643
rect 25053 16609 25087 16643
rect 25087 16609 25096 16643
rect 25044 16600 25096 16609
rect 25136 16643 25188 16652
rect 25136 16609 25145 16643
rect 25145 16609 25179 16643
rect 25179 16609 25188 16643
rect 25136 16600 25188 16609
rect 25228 16532 25280 16584
rect 26240 16532 26292 16584
rect 27068 16532 27120 16584
rect 27804 16532 27856 16584
rect 29460 16600 29512 16652
rect 30288 16600 30340 16652
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 17960 16464 18012 16516
rect 20076 16396 20128 16448
rect 21640 16464 21692 16516
rect 22652 16464 22704 16516
rect 22192 16396 22244 16448
rect 24584 16464 24636 16516
rect 27528 16464 27580 16516
rect 27436 16396 27488 16448
rect 27620 16396 27672 16448
rect 28356 16464 28408 16516
rect 28632 16575 28684 16584
rect 28632 16541 28641 16575
rect 28641 16541 28675 16575
rect 28675 16541 28684 16575
rect 28632 16532 28684 16541
rect 29644 16532 29696 16584
rect 32956 16668 33008 16720
rect 36452 16736 36504 16788
rect 35348 16668 35400 16720
rect 37464 16736 37516 16788
rect 38016 16736 38068 16788
rect 38292 16736 38344 16788
rect 39396 16779 39448 16788
rect 39396 16745 39405 16779
rect 39405 16745 39439 16779
rect 39439 16745 39448 16779
rect 39396 16736 39448 16745
rect 41236 16736 41288 16788
rect 41512 16736 41564 16788
rect 53472 16736 53524 16788
rect 54208 16779 54260 16788
rect 54208 16745 54217 16779
rect 54217 16745 54251 16779
rect 54251 16745 54260 16779
rect 54208 16736 54260 16745
rect 41880 16711 41932 16720
rect 32312 16600 32364 16652
rect 33048 16600 33100 16652
rect 33416 16600 33468 16652
rect 33508 16600 33560 16652
rect 34888 16643 34940 16652
rect 34888 16609 34897 16643
rect 34897 16609 34931 16643
rect 34931 16609 34940 16643
rect 34888 16600 34940 16609
rect 35164 16600 35216 16652
rect 35900 16600 35952 16652
rect 36636 16600 36688 16652
rect 41880 16677 41889 16711
rect 41889 16677 41923 16711
rect 41923 16677 41932 16711
rect 41880 16668 41932 16677
rect 42892 16668 42944 16720
rect 53564 16711 53616 16720
rect 53564 16677 53573 16711
rect 53573 16677 53607 16711
rect 53607 16677 53616 16711
rect 53564 16668 53616 16677
rect 37832 16600 37884 16652
rect 40408 16600 40460 16652
rect 41420 16643 41472 16652
rect 41420 16609 41429 16643
rect 41429 16609 41463 16643
rect 41463 16609 41472 16643
rect 41420 16600 41472 16609
rect 43628 16643 43680 16652
rect 43628 16609 43637 16643
rect 43637 16609 43671 16643
rect 43671 16609 43680 16643
rect 43628 16600 43680 16609
rect 29920 16439 29972 16448
rect 29920 16405 29929 16439
rect 29929 16405 29963 16439
rect 29963 16405 29972 16439
rect 29920 16396 29972 16405
rect 30012 16396 30064 16448
rect 33600 16532 33652 16584
rect 34796 16532 34848 16584
rect 36360 16575 36412 16584
rect 36360 16541 36369 16575
rect 36369 16541 36403 16575
rect 36403 16541 36412 16575
rect 36360 16532 36412 16541
rect 37280 16575 37332 16584
rect 37280 16541 37289 16575
rect 37289 16541 37323 16575
rect 37323 16541 37332 16575
rect 37280 16532 37332 16541
rect 37464 16575 37516 16584
rect 37464 16541 37473 16575
rect 37473 16541 37507 16575
rect 37507 16541 37516 16575
rect 37464 16532 37516 16541
rect 38660 16532 38712 16584
rect 39304 16532 39356 16584
rect 41880 16532 41932 16584
rect 42064 16575 42116 16584
rect 42064 16541 42073 16575
rect 42073 16541 42107 16575
rect 42107 16541 42116 16575
rect 42064 16532 42116 16541
rect 42524 16575 42576 16584
rect 42524 16541 42533 16575
rect 42533 16541 42567 16575
rect 42567 16541 42576 16575
rect 42524 16532 42576 16541
rect 33692 16464 33744 16516
rect 36544 16507 36596 16516
rect 36544 16473 36553 16507
rect 36553 16473 36587 16507
rect 36587 16473 36596 16507
rect 36544 16464 36596 16473
rect 37372 16464 37424 16516
rect 37648 16464 37700 16516
rect 38108 16464 38160 16516
rect 39028 16507 39080 16516
rect 39028 16473 39037 16507
rect 39037 16473 39071 16507
rect 39071 16473 39080 16507
rect 39028 16464 39080 16473
rect 38752 16396 38804 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 14556 16235 14608 16244
rect 14556 16201 14565 16235
rect 14565 16201 14599 16235
rect 14599 16201 14608 16235
rect 14556 16192 14608 16201
rect 15384 16192 15436 16244
rect 17316 16192 17368 16244
rect 20628 16192 20680 16244
rect 22100 16192 22152 16244
rect 24400 16192 24452 16244
rect 28172 16235 28224 16244
rect 28172 16201 28181 16235
rect 28181 16201 28215 16235
rect 28215 16201 28224 16235
rect 28172 16192 28224 16201
rect 28540 16192 28592 16244
rect 30288 16235 30340 16244
rect 15108 16167 15160 16176
rect 15108 16133 15117 16167
rect 15117 16133 15151 16167
rect 15151 16133 15160 16167
rect 15108 16124 15160 16133
rect 16856 16056 16908 16108
rect 17500 16124 17552 16176
rect 18328 16124 18380 16176
rect 17408 16056 17460 16108
rect 18420 16056 18472 16108
rect 20628 16056 20680 16108
rect 20904 16099 20956 16108
rect 20904 16065 20913 16099
rect 20913 16065 20947 16099
rect 20947 16065 20956 16099
rect 22836 16124 22888 16176
rect 23480 16167 23532 16176
rect 23480 16133 23489 16167
rect 23489 16133 23523 16167
rect 23523 16133 23532 16167
rect 23480 16124 23532 16133
rect 25872 16124 25924 16176
rect 29000 16124 29052 16176
rect 22744 16099 22796 16108
rect 20904 16056 20956 16065
rect 22744 16065 22753 16099
rect 22753 16065 22787 16099
rect 22787 16065 22796 16099
rect 22744 16056 22796 16065
rect 27160 16099 27212 16108
rect 27160 16065 27169 16099
rect 27169 16065 27203 16099
rect 27203 16065 27212 16099
rect 27160 16056 27212 16065
rect 27344 16099 27396 16108
rect 27344 16065 27353 16099
rect 27353 16065 27387 16099
rect 27387 16065 27396 16099
rect 27344 16056 27396 16065
rect 16764 15988 16816 16040
rect 16948 15988 17000 16040
rect 17224 16031 17276 16040
rect 17224 15997 17233 16031
rect 17233 15997 17267 16031
rect 17267 15997 17276 16031
rect 17224 15988 17276 15997
rect 17592 15988 17644 16040
rect 19984 16031 20036 16040
rect 19984 15997 19993 16031
rect 19993 15997 20027 16031
rect 20027 15997 20036 16031
rect 19984 15988 20036 15997
rect 21088 15988 21140 16040
rect 22008 15988 22060 16040
rect 20536 15920 20588 15972
rect 20628 15920 20680 15972
rect 22836 15920 22888 15972
rect 23388 15988 23440 16040
rect 26240 16031 26292 16040
rect 26240 15997 26249 16031
rect 26249 15997 26283 16031
rect 26283 15997 26292 16031
rect 26240 15988 26292 15997
rect 26332 15988 26384 16040
rect 25504 15920 25556 15972
rect 27344 15920 27396 15972
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 14280 15852 14332 15904
rect 15568 15895 15620 15904
rect 15568 15861 15577 15895
rect 15577 15861 15611 15895
rect 15611 15861 15620 15895
rect 15568 15852 15620 15861
rect 17868 15852 17920 15904
rect 17960 15852 18012 15904
rect 20812 15852 20864 15904
rect 24124 15852 24176 15904
rect 24216 15852 24268 15904
rect 28816 16056 28868 16108
rect 29092 16099 29144 16108
rect 29092 16065 29101 16099
rect 29101 16065 29135 16099
rect 29135 16065 29144 16099
rect 30288 16201 30297 16235
rect 30297 16201 30331 16235
rect 30331 16201 30340 16235
rect 30288 16192 30340 16201
rect 36360 16192 36412 16244
rect 37280 16192 37332 16244
rect 41512 16192 41564 16244
rect 41604 16192 41656 16244
rect 42892 16192 42944 16244
rect 54208 16235 54260 16244
rect 54208 16201 54217 16235
rect 54217 16201 54251 16235
rect 54251 16201 54260 16235
rect 54208 16192 54260 16201
rect 35164 16167 35216 16176
rect 29092 16056 29144 16065
rect 30012 16056 30064 16108
rect 31116 16099 31168 16108
rect 31116 16065 31125 16099
rect 31125 16065 31159 16099
rect 31159 16065 31168 16099
rect 31116 16056 31168 16065
rect 31852 16056 31904 16108
rect 32312 16099 32364 16108
rect 32312 16065 32321 16099
rect 32321 16065 32355 16099
rect 32355 16065 32364 16099
rect 32312 16056 32364 16065
rect 32496 16099 32548 16108
rect 32496 16065 32505 16099
rect 32505 16065 32539 16099
rect 32539 16065 32548 16099
rect 32496 16056 32548 16065
rect 32956 16099 33008 16108
rect 32956 16065 32965 16099
rect 32965 16065 32999 16099
rect 32999 16065 33008 16099
rect 32956 16056 33008 16065
rect 33048 16056 33100 16108
rect 28264 15963 28316 15972
rect 28264 15929 28273 15963
rect 28273 15929 28307 15963
rect 28307 15929 28316 15963
rect 28264 15920 28316 15929
rect 28448 15852 28500 15904
rect 32036 15988 32088 16040
rect 28816 15920 28868 15972
rect 33140 15852 33192 15904
rect 33324 15852 33376 15904
rect 35164 16133 35173 16167
rect 35173 16133 35207 16167
rect 35207 16133 35216 16167
rect 35164 16124 35216 16133
rect 36452 16124 36504 16176
rect 38200 16124 38252 16176
rect 42800 16124 42852 16176
rect 36912 16099 36964 16108
rect 36912 16065 36921 16099
rect 36921 16065 36955 16099
rect 36955 16065 36964 16099
rect 36912 16056 36964 16065
rect 34704 15988 34756 16040
rect 38108 15920 38160 15972
rect 38568 16056 38620 16108
rect 41328 16056 41380 16108
rect 54024 16099 54076 16108
rect 41420 15988 41472 16040
rect 42524 15988 42576 16040
rect 43812 15988 43864 16040
rect 43720 15963 43772 15972
rect 43720 15929 43729 15963
rect 43729 15929 43763 15963
rect 43763 15929 43772 15963
rect 43720 15920 43772 15929
rect 34428 15852 34480 15904
rect 34520 15852 34572 15904
rect 35992 15852 36044 15904
rect 37464 15895 37516 15904
rect 37464 15861 37473 15895
rect 37473 15861 37507 15895
rect 37507 15861 37516 15895
rect 37464 15852 37516 15861
rect 38200 15895 38252 15904
rect 38200 15861 38209 15895
rect 38209 15861 38243 15895
rect 38243 15861 38252 15895
rect 38200 15852 38252 15861
rect 38292 15852 38344 15904
rect 41236 15852 41288 15904
rect 41328 15852 41380 15904
rect 42616 15895 42668 15904
rect 42616 15861 42625 15895
rect 42625 15861 42659 15895
rect 42659 15861 42668 15895
rect 42616 15852 42668 15861
rect 42984 15852 43036 15904
rect 54024 16065 54033 16099
rect 54033 16065 54067 16099
rect 54067 16065 54076 16099
rect 54024 16056 54076 16065
rect 53288 15920 53340 15972
rect 53656 15852 53708 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 16488 15648 16540 15700
rect 16856 15648 16908 15700
rect 17776 15648 17828 15700
rect 20628 15648 20680 15700
rect 21640 15691 21692 15700
rect 21640 15657 21649 15691
rect 21649 15657 21683 15691
rect 21683 15657 21692 15691
rect 21640 15648 21692 15657
rect 24768 15648 24820 15700
rect 26332 15648 26384 15700
rect 28632 15648 28684 15700
rect 20812 15623 20864 15632
rect 15936 15512 15988 15564
rect 15568 15444 15620 15496
rect 20812 15589 20821 15623
rect 20821 15589 20855 15623
rect 20855 15589 20864 15623
rect 20812 15580 20864 15589
rect 21732 15580 21784 15632
rect 33692 15648 33744 15700
rect 34704 15648 34756 15700
rect 17960 15512 18012 15564
rect 18788 15555 18840 15564
rect 18788 15521 18797 15555
rect 18797 15521 18831 15555
rect 18831 15521 18840 15555
rect 18788 15512 18840 15521
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 26240 15512 26292 15564
rect 28908 15512 28960 15564
rect 29368 15512 29420 15564
rect 33600 15580 33652 15632
rect 16948 15487 17000 15496
rect 16948 15453 16957 15487
rect 16957 15453 16991 15487
rect 16991 15453 17000 15487
rect 16948 15444 17000 15453
rect 17132 15487 17184 15496
rect 17132 15453 17141 15487
rect 17141 15453 17175 15487
rect 17175 15453 17184 15487
rect 17132 15444 17184 15453
rect 17224 15487 17276 15496
rect 17224 15453 17233 15487
rect 17233 15453 17267 15487
rect 17267 15453 17276 15487
rect 19432 15487 19484 15496
rect 17224 15444 17276 15453
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 19524 15444 19576 15496
rect 21824 15487 21876 15496
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 14740 15376 14792 15428
rect 15108 15376 15160 15428
rect 17592 15376 17644 15428
rect 1676 15351 1728 15360
rect 1676 15317 1685 15351
rect 1685 15317 1719 15351
rect 1719 15317 1728 15351
rect 1676 15308 1728 15317
rect 15016 15351 15068 15360
rect 15016 15317 15025 15351
rect 15025 15317 15059 15351
rect 15059 15317 15068 15351
rect 15016 15308 15068 15317
rect 20352 15376 20404 15428
rect 18144 15351 18196 15360
rect 18144 15317 18153 15351
rect 18153 15317 18187 15351
rect 18187 15317 18196 15351
rect 18144 15308 18196 15317
rect 18236 15308 18288 15360
rect 18604 15351 18656 15360
rect 18604 15317 18613 15351
rect 18613 15317 18647 15351
rect 18647 15317 18656 15351
rect 18604 15308 18656 15317
rect 19984 15308 20036 15360
rect 24676 15444 24728 15496
rect 26516 15487 26568 15496
rect 26516 15453 26525 15487
rect 26525 15453 26559 15487
rect 26559 15453 26568 15487
rect 26516 15444 26568 15453
rect 27896 15444 27948 15496
rect 28080 15487 28132 15496
rect 28080 15453 28089 15487
rect 28089 15453 28123 15487
rect 28123 15453 28132 15487
rect 28080 15444 28132 15453
rect 28540 15444 28592 15496
rect 29460 15444 29512 15496
rect 29920 15487 29972 15496
rect 29920 15453 29929 15487
rect 29929 15453 29963 15487
rect 29963 15453 29972 15487
rect 29920 15444 29972 15453
rect 22192 15376 22244 15428
rect 24032 15376 24084 15428
rect 29184 15376 29236 15428
rect 29276 15376 29328 15428
rect 31300 15444 31352 15496
rect 33140 15512 33192 15564
rect 35532 15512 35584 15564
rect 37556 15648 37608 15700
rect 37924 15691 37976 15700
rect 37924 15657 37933 15691
rect 37933 15657 37967 15691
rect 37967 15657 37976 15691
rect 37924 15648 37976 15657
rect 36544 15580 36596 15632
rect 38384 15580 38436 15632
rect 39028 15580 39080 15632
rect 32220 15444 32272 15496
rect 30932 15419 30984 15428
rect 30932 15385 30941 15419
rect 30941 15385 30975 15419
rect 30975 15385 30984 15419
rect 30932 15376 30984 15385
rect 31116 15376 31168 15428
rect 34520 15444 34572 15496
rect 35164 15487 35216 15496
rect 35164 15453 35173 15487
rect 35173 15453 35207 15487
rect 35207 15453 35216 15487
rect 35164 15444 35216 15453
rect 35716 15444 35768 15496
rect 36452 15487 36504 15496
rect 36452 15453 36461 15487
rect 36461 15453 36495 15487
rect 36495 15453 36504 15487
rect 36452 15444 36504 15453
rect 39672 15580 39724 15632
rect 41512 15580 41564 15632
rect 42800 15648 42852 15700
rect 43168 15648 43220 15700
rect 54024 15648 54076 15700
rect 53288 15623 53340 15632
rect 41420 15555 41472 15564
rect 41420 15521 41429 15555
rect 41429 15521 41463 15555
rect 41463 15521 41472 15555
rect 41420 15512 41472 15521
rect 53288 15589 53297 15623
rect 53297 15589 53331 15623
rect 53331 15589 53340 15623
rect 53288 15580 53340 15589
rect 39304 15487 39356 15496
rect 39304 15453 39313 15487
rect 39313 15453 39347 15487
rect 39347 15453 39356 15487
rect 39304 15444 39356 15453
rect 41512 15444 41564 15496
rect 42064 15487 42116 15496
rect 42064 15453 42073 15487
rect 42073 15453 42107 15487
rect 42107 15453 42116 15487
rect 42064 15444 42116 15453
rect 42524 15487 42576 15496
rect 42524 15453 42533 15487
rect 42533 15453 42567 15487
rect 42567 15453 42576 15487
rect 42524 15444 42576 15453
rect 42892 15444 42944 15496
rect 43352 15487 43404 15496
rect 43352 15453 43361 15487
rect 43361 15453 43395 15487
rect 43395 15453 43404 15487
rect 43352 15444 43404 15453
rect 53564 15444 53616 15496
rect 54208 15487 54260 15496
rect 54208 15453 54217 15487
rect 54217 15453 54251 15487
rect 54251 15453 54260 15487
rect 54208 15444 54260 15453
rect 37464 15376 37516 15428
rect 23664 15351 23716 15360
rect 23664 15317 23673 15351
rect 23673 15317 23707 15351
rect 23707 15317 23716 15351
rect 23664 15308 23716 15317
rect 24124 15308 24176 15360
rect 26792 15308 26844 15360
rect 27620 15308 27672 15360
rect 28632 15308 28684 15360
rect 28816 15308 28868 15360
rect 30380 15308 30432 15360
rect 30840 15308 30892 15360
rect 34796 15308 34848 15360
rect 35348 15308 35400 15360
rect 38844 15308 38896 15360
rect 39396 15308 39448 15360
rect 40500 15376 40552 15428
rect 39672 15308 39724 15360
rect 41328 15308 41380 15360
rect 41696 15308 41748 15360
rect 42616 15351 42668 15360
rect 42616 15317 42625 15351
rect 42625 15317 42659 15351
rect 42659 15317 42668 15351
rect 42616 15308 42668 15317
rect 43444 15376 43496 15428
rect 53472 15419 53524 15428
rect 53472 15385 53481 15419
rect 53481 15385 53515 15419
rect 53515 15385 53524 15419
rect 53472 15376 53524 15385
rect 44456 15351 44508 15360
rect 44456 15317 44465 15351
rect 44465 15317 44499 15351
rect 44499 15317 44508 15351
rect 44456 15308 44508 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 18696 15104 18748 15156
rect 19340 15104 19392 15156
rect 20812 15147 20864 15156
rect 20812 15113 20821 15147
rect 20821 15113 20855 15147
rect 20855 15113 20864 15147
rect 20812 15104 20864 15113
rect 22744 15104 22796 15156
rect 14280 15079 14332 15088
rect 14280 15045 14289 15079
rect 14289 15045 14323 15079
rect 14323 15045 14332 15079
rect 14280 15036 14332 15045
rect 15936 15079 15988 15088
rect 15936 15045 15945 15079
rect 15945 15045 15979 15079
rect 15979 15045 15988 15079
rect 15936 15036 15988 15045
rect 17684 15036 17736 15088
rect 18328 15036 18380 15088
rect 18420 15036 18472 15088
rect 26056 15104 26108 15156
rect 26516 15104 26568 15156
rect 27436 15104 27488 15156
rect 23756 15079 23808 15088
rect 23756 15045 23765 15079
rect 23765 15045 23799 15079
rect 23799 15045 23808 15079
rect 23756 15036 23808 15045
rect 25136 15036 25188 15088
rect 28356 15104 28408 15156
rect 29000 15104 29052 15156
rect 41328 15147 41380 15156
rect 4620 14968 4672 15020
rect 14740 15011 14792 15020
rect 14740 14977 14749 15011
rect 14749 14977 14783 15011
rect 14783 14977 14792 15011
rect 14740 14968 14792 14977
rect 15384 14968 15436 15020
rect 16672 14968 16724 15020
rect 20076 14968 20128 15020
rect 11704 14900 11756 14952
rect 17132 14832 17184 14884
rect 17316 14943 17368 14952
rect 17316 14909 17325 14943
rect 17325 14909 17359 14943
rect 17359 14909 17368 14943
rect 17316 14900 17368 14909
rect 17592 14900 17644 14952
rect 20536 14900 20588 14952
rect 22560 14968 22612 15020
rect 23388 14968 23440 15020
rect 23664 15011 23716 15020
rect 23664 14977 23673 15011
rect 23673 14977 23707 15011
rect 23707 14977 23716 15011
rect 24768 15011 24820 15020
rect 23664 14968 23716 14977
rect 24768 14977 24777 15011
rect 24777 14977 24811 15011
rect 24811 14977 24820 15011
rect 24768 14968 24820 14977
rect 17776 14832 17828 14884
rect 20812 14832 20864 14884
rect 21180 14900 21232 14952
rect 22836 14943 22888 14952
rect 22836 14909 22845 14943
rect 22845 14909 22879 14943
rect 22879 14909 22888 14943
rect 22836 14900 22888 14909
rect 23848 14943 23900 14952
rect 23848 14909 23857 14943
rect 23857 14909 23891 14943
rect 23891 14909 23900 14943
rect 23848 14900 23900 14909
rect 25320 14943 25372 14952
rect 25320 14909 25329 14943
rect 25329 14909 25363 14943
rect 25363 14909 25372 14943
rect 25320 14900 25372 14909
rect 25780 14943 25832 14952
rect 25780 14909 25789 14943
rect 25789 14909 25823 14943
rect 25823 14909 25832 14943
rect 25780 14900 25832 14909
rect 26332 14943 26384 14952
rect 26332 14909 26341 14943
rect 26341 14909 26375 14943
rect 26375 14909 26384 14943
rect 26332 14900 26384 14909
rect 26884 14900 26936 14952
rect 27068 14900 27120 14952
rect 27436 14943 27488 14952
rect 27436 14909 27445 14943
rect 27445 14909 27479 14943
rect 27479 14909 27488 14943
rect 27620 14943 27672 14952
rect 27436 14900 27488 14909
rect 27620 14909 27629 14943
rect 27629 14909 27663 14943
rect 27663 14909 27672 14943
rect 27620 14900 27672 14909
rect 21640 14832 21692 14884
rect 23204 14832 23256 14884
rect 24768 14832 24820 14884
rect 27160 14832 27212 14884
rect 28264 14968 28316 15020
rect 27804 14900 27856 14952
rect 28540 15011 28592 15020
rect 28540 14977 28554 15011
rect 28554 14977 28588 15011
rect 28588 14977 28592 15011
rect 28908 15036 28960 15088
rect 29552 15079 29604 15088
rect 29552 15045 29561 15079
rect 29561 15045 29595 15079
rect 29595 15045 29604 15079
rect 29552 15036 29604 15045
rect 28540 14968 28592 14977
rect 30472 14900 30524 14952
rect 35164 14968 35216 15020
rect 35440 14968 35492 15020
rect 37832 14968 37884 15020
rect 38016 15036 38068 15088
rect 38476 15036 38528 15088
rect 39672 15079 39724 15088
rect 38200 14968 38252 15020
rect 39672 15045 39681 15079
rect 39681 15045 39715 15079
rect 39715 15045 39724 15079
rect 39672 15036 39724 15045
rect 31668 14943 31720 14952
rect 29184 14875 29236 14884
rect 1676 14807 1728 14816
rect 1676 14773 1685 14807
rect 1685 14773 1719 14807
rect 1719 14773 1728 14807
rect 1676 14764 1728 14773
rect 13176 14807 13228 14816
rect 13176 14773 13185 14807
rect 13185 14773 13219 14807
rect 13219 14773 13228 14807
rect 13176 14764 13228 14773
rect 15384 14807 15436 14816
rect 15384 14773 15393 14807
rect 15393 14773 15427 14807
rect 15427 14773 15436 14807
rect 15384 14764 15436 14773
rect 15936 14764 15988 14816
rect 16488 14764 16540 14816
rect 17408 14764 17460 14816
rect 20720 14764 20772 14816
rect 20904 14764 20956 14816
rect 22560 14764 22612 14816
rect 23940 14764 23992 14816
rect 29184 14841 29193 14875
rect 29193 14841 29227 14875
rect 29227 14841 29236 14875
rect 29184 14832 29236 14841
rect 31668 14909 31677 14943
rect 31677 14909 31711 14943
rect 31711 14909 31720 14943
rect 31668 14900 31720 14909
rect 33692 14943 33744 14952
rect 33692 14909 33701 14943
rect 33701 14909 33735 14943
rect 33735 14909 33744 14943
rect 33692 14900 33744 14909
rect 34704 14943 34756 14952
rect 34704 14909 34713 14943
rect 34713 14909 34747 14943
rect 34747 14909 34756 14943
rect 34704 14900 34756 14909
rect 39488 15011 39540 15020
rect 39488 14977 39497 15011
rect 39497 14977 39531 15011
rect 39531 14977 39540 15011
rect 39488 14968 39540 14977
rect 41328 15113 41355 15147
rect 41355 15113 41380 15147
rect 41328 15104 41380 15113
rect 43168 15147 43220 15156
rect 43168 15113 43177 15147
rect 43177 15113 43211 15147
rect 43211 15113 43220 15147
rect 43168 15104 43220 15113
rect 53564 15147 53616 15156
rect 53564 15113 53573 15147
rect 53573 15113 53607 15147
rect 53607 15113 53616 15147
rect 53564 15104 53616 15113
rect 54208 15147 54260 15156
rect 54208 15113 54217 15147
rect 54217 15113 54251 15147
rect 54251 15113 54260 15147
rect 54208 15104 54260 15113
rect 41880 15036 41932 15088
rect 42064 15036 42116 15088
rect 42524 15036 42576 15088
rect 43444 15036 43496 15088
rect 40500 15011 40552 15020
rect 40500 14977 40509 15011
rect 40509 14977 40543 15011
rect 40543 14977 40552 15011
rect 40500 14968 40552 14977
rect 43352 14968 43404 15020
rect 54024 15011 54076 15020
rect 54024 14977 54033 15011
rect 54033 14977 54067 15011
rect 54067 14977 54076 15011
rect 54024 14968 54076 14977
rect 32680 14832 32732 14884
rect 33876 14832 33928 14884
rect 37464 14875 37516 14884
rect 28172 14807 28224 14816
rect 28172 14773 28181 14807
rect 28181 14773 28215 14807
rect 28215 14773 28224 14807
rect 28172 14764 28224 14773
rect 30104 14807 30156 14816
rect 30104 14773 30113 14807
rect 30113 14773 30147 14807
rect 30147 14773 30156 14807
rect 30104 14764 30156 14773
rect 33508 14764 33560 14816
rect 33784 14764 33836 14816
rect 37096 14764 37148 14816
rect 37464 14841 37473 14875
rect 37473 14841 37507 14875
rect 37507 14841 37516 14875
rect 37464 14832 37516 14841
rect 40040 14900 40092 14952
rect 40224 14900 40276 14952
rect 40408 14900 40460 14952
rect 41696 14832 41748 14884
rect 39120 14764 39172 14816
rect 39304 14807 39356 14816
rect 39304 14773 39313 14807
rect 39313 14773 39347 14807
rect 39347 14773 39356 14807
rect 39304 14764 39356 14773
rect 39396 14764 39448 14816
rect 40224 14764 40276 14816
rect 41052 14764 41104 14816
rect 42616 14900 42668 14952
rect 41880 14832 41932 14884
rect 42064 14832 42116 14884
rect 41972 14807 42024 14816
rect 41972 14773 41981 14807
rect 41981 14773 42015 14807
rect 42015 14773 42024 14807
rect 41972 14764 42024 14773
rect 42616 14807 42668 14816
rect 42616 14773 42625 14807
rect 42625 14773 42659 14807
rect 42659 14773 42668 14807
rect 42616 14764 42668 14773
rect 43260 14764 43312 14816
rect 44272 14807 44324 14816
rect 44272 14773 44281 14807
rect 44281 14773 44315 14807
rect 44315 14773 44324 14807
rect 44272 14764 44324 14773
rect 53748 14764 53800 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 15108 14603 15160 14612
rect 15108 14569 15117 14603
rect 15117 14569 15151 14603
rect 15151 14569 15160 14603
rect 15108 14560 15160 14569
rect 15568 14603 15620 14612
rect 15568 14569 15577 14603
rect 15577 14569 15611 14603
rect 15611 14569 15620 14603
rect 15568 14560 15620 14569
rect 16580 14603 16632 14612
rect 16580 14569 16589 14603
rect 16589 14569 16623 14603
rect 16623 14569 16632 14603
rect 16580 14560 16632 14569
rect 18420 14560 18472 14612
rect 4620 14424 4672 14476
rect 11704 14424 11756 14476
rect 14740 14424 14792 14476
rect 15108 14424 15160 14476
rect 15476 14424 15528 14476
rect 15660 14356 15712 14408
rect 16028 14399 16080 14408
rect 4344 14288 4396 14340
rect 15568 14288 15620 14340
rect 1676 14263 1728 14272
rect 1676 14229 1685 14263
rect 1685 14229 1719 14263
rect 1719 14229 1728 14263
rect 1676 14220 1728 14229
rect 13176 14263 13228 14272
rect 13176 14229 13185 14263
rect 13185 14229 13219 14263
rect 13219 14229 13228 14263
rect 13176 14220 13228 14229
rect 14924 14220 14976 14272
rect 15476 14220 15528 14272
rect 16028 14365 16037 14399
rect 16037 14365 16071 14399
rect 16071 14365 16080 14399
rect 16028 14356 16080 14365
rect 16488 14424 16540 14476
rect 17408 14424 17460 14476
rect 18788 14467 18840 14476
rect 18788 14433 18797 14467
rect 18797 14433 18831 14467
rect 18831 14433 18840 14467
rect 18788 14424 18840 14433
rect 16580 14288 16632 14340
rect 17684 14356 17736 14408
rect 17868 14356 17920 14408
rect 19432 14399 19484 14408
rect 17132 14288 17184 14340
rect 17960 14288 18012 14340
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 20076 14356 20128 14408
rect 20720 14560 20772 14612
rect 23756 14560 23808 14612
rect 27804 14560 27856 14612
rect 28172 14560 28224 14612
rect 31668 14603 31720 14612
rect 28908 14492 28960 14544
rect 31668 14569 31677 14603
rect 31677 14569 31711 14603
rect 31711 14569 31720 14603
rect 31668 14560 31720 14569
rect 34704 14560 34756 14612
rect 41512 14560 41564 14612
rect 43444 14560 43496 14612
rect 37832 14492 37884 14544
rect 38936 14492 38988 14544
rect 39212 14492 39264 14544
rect 39304 14492 39356 14544
rect 54208 14535 54260 14544
rect 54208 14501 54217 14535
rect 54217 14501 54251 14535
rect 54251 14501 54260 14535
rect 54208 14492 54260 14501
rect 21180 14424 21232 14476
rect 22284 14424 22336 14476
rect 24124 14424 24176 14476
rect 24308 14424 24360 14476
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 21640 14356 21692 14365
rect 24216 14356 24268 14408
rect 29276 14424 29328 14476
rect 29828 14467 29880 14476
rect 29828 14433 29837 14467
rect 29837 14433 29871 14467
rect 29871 14433 29880 14467
rect 29828 14424 29880 14433
rect 31300 14424 31352 14476
rect 31760 14424 31812 14476
rect 32036 14467 32088 14476
rect 32036 14433 32045 14467
rect 32045 14433 32079 14467
rect 32079 14433 32088 14467
rect 32956 14467 33008 14476
rect 32036 14424 32088 14433
rect 20720 14288 20772 14340
rect 27252 14356 27304 14408
rect 27712 14399 27764 14408
rect 27712 14365 27721 14399
rect 27721 14365 27755 14399
rect 27755 14365 27764 14399
rect 27712 14356 27764 14365
rect 28540 14356 28592 14408
rect 26240 14288 26292 14340
rect 26608 14288 26660 14340
rect 28448 14288 28500 14340
rect 29092 14356 29144 14408
rect 29920 14356 29972 14408
rect 30932 14356 30984 14408
rect 29184 14288 29236 14340
rect 32128 14399 32180 14408
rect 32128 14365 32137 14399
rect 32137 14365 32171 14399
rect 32171 14365 32180 14399
rect 32956 14433 32965 14467
rect 32965 14433 32999 14467
rect 32999 14433 33008 14467
rect 32956 14424 33008 14433
rect 33784 14467 33836 14476
rect 33784 14433 33793 14467
rect 33793 14433 33827 14467
rect 33827 14433 33836 14467
rect 33784 14424 33836 14433
rect 32864 14399 32916 14408
rect 32128 14356 32180 14365
rect 32864 14365 32873 14399
rect 32873 14365 32907 14399
rect 32907 14365 32916 14399
rect 32864 14356 32916 14365
rect 33600 14356 33652 14408
rect 36268 14399 36320 14408
rect 34244 14288 34296 14340
rect 34612 14288 34664 14340
rect 35256 14288 35308 14340
rect 35900 14288 35952 14340
rect 36268 14365 36277 14399
rect 36277 14365 36311 14399
rect 36311 14365 36320 14399
rect 36268 14356 36320 14365
rect 37096 14356 37148 14408
rect 37464 14399 37516 14408
rect 37464 14365 37474 14399
rect 37474 14365 37516 14399
rect 37464 14356 37516 14365
rect 39028 14424 39080 14476
rect 38292 14399 38344 14408
rect 38292 14365 38301 14399
rect 38301 14365 38335 14399
rect 38335 14365 38344 14399
rect 38292 14356 38344 14365
rect 40224 14356 40276 14408
rect 41328 14356 41380 14408
rect 41420 14399 41472 14408
rect 41420 14365 41429 14399
rect 41429 14365 41463 14399
rect 41463 14365 41472 14399
rect 41420 14356 41472 14365
rect 42708 14356 42760 14408
rect 44272 14356 44324 14408
rect 38752 14288 38804 14340
rect 40684 14288 40736 14340
rect 40776 14288 40828 14340
rect 41512 14288 41564 14340
rect 42616 14288 42668 14340
rect 15936 14220 15988 14272
rect 18144 14263 18196 14272
rect 18144 14229 18153 14263
rect 18153 14229 18187 14263
rect 18187 14229 18196 14263
rect 18144 14220 18196 14229
rect 18696 14220 18748 14272
rect 20812 14263 20864 14272
rect 20812 14229 20821 14263
rect 20821 14229 20855 14263
rect 20855 14229 20864 14263
rect 20812 14220 20864 14229
rect 21272 14263 21324 14272
rect 21272 14229 21281 14263
rect 21281 14229 21315 14263
rect 21315 14229 21324 14263
rect 21272 14220 21324 14229
rect 21732 14263 21784 14272
rect 21732 14229 21741 14263
rect 21741 14229 21775 14263
rect 21775 14229 21784 14263
rect 21732 14220 21784 14229
rect 21824 14220 21876 14272
rect 25504 14220 25556 14272
rect 28540 14220 28592 14272
rect 30748 14220 30800 14272
rect 31208 14263 31260 14272
rect 31208 14229 31217 14263
rect 31217 14229 31251 14263
rect 31251 14229 31260 14263
rect 31208 14220 31260 14229
rect 32680 14220 32732 14272
rect 33600 14220 33652 14272
rect 34428 14220 34480 14272
rect 35348 14220 35400 14272
rect 37372 14263 37424 14272
rect 37372 14229 37381 14263
rect 37381 14229 37415 14263
rect 37415 14229 37424 14263
rect 37372 14220 37424 14229
rect 38384 14220 38436 14272
rect 39120 14220 39172 14272
rect 39856 14220 39908 14272
rect 40040 14263 40092 14272
rect 40040 14229 40049 14263
rect 40049 14229 40083 14263
rect 40083 14229 40092 14263
rect 40040 14220 40092 14229
rect 43904 14220 43956 14272
rect 54024 14399 54076 14408
rect 54024 14365 54033 14399
rect 54033 14365 54067 14399
rect 54067 14365 54076 14399
rect 54024 14356 54076 14365
rect 49056 14220 49108 14272
rect 54208 14220 54260 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 14004 14016 14056 14068
rect 15016 14016 15068 14068
rect 14464 13948 14516 14000
rect 14556 13948 14608 14000
rect 15108 13991 15160 14000
rect 15108 13957 15117 13991
rect 15117 13957 15151 13991
rect 15151 13957 15160 13991
rect 15108 13948 15160 13957
rect 4344 13880 4396 13932
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 17592 14016 17644 14068
rect 18328 14059 18380 14068
rect 18328 14025 18337 14059
rect 18337 14025 18371 14059
rect 18371 14025 18380 14059
rect 18328 14016 18380 14025
rect 18604 14016 18656 14068
rect 21824 14016 21876 14068
rect 23388 14059 23440 14068
rect 23388 14025 23397 14059
rect 23397 14025 23431 14059
rect 23431 14025 23440 14059
rect 23388 14016 23440 14025
rect 23756 14059 23808 14068
rect 23756 14025 23765 14059
rect 23765 14025 23799 14059
rect 23799 14025 23808 14059
rect 23756 14016 23808 14025
rect 23940 14016 23992 14068
rect 15844 13880 15896 13932
rect 15936 13855 15988 13864
rect 15936 13821 15945 13855
rect 15945 13821 15979 13855
rect 15979 13821 15988 13855
rect 15936 13812 15988 13821
rect 16580 13880 16632 13932
rect 16856 13880 16908 13932
rect 18236 13948 18288 14000
rect 21732 13948 21784 14000
rect 22100 13948 22152 14000
rect 31300 14059 31352 14068
rect 31300 14025 31309 14059
rect 31309 14025 31343 14059
rect 31343 14025 31352 14059
rect 31300 14016 31352 14025
rect 32036 14016 32088 14068
rect 35808 14016 35860 14068
rect 24676 13948 24728 14000
rect 17592 13880 17644 13932
rect 19616 13880 19668 13932
rect 20996 13880 21048 13932
rect 21456 13880 21508 13932
rect 24216 13880 24268 13932
rect 16396 13812 16448 13864
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 17408 13812 17460 13864
rect 20076 13812 20128 13864
rect 19892 13744 19944 13796
rect 20904 13744 20956 13796
rect 21180 13744 21232 13796
rect 23940 13855 23992 13864
rect 23940 13821 23949 13855
rect 23949 13821 23983 13855
rect 23983 13821 23992 13855
rect 23940 13812 23992 13821
rect 24308 13812 24360 13864
rect 24492 13812 24544 13864
rect 25780 13880 25832 13932
rect 26056 13880 26108 13932
rect 26700 13880 26752 13932
rect 24768 13787 24820 13796
rect 24768 13753 24777 13787
rect 24777 13753 24811 13787
rect 24811 13753 24820 13787
rect 24768 13744 24820 13753
rect 26608 13787 26660 13796
rect 26608 13753 26617 13787
rect 26617 13753 26651 13787
rect 26651 13753 26660 13787
rect 26608 13744 26660 13753
rect 27712 13880 27764 13932
rect 27988 13880 28040 13932
rect 29276 13948 29328 14000
rect 30472 13948 30524 14000
rect 33692 13948 33744 14000
rect 39948 14016 40000 14068
rect 43260 14059 43312 14068
rect 43260 14025 43269 14059
rect 43269 14025 43303 14059
rect 43303 14025 43312 14059
rect 43260 14016 43312 14025
rect 43812 14059 43864 14068
rect 43812 14025 43821 14059
rect 43821 14025 43855 14059
rect 43855 14025 43864 14059
rect 43812 14016 43864 14025
rect 43904 14016 43956 14068
rect 54024 14016 54076 14068
rect 29092 13880 29144 13932
rect 30012 13923 30064 13932
rect 30012 13889 30021 13923
rect 30021 13889 30055 13923
rect 30055 13889 30064 13923
rect 30012 13880 30064 13889
rect 30932 13880 30984 13932
rect 32128 13880 32180 13932
rect 54208 13991 54260 14000
rect 34428 13923 34480 13932
rect 34428 13889 34462 13923
rect 34462 13889 34480 13923
rect 34428 13880 34480 13889
rect 36268 13880 36320 13932
rect 38200 13880 38252 13932
rect 32956 13855 33008 13864
rect 32956 13821 32965 13855
rect 32965 13821 32999 13855
rect 32999 13821 33008 13855
rect 32956 13812 33008 13821
rect 33600 13812 33652 13864
rect 36544 13855 36596 13864
rect 36544 13821 36553 13855
rect 36553 13821 36587 13855
rect 36587 13821 36596 13855
rect 36544 13812 36596 13821
rect 38936 13880 38988 13932
rect 39764 13880 39816 13932
rect 39856 13880 39908 13932
rect 40500 13880 40552 13932
rect 41052 13923 41104 13932
rect 41052 13889 41061 13923
rect 41061 13889 41095 13923
rect 41095 13889 41104 13923
rect 41052 13880 41104 13889
rect 41144 13880 41196 13932
rect 54208 13957 54217 13991
rect 54217 13957 54251 13991
rect 54251 13957 54260 13991
rect 54208 13948 54260 13957
rect 53564 13880 53616 13932
rect 39120 13812 39172 13864
rect 41420 13812 41472 13864
rect 53840 13812 53892 13864
rect 1676 13719 1728 13728
rect 1676 13685 1685 13719
rect 1685 13685 1719 13719
rect 1719 13685 1728 13719
rect 1676 13676 1728 13685
rect 13176 13676 13228 13728
rect 15292 13719 15344 13728
rect 15292 13685 15301 13719
rect 15301 13685 15335 13719
rect 15335 13685 15344 13719
rect 15292 13676 15344 13685
rect 15660 13676 15712 13728
rect 16764 13676 16816 13728
rect 18420 13676 18472 13728
rect 18972 13676 19024 13728
rect 20628 13676 20680 13728
rect 22652 13676 22704 13728
rect 27160 13719 27212 13728
rect 27160 13685 27169 13719
rect 27169 13685 27203 13719
rect 27203 13685 27212 13719
rect 27160 13676 27212 13685
rect 27344 13676 27396 13728
rect 28908 13676 28960 13728
rect 30932 13744 30984 13796
rect 31484 13744 31536 13796
rect 35532 13744 35584 13796
rect 36360 13744 36412 13796
rect 53288 13787 53340 13796
rect 29920 13719 29972 13728
rect 29920 13685 29929 13719
rect 29929 13685 29963 13719
rect 29963 13685 29972 13719
rect 29920 13676 29972 13685
rect 33692 13676 33744 13728
rect 35440 13676 35492 13728
rect 35992 13719 36044 13728
rect 35992 13685 36001 13719
rect 36001 13685 36035 13719
rect 36035 13685 36044 13719
rect 35992 13676 36044 13685
rect 37556 13676 37608 13728
rect 39488 13719 39540 13728
rect 39488 13685 39497 13719
rect 39497 13685 39531 13719
rect 39531 13685 39540 13719
rect 39488 13676 39540 13685
rect 39856 13676 39908 13728
rect 40868 13719 40920 13728
rect 40868 13685 40877 13719
rect 40877 13685 40911 13719
rect 40911 13685 40920 13719
rect 40868 13676 40920 13685
rect 41512 13719 41564 13728
rect 41512 13685 41521 13719
rect 41521 13685 41555 13719
rect 41555 13685 41564 13719
rect 41512 13676 41564 13685
rect 53288 13753 53297 13787
rect 53297 13753 53331 13787
rect 53331 13753 53340 13787
rect 53288 13744 53340 13753
rect 54024 13676 54076 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 14924 13472 14976 13524
rect 15568 13472 15620 13524
rect 16120 13472 16172 13524
rect 22284 13515 22336 13524
rect 13728 13404 13780 13456
rect 17132 13404 17184 13456
rect 20076 13404 20128 13456
rect 15384 13336 15436 13388
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 14648 13311 14700 13320
rect 14648 13277 14657 13311
rect 14657 13277 14691 13311
rect 14691 13277 14700 13311
rect 14648 13268 14700 13277
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 15936 13268 15988 13320
rect 1676 13175 1728 13184
rect 1676 13141 1685 13175
rect 1685 13141 1719 13175
rect 1719 13141 1728 13175
rect 1676 13132 1728 13141
rect 13176 13175 13228 13184
rect 13176 13141 13185 13175
rect 13185 13141 13219 13175
rect 13219 13141 13228 13175
rect 13176 13132 13228 13141
rect 14832 13132 14884 13184
rect 16304 13132 16356 13184
rect 16488 13311 16540 13320
rect 16488 13277 16497 13311
rect 16497 13277 16531 13311
rect 16531 13277 16540 13311
rect 16488 13268 16540 13277
rect 16672 13268 16724 13320
rect 17592 13268 17644 13320
rect 22284 13481 22293 13515
rect 22293 13481 22327 13515
rect 22327 13481 22336 13515
rect 22284 13472 22336 13481
rect 23664 13472 23716 13524
rect 24584 13515 24636 13524
rect 24032 13404 24084 13456
rect 24584 13481 24593 13515
rect 24593 13481 24627 13515
rect 24627 13481 24636 13515
rect 24584 13472 24636 13481
rect 26240 13472 26292 13524
rect 26792 13472 26844 13524
rect 27344 13472 27396 13524
rect 29092 13515 29144 13524
rect 29092 13481 29101 13515
rect 29101 13481 29135 13515
rect 29135 13481 29144 13515
rect 29092 13472 29144 13481
rect 31116 13472 31168 13524
rect 32128 13472 32180 13524
rect 32864 13472 32916 13524
rect 18328 13268 18380 13320
rect 19892 13268 19944 13320
rect 19984 13268 20036 13320
rect 23756 13336 23808 13388
rect 23388 13268 23440 13320
rect 37280 13472 37332 13524
rect 37740 13472 37792 13524
rect 38476 13472 38528 13524
rect 39856 13472 39908 13524
rect 40776 13515 40828 13524
rect 40776 13481 40785 13515
rect 40785 13481 40819 13515
rect 40819 13481 40828 13515
rect 40776 13472 40828 13481
rect 41512 13515 41564 13524
rect 41512 13481 41521 13515
rect 41521 13481 41555 13515
rect 41555 13481 41564 13515
rect 41512 13472 41564 13481
rect 42524 13515 42576 13524
rect 42524 13481 42533 13515
rect 42533 13481 42567 13515
rect 42567 13481 42576 13515
rect 42524 13472 42576 13481
rect 53288 13472 53340 13524
rect 54208 13515 54260 13524
rect 54208 13481 54217 13515
rect 54217 13481 54251 13515
rect 54251 13481 54260 13515
rect 54208 13472 54260 13481
rect 53564 13447 53616 13456
rect 25320 13336 25372 13388
rect 25136 13268 25188 13320
rect 25412 13311 25464 13320
rect 25412 13277 25421 13311
rect 25421 13277 25455 13311
rect 25455 13277 25464 13311
rect 25412 13268 25464 13277
rect 27068 13268 27120 13320
rect 30472 13336 30524 13388
rect 31208 13336 31260 13388
rect 17040 13200 17092 13252
rect 17960 13132 18012 13184
rect 20168 13175 20220 13184
rect 20168 13141 20177 13175
rect 20177 13141 20211 13175
rect 20211 13141 20220 13175
rect 20168 13132 20220 13141
rect 25044 13200 25096 13252
rect 28356 13268 28408 13320
rect 29552 13268 29604 13320
rect 30380 13268 30432 13320
rect 30748 13311 30800 13320
rect 30748 13277 30757 13311
rect 30757 13277 30791 13311
rect 30791 13277 30800 13311
rect 30748 13268 30800 13277
rect 30840 13311 30892 13320
rect 30840 13277 30849 13311
rect 30849 13277 30883 13311
rect 30883 13277 30892 13311
rect 30840 13268 30892 13277
rect 29000 13200 29052 13252
rect 29920 13200 29972 13252
rect 31484 13268 31536 13320
rect 33140 13336 33192 13388
rect 33508 13379 33560 13388
rect 33508 13345 33517 13379
rect 33517 13345 33551 13379
rect 33551 13345 33560 13379
rect 33508 13336 33560 13345
rect 36268 13379 36320 13388
rect 36268 13345 36277 13379
rect 36277 13345 36311 13379
rect 36311 13345 36320 13379
rect 36268 13336 36320 13345
rect 31852 13268 31904 13320
rect 53564 13413 53573 13447
rect 53573 13413 53607 13447
rect 53607 13413 53616 13447
rect 53564 13404 53616 13413
rect 37372 13336 37424 13388
rect 37832 13336 37884 13388
rect 37096 13311 37148 13320
rect 37096 13277 37105 13311
rect 37105 13277 37139 13311
rect 37139 13277 37148 13311
rect 37096 13268 37148 13277
rect 37556 13311 37608 13320
rect 37556 13277 37568 13311
rect 37568 13277 37602 13311
rect 37602 13277 37608 13311
rect 37556 13268 37608 13277
rect 38108 13268 38160 13320
rect 38476 13268 38528 13320
rect 39488 13336 39540 13388
rect 39396 13311 39448 13320
rect 39396 13277 39405 13311
rect 39405 13277 39439 13311
rect 39439 13277 39448 13311
rect 39396 13268 39448 13277
rect 40040 13311 40092 13320
rect 40040 13277 40049 13311
rect 40049 13277 40083 13311
rect 40083 13277 40092 13311
rect 40040 13268 40092 13277
rect 40684 13268 40736 13320
rect 54024 13311 54076 13320
rect 54024 13277 54033 13311
rect 54033 13277 54067 13311
rect 54067 13277 54076 13311
rect 54024 13268 54076 13277
rect 32680 13200 32732 13252
rect 34428 13200 34480 13252
rect 35992 13243 36044 13252
rect 35992 13209 36010 13243
rect 36010 13209 36044 13243
rect 35992 13200 36044 13209
rect 20720 13132 20772 13184
rect 24124 13132 24176 13184
rect 24400 13132 24452 13184
rect 27252 13175 27304 13184
rect 27252 13141 27261 13175
rect 27261 13141 27295 13175
rect 27295 13141 27304 13175
rect 27252 13132 27304 13141
rect 28816 13132 28868 13184
rect 28908 13132 28960 13184
rect 30380 13132 30432 13184
rect 30656 13132 30708 13184
rect 31208 13175 31260 13184
rect 31208 13141 31217 13175
rect 31217 13141 31251 13175
rect 31251 13141 31260 13175
rect 31208 13132 31260 13141
rect 33048 13132 33100 13184
rect 35532 13132 35584 13184
rect 37372 13132 37424 13184
rect 40132 13200 40184 13252
rect 39028 13175 39080 13184
rect 39028 13141 39037 13175
rect 39037 13141 39071 13175
rect 39071 13141 39080 13175
rect 39028 13132 39080 13141
rect 39764 13132 39816 13184
rect 41144 13132 41196 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 1860 12928 1912 12980
rect 14188 12928 14240 12980
rect 16120 12928 16172 12980
rect 17040 12971 17092 12980
rect 17040 12937 17049 12971
rect 17049 12937 17083 12971
rect 17083 12937 17092 12971
rect 17040 12928 17092 12937
rect 17132 12928 17184 12980
rect 18236 12971 18288 12980
rect 18236 12937 18245 12971
rect 18245 12937 18279 12971
rect 18279 12937 18288 12971
rect 18236 12928 18288 12937
rect 15108 12903 15160 12912
rect 15108 12869 15117 12903
rect 15117 12869 15151 12903
rect 15151 12869 15160 12903
rect 15108 12860 15160 12869
rect 13176 12792 13228 12844
rect 13360 12792 13412 12844
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13728 12835 13780 12844
rect 13544 12792 13596 12801
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 14188 12792 14240 12844
rect 14740 12792 14792 12844
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 16304 12792 16356 12844
rect 17592 12860 17644 12912
rect 19984 12928 20036 12980
rect 20168 12928 20220 12980
rect 15936 12767 15988 12776
rect 15936 12733 15945 12767
rect 15945 12733 15979 12767
rect 15979 12733 15988 12767
rect 15936 12724 15988 12733
rect 15844 12656 15896 12708
rect 16212 12767 16264 12776
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 19984 12792 20036 12844
rect 20076 12835 20128 12844
rect 20076 12801 20085 12835
rect 20085 12801 20119 12835
rect 20119 12801 20128 12835
rect 22284 12860 22336 12912
rect 22560 12860 22612 12912
rect 23020 12903 23072 12912
rect 23020 12869 23029 12903
rect 23029 12869 23063 12903
rect 23063 12869 23072 12903
rect 23020 12860 23072 12869
rect 26608 12928 26660 12980
rect 27988 12971 28040 12980
rect 27988 12937 27997 12971
rect 27997 12937 28031 12971
rect 28031 12937 28040 12971
rect 27988 12928 28040 12937
rect 29736 12928 29788 12980
rect 26240 12860 26292 12912
rect 27160 12860 27212 12912
rect 27436 12860 27488 12912
rect 28448 12860 28500 12912
rect 20352 12835 20404 12844
rect 20076 12792 20128 12801
rect 20352 12801 20386 12835
rect 20386 12801 20404 12835
rect 20352 12792 20404 12801
rect 20720 12792 20772 12844
rect 21456 12792 21508 12844
rect 22100 12792 22152 12844
rect 24032 12835 24084 12844
rect 24032 12801 24041 12835
rect 24041 12801 24075 12835
rect 24075 12801 24084 12835
rect 24032 12792 24084 12801
rect 25320 12792 25372 12844
rect 16212 12724 16264 12733
rect 18144 12724 18196 12776
rect 17960 12656 18012 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 19340 12588 19392 12640
rect 20720 12588 20772 12640
rect 23848 12724 23900 12776
rect 21456 12699 21508 12708
rect 21456 12665 21465 12699
rect 21465 12665 21499 12699
rect 21499 12665 21508 12699
rect 21456 12656 21508 12665
rect 22744 12656 22796 12708
rect 21180 12588 21232 12640
rect 24952 12588 25004 12640
rect 26148 12656 26200 12708
rect 28816 12835 28868 12844
rect 28816 12801 28825 12835
rect 28825 12801 28859 12835
rect 28859 12801 28868 12835
rect 28816 12792 28868 12801
rect 29828 12860 29880 12912
rect 30564 12928 30616 12980
rect 32128 12928 32180 12980
rect 29736 12835 29788 12844
rect 29736 12801 29746 12835
rect 29746 12801 29780 12835
rect 29780 12801 29788 12835
rect 29736 12792 29788 12801
rect 30656 12860 30708 12912
rect 30012 12835 30064 12844
rect 30012 12801 30021 12835
rect 30021 12801 30055 12835
rect 30055 12801 30064 12835
rect 30012 12792 30064 12801
rect 30748 12792 30800 12844
rect 31392 12860 31444 12912
rect 31024 12835 31076 12844
rect 31024 12801 31033 12835
rect 31033 12801 31067 12835
rect 31067 12801 31076 12835
rect 31024 12792 31076 12801
rect 31208 12835 31260 12844
rect 31208 12801 31217 12835
rect 31217 12801 31251 12835
rect 31251 12801 31260 12835
rect 31208 12792 31260 12801
rect 32772 12860 32824 12912
rect 35716 12860 35768 12912
rect 36544 12928 36596 12980
rect 32588 12835 32640 12844
rect 32588 12801 32597 12835
rect 32597 12801 32631 12835
rect 32631 12801 32640 12835
rect 32588 12792 32640 12801
rect 33140 12792 33192 12844
rect 33784 12792 33836 12844
rect 35348 12835 35400 12844
rect 35348 12801 35357 12835
rect 35357 12801 35391 12835
rect 35391 12801 35400 12835
rect 35348 12792 35400 12801
rect 36360 12835 36412 12844
rect 32404 12724 32456 12776
rect 26516 12588 26568 12640
rect 27344 12588 27396 12640
rect 30288 12631 30340 12640
rect 30288 12597 30297 12631
rect 30297 12597 30331 12631
rect 30331 12597 30340 12631
rect 30288 12588 30340 12597
rect 31208 12656 31260 12708
rect 31392 12656 31444 12708
rect 32220 12656 32272 12708
rect 32772 12767 32824 12776
rect 32772 12733 32781 12767
rect 32781 12733 32815 12767
rect 32815 12733 32824 12767
rect 32772 12724 32824 12733
rect 33692 12724 33744 12776
rect 36360 12801 36369 12835
rect 36369 12801 36403 12835
rect 36403 12801 36412 12835
rect 36360 12792 36412 12801
rect 37740 12860 37792 12912
rect 38844 12928 38896 12980
rect 39948 12928 40000 12980
rect 41420 12928 41472 12980
rect 53840 12928 53892 12980
rect 54208 12971 54260 12980
rect 54208 12937 54217 12971
rect 54217 12937 54251 12971
rect 54251 12937 54260 12971
rect 54208 12928 54260 12937
rect 38384 12792 38436 12844
rect 40132 12835 40184 12844
rect 40132 12801 40141 12835
rect 40141 12801 40175 12835
rect 40175 12801 40184 12835
rect 40132 12792 40184 12801
rect 40500 12792 40552 12844
rect 41788 12792 41840 12844
rect 36268 12767 36320 12776
rect 36268 12733 36277 12767
rect 36277 12733 36311 12767
rect 36311 12733 36320 12767
rect 36268 12724 36320 12733
rect 38200 12724 38252 12776
rect 32128 12588 32180 12640
rect 32312 12631 32364 12640
rect 32312 12597 32321 12631
rect 32321 12597 32355 12631
rect 32355 12597 32364 12631
rect 32312 12588 32364 12597
rect 34244 12631 34296 12640
rect 34244 12597 34253 12631
rect 34253 12597 34287 12631
rect 34287 12597 34296 12631
rect 34244 12588 34296 12597
rect 34520 12588 34572 12640
rect 37648 12631 37700 12640
rect 37648 12597 37657 12631
rect 37657 12597 37691 12631
rect 37691 12597 37700 12631
rect 37648 12588 37700 12597
rect 39396 12656 39448 12708
rect 41788 12588 41840 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 13544 12384 13596 12436
rect 15844 12427 15896 12436
rect 15844 12393 15853 12427
rect 15853 12393 15887 12427
rect 15887 12393 15896 12427
rect 15844 12384 15896 12393
rect 17316 12427 17368 12436
rect 17316 12393 17325 12427
rect 17325 12393 17359 12427
rect 17359 12393 17368 12427
rect 17316 12384 17368 12393
rect 17592 12384 17644 12436
rect 20812 12384 20864 12436
rect 22560 12384 22612 12436
rect 16672 12316 16724 12368
rect 17040 12316 17092 12368
rect 17868 12316 17920 12368
rect 19800 12316 19852 12368
rect 15752 12248 15804 12300
rect 18236 12248 18288 12300
rect 18880 12248 18932 12300
rect 13912 12180 13964 12232
rect 15936 12180 15988 12232
rect 14004 12112 14056 12164
rect 15200 12112 15252 12164
rect 16120 12112 16172 12164
rect 16580 12180 16632 12232
rect 16672 12180 16724 12232
rect 17132 12180 17184 12232
rect 17868 12180 17920 12232
rect 18144 12180 18196 12232
rect 19248 12180 19300 12232
rect 20628 12248 20680 12300
rect 21180 12291 21232 12300
rect 21180 12257 21189 12291
rect 21189 12257 21223 12291
rect 21223 12257 21232 12291
rect 21180 12248 21232 12257
rect 23204 12316 23256 12368
rect 23940 12248 23992 12300
rect 26608 12384 26660 12436
rect 29092 12384 29144 12436
rect 29736 12384 29788 12436
rect 30012 12384 30064 12436
rect 31116 12427 31168 12436
rect 31116 12393 31125 12427
rect 31125 12393 31159 12427
rect 31159 12393 31168 12427
rect 31116 12384 31168 12393
rect 31484 12384 31536 12436
rect 20720 12180 20772 12232
rect 23664 12223 23716 12232
rect 23664 12189 23673 12223
rect 23673 12189 23707 12223
rect 23707 12189 23716 12223
rect 23664 12180 23716 12189
rect 25412 12180 25464 12232
rect 22192 12155 22244 12164
rect 1676 12087 1728 12096
rect 1676 12053 1685 12087
rect 1685 12053 1719 12087
rect 1719 12053 1728 12087
rect 1676 12044 1728 12053
rect 12624 12087 12676 12096
rect 12624 12053 12633 12087
rect 12633 12053 12667 12087
rect 12667 12053 12676 12087
rect 12624 12044 12676 12053
rect 13728 12044 13780 12096
rect 14832 12044 14884 12096
rect 15016 12044 15068 12096
rect 15844 12044 15896 12096
rect 22192 12121 22201 12155
rect 22201 12121 22235 12155
rect 22235 12121 22244 12155
rect 22192 12112 22244 12121
rect 22468 12155 22520 12164
rect 22468 12121 22477 12155
rect 22477 12121 22511 12155
rect 22511 12121 22520 12155
rect 22468 12112 22520 12121
rect 24032 12112 24084 12164
rect 25044 12112 25096 12164
rect 27160 12248 27212 12300
rect 29000 12316 29052 12368
rect 34060 12316 34112 12368
rect 34244 12316 34296 12368
rect 34520 12316 34572 12368
rect 34704 12316 34756 12368
rect 34796 12316 34848 12368
rect 36360 12384 36412 12436
rect 37556 12384 37608 12436
rect 37740 12384 37792 12436
rect 38384 12384 38436 12436
rect 40040 12427 40092 12436
rect 40040 12393 40049 12427
rect 40049 12393 40083 12427
rect 40083 12393 40092 12427
rect 40040 12384 40092 12393
rect 38844 12316 38896 12368
rect 28540 12248 28592 12300
rect 30840 12248 30892 12300
rect 32128 12291 32180 12300
rect 32128 12257 32137 12291
rect 32137 12257 32171 12291
rect 32171 12257 32180 12291
rect 32128 12248 32180 12257
rect 18052 12044 18104 12096
rect 18512 12087 18564 12096
rect 18512 12053 18521 12087
rect 18521 12053 18555 12087
rect 18555 12053 18564 12087
rect 18512 12044 18564 12053
rect 20076 12044 20128 12096
rect 20168 12044 20220 12096
rect 20904 12087 20956 12096
rect 20904 12053 20913 12087
rect 20913 12053 20947 12087
rect 20947 12053 20956 12087
rect 20904 12044 20956 12053
rect 20996 12087 21048 12096
rect 20996 12053 21005 12087
rect 21005 12053 21039 12087
rect 21039 12053 21048 12087
rect 20996 12044 21048 12053
rect 22376 12044 22428 12096
rect 22836 12044 22888 12096
rect 23020 12044 23072 12096
rect 24216 12044 24268 12096
rect 26332 12044 26384 12096
rect 26884 12044 26936 12096
rect 29644 12180 29696 12232
rect 29828 12180 29880 12232
rect 30748 12180 30800 12232
rect 33140 12180 33192 12232
rect 37096 12248 37148 12300
rect 37740 12291 37792 12300
rect 37740 12257 37749 12291
rect 37749 12257 37783 12291
rect 37783 12257 37792 12291
rect 37740 12248 37792 12257
rect 38292 12248 38344 12300
rect 28908 12112 28960 12164
rect 28264 12044 28316 12096
rect 29276 12112 29328 12164
rect 30656 12112 30708 12164
rect 31668 12112 31720 12164
rect 33508 12112 33560 12164
rect 36544 12180 36596 12232
rect 36728 12180 36780 12232
rect 36912 12180 36964 12232
rect 37004 12180 37056 12232
rect 35348 12155 35400 12164
rect 35348 12121 35357 12155
rect 35357 12121 35391 12155
rect 35391 12121 35400 12155
rect 35348 12112 35400 12121
rect 37188 12112 37240 12164
rect 38476 12223 38528 12232
rect 38476 12189 38485 12223
rect 38485 12189 38519 12223
rect 38519 12189 38528 12223
rect 38476 12180 38528 12189
rect 39028 12248 39080 12300
rect 39304 12180 39356 12232
rect 49700 12180 49752 12232
rect 54208 12223 54260 12232
rect 54208 12189 54217 12223
rect 54217 12189 54251 12223
rect 54251 12189 54260 12223
rect 54208 12180 54260 12189
rect 39764 12112 39816 12164
rect 53196 12112 53248 12164
rect 53472 12155 53524 12164
rect 53472 12121 53481 12155
rect 53481 12121 53515 12155
rect 53515 12121 53524 12155
rect 53472 12112 53524 12121
rect 53564 12112 53616 12164
rect 31576 12087 31628 12096
rect 31576 12053 31585 12087
rect 31585 12053 31619 12087
rect 31619 12053 31628 12087
rect 31576 12044 31628 12053
rect 31760 12044 31812 12096
rect 33600 12044 33652 12096
rect 34704 12044 34756 12096
rect 34796 12044 34848 12096
rect 36636 12044 36688 12096
rect 37372 12044 37424 12096
rect 37648 12044 37700 12096
rect 39396 12044 39448 12096
rect 41236 12044 41288 12096
rect 41788 12087 41840 12096
rect 41788 12053 41797 12087
rect 41797 12053 41831 12087
rect 41831 12053 41840 12087
rect 41788 12044 41840 12053
rect 42524 12044 42576 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 13360 11840 13412 11892
rect 15752 11883 15804 11892
rect 15752 11849 15761 11883
rect 15761 11849 15795 11883
rect 15795 11849 15804 11883
rect 15752 11840 15804 11849
rect 18512 11840 18564 11892
rect 18788 11840 18840 11892
rect 16948 11772 17000 11824
rect 20904 11840 20956 11892
rect 15844 11704 15896 11756
rect 17592 11704 17644 11756
rect 17960 11704 18012 11756
rect 22284 11772 22336 11824
rect 22652 11772 22704 11824
rect 23572 11772 23624 11824
rect 23756 11772 23808 11824
rect 26240 11840 26292 11892
rect 27344 11840 27396 11892
rect 29644 11883 29696 11892
rect 28908 11772 28960 11824
rect 29092 11815 29144 11824
rect 29092 11781 29101 11815
rect 29101 11781 29135 11815
rect 29135 11781 29144 11815
rect 29092 11772 29144 11781
rect 19432 11704 19484 11756
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 15108 11679 15160 11688
rect 15108 11645 15117 11679
rect 15117 11645 15151 11679
rect 15151 11645 15160 11679
rect 15108 11636 15160 11645
rect 15200 11679 15252 11688
rect 15200 11645 15209 11679
rect 15209 11645 15243 11679
rect 15243 11645 15252 11679
rect 15936 11679 15988 11688
rect 15200 11636 15252 11645
rect 15936 11645 15945 11679
rect 15945 11645 15979 11679
rect 15979 11645 15988 11679
rect 15936 11636 15988 11645
rect 16120 11679 16172 11688
rect 16120 11645 16129 11679
rect 16129 11645 16163 11679
rect 16163 11645 16172 11679
rect 16120 11636 16172 11645
rect 15292 11568 15344 11620
rect 19340 11636 19392 11688
rect 20996 11704 21048 11756
rect 24860 11704 24912 11756
rect 22284 11636 22336 11688
rect 22836 11679 22888 11688
rect 22836 11645 22845 11679
rect 22845 11645 22879 11679
rect 22879 11645 22888 11679
rect 22836 11636 22888 11645
rect 23664 11636 23716 11688
rect 24216 11636 24268 11688
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 28540 11679 28592 11688
rect 28540 11645 28549 11679
rect 28549 11645 28583 11679
rect 28583 11645 28592 11679
rect 28540 11636 28592 11645
rect 1676 11543 1728 11552
rect 1676 11509 1685 11543
rect 1685 11509 1719 11543
rect 1719 11509 1728 11543
rect 1676 11500 1728 11509
rect 13176 11543 13228 11552
rect 13176 11509 13185 11543
rect 13185 11509 13219 11543
rect 13219 11509 13228 11543
rect 13176 11500 13228 11509
rect 13728 11500 13780 11552
rect 17776 11500 17828 11552
rect 19248 11543 19300 11552
rect 19248 11509 19257 11543
rect 19257 11509 19291 11543
rect 19291 11509 19300 11543
rect 22376 11611 22428 11620
rect 22376 11577 22385 11611
rect 22385 11577 22419 11611
rect 22419 11577 22428 11611
rect 22376 11568 22428 11577
rect 19248 11500 19300 11509
rect 20904 11500 20956 11552
rect 22192 11500 22244 11552
rect 27160 11543 27212 11552
rect 27160 11509 27169 11543
rect 27169 11509 27203 11543
rect 27203 11509 27212 11543
rect 27160 11500 27212 11509
rect 27620 11500 27672 11552
rect 29644 11849 29653 11883
rect 29653 11849 29687 11883
rect 29687 11849 29696 11883
rect 29644 11840 29696 11849
rect 30012 11883 30064 11892
rect 30012 11849 30021 11883
rect 30021 11849 30055 11883
rect 30055 11849 30064 11883
rect 30012 11840 30064 11849
rect 31484 11883 31536 11892
rect 31484 11849 31493 11883
rect 31493 11849 31527 11883
rect 31527 11849 31536 11883
rect 31484 11840 31536 11849
rect 31668 11840 31720 11892
rect 33508 11840 33560 11892
rect 35900 11840 35952 11892
rect 37740 11840 37792 11892
rect 29920 11772 29972 11824
rect 30748 11772 30800 11824
rect 29092 11636 29144 11688
rect 30288 11704 30340 11756
rect 31760 11772 31812 11824
rect 39212 11840 39264 11892
rect 39304 11840 39356 11892
rect 41144 11883 41196 11892
rect 41144 11849 41153 11883
rect 41153 11849 41187 11883
rect 41187 11849 41196 11883
rect 41144 11840 41196 11849
rect 41236 11840 41288 11892
rect 53564 11883 53616 11892
rect 53564 11849 53573 11883
rect 53573 11849 53607 11883
rect 53607 11849 53616 11883
rect 53564 11840 53616 11849
rect 54208 11883 54260 11892
rect 54208 11849 54217 11883
rect 54217 11849 54251 11883
rect 54251 11849 54260 11883
rect 54208 11840 54260 11849
rect 31208 11747 31260 11756
rect 31208 11713 31217 11747
rect 31217 11713 31251 11747
rect 31251 11713 31260 11747
rect 34796 11747 34848 11756
rect 31208 11704 31260 11713
rect 34796 11713 34805 11747
rect 34805 11713 34839 11747
rect 34839 11713 34848 11747
rect 34796 11704 34848 11713
rect 35992 11704 36044 11756
rect 29460 11568 29512 11620
rect 30656 11568 30708 11620
rect 32588 11636 32640 11688
rect 35348 11636 35400 11688
rect 32864 11568 32916 11620
rect 33232 11568 33284 11620
rect 36820 11704 36872 11756
rect 37648 11747 37700 11756
rect 37648 11713 37657 11747
rect 37657 11713 37691 11747
rect 37691 11713 37700 11747
rect 37648 11704 37700 11713
rect 38200 11704 38252 11756
rect 39120 11772 39172 11824
rect 40960 11772 41012 11824
rect 40040 11704 40092 11756
rect 40224 11704 40276 11756
rect 51080 11772 51132 11824
rect 46940 11704 46992 11756
rect 38384 11568 38436 11620
rect 41144 11636 41196 11688
rect 43628 11636 43680 11688
rect 29644 11500 29696 11552
rect 31852 11500 31904 11552
rect 33876 11500 33928 11552
rect 37648 11500 37700 11552
rect 39212 11500 39264 11552
rect 40500 11500 40552 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 15292 11296 15344 11348
rect 16212 11296 16264 11348
rect 14464 11228 14516 11280
rect 15936 11271 15988 11280
rect 15936 11237 15945 11271
rect 15945 11237 15979 11271
rect 15979 11237 15988 11271
rect 15936 11228 15988 11237
rect 15292 11160 15344 11212
rect 16120 11160 16172 11212
rect 11060 11092 11112 11144
rect 15016 11092 15068 11144
rect 23848 11296 23900 11348
rect 25044 11339 25096 11348
rect 25044 11305 25053 11339
rect 25053 11305 25087 11339
rect 25087 11305 25096 11339
rect 25044 11296 25096 11305
rect 27160 11296 27212 11348
rect 35992 11339 36044 11348
rect 18696 11228 18748 11280
rect 20168 11228 20220 11280
rect 23940 11228 23992 11280
rect 13820 11024 13872 11076
rect 14004 11024 14056 11076
rect 1676 10999 1728 11008
rect 1676 10965 1685 10999
rect 1685 10965 1719 10999
rect 1719 10965 1728 10999
rect 1676 10956 1728 10965
rect 13728 10999 13780 11008
rect 13728 10965 13737 10999
rect 13737 10965 13771 10999
rect 13771 10965 13780 10999
rect 13728 10956 13780 10965
rect 15844 10956 15896 11008
rect 16672 11024 16724 11076
rect 16856 11024 16908 11076
rect 19340 11092 19392 11144
rect 22284 11135 22336 11144
rect 22284 11101 22293 11135
rect 22293 11101 22327 11135
rect 22327 11101 22336 11135
rect 22284 11092 22336 11101
rect 26608 11160 26660 11212
rect 29460 11228 29512 11280
rect 32036 11228 32088 11280
rect 33416 11228 33468 11280
rect 33876 11228 33928 11280
rect 35992 11305 36001 11339
rect 36001 11305 36035 11339
rect 36035 11305 36044 11339
rect 35992 11296 36044 11305
rect 27988 11160 28040 11212
rect 24952 11092 25004 11144
rect 26332 11135 26384 11144
rect 26332 11101 26341 11135
rect 26341 11101 26375 11135
rect 26375 11101 26384 11135
rect 26332 11092 26384 11101
rect 27068 11092 27120 11144
rect 27436 11092 27488 11144
rect 17776 11067 17828 11076
rect 17776 11033 17810 11067
rect 17810 11033 17828 11067
rect 17776 11024 17828 11033
rect 20812 11024 20864 11076
rect 21456 11024 21508 11076
rect 22836 11024 22888 11076
rect 24768 11024 24820 11076
rect 26148 11024 26200 11076
rect 17316 10956 17368 11008
rect 18604 10956 18656 11008
rect 20076 10956 20128 11008
rect 23664 10999 23716 11008
rect 23664 10965 23673 10999
rect 23673 10965 23707 10999
rect 23707 10965 23716 10999
rect 23664 10956 23716 10965
rect 27344 10956 27396 11008
rect 28632 11092 28684 11144
rect 30564 11135 30616 11144
rect 28724 11067 28776 11076
rect 28724 11033 28733 11067
rect 28733 11033 28767 11067
rect 28767 11033 28776 11067
rect 28724 11024 28776 11033
rect 29644 11024 29696 11076
rect 30196 11024 30248 11076
rect 30564 11101 30573 11135
rect 30573 11101 30607 11135
rect 30607 11101 30616 11135
rect 30564 11092 30616 11101
rect 30748 11135 30800 11144
rect 30748 11101 30752 11135
rect 30752 11101 30786 11135
rect 30786 11101 30800 11135
rect 30748 11092 30800 11101
rect 30840 11135 30892 11144
rect 30840 11101 30849 11135
rect 30849 11101 30883 11135
rect 30883 11101 30892 11135
rect 30840 11092 30892 11101
rect 31024 11092 31076 11144
rect 32864 11160 32916 11212
rect 31484 11092 31536 11144
rect 31668 11135 31720 11144
rect 31668 11101 31677 11135
rect 31677 11101 31711 11135
rect 31711 11101 31720 11135
rect 31668 11092 31720 11101
rect 31852 11135 31904 11144
rect 31852 11101 31861 11135
rect 31861 11101 31895 11135
rect 31895 11101 31904 11135
rect 31852 11092 31904 11101
rect 32036 11135 32088 11144
rect 32036 11101 32045 11135
rect 32045 11101 32079 11135
rect 32079 11101 32088 11135
rect 32036 11092 32088 11101
rect 33508 11092 33560 11144
rect 33600 11092 33652 11144
rect 34336 11135 34388 11144
rect 34336 11101 34345 11135
rect 34345 11101 34379 11135
rect 34379 11101 34388 11135
rect 34336 11092 34388 11101
rect 34796 11092 34848 11144
rect 35808 11092 35860 11144
rect 36084 11228 36136 11280
rect 37280 11296 37332 11348
rect 37372 11296 37424 11348
rect 37832 11296 37884 11348
rect 38384 11296 38436 11348
rect 40040 11339 40092 11348
rect 40040 11305 40049 11339
rect 40049 11305 40083 11339
rect 40083 11305 40092 11339
rect 40040 11296 40092 11305
rect 40960 11339 41012 11348
rect 40960 11305 40969 11339
rect 40969 11305 41003 11339
rect 41003 11305 41012 11339
rect 40960 11296 41012 11305
rect 36452 11228 36504 11280
rect 54208 11271 54260 11280
rect 54208 11237 54217 11271
rect 54217 11237 54251 11271
rect 54251 11237 54260 11271
rect 54208 11228 54260 11237
rect 37372 11160 37424 11212
rect 32588 11024 32640 11076
rect 32956 11024 33008 11076
rect 34704 11024 34756 11076
rect 36636 11135 36688 11144
rect 36636 11101 36645 11135
rect 36645 11101 36679 11135
rect 36679 11101 36688 11135
rect 36636 11092 36688 11101
rect 37188 11092 37240 11144
rect 40316 11160 40368 11212
rect 40500 11203 40552 11212
rect 40500 11169 40509 11203
rect 40509 11169 40543 11203
rect 40543 11169 40552 11203
rect 40500 11160 40552 11169
rect 37004 11024 37056 11076
rect 37372 11067 37424 11076
rect 32680 10956 32732 11008
rect 33232 10999 33284 11008
rect 33232 10965 33241 10999
rect 33241 10965 33275 10999
rect 33275 10965 33284 10999
rect 33232 10956 33284 10965
rect 33692 10956 33744 11008
rect 35624 10956 35676 11008
rect 36452 10956 36504 11008
rect 37372 11033 37381 11067
rect 37381 11033 37415 11067
rect 37415 11033 37424 11067
rect 37372 11024 37424 11033
rect 37832 11092 37884 11144
rect 38108 11024 38160 11076
rect 38384 11135 38436 11144
rect 38384 11101 38393 11135
rect 38393 11101 38427 11135
rect 38427 11101 38436 11135
rect 38568 11135 38620 11144
rect 38384 11092 38436 11101
rect 38568 11101 38577 11135
rect 38577 11101 38611 11135
rect 38611 11101 38620 11135
rect 38568 11092 38620 11101
rect 38660 11135 38712 11144
rect 38660 11101 38669 11135
rect 38669 11101 38703 11135
rect 38703 11101 38712 11135
rect 38660 11092 38712 11101
rect 39212 11092 39264 11144
rect 39764 11092 39816 11144
rect 51080 11092 51132 11144
rect 40224 10956 40276 11008
rect 54208 10956 54260 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 11060 10752 11112 10804
rect 14004 10727 14056 10736
rect 14004 10693 14013 10727
rect 14013 10693 14047 10727
rect 14047 10693 14056 10727
rect 14004 10684 14056 10693
rect 16580 10752 16632 10804
rect 20996 10752 21048 10804
rect 17960 10684 18012 10736
rect 15016 10616 15068 10668
rect 13820 10548 13872 10600
rect 14924 10548 14976 10600
rect 15292 10591 15344 10600
rect 15292 10557 15301 10591
rect 15301 10557 15335 10591
rect 15335 10557 15344 10591
rect 15292 10548 15344 10557
rect 18052 10616 18104 10668
rect 18236 10616 18288 10668
rect 22836 10684 22888 10736
rect 20996 10659 21048 10668
rect 20996 10625 21005 10659
rect 21005 10625 21039 10659
rect 21039 10625 21048 10659
rect 20996 10616 21048 10625
rect 22744 10659 22796 10668
rect 22744 10625 22753 10659
rect 22753 10625 22787 10659
rect 22787 10625 22796 10659
rect 22744 10616 22796 10625
rect 23388 10659 23440 10668
rect 23388 10625 23397 10659
rect 23397 10625 23431 10659
rect 23431 10625 23440 10659
rect 23388 10616 23440 10625
rect 14280 10523 14332 10532
rect 14280 10489 14289 10523
rect 14289 10489 14323 10523
rect 14323 10489 14332 10523
rect 14280 10480 14332 10489
rect 14372 10480 14424 10532
rect 15568 10480 15620 10532
rect 17316 10591 17368 10600
rect 17316 10557 17325 10591
rect 17325 10557 17359 10591
rect 17359 10557 17368 10591
rect 17316 10548 17368 10557
rect 18052 10480 18104 10532
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 15200 10412 15252 10464
rect 20076 10548 20128 10600
rect 21180 10591 21232 10600
rect 21180 10557 21189 10591
rect 21189 10557 21223 10591
rect 21223 10557 21232 10591
rect 21180 10548 21232 10557
rect 23020 10548 23072 10600
rect 19248 10480 19300 10532
rect 22468 10480 22520 10532
rect 19340 10412 19392 10464
rect 20628 10455 20680 10464
rect 20628 10421 20637 10455
rect 20637 10421 20671 10455
rect 20671 10421 20680 10455
rect 20628 10412 20680 10421
rect 22560 10412 22612 10464
rect 23848 10412 23900 10464
rect 24768 10752 24820 10804
rect 26424 10752 26476 10804
rect 29184 10795 29236 10804
rect 29184 10761 29193 10795
rect 29193 10761 29227 10795
rect 29227 10761 29236 10795
rect 29184 10752 29236 10761
rect 27160 10684 27212 10736
rect 26240 10659 26292 10668
rect 26240 10625 26249 10659
rect 26249 10625 26283 10659
rect 26283 10625 26292 10659
rect 26240 10616 26292 10625
rect 27344 10659 27396 10668
rect 27344 10625 27353 10659
rect 27353 10625 27387 10659
rect 27387 10625 27396 10659
rect 27344 10616 27396 10625
rect 28172 10659 28224 10668
rect 28172 10625 28181 10659
rect 28181 10625 28215 10659
rect 28215 10625 28224 10659
rect 28172 10616 28224 10625
rect 30104 10752 30156 10804
rect 31668 10752 31720 10804
rect 32772 10752 32824 10804
rect 34060 10752 34112 10804
rect 35532 10752 35584 10804
rect 37556 10795 37608 10804
rect 37556 10761 37565 10795
rect 37565 10761 37599 10795
rect 37599 10761 37608 10795
rect 37556 10752 37608 10761
rect 37740 10752 37792 10804
rect 38936 10752 38988 10804
rect 41420 10752 41472 10804
rect 42064 10752 42116 10804
rect 29644 10684 29696 10736
rect 29920 10684 29972 10736
rect 29828 10659 29880 10668
rect 29828 10625 29837 10659
rect 29837 10625 29871 10659
rect 29871 10625 29880 10659
rect 29828 10616 29880 10625
rect 31392 10684 31444 10736
rect 31852 10684 31904 10736
rect 26332 10548 26384 10600
rect 29184 10548 29236 10600
rect 29736 10591 29788 10600
rect 29736 10557 29745 10591
rect 29745 10557 29779 10591
rect 29779 10557 29788 10591
rect 29736 10548 29788 10557
rect 29920 10591 29972 10600
rect 29920 10557 29929 10591
rect 29929 10557 29963 10591
rect 29963 10557 29972 10591
rect 30748 10616 30800 10668
rect 30932 10659 30984 10668
rect 30932 10625 30941 10659
rect 30941 10625 30975 10659
rect 30975 10625 30984 10659
rect 30932 10616 30984 10625
rect 31484 10616 31536 10668
rect 32772 10659 32824 10668
rect 32772 10625 32781 10659
rect 32781 10625 32815 10659
rect 32815 10625 32824 10659
rect 32772 10616 32824 10625
rect 29920 10548 29972 10557
rect 32312 10548 32364 10600
rect 33140 10616 33192 10668
rect 34796 10616 34848 10668
rect 35808 10616 35860 10668
rect 36360 10659 36412 10668
rect 35348 10591 35400 10600
rect 35348 10557 35357 10591
rect 35357 10557 35391 10591
rect 35391 10557 35400 10591
rect 35348 10548 35400 10557
rect 32496 10480 32548 10532
rect 36360 10625 36369 10659
rect 36369 10625 36403 10659
rect 36403 10625 36412 10659
rect 36360 10616 36412 10625
rect 36452 10659 36504 10668
rect 36452 10625 36461 10659
rect 36461 10625 36495 10659
rect 36495 10625 36504 10659
rect 36452 10616 36504 10625
rect 37740 10659 37792 10668
rect 37740 10625 37749 10659
rect 37749 10625 37783 10659
rect 37783 10625 37792 10659
rect 37740 10616 37792 10625
rect 38476 10659 38528 10668
rect 38476 10625 38510 10659
rect 38510 10625 38528 10659
rect 48964 10684 49016 10736
rect 54208 10727 54260 10736
rect 54208 10693 54217 10727
rect 54217 10693 54251 10727
rect 54251 10693 54260 10727
rect 54208 10684 54260 10693
rect 38476 10616 38528 10625
rect 40316 10616 40368 10668
rect 41420 10659 41472 10668
rect 41420 10625 41429 10659
rect 41429 10625 41463 10659
rect 41463 10625 41472 10659
rect 53472 10659 53524 10668
rect 41420 10616 41472 10625
rect 53472 10625 53481 10659
rect 53481 10625 53515 10659
rect 53515 10625 53524 10659
rect 53472 10616 53524 10625
rect 37924 10548 37976 10600
rect 38200 10591 38252 10600
rect 38200 10557 38209 10591
rect 38209 10557 38243 10591
rect 38243 10557 38252 10591
rect 38200 10548 38252 10557
rect 25872 10412 25924 10464
rect 27528 10455 27580 10464
rect 27528 10421 27537 10455
rect 27537 10421 27571 10455
rect 27571 10421 27580 10455
rect 27528 10412 27580 10421
rect 27988 10455 28040 10464
rect 27988 10421 27997 10455
rect 27997 10421 28031 10455
rect 28031 10421 28040 10455
rect 27988 10412 28040 10421
rect 30748 10412 30800 10464
rect 36360 10412 36412 10464
rect 36912 10455 36964 10464
rect 36912 10421 36921 10455
rect 36921 10421 36955 10455
rect 36955 10421 36964 10455
rect 36912 10412 36964 10421
rect 53288 10480 53340 10532
rect 38384 10412 38436 10464
rect 39580 10455 39632 10464
rect 39580 10421 39589 10455
rect 39589 10421 39623 10455
rect 39623 10421 39632 10455
rect 39580 10412 39632 10421
rect 41328 10455 41380 10464
rect 41328 10421 41337 10455
rect 41337 10421 41371 10455
rect 41371 10421 41380 10455
rect 41328 10412 41380 10421
rect 53380 10455 53432 10464
rect 53380 10421 53389 10455
rect 53389 10421 53423 10455
rect 53423 10421 53432 10455
rect 53380 10412 53432 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 14372 10208 14424 10260
rect 15016 10251 15068 10260
rect 15016 10217 15025 10251
rect 15025 10217 15059 10251
rect 15059 10217 15068 10251
rect 15016 10208 15068 10217
rect 16028 10208 16080 10260
rect 13176 10140 13228 10192
rect 15292 10140 15344 10192
rect 14004 10072 14056 10124
rect 15660 10072 15712 10124
rect 15016 10004 15068 10056
rect 15200 10047 15252 10056
rect 15200 10013 15209 10047
rect 15209 10013 15243 10047
rect 15243 10013 15252 10047
rect 15200 10004 15252 10013
rect 15476 10047 15528 10056
rect 15476 10013 15485 10047
rect 15485 10013 15519 10047
rect 15519 10013 15528 10047
rect 15476 10004 15528 10013
rect 16856 10140 16908 10192
rect 17776 10208 17828 10260
rect 17868 10208 17920 10260
rect 19432 10208 19484 10260
rect 19984 10208 20036 10260
rect 21640 10208 21692 10260
rect 23572 10251 23624 10260
rect 20996 10140 21048 10192
rect 23572 10217 23581 10251
rect 23581 10217 23615 10251
rect 23615 10217 23624 10251
rect 23572 10208 23624 10217
rect 28356 10251 28408 10260
rect 28356 10217 28365 10251
rect 28365 10217 28399 10251
rect 28399 10217 28408 10251
rect 28356 10208 28408 10217
rect 29276 10208 29328 10260
rect 29736 10208 29788 10260
rect 33692 10208 33744 10260
rect 18880 10072 18932 10124
rect 21180 10072 21232 10124
rect 17132 10004 17184 10056
rect 17868 10004 17920 10056
rect 17960 10004 18012 10056
rect 19248 10004 19300 10056
rect 1676 9911 1728 9920
rect 1676 9877 1685 9911
rect 1685 9877 1719 9911
rect 1719 9877 1728 9911
rect 1676 9868 1728 9877
rect 19064 9936 19116 9988
rect 21272 10004 21324 10056
rect 22100 10072 22152 10124
rect 22284 10004 22336 10056
rect 22468 10047 22520 10056
rect 22468 10013 22502 10047
rect 22502 10013 22520 10047
rect 22468 10004 22520 10013
rect 23664 10004 23716 10056
rect 22560 9936 22612 9988
rect 23940 9936 23992 9988
rect 29828 10140 29880 10192
rect 30380 10140 30432 10192
rect 30564 10140 30616 10192
rect 30656 10140 30708 10192
rect 33048 10140 33100 10192
rect 25228 10115 25280 10124
rect 25228 10081 25237 10115
rect 25237 10081 25271 10115
rect 25271 10081 25280 10115
rect 25228 10072 25280 10081
rect 27528 10072 27580 10124
rect 31852 10115 31904 10124
rect 25872 10004 25924 10056
rect 26056 10047 26108 10056
rect 26056 10013 26065 10047
rect 26065 10013 26099 10047
rect 26099 10013 26108 10047
rect 26056 10004 26108 10013
rect 28264 10047 28316 10056
rect 28264 10013 28273 10047
rect 28273 10013 28307 10047
rect 28307 10013 28316 10047
rect 28264 10004 28316 10013
rect 29000 10047 29052 10056
rect 29000 10013 29009 10047
rect 29009 10013 29043 10047
rect 29043 10013 29052 10047
rect 29000 10004 29052 10013
rect 30840 10004 30892 10056
rect 31852 10081 31861 10115
rect 31861 10081 31895 10115
rect 31895 10081 31904 10115
rect 31852 10072 31904 10081
rect 34520 10140 34572 10192
rect 35256 10140 35308 10192
rect 36268 10208 36320 10260
rect 38476 10208 38528 10260
rect 41328 10208 41380 10260
rect 48320 10208 48372 10260
rect 54208 10251 54260 10260
rect 54208 10217 54217 10251
rect 54217 10217 54251 10251
rect 54251 10217 54260 10251
rect 54208 10208 54260 10217
rect 53472 10183 53524 10192
rect 53472 10149 53481 10183
rect 53481 10149 53515 10183
rect 53515 10149 53524 10183
rect 53472 10140 53524 10149
rect 32772 10004 32824 10056
rect 33140 10047 33192 10056
rect 33140 10013 33149 10047
rect 33149 10013 33183 10047
rect 33183 10013 33192 10047
rect 33140 10004 33192 10013
rect 33324 10004 33376 10056
rect 33784 10004 33836 10056
rect 39580 10072 39632 10124
rect 26332 9936 26384 9988
rect 27896 9936 27948 9988
rect 29920 9936 29972 9988
rect 30288 9936 30340 9988
rect 30472 9979 30524 9988
rect 30472 9945 30481 9979
rect 30481 9945 30515 9979
rect 30515 9945 30524 9979
rect 30472 9936 30524 9945
rect 30748 9979 30800 9988
rect 30748 9945 30757 9979
rect 30757 9945 30791 9979
rect 30791 9945 30800 9979
rect 30748 9936 30800 9945
rect 34060 10004 34112 10056
rect 34980 10047 35032 10056
rect 34980 10013 34989 10047
rect 34989 10013 35023 10047
rect 35023 10013 35032 10047
rect 34980 10004 35032 10013
rect 34520 9936 34572 9988
rect 35624 10004 35676 10056
rect 18604 9911 18656 9920
rect 18604 9877 18613 9911
rect 18613 9877 18647 9911
rect 18647 9877 18656 9911
rect 19432 9911 19484 9920
rect 18604 9868 18656 9877
rect 19432 9877 19441 9911
rect 19441 9877 19475 9911
rect 19475 9877 19484 9911
rect 19432 9868 19484 9877
rect 19984 9868 20036 9920
rect 20260 9868 20312 9920
rect 21548 9911 21600 9920
rect 21548 9877 21557 9911
rect 21557 9877 21591 9911
rect 21591 9877 21600 9911
rect 21548 9868 21600 9877
rect 22100 9868 22152 9920
rect 25044 9911 25096 9920
rect 25044 9877 25053 9911
rect 25053 9877 25087 9911
rect 25087 9877 25096 9911
rect 25044 9868 25096 9877
rect 27620 9868 27672 9920
rect 30380 9868 30432 9920
rect 32956 9868 33008 9920
rect 34060 9911 34112 9920
rect 34060 9877 34069 9911
rect 34069 9877 34103 9911
rect 34103 9877 34112 9911
rect 35532 9936 35584 9988
rect 34060 9868 34112 9877
rect 35440 9868 35492 9920
rect 38200 10004 38252 10056
rect 38384 10004 38436 10056
rect 40224 10047 40276 10056
rect 40224 10013 40233 10047
rect 40233 10013 40267 10047
rect 40267 10013 40276 10047
rect 40224 10004 40276 10013
rect 53564 10072 53616 10124
rect 36912 9936 36964 9988
rect 39304 9979 39356 9988
rect 39304 9945 39313 9979
rect 39313 9945 39347 9979
rect 39347 9945 39356 9979
rect 39304 9936 39356 9945
rect 37924 9911 37976 9920
rect 37924 9877 37933 9911
rect 37933 9877 37967 9911
rect 37967 9877 37976 9911
rect 37924 9868 37976 9877
rect 38016 9868 38068 9920
rect 53380 9936 53432 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 15200 9664 15252 9716
rect 15384 9664 15436 9716
rect 17132 9664 17184 9716
rect 20168 9664 20220 9716
rect 20536 9664 20588 9716
rect 22836 9707 22888 9716
rect 22836 9673 22845 9707
rect 22845 9673 22879 9707
rect 22879 9673 22888 9707
rect 22836 9664 22888 9673
rect 14004 9596 14056 9648
rect 16212 9596 16264 9648
rect 17316 9639 17368 9648
rect 14556 9528 14608 9580
rect 15108 9571 15160 9580
rect 15108 9537 15117 9571
rect 15117 9537 15151 9571
rect 15151 9537 15160 9571
rect 15108 9528 15160 9537
rect 14096 9460 14148 9512
rect 14648 9460 14700 9512
rect 13360 9435 13412 9444
rect 13360 9401 13369 9435
rect 13369 9401 13403 9435
rect 13403 9401 13412 9435
rect 13360 9392 13412 9401
rect 15108 9392 15160 9444
rect 15752 9460 15804 9512
rect 16396 9460 16448 9512
rect 15660 9392 15712 9444
rect 16580 9392 16632 9444
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 15016 9324 15068 9376
rect 17316 9605 17325 9639
rect 17325 9605 17359 9639
rect 17359 9605 17368 9639
rect 17316 9596 17368 9605
rect 23572 9596 23624 9648
rect 25044 9664 25096 9716
rect 17776 9571 17828 9580
rect 17776 9537 17785 9571
rect 17785 9537 17819 9571
rect 17819 9537 17828 9571
rect 17776 9528 17828 9537
rect 18696 9528 18748 9580
rect 19984 9528 20036 9580
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 22100 9528 22152 9580
rect 22192 9571 22244 9580
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 23480 9528 23532 9580
rect 26332 9596 26384 9648
rect 24768 9571 24820 9580
rect 24768 9537 24777 9571
rect 24777 9537 24811 9571
rect 24811 9537 24820 9571
rect 24768 9528 24820 9537
rect 25872 9528 25924 9580
rect 26148 9571 26200 9580
rect 26148 9537 26157 9571
rect 26157 9537 26191 9571
rect 26191 9537 26200 9571
rect 26148 9528 26200 9537
rect 27160 9528 27212 9580
rect 28356 9596 28408 9648
rect 19524 9460 19576 9512
rect 19616 9460 19668 9512
rect 23112 9460 23164 9512
rect 23572 9460 23624 9512
rect 26332 9503 26384 9512
rect 18788 9435 18840 9444
rect 18788 9401 18797 9435
rect 18797 9401 18831 9435
rect 18831 9401 18840 9435
rect 18788 9392 18840 9401
rect 20076 9392 20128 9444
rect 20812 9435 20864 9444
rect 20812 9401 20821 9435
rect 20821 9401 20855 9435
rect 20855 9401 20864 9435
rect 20812 9392 20864 9401
rect 21456 9435 21508 9444
rect 21456 9401 21465 9435
rect 21465 9401 21499 9435
rect 21499 9401 21508 9435
rect 21456 9392 21508 9401
rect 23756 9392 23808 9444
rect 18972 9324 19024 9376
rect 19800 9324 19852 9376
rect 20720 9324 20772 9376
rect 21916 9324 21968 9376
rect 24124 9324 24176 9376
rect 26332 9469 26341 9503
rect 26341 9469 26375 9503
rect 26375 9469 26384 9503
rect 26332 9460 26384 9469
rect 27896 9528 27948 9580
rect 29460 9596 29512 9648
rect 28448 9503 28500 9512
rect 28448 9469 28457 9503
rect 28457 9469 28491 9503
rect 28491 9469 28500 9503
rect 28448 9460 28500 9469
rect 28908 9528 28960 9580
rect 29460 9503 29512 9512
rect 25964 9392 26016 9444
rect 26976 9392 27028 9444
rect 29460 9469 29469 9503
rect 29469 9469 29503 9503
rect 29503 9469 29512 9503
rect 29460 9460 29512 9469
rect 29736 9571 29788 9580
rect 29736 9537 29745 9571
rect 29745 9537 29779 9571
rect 29779 9537 29788 9571
rect 29736 9528 29788 9537
rect 30380 9528 30432 9580
rect 30932 9596 30984 9648
rect 31116 9596 31168 9648
rect 30656 9571 30708 9580
rect 30656 9537 30665 9571
rect 30665 9537 30699 9571
rect 30699 9537 30708 9571
rect 31852 9596 31904 9648
rect 33140 9664 33192 9716
rect 34060 9596 34112 9648
rect 30656 9528 30708 9537
rect 31668 9528 31720 9580
rect 31760 9528 31812 9580
rect 32036 9528 32088 9580
rect 32496 9528 32548 9580
rect 31116 9460 31168 9512
rect 33692 9503 33744 9512
rect 33692 9469 33701 9503
rect 33701 9469 33735 9503
rect 33735 9469 33744 9503
rect 35348 9596 35400 9648
rect 34704 9528 34756 9580
rect 35532 9664 35584 9716
rect 38016 9664 38068 9716
rect 38292 9664 38344 9716
rect 36544 9639 36596 9648
rect 36544 9605 36553 9639
rect 36553 9605 36587 9639
rect 36587 9605 36596 9639
rect 36544 9596 36596 9605
rect 37556 9528 37608 9580
rect 44456 9596 44508 9648
rect 38108 9528 38160 9580
rect 48412 9596 48464 9648
rect 53380 9596 53432 9648
rect 48780 9571 48832 9580
rect 48780 9537 48789 9571
rect 48789 9537 48823 9571
rect 48823 9537 48832 9571
rect 48780 9528 48832 9537
rect 49056 9571 49108 9580
rect 49056 9537 49090 9571
rect 49090 9537 49108 9571
rect 49056 9528 49108 9537
rect 33692 9460 33744 9469
rect 31576 9392 31628 9444
rect 32128 9392 32180 9444
rect 25780 9324 25832 9376
rect 28724 9324 28776 9376
rect 29828 9324 29880 9376
rect 30104 9367 30156 9376
rect 30104 9333 30113 9367
rect 30113 9333 30147 9367
rect 30147 9333 30156 9367
rect 30104 9324 30156 9333
rect 31760 9367 31812 9376
rect 31760 9333 31769 9367
rect 31769 9333 31803 9367
rect 31803 9333 31812 9367
rect 31760 9324 31812 9333
rect 32036 9324 32088 9376
rect 37372 9392 37424 9444
rect 50896 9528 50948 9580
rect 53564 9528 53616 9580
rect 35992 9367 36044 9376
rect 35992 9333 36001 9367
rect 36001 9333 36035 9367
rect 36035 9333 36044 9367
rect 35992 9324 36044 9333
rect 37004 9324 37056 9376
rect 37648 9324 37700 9376
rect 39120 9324 39172 9376
rect 43628 9324 43680 9376
rect 50436 9324 50488 9376
rect 54208 9435 54260 9444
rect 54208 9401 54217 9435
rect 54217 9401 54251 9435
rect 54251 9401 54260 9435
rect 54208 9392 54260 9401
rect 51632 9324 51684 9376
rect 52276 9367 52328 9376
rect 52276 9333 52285 9367
rect 52285 9333 52319 9367
rect 52319 9333 52328 9367
rect 52276 9324 52328 9333
rect 52460 9324 52512 9376
rect 53104 9324 53156 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 14556 9120 14608 9172
rect 13268 9052 13320 9104
rect 16212 9095 16264 9104
rect 16212 9061 16221 9095
rect 16221 9061 16255 9095
rect 16255 9061 16264 9095
rect 16212 9052 16264 9061
rect 16488 9120 16540 9172
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 17316 9120 17368 9172
rect 18236 9163 18288 9172
rect 18236 9129 18245 9163
rect 18245 9129 18279 9163
rect 18279 9129 18288 9163
rect 18236 9120 18288 9129
rect 21364 9120 21416 9172
rect 24032 9163 24084 9172
rect 24032 9129 24041 9163
rect 24041 9129 24075 9163
rect 24075 9129 24084 9163
rect 24032 9120 24084 9129
rect 24768 9120 24820 9172
rect 18328 9052 18380 9104
rect 18420 9052 18472 9104
rect 25780 9052 25832 9104
rect 17960 8984 18012 9036
rect 14096 8916 14148 8968
rect 14648 8959 14700 8968
rect 14648 8925 14657 8959
rect 14657 8925 14691 8959
rect 14691 8925 14700 8959
rect 14648 8916 14700 8925
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 19432 8984 19484 9036
rect 19524 8984 19576 9036
rect 21548 9027 21600 9036
rect 21548 8993 21557 9027
rect 21557 8993 21591 9027
rect 21591 8993 21600 9027
rect 21548 8984 21600 8993
rect 22836 8984 22888 9036
rect 25136 9027 25188 9036
rect 25136 8993 25145 9027
rect 25145 8993 25179 9027
rect 25179 8993 25188 9027
rect 25136 8984 25188 8993
rect 14740 8916 14792 8925
rect 1676 8823 1728 8832
rect 1676 8789 1685 8823
rect 1685 8789 1719 8823
rect 1719 8789 1728 8823
rect 1676 8780 1728 8789
rect 14556 8848 14608 8900
rect 14464 8780 14516 8832
rect 16948 8848 17000 8900
rect 17316 8848 17368 8900
rect 19800 8891 19852 8900
rect 18880 8823 18932 8832
rect 18880 8789 18889 8823
rect 18889 8789 18923 8823
rect 18923 8789 18932 8823
rect 18880 8780 18932 8789
rect 19800 8857 19809 8891
rect 19809 8857 19843 8891
rect 19843 8857 19852 8891
rect 19800 8848 19852 8857
rect 20076 8780 20128 8832
rect 21456 8916 21508 8968
rect 21640 8916 21692 8968
rect 23204 8959 23256 8968
rect 23204 8925 23213 8959
rect 23213 8925 23247 8959
rect 23247 8925 23256 8959
rect 23204 8916 23256 8925
rect 23848 8959 23900 8968
rect 23848 8925 23857 8959
rect 23857 8925 23891 8959
rect 23891 8925 23900 8959
rect 23848 8916 23900 8925
rect 26424 8984 26476 9036
rect 28172 9120 28224 9172
rect 28356 9120 28408 9172
rect 28540 9120 28592 9172
rect 31208 9120 31260 9172
rect 31668 9163 31720 9172
rect 31668 9129 31677 9163
rect 31677 9129 31711 9163
rect 31711 9129 31720 9163
rect 31668 9120 31720 9129
rect 34520 9120 34572 9172
rect 35808 9120 35860 9172
rect 38660 9120 38712 9172
rect 49056 9120 49108 9172
rect 49148 9120 49200 9172
rect 28448 9027 28500 9036
rect 28448 8993 28457 9027
rect 28457 8993 28491 9027
rect 28491 8993 28500 9027
rect 28448 8984 28500 8993
rect 29092 8984 29144 9036
rect 29460 8984 29512 9036
rect 31852 8984 31904 9036
rect 32312 9027 32364 9036
rect 32312 8993 32321 9027
rect 32321 8993 32355 9027
rect 32355 8993 32364 9027
rect 32312 8984 32364 8993
rect 32956 8984 33008 9036
rect 23756 8848 23808 8900
rect 21364 8780 21416 8832
rect 22560 8823 22612 8832
rect 22560 8789 22569 8823
rect 22569 8789 22603 8823
rect 22603 8789 22612 8823
rect 22560 8780 22612 8789
rect 23112 8780 23164 8832
rect 27436 8916 27488 8968
rect 27620 8916 27672 8968
rect 29736 8959 29788 8968
rect 29736 8925 29745 8959
rect 29745 8925 29779 8959
rect 29779 8925 29788 8959
rect 29736 8916 29788 8925
rect 29828 8916 29880 8968
rect 33324 8916 33376 8968
rect 33600 8984 33652 9036
rect 33784 8984 33836 9036
rect 35624 9052 35676 9104
rect 35900 9052 35952 9104
rect 42984 9052 43036 9104
rect 46204 9052 46256 9104
rect 52460 9052 52512 9104
rect 52736 9120 52788 9172
rect 37924 9027 37976 9036
rect 37924 8993 37933 9027
rect 37933 8993 37967 9027
rect 37967 8993 37976 9027
rect 37924 8984 37976 8993
rect 52276 8984 52328 9036
rect 36728 8959 36780 8968
rect 36728 8925 36737 8959
rect 36737 8925 36771 8959
rect 36771 8925 36780 8959
rect 36728 8916 36780 8925
rect 39120 8959 39172 8968
rect 27252 8891 27304 8900
rect 27252 8857 27270 8891
rect 27270 8857 27304 8891
rect 27252 8848 27304 8857
rect 24584 8823 24636 8832
rect 24584 8789 24593 8823
rect 24593 8789 24627 8823
rect 24627 8789 24636 8823
rect 24584 8780 24636 8789
rect 25964 8780 26016 8832
rect 26332 8780 26384 8832
rect 26424 8780 26476 8832
rect 31024 8848 31076 8900
rect 38660 8848 38712 8900
rect 39120 8925 39129 8959
rect 39129 8925 39163 8959
rect 39163 8925 39172 8959
rect 39120 8916 39172 8925
rect 42524 8916 42576 8968
rect 48964 8959 49016 8968
rect 40224 8848 40276 8900
rect 48964 8925 48973 8959
rect 48973 8925 49007 8959
rect 49007 8925 49016 8959
rect 51632 8959 51684 8968
rect 48964 8916 49016 8925
rect 50436 8891 50488 8900
rect 28632 8780 28684 8832
rect 28724 8780 28776 8832
rect 31852 8780 31904 8832
rect 32128 8780 32180 8832
rect 33508 8780 33560 8832
rect 33876 8823 33928 8832
rect 33876 8789 33885 8823
rect 33885 8789 33919 8823
rect 33919 8789 33928 8823
rect 33876 8780 33928 8789
rect 34428 8780 34480 8832
rect 34520 8780 34572 8832
rect 34980 8780 35032 8832
rect 36636 8780 36688 8832
rect 36728 8780 36780 8832
rect 48412 8780 48464 8832
rect 50436 8857 50445 8891
rect 50445 8857 50479 8891
rect 50479 8857 50488 8891
rect 50436 8848 50488 8857
rect 51632 8925 51641 8959
rect 51641 8925 51675 8959
rect 51675 8925 51684 8959
rect 51632 8916 51684 8925
rect 52460 8916 52512 8968
rect 52736 8959 52788 8968
rect 52736 8925 52745 8959
rect 52745 8925 52779 8959
rect 52779 8925 52788 8959
rect 52736 8916 52788 8925
rect 53196 8848 53248 8900
rect 49700 8780 49752 8832
rect 52736 8780 52788 8832
rect 53564 8823 53616 8832
rect 53564 8789 53573 8823
rect 53573 8789 53607 8823
rect 53607 8789 53616 8823
rect 53564 8780 53616 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 15476 8576 15528 8628
rect 17408 8576 17460 8628
rect 18880 8576 18932 8628
rect 14464 8508 14516 8560
rect 11060 8440 11112 8492
rect 14648 8440 14700 8492
rect 17132 8508 17184 8560
rect 19340 8508 19392 8560
rect 15108 8372 15160 8424
rect 1676 8347 1728 8356
rect 1676 8313 1685 8347
rect 1685 8313 1719 8347
rect 1719 8313 1728 8347
rect 1676 8304 1728 8313
rect 13636 8304 13688 8356
rect 15292 8304 15344 8356
rect 16672 8304 16724 8356
rect 17592 8304 17644 8356
rect 18512 8483 18564 8492
rect 18512 8449 18546 8483
rect 18546 8449 18564 8483
rect 18512 8440 18564 8449
rect 18788 8440 18840 8492
rect 23112 8576 23164 8628
rect 22284 8440 22336 8492
rect 22652 8440 22704 8492
rect 19340 8372 19392 8424
rect 19984 8372 20036 8424
rect 21272 8372 21324 8424
rect 25136 8576 25188 8628
rect 25688 8576 25740 8628
rect 23572 8483 23624 8492
rect 23572 8449 23606 8483
rect 23606 8449 23624 8483
rect 23572 8440 23624 8449
rect 27988 8576 28040 8628
rect 28448 8576 28500 8628
rect 32036 8576 32088 8628
rect 32496 8619 32548 8628
rect 32496 8585 32505 8619
rect 32505 8585 32539 8619
rect 32539 8585 32548 8619
rect 32496 8576 32548 8585
rect 26424 8508 26476 8560
rect 27620 8508 27672 8560
rect 29736 8508 29788 8560
rect 33692 8576 33744 8628
rect 34704 8576 34756 8628
rect 36820 8576 36872 8628
rect 38292 8576 38344 8628
rect 38660 8576 38712 8628
rect 50896 8576 50948 8628
rect 19616 8347 19668 8356
rect 19616 8313 19625 8347
rect 19625 8313 19659 8347
rect 19659 8313 19668 8347
rect 19616 8304 19668 8313
rect 19892 8304 19944 8356
rect 21364 8304 21416 8356
rect 21548 8304 21600 8356
rect 22008 8304 22060 8356
rect 25412 8372 25464 8424
rect 26424 8415 26476 8424
rect 26424 8381 26433 8415
rect 26433 8381 26467 8415
rect 26467 8381 26476 8415
rect 26424 8372 26476 8381
rect 29460 8440 29512 8492
rect 30104 8440 30156 8492
rect 31760 8440 31812 8492
rect 34428 8508 34480 8560
rect 35992 8508 36044 8560
rect 36636 8508 36688 8560
rect 54208 8619 54260 8628
rect 54208 8585 54217 8619
rect 54217 8585 54251 8619
rect 54251 8585 54260 8619
rect 54208 8576 54260 8585
rect 33508 8440 33560 8492
rect 35440 8483 35492 8492
rect 35440 8449 35449 8483
rect 35449 8449 35483 8483
rect 35483 8449 35492 8483
rect 35440 8440 35492 8449
rect 39120 8440 39172 8492
rect 52184 8483 52236 8492
rect 52184 8449 52193 8483
rect 52193 8449 52227 8483
rect 52227 8449 52236 8483
rect 52184 8440 52236 8449
rect 53472 8483 53524 8492
rect 53472 8449 53481 8483
rect 53481 8449 53515 8483
rect 53515 8449 53524 8483
rect 53472 8440 53524 8449
rect 24492 8304 24544 8356
rect 30380 8372 30432 8424
rect 31576 8415 31628 8424
rect 31024 8304 31076 8356
rect 31576 8381 31585 8415
rect 31585 8381 31619 8415
rect 31619 8381 31628 8415
rect 31576 8372 31628 8381
rect 31484 8304 31536 8356
rect 33232 8304 33284 8356
rect 37648 8372 37700 8424
rect 46204 8372 46256 8424
rect 34796 8347 34848 8356
rect 28632 8236 28684 8288
rect 30932 8236 30984 8288
rect 31208 8279 31260 8288
rect 31208 8245 31217 8279
rect 31217 8245 31251 8279
rect 31251 8245 31260 8279
rect 31208 8236 31260 8245
rect 34796 8313 34805 8347
rect 34805 8313 34839 8347
rect 34839 8313 34848 8347
rect 34796 8304 34848 8313
rect 37556 8347 37608 8356
rect 37556 8313 37565 8347
rect 37565 8313 37599 8347
rect 37599 8313 37608 8347
rect 37556 8304 37608 8313
rect 48320 8304 48372 8356
rect 53564 8304 53616 8356
rect 35624 8236 35676 8288
rect 35900 8279 35952 8288
rect 35900 8245 35909 8279
rect 35909 8245 35943 8279
rect 35943 8245 35952 8279
rect 35900 8236 35952 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 14648 8075 14700 8084
rect 12992 7896 13044 7948
rect 14648 8041 14657 8075
rect 14657 8041 14691 8075
rect 14691 8041 14700 8075
rect 14648 8032 14700 8041
rect 15200 8032 15252 8084
rect 17132 8032 17184 8084
rect 17500 8032 17552 8084
rect 18052 7964 18104 8016
rect 13728 7896 13780 7948
rect 19432 7896 19484 7948
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 19616 7828 19668 7880
rect 19984 7828 20036 7880
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 17132 7692 17184 7744
rect 19248 7760 19300 7812
rect 19432 7760 19484 7812
rect 23572 8032 23624 8084
rect 24676 8075 24728 8084
rect 24676 8041 24685 8075
rect 24685 8041 24719 8075
rect 24719 8041 24728 8075
rect 24676 8032 24728 8041
rect 23756 7964 23808 8016
rect 25228 8032 25280 8084
rect 31116 8075 31168 8084
rect 22652 7939 22704 7948
rect 22652 7905 22661 7939
rect 22661 7905 22695 7939
rect 22695 7905 22704 7939
rect 22652 7896 22704 7905
rect 25136 7896 25188 7948
rect 26424 7896 26476 7948
rect 22468 7828 22520 7880
rect 22560 7828 22612 7880
rect 23204 7828 23256 7880
rect 27620 7964 27672 8016
rect 31116 8041 31125 8075
rect 31125 8041 31159 8075
rect 31159 8041 31168 8075
rect 31116 8032 31168 8041
rect 32220 8075 32272 8084
rect 32220 8041 32229 8075
rect 32229 8041 32263 8075
rect 32263 8041 32272 8075
rect 32220 8032 32272 8041
rect 32312 8032 32364 8084
rect 33324 8075 33376 8084
rect 33324 8041 33333 8075
rect 33333 8041 33367 8075
rect 33367 8041 33376 8075
rect 33324 8032 33376 8041
rect 35532 8075 35584 8084
rect 35532 8041 35541 8075
rect 35541 8041 35575 8075
rect 35575 8041 35584 8075
rect 35532 8032 35584 8041
rect 35900 8032 35952 8084
rect 36636 8075 36688 8084
rect 36636 8041 36645 8075
rect 36645 8041 36679 8075
rect 36679 8041 36688 8075
rect 36636 8032 36688 8041
rect 52460 8075 52512 8084
rect 52460 8041 52469 8075
rect 52469 8041 52503 8075
rect 52503 8041 52512 8075
rect 52460 8032 52512 8041
rect 29092 7896 29144 7948
rect 29184 7939 29236 7948
rect 29184 7905 29193 7939
rect 29193 7905 29227 7939
rect 29227 7905 29236 7939
rect 29736 7939 29788 7948
rect 29184 7896 29236 7905
rect 29736 7905 29745 7939
rect 29745 7905 29779 7939
rect 29779 7905 29788 7939
rect 29736 7896 29788 7905
rect 28632 7828 28684 7880
rect 29000 7871 29052 7880
rect 29000 7837 29009 7871
rect 29009 7837 29043 7871
rect 29043 7837 29052 7871
rect 29000 7828 29052 7837
rect 31576 7828 31628 7880
rect 34520 7896 34572 7948
rect 24308 7760 24360 7812
rect 24768 7760 24820 7812
rect 18604 7692 18656 7744
rect 19340 7692 19392 7744
rect 21272 7735 21324 7744
rect 21272 7701 21281 7735
rect 21281 7701 21315 7735
rect 21315 7701 21324 7735
rect 21272 7692 21324 7701
rect 24860 7692 24912 7744
rect 28724 7760 28776 7812
rect 30380 7760 30432 7812
rect 33876 7828 33928 7880
rect 37464 7896 37516 7948
rect 52276 7871 52328 7880
rect 52276 7837 52285 7871
rect 52285 7837 52319 7871
rect 52319 7837 52328 7871
rect 52276 7828 52328 7837
rect 52920 7871 52972 7880
rect 52920 7837 52929 7871
rect 52929 7837 52963 7871
rect 52963 7837 52972 7871
rect 52920 7828 52972 7837
rect 52736 7760 52788 7812
rect 26424 7735 26476 7744
rect 26424 7701 26433 7735
rect 26433 7701 26467 7735
rect 26467 7701 26476 7735
rect 26424 7692 26476 7701
rect 26884 7735 26936 7744
rect 26884 7701 26893 7735
rect 26893 7701 26927 7735
rect 26927 7701 26936 7735
rect 26884 7692 26936 7701
rect 28356 7692 28408 7744
rect 30196 7692 30248 7744
rect 30564 7692 30616 7744
rect 34060 7692 34112 7744
rect 34244 7692 34296 7744
rect 39672 7692 39724 7744
rect 51080 7692 51132 7744
rect 54300 7735 54352 7744
rect 54300 7701 54309 7735
rect 54309 7701 54343 7735
rect 54343 7701 54352 7735
rect 54300 7692 54352 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 11060 7488 11112 7540
rect 13728 7531 13780 7540
rect 13728 7497 13737 7531
rect 13737 7497 13771 7531
rect 13771 7497 13780 7531
rect 13728 7488 13780 7497
rect 15752 7531 15804 7540
rect 15752 7497 15761 7531
rect 15761 7497 15795 7531
rect 15795 7497 15804 7531
rect 15752 7488 15804 7497
rect 17224 7531 17276 7540
rect 17224 7497 17233 7531
rect 17233 7497 17267 7531
rect 17267 7497 17276 7531
rect 17224 7488 17276 7497
rect 18604 7488 18656 7540
rect 22192 7488 22244 7540
rect 23204 7488 23256 7540
rect 27252 7488 27304 7540
rect 29000 7488 29052 7540
rect 30380 7531 30432 7540
rect 30380 7497 30389 7531
rect 30389 7497 30423 7531
rect 30423 7497 30432 7531
rect 30380 7488 30432 7497
rect 30932 7488 30984 7540
rect 33784 7488 33836 7540
rect 35900 7488 35952 7540
rect 48780 7488 48832 7540
rect 52920 7488 52972 7540
rect 53196 7531 53248 7540
rect 53196 7497 53205 7531
rect 53205 7497 53239 7531
rect 53239 7497 53248 7531
rect 53196 7488 53248 7497
rect 11060 7352 11112 7404
rect 12532 7352 12584 7404
rect 17132 7352 17184 7404
rect 17500 7352 17552 7404
rect 19984 7420 20036 7472
rect 18328 7352 18380 7404
rect 19064 7352 19116 7404
rect 1676 7191 1728 7200
rect 1676 7157 1685 7191
rect 1685 7157 1719 7191
rect 1719 7157 1728 7191
rect 1676 7148 1728 7157
rect 12992 7327 13044 7336
rect 12992 7293 13001 7327
rect 13001 7293 13035 7327
rect 13035 7293 13044 7327
rect 12992 7284 13044 7293
rect 13452 7284 13504 7336
rect 17960 7216 18012 7268
rect 21364 7352 21416 7404
rect 22284 7420 22336 7472
rect 22008 7352 22060 7404
rect 22284 7284 22336 7336
rect 24952 7352 25004 7404
rect 26884 7420 26936 7472
rect 30656 7420 30708 7472
rect 30748 7420 30800 7472
rect 49700 7420 49752 7472
rect 28356 7352 28408 7404
rect 28540 7395 28592 7404
rect 28540 7361 28549 7395
rect 28549 7361 28583 7395
rect 28583 7361 28592 7395
rect 28540 7352 28592 7361
rect 29184 7352 29236 7404
rect 29368 7352 29420 7404
rect 29092 7284 29144 7336
rect 19984 7148 20036 7200
rect 21640 7148 21692 7200
rect 23572 7148 23624 7200
rect 24768 7148 24820 7200
rect 27988 7216 28040 7268
rect 29460 7216 29512 7268
rect 31208 7352 31260 7404
rect 53380 7395 53432 7404
rect 53380 7361 53389 7395
rect 53389 7361 53423 7395
rect 53423 7361 53432 7395
rect 53380 7352 53432 7361
rect 54392 7352 54444 7404
rect 31024 7284 31076 7336
rect 30288 7216 30340 7268
rect 26424 7148 26476 7200
rect 30840 7148 30892 7200
rect 31576 7191 31628 7200
rect 31576 7157 31585 7191
rect 31585 7157 31619 7191
rect 31619 7157 31628 7191
rect 31576 7148 31628 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 18604 6944 18656 6996
rect 21364 6944 21416 6996
rect 22192 6944 22244 6996
rect 24952 6944 25004 6996
rect 33876 6987 33928 6996
rect 33876 6953 33885 6987
rect 33885 6953 33919 6987
rect 33919 6953 33928 6987
rect 33876 6944 33928 6953
rect 53380 6944 53432 6996
rect 54116 6987 54168 6996
rect 54116 6953 54125 6987
rect 54125 6953 54159 6987
rect 54159 6953 54168 6987
rect 54116 6944 54168 6953
rect 11060 6808 11112 6860
rect 29368 6876 29420 6928
rect 12992 6740 13044 6792
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 13084 6672 13136 6724
rect 1676 6647 1728 6656
rect 1676 6613 1685 6647
rect 1685 6613 1719 6647
rect 1719 6613 1728 6647
rect 1676 6604 1728 6613
rect 12072 6604 12124 6656
rect 17408 6808 17460 6860
rect 17500 6851 17552 6860
rect 17500 6817 17509 6851
rect 17509 6817 17543 6851
rect 17543 6817 17552 6851
rect 17500 6808 17552 6817
rect 18788 6740 18840 6792
rect 19432 6740 19484 6792
rect 22284 6808 22336 6860
rect 25136 6808 25188 6860
rect 26516 6851 26568 6860
rect 21640 6783 21692 6792
rect 17684 6604 17736 6656
rect 19984 6672 20036 6724
rect 21640 6749 21649 6783
rect 21649 6749 21683 6783
rect 21683 6749 21692 6783
rect 21640 6740 21692 6749
rect 25320 6740 25372 6792
rect 23572 6672 23624 6724
rect 23664 6672 23716 6724
rect 24676 6672 24728 6724
rect 19248 6604 19300 6656
rect 22192 6647 22244 6656
rect 22192 6613 22201 6647
rect 22201 6613 22235 6647
rect 22235 6613 22244 6647
rect 22192 6604 22244 6613
rect 22376 6604 22428 6656
rect 22836 6604 22888 6656
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 27344 6808 27396 6860
rect 27896 6808 27948 6860
rect 29552 6808 29604 6860
rect 30472 6808 30524 6860
rect 31392 6808 31444 6860
rect 33048 6851 33100 6860
rect 33048 6817 33057 6851
rect 33057 6817 33091 6851
rect 33091 6817 33100 6851
rect 33048 6808 33100 6817
rect 43720 6808 43772 6860
rect 51264 6808 51316 6860
rect 30380 6783 30432 6792
rect 30380 6749 30389 6783
rect 30389 6749 30423 6783
rect 30423 6749 30432 6783
rect 30380 6740 30432 6749
rect 31300 6740 31352 6792
rect 44916 6740 44968 6792
rect 49976 6740 50028 6792
rect 54300 6783 54352 6792
rect 54300 6749 54309 6783
rect 54309 6749 54343 6783
rect 54343 6749 54352 6783
rect 54300 6740 54352 6749
rect 27068 6672 27120 6724
rect 29368 6672 29420 6724
rect 30012 6672 30064 6724
rect 31576 6672 31628 6724
rect 29000 6604 29052 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 12532 6443 12584 6452
rect 12532 6409 12541 6443
rect 12541 6409 12575 6443
rect 12575 6409 12584 6443
rect 12532 6400 12584 6409
rect 12992 6443 13044 6452
rect 12992 6409 13001 6443
rect 13001 6409 13035 6443
rect 13035 6409 13044 6443
rect 12992 6400 13044 6409
rect 13084 6400 13136 6452
rect 8300 6332 8352 6384
rect 12440 6332 12492 6384
rect 13084 6264 13136 6316
rect 14188 6400 14240 6452
rect 17500 6400 17552 6452
rect 18512 6400 18564 6452
rect 19984 6400 20036 6452
rect 20168 6443 20220 6452
rect 20168 6409 20177 6443
rect 20177 6409 20211 6443
rect 20211 6409 20220 6443
rect 20168 6400 20220 6409
rect 20720 6443 20772 6452
rect 20720 6409 20729 6443
rect 20729 6409 20763 6443
rect 20763 6409 20772 6443
rect 20720 6400 20772 6409
rect 21456 6443 21508 6452
rect 21456 6409 21465 6443
rect 21465 6409 21499 6443
rect 21499 6409 21508 6443
rect 21456 6400 21508 6409
rect 23112 6400 23164 6452
rect 23664 6443 23716 6452
rect 23664 6409 23673 6443
rect 23673 6409 23707 6443
rect 23707 6409 23716 6443
rect 23664 6400 23716 6409
rect 25044 6400 25096 6452
rect 25320 6400 25372 6452
rect 25780 6443 25832 6452
rect 25780 6409 25789 6443
rect 25789 6409 25823 6443
rect 25823 6409 25832 6443
rect 25780 6400 25832 6409
rect 27068 6400 27120 6452
rect 29184 6400 29236 6452
rect 30472 6400 30524 6452
rect 31484 6443 31536 6452
rect 31484 6409 31493 6443
rect 31493 6409 31527 6443
rect 31527 6409 31536 6443
rect 31484 6400 31536 6409
rect 12072 6239 12124 6248
rect 12072 6205 12081 6239
rect 12081 6205 12115 6239
rect 12115 6205 12124 6239
rect 12072 6196 12124 6205
rect 10876 6128 10928 6180
rect 12992 6196 13044 6248
rect 31576 6332 31628 6384
rect 18972 6264 19024 6316
rect 19340 6307 19392 6316
rect 19340 6273 19349 6307
rect 19349 6273 19383 6307
rect 19383 6273 19392 6307
rect 19340 6264 19392 6273
rect 24584 6264 24636 6316
rect 27436 6264 27488 6316
rect 29736 6264 29788 6316
rect 30288 6264 30340 6316
rect 30564 6264 30616 6316
rect 12716 6128 12768 6180
rect 12808 6128 12860 6180
rect 24492 6196 24544 6248
rect 25136 6239 25188 6248
rect 25136 6205 25145 6239
rect 25145 6205 25179 6239
rect 25179 6205 25188 6239
rect 25136 6196 25188 6205
rect 33048 6400 33100 6452
rect 54392 6400 54444 6452
rect 22468 6128 22520 6180
rect 24676 6128 24728 6180
rect 44824 6128 44876 6180
rect 51540 6128 51592 6180
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 12440 6060 12492 6112
rect 17224 6060 17276 6112
rect 24216 6060 24268 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 12900 5856 12952 5908
rect 13084 5899 13136 5908
rect 13084 5865 13093 5899
rect 13093 5865 13127 5899
rect 13127 5865 13136 5899
rect 13084 5856 13136 5865
rect 11520 5831 11572 5840
rect 11520 5797 11529 5831
rect 11529 5797 11563 5831
rect 11563 5797 11572 5831
rect 11520 5788 11572 5797
rect 12532 5831 12584 5840
rect 12532 5797 12541 5831
rect 12541 5797 12575 5831
rect 12575 5797 12584 5831
rect 12532 5788 12584 5797
rect 12992 5788 13044 5840
rect 13452 5856 13504 5908
rect 13544 5788 13596 5840
rect 23204 5856 23256 5908
rect 24124 5856 24176 5908
rect 24676 5899 24728 5908
rect 24676 5865 24685 5899
rect 24685 5865 24719 5899
rect 24719 5865 24728 5899
rect 24676 5856 24728 5865
rect 26056 5856 26108 5908
rect 28724 5856 28776 5908
rect 30472 5856 30524 5908
rect 21456 5788 21508 5840
rect 12440 5652 12492 5704
rect 12624 5652 12676 5704
rect 13544 5695 13596 5704
rect 11704 5584 11756 5636
rect 12072 5584 12124 5636
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 11152 5516 11204 5568
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 17224 5652 17276 5704
rect 27160 5720 27212 5772
rect 23112 5652 23164 5704
rect 24308 5652 24360 5704
rect 26148 5652 26200 5704
rect 19248 5584 19300 5636
rect 29000 5652 29052 5704
rect 30472 5652 30524 5704
rect 26332 5584 26384 5636
rect 37464 5584 37516 5636
rect 25780 5516 25832 5568
rect 32772 5516 32824 5568
rect 34612 5516 34664 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 12440 5355 12492 5364
rect 12440 5321 12449 5355
rect 12449 5321 12483 5355
rect 12483 5321 12492 5355
rect 12440 5312 12492 5321
rect 16028 5312 16080 5364
rect 22836 5312 22888 5364
rect 25044 5312 25096 5364
rect 25872 5312 25924 5364
rect 25964 5312 26016 5364
rect 27620 5312 27672 5364
rect 28632 5312 28684 5364
rect 30012 5355 30064 5364
rect 30012 5321 30021 5355
rect 30021 5321 30055 5355
rect 30055 5321 30064 5355
rect 30012 5312 30064 5321
rect 30472 5312 30524 5364
rect 10508 5176 10560 5228
rect 12900 5219 12952 5228
rect 12900 5185 12910 5219
rect 12910 5185 12944 5219
rect 12944 5185 12952 5219
rect 14832 5244 14884 5296
rect 37556 5244 37608 5296
rect 38384 5244 38436 5296
rect 12900 5176 12952 5185
rect 14188 5176 14240 5228
rect 29184 5176 29236 5228
rect 7104 5108 7156 5160
rect 12440 5108 12492 5160
rect 13452 5151 13504 5160
rect 11796 5040 11848 5092
rect 1676 5015 1728 5024
rect 1676 4981 1685 5015
rect 1685 4981 1719 5015
rect 1719 4981 1728 5015
rect 1676 4972 1728 4981
rect 9588 4972 9640 5024
rect 9864 5015 9916 5024
rect 9864 4981 9873 5015
rect 9873 4981 9907 5015
rect 9907 4981 9916 5015
rect 9864 4972 9916 4981
rect 10692 4972 10744 5024
rect 12348 4972 12400 5024
rect 13452 5117 13461 5151
rect 13461 5117 13495 5151
rect 13495 5117 13504 5151
rect 13452 5108 13504 5117
rect 13820 5108 13872 5160
rect 25872 5108 25924 5160
rect 12992 5040 13044 5092
rect 13728 5083 13780 5092
rect 13728 5049 13737 5083
rect 13737 5049 13771 5083
rect 13771 5049 13780 5083
rect 13728 5040 13780 5049
rect 14740 5040 14792 5092
rect 18144 5040 18196 5092
rect 26884 5040 26936 5092
rect 16028 4972 16080 5024
rect 24952 5015 25004 5024
rect 24952 4981 24961 5015
rect 24961 4981 24995 5015
rect 24995 4981 25004 5015
rect 24952 4972 25004 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 10508 4811 10560 4820
rect 10508 4777 10517 4811
rect 10517 4777 10551 4811
rect 10551 4777 10560 4811
rect 10508 4768 10560 4777
rect 12808 4768 12860 4820
rect 12900 4768 12952 4820
rect 25780 4768 25832 4820
rect 28724 4768 28776 4820
rect 38384 4811 38436 4820
rect 38384 4777 38393 4811
rect 38393 4777 38427 4811
rect 38427 4777 38436 4811
rect 38384 4768 38436 4777
rect 41696 4768 41748 4820
rect 42432 4811 42484 4820
rect 42432 4777 42441 4811
rect 42441 4777 42475 4811
rect 42475 4777 42484 4811
rect 42432 4768 42484 4777
rect 42984 4811 43036 4820
rect 42984 4777 42993 4811
rect 42993 4777 43027 4811
rect 43027 4777 43036 4811
rect 42984 4768 43036 4777
rect 11244 4700 11296 4752
rect 13084 4743 13136 4752
rect 13084 4709 13093 4743
rect 13093 4709 13127 4743
rect 13127 4709 13136 4743
rect 13084 4700 13136 4709
rect 26884 4700 26936 4752
rect 46940 4700 46992 4752
rect 21272 4632 21324 4684
rect 23296 4632 23348 4684
rect 27436 4632 27488 4684
rect 10508 4564 10560 4616
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 10968 4607 11020 4616
rect 10968 4573 10977 4607
rect 10977 4573 11011 4607
rect 11011 4573 11020 4607
rect 10968 4564 11020 4573
rect 8668 4496 8720 4548
rect 12808 4564 12860 4616
rect 15200 4564 15252 4616
rect 45560 4607 45612 4616
rect 45560 4573 45569 4607
rect 45569 4573 45603 4607
rect 45603 4573 45612 4607
rect 45560 4564 45612 4573
rect 11704 4496 11756 4548
rect 13452 4539 13504 4548
rect 13452 4505 13461 4539
rect 13461 4505 13495 4539
rect 13495 4505 13504 4539
rect 13452 4496 13504 4505
rect 13912 4496 13964 4548
rect 22560 4496 22612 4548
rect 32404 4496 32456 4548
rect 1676 4471 1728 4480
rect 1676 4437 1685 4471
rect 1685 4437 1719 4471
rect 1719 4437 1728 4471
rect 1676 4428 1728 4437
rect 7748 4428 7800 4480
rect 10784 4428 10836 4480
rect 11612 4471 11664 4480
rect 11612 4437 11621 4471
rect 11621 4437 11655 4471
rect 11655 4437 11664 4471
rect 11612 4428 11664 4437
rect 12992 4428 13044 4480
rect 14556 4428 14608 4480
rect 23296 4471 23348 4480
rect 23296 4437 23305 4471
rect 23305 4437 23339 4471
rect 23339 4437 23348 4471
rect 23296 4428 23348 4437
rect 23664 4428 23716 4480
rect 25412 4428 25464 4480
rect 38660 4428 38712 4480
rect 43628 4471 43680 4480
rect 43628 4437 43637 4471
rect 43637 4437 43671 4471
rect 43671 4437 43680 4471
rect 43628 4428 43680 4437
rect 45928 4428 45980 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 10968 4224 11020 4276
rect 25320 4224 25372 4276
rect 10324 4156 10376 4208
rect 10416 4088 10468 4140
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 10508 4063 10560 4072
rect 10508 4029 10517 4063
rect 10517 4029 10551 4063
rect 10551 4029 10560 4063
rect 10508 4020 10560 4029
rect 12992 4156 13044 4208
rect 13728 4156 13780 4208
rect 10692 4063 10744 4072
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 10876 4063 10928 4072
rect 10876 4029 10885 4063
rect 10885 4029 10919 4063
rect 10919 4029 10928 4063
rect 10876 4020 10928 4029
rect 10968 4063 11020 4072
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 11704 4020 11756 4072
rect 12348 4088 12400 4140
rect 22100 4088 22152 4140
rect 26332 4156 26384 4208
rect 26240 4088 26292 4140
rect 26700 4088 26752 4140
rect 32404 4224 32456 4276
rect 35716 4224 35768 4276
rect 32772 4199 32824 4208
rect 32772 4165 32781 4199
rect 32781 4165 32815 4199
rect 32815 4165 32824 4199
rect 32772 4156 32824 4165
rect 32864 4156 32916 4208
rect 36176 4156 36228 4208
rect 36636 4156 36688 4208
rect 30380 4088 30432 4140
rect 30932 4088 30984 4140
rect 32496 4088 32548 4140
rect 9772 3952 9824 4004
rect 11060 3952 11112 4004
rect 13544 4020 13596 4072
rect 14648 4020 14700 4072
rect 23112 4020 23164 4072
rect 23940 4020 23992 4072
rect 25136 4020 25188 4072
rect 25504 4020 25556 4072
rect 25872 4020 25924 4072
rect 27988 4020 28040 4072
rect 40040 4088 40092 4140
rect 42708 4131 42760 4140
rect 42708 4097 42717 4131
rect 42717 4097 42751 4131
rect 42751 4097 42760 4131
rect 42708 4088 42760 4097
rect 45560 4088 45612 4140
rect 15108 3952 15160 4004
rect 37464 3995 37516 4004
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 6828 3927 6880 3936
rect 6828 3893 6837 3927
rect 6837 3893 6871 3927
rect 6871 3893 6880 3927
rect 6828 3884 6880 3893
rect 7656 3884 7708 3936
rect 8392 3884 8444 3936
rect 10048 3884 10100 3936
rect 10784 3884 10836 3936
rect 11428 3884 11480 3936
rect 12532 3884 12584 3936
rect 12900 3884 12952 3936
rect 13728 3884 13780 3936
rect 14096 3927 14148 3936
rect 14096 3893 14105 3927
rect 14105 3893 14139 3927
rect 14139 3893 14148 3927
rect 14096 3884 14148 3893
rect 14832 3884 14884 3936
rect 14924 3884 14976 3936
rect 37464 3961 37473 3995
rect 37473 3961 37507 3995
rect 37507 3961 37516 3995
rect 37464 3952 37516 3961
rect 38660 3952 38712 4004
rect 15384 3884 15436 3936
rect 17868 3884 17920 3936
rect 23480 3884 23532 3936
rect 23756 3927 23808 3936
rect 23756 3893 23765 3927
rect 23765 3893 23799 3927
rect 23799 3893 23808 3927
rect 23756 3884 23808 3893
rect 25044 3884 25096 3936
rect 27896 3884 27948 3936
rect 30932 3927 30984 3936
rect 30932 3893 30941 3927
rect 30941 3893 30975 3927
rect 30975 3893 30984 3927
rect 30932 3884 30984 3893
rect 32680 3884 32732 3936
rect 34152 3884 34204 3936
rect 38936 3884 38988 3936
rect 39304 3927 39356 3936
rect 39304 3893 39313 3927
rect 39313 3893 39347 3927
rect 39347 3893 39356 3927
rect 39304 3884 39356 3893
rect 43904 3952 43956 4004
rect 45744 3952 45796 4004
rect 41788 3927 41840 3936
rect 41788 3893 41797 3927
rect 41797 3893 41831 3927
rect 41831 3893 41840 3927
rect 41788 3884 41840 3893
rect 43076 3884 43128 3936
rect 44640 3884 44692 3936
rect 45652 3884 45704 3936
rect 46296 3884 46348 3936
rect 47768 3884 47820 3936
rect 49056 3927 49108 3936
rect 49056 3893 49065 3927
rect 49065 3893 49099 3927
rect 49099 3893 49108 3927
rect 49056 3884 49108 3893
rect 50160 3927 50212 3936
rect 50160 3893 50169 3927
rect 50169 3893 50203 3927
rect 50203 3893 50212 3927
rect 50160 3884 50212 3893
rect 50988 3927 51040 3936
rect 50988 3893 50997 3927
rect 50997 3893 51031 3927
rect 51031 3893 51040 3927
rect 50988 3884 51040 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 7104 3723 7156 3732
rect 7104 3689 7113 3723
rect 7113 3689 7147 3723
rect 7147 3689 7156 3723
rect 7104 3680 7156 3689
rect 8300 3680 8352 3732
rect 9588 3680 9640 3732
rect 10232 3680 10284 3732
rect 10416 3723 10468 3732
rect 10416 3689 10425 3723
rect 10425 3689 10459 3723
rect 10459 3689 10468 3723
rect 10416 3680 10468 3689
rect 12716 3680 12768 3732
rect 13360 3680 13412 3732
rect 15844 3680 15896 3732
rect 26792 3723 26844 3732
rect 8484 3612 8536 3664
rect 10324 3612 10376 3664
rect 10140 3544 10192 3596
rect 10876 3612 10928 3664
rect 13084 3612 13136 3664
rect 14464 3587 14516 3596
rect 14464 3553 14473 3587
rect 14473 3553 14507 3587
rect 14507 3553 14516 3587
rect 14464 3544 14516 3553
rect 14648 3587 14700 3596
rect 14648 3553 14657 3587
rect 14657 3553 14691 3587
rect 14691 3553 14700 3587
rect 14648 3544 14700 3553
rect 19064 3544 19116 3596
rect 26792 3689 26801 3723
rect 26801 3689 26835 3723
rect 26835 3689 26844 3723
rect 26792 3680 26844 3689
rect 27804 3680 27856 3732
rect 27896 3680 27948 3732
rect 28080 3680 28132 3732
rect 28632 3723 28684 3732
rect 28632 3689 28641 3723
rect 28641 3689 28675 3723
rect 28675 3689 28684 3723
rect 28632 3680 28684 3689
rect 31760 3680 31812 3732
rect 32404 3680 32456 3732
rect 32864 3680 32916 3732
rect 33324 3723 33376 3732
rect 33324 3689 33333 3723
rect 33333 3689 33367 3723
rect 33367 3689 33376 3723
rect 33324 3680 33376 3689
rect 33784 3680 33836 3732
rect 33968 3680 34020 3732
rect 34520 3680 34572 3732
rect 41696 3680 41748 3732
rect 42708 3680 42760 3732
rect 51172 3723 51224 3732
rect 23112 3612 23164 3664
rect 30288 3612 30340 3664
rect 30380 3612 30432 3664
rect 31668 3612 31720 3664
rect 31852 3655 31904 3664
rect 31852 3621 31861 3655
rect 31861 3621 31895 3655
rect 31895 3621 31904 3655
rect 31852 3612 31904 3621
rect 35348 3612 35400 3664
rect 41512 3612 41564 3664
rect 51172 3689 51181 3723
rect 51181 3689 51215 3723
rect 51215 3689 51224 3723
rect 51172 3680 51224 3689
rect 6828 3476 6880 3528
rect 7748 3519 7800 3528
rect 7748 3485 7757 3519
rect 7757 3485 7791 3519
rect 7791 3485 7800 3519
rect 7748 3476 7800 3485
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 7012 3340 7064 3392
rect 9588 3408 9640 3460
rect 8944 3340 8996 3392
rect 9680 3340 9732 3392
rect 9956 3383 10008 3392
rect 9956 3349 9965 3383
rect 9965 3349 9999 3383
rect 9999 3349 10008 3383
rect 9956 3340 10008 3349
rect 10692 3485 10724 3504
rect 10724 3485 10744 3504
rect 10692 3452 10744 3485
rect 10876 3519 10928 3528
rect 10876 3485 10886 3519
rect 10886 3485 10920 3519
rect 10920 3485 10928 3519
rect 11428 3519 11480 3528
rect 10876 3476 10928 3485
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 11612 3476 11664 3528
rect 12348 3476 12400 3528
rect 13452 3476 13504 3528
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 14556 3476 14608 3528
rect 14924 3519 14976 3528
rect 14924 3485 14933 3519
rect 14933 3485 14967 3519
rect 14967 3485 14976 3519
rect 14924 3476 14976 3485
rect 19984 3476 20036 3528
rect 22100 3451 22152 3460
rect 22100 3417 22109 3451
rect 22109 3417 22143 3451
rect 22143 3417 22152 3451
rect 22100 3408 22152 3417
rect 22744 3408 22796 3460
rect 14648 3340 14700 3392
rect 16120 3340 16172 3392
rect 16396 3383 16448 3392
rect 16396 3349 16405 3383
rect 16405 3349 16439 3383
rect 16439 3349 16448 3383
rect 16396 3340 16448 3349
rect 17776 3340 17828 3392
rect 18512 3340 18564 3392
rect 18604 3340 18656 3392
rect 24952 3476 25004 3528
rect 25320 3476 25372 3528
rect 23480 3408 23532 3460
rect 34060 3476 34112 3528
rect 37464 3476 37516 3528
rect 38936 3519 38988 3528
rect 38936 3485 38945 3519
rect 38945 3485 38979 3519
rect 38979 3485 38988 3519
rect 38936 3476 38988 3485
rect 40040 3519 40092 3528
rect 40040 3485 40049 3519
rect 40049 3485 40083 3519
rect 40083 3485 40092 3519
rect 40040 3476 40092 3485
rect 41696 3476 41748 3528
rect 41788 3476 41840 3528
rect 43076 3519 43128 3528
rect 26332 3408 26384 3460
rect 27712 3408 27764 3460
rect 29000 3408 29052 3460
rect 39304 3408 39356 3460
rect 43076 3485 43085 3519
rect 43085 3485 43119 3519
rect 43119 3485 43128 3519
rect 43076 3476 43128 3485
rect 45928 3519 45980 3528
rect 45928 3485 45937 3519
rect 45937 3485 45971 3519
rect 45971 3485 45980 3519
rect 45928 3476 45980 3485
rect 46940 3519 46992 3528
rect 46940 3485 46949 3519
rect 46949 3485 46983 3519
rect 46983 3485 46992 3519
rect 46940 3476 46992 3485
rect 50988 3408 51040 3460
rect 24860 3340 24912 3392
rect 35900 3340 35952 3392
rect 36268 3340 36320 3392
rect 37924 3340 37976 3392
rect 38108 3383 38160 3392
rect 38108 3349 38117 3383
rect 38117 3349 38151 3383
rect 38151 3349 38160 3383
rect 38108 3340 38160 3349
rect 40040 3340 40092 3392
rect 40776 3340 40828 3392
rect 42800 3340 42852 3392
rect 43628 3340 43680 3392
rect 44088 3340 44140 3392
rect 45192 3340 45244 3392
rect 45560 3340 45612 3392
rect 45836 3340 45888 3392
rect 46572 3340 46624 3392
rect 47676 3340 47728 3392
rect 48872 3383 48924 3392
rect 48872 3349 48881 3383
rect 48881 3349 48915 3383
rect 48915 3349 48924 3383
rect 48872 3340 48924 3349
rect 49424 3383 49476 3392
rect 49424 3349 49433 3383
rect 49433 3349 49467 3383
rect 49467 3349 49476 3383
rect 49424 3340 49476 3349
rect 49608 3340 49660 3392
rect 51816 3383 51868 3392
rect 51816 3349 51825 3383
rect 51825 3349 51859 3383
rect 51859 3349 51868 3383
rect 51816 3340 51868 3349
rect 52000 3340 52052 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 7656 3136 7708 3188
rect 8300 3136 8352 3188
rect 8484 3179 8536 3188
rect 8484 3145 8493 3179
rect 8493 3145 8527 3179
rect 8527 3145 8536 3179
rect 8484 3136 8536 3145
rect 8760 3136 8812 3188
rect 9404 3136 9456 3188
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 10968 3136 11020 3188
rect 12900 3136 12952 3188
rect 13636 3136 13688 3188
rect 14280 3136 14332 3188
rect 14924 3136 14976 3188
rect 15568 3179 15620 3188
rect 15568 3145 15577 3179
rect 15577 3145 15611 3179
rect 15611 3145 15620 3179
rect 15568 3136 15620 3145
rect 16580 3136 16632 3188
rect 16764 3136 16816 3188
rect 17592 3179 17644 3188
rect 17592 3145 17601 3179
rect 17601 3145 17635 3179
rect 17635 3145 17644 3179
rect 17592 3136 17644 3145
rect 17960 3136 18012 3188
rect 24400 3136 24452 3188
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 8392 3068 8444 3120
rect 9036 3068 9088 3120
rect 8760 3000 8812 3052
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 25412 3068 25464 3120
rect 28816 3136 28868 3188
rect 29644 3179 29696 3188
rect 29644 3145 29653 3179
rect 29653 3145 29687 3179
rect 29687 3145 29696 3179
rect 29644 3136 29696 3145
rect 29920 3136 29972 3188
rect 38936 3136 38988 3188
rect 40132 3136 40184 3188
rect 47860 3179 47912 3188
rect 34428 3068 34480 3120
rect 9864 3000 9916 3052
rect 10140 3000 10192 3052
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 11612 3000 11664 3052
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 10324 2932 10376 2984
rect 12900 3000 12952 3052
rect 13636 3000 13688 3052
rect 14096 3000 14148 3052
rect 14556 3000 14608 3052
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 16396 3000 16448 3052
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 17500 3000 17552 3052
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 18236 3000 18288 3052
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 23664 3043 23716 3052
rect 23664 3009 23673 3043
rect 23673 3009 23707 3043
rect 23707 3009 23716 3043
rect 23664 3000 23716 3009
rect 23756 3000 23808 3052
rect 12716 2932 12768 2984
rect 15200 2932 15252 2984
rect 12992 2864 13044 2916
rect 14648 2907 14700 2916
rect 14648 2873 14657 2907
rect 14657 2873 14691 2907
rect 14691 2873 14700 2907
rect 14648 2864 14700 2873
rect 24124 2932 24176 2984
rect 25044 3000 25096 3052
rect 26240 3000 26292 3052
rect 26792 3000 26844 3052
rect 27804 3043 27856 3052
rect 27804 3009 27813 3043
rect 27813 3009 27847 3043
rect 27847 3009 27856 3043
rect 27804 3000 27856 3009
rect 28816 3000 28868 3052
rect 30380 3043 30432 3052
rect 30380 3009 30389 3043
rect 30389 3009 30423 3043
rect 30423 3009 30432 3043
rect 30380 3000 30432 3009
rect 31760 3000 31812 3052
rect 32864 3000 32916 3052
rect 33324 3043 33376 3052
rect 33324 3009 33333 3043
rect 33333 3009 33367 3043
rect 33367 3009 33376 3043
rect 33324 3000 33376 3009
rect 35532 3000 35584 3052
rect 38108 3043 38160 3052
rect 38108 3009 38117 3043
rect 38117 3009 38151 3043
rect 38151 3009 38160 3043
rect 38108 3000 38160 3009
rect 38384 3000 38436 3052
rect 39304 3043 39356 3052
rect 39304 3009 39313 3043
rect 39313 3009 39347 3043
rect 39347 3009 39356 3043
rect 39304 3000 39356 3009
rect 47860 3145 47869 3179
rect 47869 3145 47903 3179
rect 47903 3145 47912 3179
rect 47860 3136 47912 3145
rect 48596 3179 48648 3188
rect 48596 3145 48605 3179
rect 48605 3145 48639 3179
rect 48639 3145 48648 3179
rect 48596 3136 48648 3145
rect 49332 3179 49384 3188
rect 49332 3145 49341 3179
rect 49341 3145 49375 3179
rect 49375 3145 49384 3179
rect 49332 3136 49384 3145
rect 50068 3179 50120 3188
rect 50068 3145 50077 3179
rect 50077 3145 50111 3179
rect 50111 3145 50120 3179
rect 50068 3136 50120 3145
rect 50804 3179 50856 3188
rect 50804 3145 50813 3179
rect 50813 3145 50847 3179
rect 50847 3145 50856 3179
rect 50804 3136 50856 3145
rect 51540 3179 51592 3188
rect 51540 3145 51549 3179
rect 51549 3145 51583 3179
rect 51583 3145 51592 3179
rect 51540 3136 51592 3145
rect 47676 3068 47728 3120
rect 50620 3068 50672 3120
rect 51816 3068 51868 3120
rect 41696 3000 41748 3052
rect 42432 3000 42484 3052
rect 43628 3043 43680 3052
rect 43628 3009 43637 3043
rect 43637 3009 43671 3043
rect 43671 3009 43680 3043
rect 43628 3000 43680 3009
rect 44088 3043 44140 3052
rect 44088 3009 44097 3043
rect 44097 3009 44131 3043
rect 44131 3009 44140 3043
rect 44088 3000 44140 3009
rect 44640 3000 44692 3052
rect 45560 3043 45612 3052
rect 45560 3009 45569 3043
rect 45569 3009 45603 3043
rect 45603 3009 45612 3043
rect 45560 3000 45612 3009
rect 46296 3043 46348 3052
rect 46296 3009 46305 3043
rect 46305 3009 46339 3043
rect 46339 3009 46348 3043
rect 46296 3000 46348 3009
rect 46940 3000 46992 3052
rect 48412 3000 48464 3052
rect 49424 3043 49476 3052
rect 49424 3009 49433 3043
rect 49433 3009 49467 3043
rect 49467 3009 49476 3043
rect 49424 3000 49476 3009
rect 32220 2932 32272 2984
rect 32956 2932 33008 2984
rect 31484 2864 31536 2916
rect 33692 2864 33744 2916
rect 35348 2932 35400 2984
rect 49148 2932 49200 2984
rect 49608 2932 49660 2984
rect 42524 2864 42576 2916
rect 18972 2796 19024 2848
rect 20076 2839 20128 2848
rect 20076 2805 20085 2839
rect 20085 2805 20119 2839
rect 20119 2805 20128 2839
rect 20076 2796 20128 2805
rect 20444 2796 20496 2848
rect 21548 2796 21600 2848
rect 22284 2839 22336 2848
rect 22284 2805 22293 2839
rect 22293 2805 22327 2839
rect 22327 2805 22336 2839
rect 22284 2796 22336 2805
rect 22652 2796 22704 2848
rect 23388 2796 23440 2848
rect 24124 2796 24176 2848
rect 25228 2796 25280 2848
rect 25964 2796 26016 2848
rect 26700 2796 26752 2848
rect 27436 2796 27488 2848
rect 28172 2796 28224 2848
rect 30012 2796 30064 2848
rect 30748 2796 30800 2848
rect 32220 2796 32272 2848
rect 37740 2796 37792 2848
rect 38476 2796 38528 2848
rect 38844 2796 38896 2848
rect 39580 2796 39632 2848
rect 40316 2796 40368 2848
rect 41052 2796 41104 2848
rect 41788 2796 41840 2848
rect 43260 2864 43312 2916
rect 43996 2864 44048 2916
rect 45468 2864 45520 2916
rect 49884 2864 49936 2916
rect 44732 2796 44784 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 11060 2592 11112 2644
rect 11520 2592 11572 2644
rect 12532 2592 12584 2644
rect 13084 2635 13136 2644
rect 13084 2601 13093 2635
rect 13093 2601 13127 2635
rect 13127 2601 13136 2635
rect 13084 2592 13136 2601
rect 14280 2592 14332 2644
rect 16212 2592 16264 2644
rect 17040 2592 17092 2644
rect 17408 2635 17460 2644
rect 17408 2601 17417 2635
rect 17417 2601 17451 2635
rect 17451 2601 17460 2635
rect 17408 2592 17460 2601
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 5448 2295 5500 2304
rect 5448 2261 5457 2295
rect 5457 2261 5491 2295
rect 5491 2261 5500 2295
rect 5448 2252 5500 2261
rect 6000 2295 6052 2304
rect 6000 2261 6009 2295
rect 6009 2261 6043 2295
rect 6043 2261 6052 2295
rect 6000 2252 6052 2261
rect 7564 2388 7616 2440
rect 10324 2524 10376 2576
rect 11244 2524 11296 2576
rect 15936 2524 15988 2576
rect 24308 2592 24360 2644
rect 30288 2592 30340 2644
rect 20812 2524 20864 2576
rect 28908 2524 28960 2576
rect 30380 2524 30432 2576
rect 31852 2524 31904 2576
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 10876 2388 10928 2440
rect 11612 2388 11664 2440
rect 12808 2388 12860 2440
rect 13912 2388 13964 2440
rect 14832 2431 14884 2440
rect 14832 2397 14841 2431
rect 14841 2397 14875 2431
rect 14875 2397 14884 2431
rect 14832 2388 14884 2397
rect 15384 2388 15436 2440
rect 8668 2252 8720 2304
rect 13268 2252 13320 2304
rect 14188 2320 14240 2372
rect 16028 2388 16080 2440
rect 16120 2431 16172 2440
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 16764 2388 16816 2440
rect 17868 2388 17920 2440
rect 22192 2456 22244 2508
rect 33416 2456 33468 2508
rect 18604 2388 18656 2440
rect 19340 2388 19392 2440
rect 21180 2388 21232 2440
rect 21916 2388 21968 2440
rect 22560 2431 22612 2440
rect 22560 2397 22569 2431
rect 22569 2397 22603 2431
rect 22603 2397 22612 2431
rect 22560 2388 22612 2397
rect 23296 2431 23348 2440
rect 23296 2397 23305 2431
rect 23305 2397 23339 2431
rect 23339 2397 23348 2431
rect 23296 2388 23348 2397
rect 23480 2388 23532 2440
rect 25044 2388 25096 2440
rect 25872 2388 25924 2440
rect 26332 2431 26384 2440
rect 26332 2397 26341 2431
rect 26341 2397 26375 2431
rect 26375 2397 26384 2431
rect 26332 2388 26384 2397
rect 27896 2388 27948 2440
rect 28540 2388 28592 2440
rect 29644 2388 29696 2440
rect 29920 2388 29972 2440
rect 30932 2388 30984 2440
rect 31760 2388 31812 2440
rect 32864 2388 32916 2440
rect 33784 2388 33836 2440
rect 34152 2388 34204 2440
rect 47584 2592 47636 2644
rect 37372 2524 37424 2576
rect 39948 2524 40000 2576
rect 41420 2524 41472 2576
rect 42892 2524 42944 2576
rect 44364 2524 44416 2576
rect 46204 2524 46256 2576
rect 48504 2567 48556 2576
rect 48504 2533 48513 2567
rect 48513 2533 48547 2567
rect 48547 2533 48556 2567
rect 48504 2524 48556 2533
rect 49976 2524 50028 2576
rect 51080 2567 51132 2576
rect 51080 2533 51089 2567
rect 51089 2533 51123 2567
rect 51123 2533 51132 2567
rect 51080 2524 51132 2533
rect 42800 2456 42852 2508
rect 37924 2388 37976 2440
rect 38752 2388 38804 2440
rect 40040 2431 40092 2440
rect 40040 2397 40049 2431
rect 40049 2397 40083 2431
rect 40083 2397 40092 2431
rect 40040 2388 40092 2397
rect 40776 2431 40828 2440
rect 40776 2397 40785 2431
rect 40785 2397 40819 2431
rect 40819 2397 40828 2431
rect 40776 2388 40828 2397
rect 41512 2431 41564 2440
rect 41512 2397 41521 2431
rect 41521 2397 41555 2431
rect 41555 2397 41564 2431
rect 41512 2388 41564 2397
rect 42984 2388 43036 2440
rect 45652 2456 45704 2508
rect 43904 2388 43956 2440
rect 45192 2431 45244 2440
rect 45192 2397 45201 2431
rect 45201 2397 45235 2431
rect 45235 2397 45244 2431
rect 45192 2388 45244 2397
rect 45744 2388 45796 2440
rect 47768 2431 47820 2440
rect 47768 2397 47777 2431
rect 47777 2397 47811 2431
rect 47811 2397 47820 2431
rect 47768 2388 47820 2397
rect 48044 2388 48096 2440
rect 49056 2388 49108 2440
rect 49700 2388 49752 2440
rect 34520 2320 34572 2372
rect 34796 2320 34848 2372
rect 45100 2320 45152 2372
rect 17132 2252 17184 2304
rect 23020 2252 23072 2304
rect 23756 2252 23808 2304
rect 24492 2252 24544 2304
rect 25596 2252 25648 2304
rect 26332 2252 26384 2304
rect 27068 2252 27120 2304
rect 27804 2252 27856 2304
rect 28540 2252 28592 2304
rect 29276 2252 29328 2304
rect 29644 2252 29696 2304
rect 31116 2252 31168 2304
rect 32588 2252 32640 2304
rect 37004 2252 37056 2304
rect 38108 2252 38160 2304
rect 39212 2252 39264 2304
rect 40684 2252 40736 2304
rect 42156 2252 42208 2304
rect 43628 2252 43680 2304
rect 47308 2320 47360 2372
rect 48872 2320 48924 2372
rect 48964 2320 49016 2372
rect 50160 2320 50212 2372
rect 51816 2363 51868 2372
rect 51816 2329 51825 2363
rect 51825 2329 51859 2363
rect 51859 2329 51868 2363
rect 51816 2320 51868 2329
rect 52000 2363 52052 2372
rect 52000 2329 52009 2363
rect 52009 2329 52043 2363
rect 52043 2329 52052 2363
rect 52000 2320 52052 2329
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 5448 2048 5500 2100
rect 9680 2048 9732 2100
rect 10876 2048 10928 2100
rect 13912 2048 13964 2100
rect 14924 2048 14976 2100
rect 50252 2048 50304 2100
rect 52000 2048 52052 2100
rect 6000 1980 6052 2032
rect 11612 1980 11664 2032
<< metal2 >>
rect 1674 55200 1730 56000
rect 2870 55298 2926 56000
rect 2870 55270 3188 55298
rect 2870 55200 2926 55270
rect 1688 53038 1716 55200
rect 3160 53174 3188 55270
rect 4066 55200 4122 56000
rect 5262 55298 5318 56000
rect 6458 55298 6514 56000
rect 7654 55298 7710 56000
rect 8850 55298 8906 56000
rect 5262 55270 5488 55298
rect 5262 55200 5318 55270
rect 3148 53168 3200 53174
rect 3148 53110 3200 53116
rect 1676 53032 1728 53038
rect 1676 52974 1728 52980
rect 2596 53032 2648 53038
rect 2596 52974 2648 52980
rect 1768 52488 1820 52494
rect 1768 52430 1820 52436
rect 2504 52488 2556 52494
rect 2504 52430 2556 52436
rect 1492 52352 1544 52358
rect 1492 52294 1544 52300
rect 1504 52193 1532 52294
rect 1490 52184 1546 52193
rect 1490 52119 1546 52128
rect 1676 52012 1728 52018
rect 1676 51954 1728 51960
rect 1688 51649 1716 51954
rect 1674 51640 1730 51649
rect 1674 51575 1730 51584
rect 1676 51332 1728 51338
rect 1676 51274 1728 51280
rect 1688 51105 1716 51274
rect 1674 51096 1730 51105
rect 1674 51031 1730 51040
rect 1676 49836 1728 49842
rect 1676 49778 1728 49784
rect 1688 49473 1716 49778
rect 1674 49464 1730 49473
rect 1674 49399 1730 49408
rect 1780 43178 1808 52430
rect 1860 51876 1912 51882
rect 1860 51818 1912 51824
rect 1872 43382 1900 51818
rect 2320 50856 2372 50862
rect 2320 50798 2372 50804
rect 2136 50312 2188 50318
rect 2136 50254 2188 50260
rect 2044 49768 2096 49774
rect 2044 49710 2096 49716
rect 1860 43376 1912 43382
rect 1860 43318 1912 43324
rect 1768 43172 1820 43178
rect 1768 43114 1820 43120
rect 2056 41177 2084 49710
rect 2148 48550 2176 50254
rect 2332 49314 2360 50798
rect 2332 49286 2452 49314
rect 2320 49224 2372 49230
rect 2320 49166 2372 49172
rect 2228 48680 2280 48686
rect 2228 48622 2280 48628
rect 2136 48544 2188 48550
rect 2136 48486 2188 48492
rect 2240 46442 2268 48622
rect 2332 47530 2360 49166
rect 2320 47524 2372 47530
rect 2320 47466 2372 47472
rect 2228 46436 2280 46442
rect 2228 46378 2280 46384
rect 2424 46102 2452 49286
rect 2412 46096 2464 46102
rect 2412 46038 2464 46044
rect 2320 45960 2372 45966
rect 2320 45902 2372 45908
rect 2228 44328 2280 44334
rect 2228 44270 2280 44276
rect 2136 43784 2188 43790
rect 2136 43726 2188 43732
rect 2042 41168 2098 41177
rect 2042 41103 2098 41112
rect 2148 40610 2176 43726
rect 2056 40582 2176 40610
rect 1676 38276 1728 38282
rect 1676 38218 1728 38224
rect 1688 38049 1716 38218
rect 1674 38040 1730 38049
rect 1674 37975 1730 37984
rect 1584 37868 1636 37874
rect 1584 37810 1636 37816
rect 1596 37505 1624 37810
rect 1582 37496 1638 37505
rect 1582 37431 1638 37440
rect 2056 36106 2084 40582
rect 2136 40520 2188 40526
rect 2136 40462 2188 40468
rect 2148 37942 2176 40462
rect 2136 37936 2188 37942
rect 2136 37878 2188 37884
rect 2240 36689 2268 44270
rect 2332 43858 2360 45902
rect 2516 44305 2544 52430
rect 2608 52086 2636 52974
rect 2778 52728 2834 52737
rect 3160 52698 3188 53110
rect 4080 53106 4108 55200
rect 5460 53174 5488 55270
rect 6458 55270 6684 55298
rect 6458 55200 6514 55270
rect 6656 53174 6684 55270
rect 7654 55270 7788 55298
rect 7654 55200 7710 55270
rect 5448 53168 5500 53174
rect 5448 53110 5500 53116
rect 6644 53168 6696 53174
rect 6644 53110 6696 53116
rect 4068 53100 4120 53106
rect 4068 53042 4120 53048
rect 3240 52896 3292 52902
rect 3240 52838 3292 52844
rect 2778 52663 2834 52672
rect 3148 52692 3200 52698
rect 2792 52426 2820 52663
rect 3148 52634 3200 52640
rect 2780 52420 2832 52426
rect 2780 52362 2832 52368
rect 2792 52154 2820 52362
rect 2872 52352 2924 52358
rect 2872 52294 2924 52300
rect 2780 52148 2832 52154
rect 2780 52090 2832 52096
rect 2596 52080 2648 52086
rect 2596 52022 2648 52028
rect 2884 51610 2912 52294
rect 2872 51604 2924 51610
rect 2872 51546 2924 51552
rect 2688 51264 2740 51270
rect 2688 51206 2740 51212
rect 2700 48006 2728 51206
rect 2780 50856 2832 50862
rect 2780 50798 2832 50804
rect 2792 50561 2820 50798
rect 2778 50552 2834 50561
rect 2778 50487 2834 50496
rect 2780 50312 2832 50318
rect 2780 50254 2832 50260
rect 2792 50017 2820 50254
rect 2778 50008 2834 50017
rect 2778 49943 2834 49952
rect 2780 49224 2832 49230
rect 2780 49166 2832 49172
rect 2792 48929 2820 49166
rect 2778 48920 2834 48929
rect 2778 48855 2834 48864
rect 2780 48680 2832 48686
rect 2780 48622 2832 48628
rect 2792 48385 2820 48622
rect 2778 48376 2834 48385
rect 2778 48311 2834 48320
rect 2780 48136 2832 48142
rect 2780 48078 2832 48084
rect 2688 48000 2740 48006
rect 2688 47942 2740 47948
rect 2792 47841 2820 48078
rect 2778 47832 2834 47841
rect 2778 47767 2834 47776
rect 2780 47592 2832 47598
rect 2780 47534 2832 47540
rect 2792 47297 2820 47534
rect 2778 47288 2834 47297
rect 2778 47223 2834 47232
rect 2688 47116 2740 47122
rect 2688 47058 2740 47064
rect 2596 46572 2648 46578
rect 2596 46514 2648 46520
rect 2502 44296 2558 44305
rect 2502 44231 2558 44240
rect 2320 43852 2372 43858
rect 2320 43794 2372 43800
rect 2504 43308 2556 43314
rect 2504 43250 2556 43256
rect 2320 42152 2372 42158
rect 2320 42094 2372 42100
rect 2332 37466 2360 42094
rect 2320 37460 2372 37466
rect 2320 37402 2372 37408
rect 2226 36680 2282 36689
rect 2226 36615 2282 36624
rect 2044 36100 2096 36106
rect 2044 36042 2096 36048
rect 2516 35494 2544 43250
rect 2608 42770 2636 46514
rect 2700 43314 2728 47058
rect 2780 47048 2832 47054
rect 2780 46990 2832 46996
rect 2792 46753 2820 46990
rect 2778 46744 2834 46753
rect 2778 46679 2834 46688
rect 2780 46504 2832 46510
rect 2780 46446 2832 46452
rect 2792 46209 2820 46446
rect 2778 46200 2834 46209
rect 2778 46135 2834 46144
rect 2780 45960 2832 45966
rect 2780 45902 2832 45908
rect 2792 45665 2820 45902
rect 2778 45656 2834 45665
rect 2778 45591 2834 45600
rect 2780 45416 2832 45422
rect 2780 45358 2832 45364
rect 2792 45121 2820 45358
rect 2778 45112 2834 45121
rect 2778 45047 2834 45056
rect 2780 44872 2832 44878
rect 2780 44814 2832 44820
rect 2792 44577 2820 44814
rect 2778 44568 2834 44577
rect 2778 44503 2834 44512
rect 2780 44328 2832 44334
rect 2780 44270 2832 44276
rect 2792 44033 2820 44270
rect 2778 44024 2834 44033
rect 2778 43959 2834 43968
rect 2780 43784 2832 43790
rect 2780 43726 2832 43732
rect 2792 43489 2820 43726
rect 2778 43480 2834 43489
rect 2778 43415 2834 43424
rect 2688 43308 2740 43314
rect 2688 43250 2740 43256
rect 2780 43240 2832 43246
rect 2780 43182 2832 43188
rect 2792 42945 2820 43182
rect 2778 42936 2834 42945
rect 2778 42871 2834 42880
rect 2596 42764 2648 42770
rect 2596 42706 2648 42712
rect 2780 42696 2832 42702
rect 2780 42638 2832 42644
rect 2792 42401 2820 42638
rect 2778 42392 2834 42401
rect 2778 42327 2834 42336
rect 2780 42152 2832 42158
rect 2780 42094 2832 42100
rect 2792 41857 2820 42094
rect 2778 41848 2834 41857
rect 2778 41783 2834 41792
rect 2780 41608 2832 41614
rect 2780 41550 2832 41556
rect 2792 41313 2820 41550
rect 2778 41304 2834 41313
rect 2778 41239 2834 41248
rect 2780 41064 2832 41070
rect 2780 41006 2832 41012
rect 2792 40769 2820 41006
rect 2778 40760 2834 40769
rect 2778 40695 2834 40704
rect 2780 40520 2832 40526
rect 2780 40462 2832 40468
rect 2792 40225 2820 40462
rect 2778 40216 2834 40225
rect 2778 40151 2834 40160
rect 2780 39976 2832 39982
rect 2780 39918 2832 39924
rect 2792 39681 2820 39918
rect 2778 39672 2834 39681
rect 2778 39607 2834 39616
rect 2780 39432 2832 39438
rect 2780 39374 2832 39380
rect 2792 39137 2820 39374
rect 2778 39128 2834 39137
rect 2778 39063 2834 39072
rect 2780 38888 2832 38894
rect 2780 38830 2832 38836
rect 2792 38593 2820 38830
rect 2778 38584 2834 38593
rect 2778 38519 2834 38528
rect 2780 37664 2832 37670
rect 2780 37606 2832 37612
rect 2792 37330 2820 37606
rect 2780 37324 2832 37330
rect 2780 37266 2832 37272
rect 2792 36961 2820 37266
rect 2778 36952 2834 36961
rect 2778 36887 2834 36896
rect 2780 36712 2832 36718
rect 2780 36654 2832 36660
rect 2792 36417 2820 36654
rect 2778 36408 2834 36417
rect 2778 36343 2834 36352
rect 2780 36168 2832 36174
rect 2780 36110 2832 36116
rect 2792 35873 2820 36110
rect 2778 35864 2834 35873
rect 2778 35799 2834 35808
rect 2780 35624 2832 35630
rect 2780 35566 2832 35572
rect 2504 35488 2556 35494
rect 2504 35430 2556 35436
rect 2792 35329 2820 35566
rect 2778 35320 2834 35329
rect 2778 35255 2834 35264
rect 1584 35080 1636 35086
rect 3252 35057 3280 52838
rect 4080 52698 4108 53042
rect 5540 52896 5592 52902
rect 5540 52838 5592 52844
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4068 52692 4120 52698
rect 4068 52634 4120 52640
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 5552 38282 5580 52838
rect 6656 52698 6684 53110
rect 7760 53106 7788 55270
rect 8588 55270 8906 55298
rect 8588 53242 8616 55270
rect 8850 55200 8906 55270
rect 10046 55298 10102 56000
rect 11242 55298 11298 56000
rect 12438 55298 12494 56000
rect 10046 55270 10180 55298
rect 10046 55200 10102 55270
rect 8576 53236 8628 53242
rect 8576 53178 8628 53184
rect 9312 53236 9364 53242
rect 9312 53178 9364 53184
rect 7748 53100 7800 53106
rect 7748 53042 7800 53048
rect 6736 52896 6788 52902
rect 6736 52838 6788 52844
rect 6644 52692 6696 52698
rect 6644 52634 6696 52640
rect 5540 38276 5592 38282
rect 5540 38218 5592 38224
rect 4344 38208 4396 38214
rect 4344 38150 4396 38156
rect 4356 37806 4384 38150
rect 4344 37800 4396 37806
rect 4344 37742 4396 37748
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 1584 35022 1636 35028
rect 3238 35048 3294 35057
rect 1596 34785 1624 35022
rect 3238 34983 3294 34992
rect 1768 34944 1820 34950
rect 1768 34886 1820 34892
rect 2780 34944 2832 34950
rect 2780 34886 2832 34892
rect 1582 34776 1638 34785
rect 1780 34746 1808 34886
rect 1582 34711 1638 34720
rect 1768 34740 1820 34746
rect 1768 34682 1820 34688
rect 2792 34542 2820 34886
rect 2780 34536 2832 34542
rect 2780 34478 2832 34484
rect 2792 34241 2820 34478
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 2778 34232 2834 34241
rect 4214 34235 4522 34244
rect 2778 34167 2834 34176
rect 2780 33992 2832 33998
rect 2780 33934 2832 33940
rect 2792 33697 2820 33934
rect 2778 33688 2834 33697
rect 2778 33623 2834 33632
rect 6748 33522 6776 52838
rect 7760 52698 7788 53042
rect 8208 53032 8260 53038
rect 8208 52974 8260 52980
rect 7748 52692 7800 52698
rect 7748 52634 7800 52640
rect 8220 50386 8248 52974
rect 9324 51950 9352 53178
rect 10152 53106 10180 55270
rect 11242 55270 11376 55298
rect 11242 55200 11298 55270
rect 10140 53100 10192 53106
rect 10140 53042 10192 53048
rect 10152 52698 10180 53042
rect 10416 53032 10468 53038
rect 10416 52974 10468 52980
rect 10140 52692 10192 52698
rect 10140 52634 10192 52640
rect 9312 51944 9364 51950
rect 9312 51886 9364 51892
rect 8208 50380 8260 50386
rect 8208 50322 8260 50328
rect 10428 44334 10456 52974
rect 11348 52562 11376 55270
rect 12438 55270 12572 55298
rect 12438 55200 12494 55270
rect 12544 53106 12572 55270
rect 13634 55200 13690 56000
rect 14830 55200 14886 56000
rect 16026 55298 16082 56000
rect 17222 55298 17278 56000
rect 16026 55270 16344 55298
rect 16026 55200 16082 55270
rect 12532 53100 12584 53106
rect 12532 53042 12584 53048
rect 12808 53032 12860 53038
rect 12808 52974 12860 52980
rect 11704 52896 11756 52902
rect 11704 52838 11756 52844
rect 11336 52556 11388 52562
rect 11336 52498 11388 52504
rect 11612 52488 11664 52494
rect 11612 52430 11664 52436
rect 10416 44328 10468 44334
rect 10416 44270 10468 44276
rect 11624 43217 11652 52430
rect 11610 43208 11666 43217
rect 11610 43143 11666 43152
rect 11716 39098 11744 52838
rect 12820 43926 12848 52974
rect 13648 52698 13676 55200
rect 14844 53106 14872 55200
rect 16316 53106 16344 55270
rect 17222 55270 17356 55298
rect 17222 55200 17278 55270
rect 14832 53100 14884 53106
rect 14832 53042 14884 53048
rect 16304 53100 16356 53106
rect 16304 53042 16356 53048
rect 14844 52698 14872 53042
rect 16028 53032 16080 53038
rect 16028 52974 16080 52980
rect 15016 52896 15068 52902
rect 15016 52838 15068 52844
rect 13636 52692 13688 52698
rect 13636 52634 13688 52640
rect 14832 52692 14884 52698
rect 14832 52634 14884 52640
rect 13648 52494 13676 52634
rect 13636 52488 13688 52494
rect 13636 52430 13688 52436
rect 14280 52352 14332 52358
rect 14280 52294 14332 52300
rect 12808 43920 12860 43926
rect 12808 43862 12860 43868
rect 11704 39092 11756 39098
rect 11704 39034 11756 39040
rect 13452 36576 13504 36582
rect 13452 36518 13504 36524
rect 13464 36310 13492 36518
rect 13452 36304 13504 36310
rect 13452 36246 13504 36252
rect 14292 34610 14320 52294
rect 14832 38888 14884 38894
rect 14832 38830 14884 38836
rect 14844 37738 14872 38830
rect 14832 37732 14884 37738
rect 14832 37674 14884 37680
rect 15028 35222 15056 52838
rect 16040 50454 16068 52974
rect 17328 52562 17356 55270
rect 18418 55200 18474 56000
rect 19614 55298 19670 56000
rect 19444 55270 19670 55298
rect 18432 53106 18460 55200
rect 19444 53106 19472 55270
rect 19614 55200 19670 55270
rect 20810 55298 20866 56000
rect 20810 55270 20944 55298
rect 20810 55200 20866 55270
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 20916 53106 20944 55270
rect 22006 55200 22062 56000
rect 23202 55298 23258 56000
rect 24398 55298 24454 56000
rect 25594 55298 25650 56000
rect 26790 55298 26846 56000
rect 23202 55270 23336 55298
rect 23202 55200 23258 55270
rect 22020 53106 22048 55200
rect 23308 53106 23336 55270
rect 24398 55270 24624 55298
rect 24398 55200 24454 55270
rect 24492 53168 24544 53174
rect 24492 53110 24544 53116
rect 18420 53100 18472 53106
rect 18420 53042 18472 53048
rect 18788 53100 18840 53106
rect 18788 53042 18840 53048
rect 19432 53100 19484 53106
rect 19432 53042 19484 53048
rect 20904 53100 20956 53106
rect 20904 53042 20956 53048
rect 22008 53100 22060 53106
rect 22008 53042 22060 53048
rect 23296 53100 23348 53106
rect 23296 53042 23348 53048
rect 18800 52698 18828 53042
rect 19444 52698 19472 53042
rect 21456 53032 21508 53038
rect 21456 52974 21508 52980
rect 18788 52692 18840 52698
rect 18788 52634 18840 52640
rect 19432 52692 19484 52698
rect 19432 52634 19484 52640
rect 17316 52556 17368 52562
rect 17316 52498 17368 52504
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 16028 50448 16080 50454
rect 16028 50390 16080 50396
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19340 39976 19392 39982
rect 19340 39918 19392 39924
rect 17224 39840 17276 39846
rect 17224 39782 17276 39788
rect 17236 36786 17264 39782
rect 17316 38956 17368 38962
rect 17316 38898 17368 38904
rect 17328 38214 17356 38898
rect 17316 38208 17368 38214
rect 17316 38150 17368 38156
rect 17224 36780 17276 36786
rect 17224 36722 17276 36728
rect 17328 36310 17356 38150
rect 17316 36304 17368 36310
rect 17316 36246 17368 36252
rect 15108 36032 15160 36038
rect 15108 35974 15160 35980
rect 15120 35698 15148 35974
rect 15108 35692 15160 35698
rect 15108 35634 15160 35640
rect 15108 35284 15160 35290
rect 15108 35226 15160 35232
rect 16672 35284 16724 35290
rect 16672 35226 16724 35232
rect 15016 35216 15068 35222
rect 15016 35158 15068 35164
rect 14556 35148 14608 35154
rect 14556 35090 14608 35096
rect 14568 34950 14596 35090
rect 15120 35034 15148 35226
rect 15028 35018 15148 35034
rect 15660 35080 15712 35086
rect 15660 35022 15712 35028
rect 15016 35012 15148 35018
rect 15068 35006 15148 35012
rect 15016 34954 15068 34960
rect 14556 34944 14608 34950
rect 14556 34886 14608 34892
rect 14280 34604 14332 34610
rect 14280 34546 14332 34552
rect 13452 34536 13504 34542
rect 13452 34478 13504 34484
rect 6736 33516 6788 33522
rect 6736 33458 6788 33464
rect 2780 33448 2832 33454
rect 2780 33390 2832 33396
rect 2792 33153 2820 33390
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 2778 33144 2834 33153
rect 4214 33147 4522 33156
rect 2778 33079 2834 33088
rect 1584 32904 1636 32910
rect 1584 32846 1636 32852
rect 1596 32609 1624 32846
rect 2780 32768 2832 32774
rect 2780 32710 2832 32716
rect 1582 32600 1638 32609
rect 1582 32535 1638 32544
rect 2792 32366 2820 32710
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2792 32065 2820 32302
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 2778 32056 2834 32065
rect 4214 32059 4522 32068
rect 2778 31991 2834 32000
rect 2136 31816 2188 31822
rect 2136 31758 2188 31764
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 2148 30394 2176 31758
rect 2792 31521 2820 31758
rect 2778 31512 2834 31521
rect 2778 31447 2834 31456
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2792 30977 2820 31214
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 2778 30968 2834 30977
rect 4214 30971 4522 30980
rect 2778 30903 2834 30912
rect 2780 30728 2832 30734
rect 2780 30670 2832 30676
rect 2792 30433 2820 30670
rect 2778 30424 2834 30433
rect 2136 30388 2188 30394
rect 2778 30359 2834 30368
rect 2136 30330 2188 30336
rect 2228 30184 2280 30190
rect 2228 30126 2280 30132
rect 2240 29889 2268 30126
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 2226 29880 2282 29889
rect 4214 29883 4522 29892
rect 2226 29815 2228 29824
rect 2280 29815 2282 29824
rect 2228 29786 2280 29792
rect 1584 29640 1636 29646
rect 1584 29582 1636 29588
rect 4528 29640 4580 29646
rect 4528 29582 4580 29588
rect 1596 29345 1624 29582
rect 1582 29336 1638 29345
rect 1582 29271 1638 29280
rect 4540 29170 4568 29582
rect 11060 29232 11112 29238
rect 11060 29174 11112 29180
rect 4528 29164 4580 29170
rect 4528 29106 4580 29112
rect 2780 29096 2832 29102
rect 2780 29038 2832 29044
rect 2792 28801 2820 29038
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 2778 28792 2834 28801
rect 4214 28795 4522 28804
rect 2778 28727 2834 28736
rect 2780 28552 2832 28558
rect 2780 28494 2832 28500
rect 2792 28257 2820 28494
rect 2778 28248 2834 28257
rect 2778 28183 2834 28192
rect 2688 28076 2740 28082
rect 2688 28018 2740 28024
rect 2228 28008 2280 28014
rect 2228 27950 2280 27956
rect 2240 27713 2268 27950
rect 2226 27704 2282 27713
rect 2226 27639 2228 27648
rect 2280 27639 2282 27648
rect 2228 27610 2280 27616
rect 1584 27464 1636 27470
rect 1584 27406 1636 27412
rect 1596 27169 1624 27406
rect 1582 27160 1638 27169
rect 1582 27095 1638 27104
rect 2700 26518 2728 28018
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 11072 27402 11100 29174
rect 13360 29096 13412 29102
rect 13360 29038 13412 29044
rect 11060 27396 11112 27402
rect 11060 27338 11112 27344
rect 2780 26920 2832 26926
rect 2780 26862 2832 26868
rect 2792 26625 2820 26862
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 2778 26616 2834 26625
rect 4214 26619 4522 26628
rect 2778 26551 2834 26560
rect 2688 26512 2740 26518
rect 2688 26454 2740 26460
rect 2228 26376 2280 26382
rect 2228 26318 2280 26324
rect 2240 26081 2268 26318
rect 2226 26072 2282 26081
rect 2226 26007 2228 26016
rect 2280 26007 2282 26016
rect 2228 25978 2280 25984
rect 2240 25947 2268 25978
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 1596 25537 1624 25842
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 1582 25528 1638 25537
rect 4214 25531 4522 25540
rect 1582 25463 1584 25472
rect 1636 25463 1638 25472
rect 1584 25434 1636 25440
rect 1596 25403 1624 25434
rect 1584 25288 1636 25294
rect 1584 25230 1636 25236
rect 1596 24993 1624 25230
rect 1582 24984 1638 24993
rect 1582 24919 1638 24928
rect 1676 24812 1728 24818
rect 1676 24754 1728 24760
rect 1688 24449 1716 24754
rect 4068 24608 4120 24614
rect 4068 24550 4120 24556
rect 1674 24440 1730 24449
rect 1674 24375 1730 24384
rect 1676 24132 1728 24138
rect 1676 24074 1728 24080
rect 1688 23905 1716 24074
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1674 23896 1730 23905
rect 1674 23831 1730 23840
rect 1780 23798 1808 24006
rect 4080 23866 4108 24550
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 1768 23792 1820 23798
rect 1768 23734 1820 23740
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1688 23361 1716 23462
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 1674 23352 1730 23361
rect 4214 23355 4522 23364
rect 1674 23287 1730 23296
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1688 22817 1716 22918
rect 1674 22808 1730 22817
rect 2332 22778 2360 23054
rect 1674 22743 1730 22752
rect 2320 22772 2372 22778
rect 2320 22714 2372 22720
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 1676 22432 1728 22438
rect 1676 22374 1728 22380
rect 1688 22273 1716 22374
rect 1674 22264 1730 22273
rect 1674 22199 1730 22208
rect 1872 22166 1900 22578
rect 2596 22568 2648 22574
rect 2596 22510 2648 22516
rect 1860 22160 1912 22166
rect 1860 22102 1912 22108
rect 2412 22024 2464 22030
rect 2412 21966 2464 21972
rect 1676 21888 1728 21894
rect 1676 21830 1728 21836
rect 1688 21729 1716 21830
rect 1674 21720 1730 21729
rect 2424 21690 2452 21966
rect 1674 21655 1730 21664
rect 2412 21684 2464 21690
rect 2412 21626 2464 21632
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 2412 21548 2464 21554
rect 2412 21490 2464 21496
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 1688 21185 1716 21286
rect 1674 21176 1730 21185
rect 2424 21146 2452 21490
rect 1674 21111 1730 21120
rect 2412 21140 2464 21146
rect 2412 21082 2464 21088
rect 1676 20800 1728 20806
rect 1676 20742 1728 20748
rect 1688 20641 1716 20742
rect 1674 20632 1730 20641
rect 1674 20567 1730 20576
rect 1676 20256 1728 20262
rect 1676 20198 1728 20204
rect 1688 20097 1716 20198
rect 1674 20088 1730 20097
rect 2516 20058 2544 21626
rect 1674 20023 1730 20032
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 19553 1716 19654
rect 1674 19544 1730 19553
rect 1674 19479 1730 19488
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 1688 19009 1716 19110
rect 1674 19000 1730 19009
rect 2608 18970 2636 22510
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 1674 18935 1730 18944
rect 2596 18964 2648 18970
rect 2596 18906 2648 18912
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1688 18465 1716 18566
rect 1674 18456 1730 18465
rect 1674 18391 1730 18400
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17921 1624 18022
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 1582 17912 1638 17921
rect 4214 17915 4522 17924
rect 1582 17847 1638 17856
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1688 17377 1716 17478
rect 1674 17368 1730 17377
rect 1674 17303 1730 17312
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 16833 1716 16934
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 1674 16824 1730 16833
rect 4214 16827 4522 16836
rect 1674 16759 1730 16768
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1688 16289 1716 16390
rect 1674 16280 1730 16289
rect 1674 16215 1730 16224
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15745 1716 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 1674 15736 1730 15745
rect 4214 15739 4522 15748
rect 1674 15671 1730 15680
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1688 15201 1716 15302
rect 1674 15192 1730 15201
rect 1674 15127 1730 15136
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1688 14657 1716 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 1674 14648 1730 14657
rect 4214 14651 4522 14660
rect 1674 14583 1730 14592
rect 4632 14482 4660 14962
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11716 14482 11744 14894
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 4344 14340 4396 14346
rect 4344 14282 4396 14288
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1688 14113 1716 14214
rect 1674 14104 1730 14113
rect 1674 14039 1730 14048
rect 4356 13938 4384 14282
rect 13188 14278 13216 14758
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 13188 13734 13216 14214
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 1688 13569 1716 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 1674 13560 1730 13569
rect 4214 13563 4522 13572
rect 1674 13495 1730 13504
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1688 13025 1716 13126
rect 1674 13016 1730 13025
rect 1872 12986 1900 13262
rect 13188 13190 13216 13670
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 1674 12951 1730 12960
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 13188 12850 13216 13126
rect 13372 12850 13400 29038
rect 13464 25226 13492 34478
rect 13544 33380 13596 33386
rect 13544 33322 13596 33328
rect 13452 25220 13504 25226
rect 13452 25162 13504 25168
rect 13556 12850 13584 33322
rect 13820 29572 13872 29578
rect 13820 29514 13872 29520
rect 13832 29170 13860 29514
rect 13820 29164 13872 29170
rect 13820 29106 13872 29112
rect 14188 29164 14240 29170
rect 14188 29106 14240 29112
rect 14200 28422 14228 29106
rect 14188 28416 14240 28422
rect 14188 28358 14240 28364
rect 14568 25770 14596 34886
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14752 34202 14780 34546
rect 15028 34542 15056 34954
rect 15672 34610 15700 35022
rect 15660 34604 15712 34610
rect 15660 34546 15712 34552
rect 16684 34542 16712 35226
rect 15016 34536 15068 34542
rect 15016 34478 15068 34484
rect 16672 34536 16724 34542
rect 16672 34478 16724 34484
rect 14740 34196 14792 34202
rect 14740 34138 14792 34144
rect 14556 25764 14608 25770
rect 14556 25706 14608 25712
rect 14648 24404 14700 24410
rect 14648 24346 14700 24352
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 14108 21554 14136 22374
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 13924 20942 13952 21286
rect 13912 20936 13964 20942
rect 13912 20878 13964 20884
rect 14476 19854 14504 24006
rect 14660 23526 14688 24346
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 14660 22982 14688 23462
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 14292 19378 14320 19654
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 14568 16250 14596 22646
rect 14660 22438 14688 22918
rect 14752 22642 14780 34138
rect 15028 31362 15056 34478
rect 15108 33312 15160 33318
rect 15108 33254 15160 33260
rect 15120 32842 15148 33254
rect 15108 32836 15160 32842
rect 15108 32778 15160 32784
rect 17328 31754 17356 36246
rect 19352 35086 19380 39918
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 21468 38214 21496 52974
rect 22020 52698 22048 53042
rect 24032 52964 24084 52970
rect 24032 52906 24084 52912
rect 22284 52896 22336 52902
rect 22284 52838 22336 52844
rect 22008 52692 22060 52698
rect 22008 52634 22060 52640
rect 22192 45348 22244 45354
rect 22192 45290 22244 45296
rect 22204 39642 22232 45290
rect 22296 44470 22324 52838
rect 22836 52488 22888 52494
rect 22836 52430 22888 52436
rect 22284 44464 22336 44470
rect 22284 44406 22336 44412
rect 22744 39908 22796 39914
rect 22744 39850 22796 39856
rect 22192 39636 22244 39642
rect 22192 39578 22244 39584
rect 22756 39030 22784 39850
rect 22744 39024 22796 39030
rect 22744 38966 22796 38972
rect 21916 38412 21968 38418
rect 21916 38354 21968 38360
rect 21456 38208 21508 38214
rect 21456 38150 21508 38156
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 21270 36136 21326 36145
rect 21270 36071 21272 36080
rect 21324 36071 21326 36080
rect 21272 36042 21324 36048
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 20812 35828 20864 35834
rect 20812 35770 20864 35776
rect 20824 35494 20852 35770
rect 20812 35488 20864 35494
rect 20812 35430 20864 35436
rect 19340 35080 19392 35086
rect 19340 35022 19392 35028
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 17868 34536 17920 34542
rect 17868 34478 17920 34484
rect 17236 31726 17356 31754
rect 15028 31334 15148 31362
rect 15120 28422 15148 31334
rect 15108 28416 15160 28422
rect 15108 28358 15160 28364
rect 15120 28014 15148 28358
rect 15108 28008 15160 28014
rect 15108 27950 15160 27956
rect 14924 25764 14976 25770
rect 14924 25706 14976 25712
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 14752 22234 14780 22578
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14292 15094 14320 15846
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13740 12850 13768 13398
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12481 1716 12582
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 1674 12472 1730 12481
rect 4214 12475 4522 12484
rect 1674 12407 1730 12416
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 1688 11937 1716 12038
rect 1674 11928 1730 11937
rect 1674 11863 1730 11872
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 11393 1716 11494
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 1674 11384 1730 11393
rect 4214 11387 4522 11396
rect 1674 11319 1730 11328
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1688 10849 1716 10950
rect 1674 10840 1730 10849
rect 11072 10810 11100 11086
rect 1674 10775 1730 10784
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10305 1716 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 1674 10296 1730 10305
rect 4214 10299 4522 10308
rect 1674 10231 1730 10240
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9761 1716 9862
rect 1674 9752 1730 9761
rect 1674 9687 1730 9696
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 9217 1716 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 1674 9208 1730 9217
rect 4214 9211 4522 9220
rect 1674 9143 1730 9152
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 8673 1716 8774
rect 1674 8664 1730 8673
rect 1674 8599 1730 8608
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1688 8129 1716 8298
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 1674 8120 1730 8129
rect 4214 8123 4522 8132
rect 1674 8055 1730 8064
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7585 1716 7686
rect 1674 7576 1730 7585
rect 11072 7546 11100 8434
rect 1674 7511 1730 7520
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 7041 1716 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 1674 7032 1730 7041
rect 4214 7035 4522 7044
rect 1674 6967 1730 6976
rect 11072 6866 11100 7346
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 1688 6497 1716 6598
rect 1674 6488 1730 6497
rect 1674 6423 1730 6432
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 5953 1716 6054
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 1674 5944 1730 5953
rect 4214 5947 4522 5956
rect 1674 5879 1730 5888
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1688 5409 1716 5510
rect 1674 5400 1730 5409
rect 1674 5335 1730 5344
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4865 1716 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 1674 4856 1730 4865
rect 4214 4859 4522 4868
rect 1674 4791 1730 4800
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1688 4321 1716 4422
rect 1674 4312 1730 4321
rect 1674 4247 1730 4256
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 1688 3777 1716 3878
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 1674 3768 1730 3777
rect 4214 3771 4522 3780
rect 1674 3703 1730 3712
rect 6840 3534 6868 3878
rect 7116 3738 7144 5102
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1688 3233 1716 3334
rect 1674 3224 1730 3233
rect 1674 3159 1730 3168
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 5460 2106 5488 2246
rect 5448 2100 5500 2106
rect 5448 2042 5500 2048
rect 6012 2038 6040 2246
rect 6000 2032 6052 2038
rect 6000 1974 6052 1980
rect 6840 800 6868 3470
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7024 3058 7052 3334
rect 7668 3194 7696 3878
rect 7760 3534 7788 4422
rect 8312 3738 8340 6326
rect 12084 6254 12112 6598
rect 12544 6458 12572 7346
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8404 3534 8432 3878
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7668 3058 7696 3130
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7024 2774 7052 2994
rect 7760 2774 7788 3470
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 7024 2746 7236 2774
rect 7760 2746 7972 2774
rect 7208 800 7236 2746
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7576 800 7604 2382
rect 7944 800 7972 2746
rect 8312 800 8340 3130
rect 8404 3126 8432 3470
rect 8496 3194 8524 3606
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 8680 2310 8708 4490
rect 9600 4162 9628 4966
rect 9600 4134 9720 4162
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9600 3738 9628 4014
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9600 3466 9628 3674
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9692 3398 9720 4134
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8772 3058 8800 3130
rect 8956 3058 8984 3334
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8680 800 8708 2246
rect 9048 800 9076 3062
rect 9416 800 9444 3130
rect 9692 2774 9720 3334
rect 9784 3194 9812 3946
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9876 3058 9904 4966
rect 10520 4826 10548 5170
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10704 4622 10732 4966
rect 10888 4622 10916 6122
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10048 3936 10100 3942
rect 10046 3904 10048 3913
rect 10100 3904 10102 3913
rect 10046 3839 10102 3848
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10138 3632 10194 3641
rect 10138 3567 10140 3576
rect 10192 3567 10194 3576
rect 10140 3538 10192 3544
rect 9956 3392 10008 3398
rect 9954 3360 9956 3369
rect 10008 3360 10010 3369
rect 9954 3295 10010 3304
rect 10244 3058 10272 3674
rect 10336 3670 10364 4150
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10428 3738 10456 4082
rect 10520 4078 10548 4558
rect 10704 4078 10732 4558
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10796 3942 10824 4422
rect 10888 4078 10916 4558
rect 10980 4282 11008 4558
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10784 3936 10836 3942
rect 10690 3904 10746 3913
rect 10784 3878 10836 3884
rect 10690 3839 10746 3848
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10704 3510 10732 3839
rect 10692 3504 10744 3510
rect 10692 3446 10744 3452
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 9692 2746 9812 2774
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9692 2106 9720 2382
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 9784 800 9812 2746
rect 10152 800 10180 2994
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 10336 2582 10364 2926
rect 10796 2774 10824 3878
rect 10888 3670 10916 4014
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 3369 10916 3470
rect 10874 3360 10930 3369
rect 10874 3295 10930 3304
rect 10980 3194 11008 4014
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10520 2746 10824 2774
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 10520 800 10548 2746
rect 11072 2650 11100 3946
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10876 2440 10928 2446
rect 11164 2428 11192 5510
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11256 2582 11284 4694
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3534 11468 3878
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11532 2650 11560 5782
rect 12084 5642 12112 6190
rect 12452 6118 12480 6326
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 11716 4554 11744 5578
rect 12452 5370 12480 5646
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12440 5160 12492 5166
rect 12438 5128 12440 5137
rect 12492 5128 12494 5137
rect 11796 5092 11848 5098
rect 12438 5063 12494 5072
rect 11796 5034 11848 5040
rect 11704 4548 11756 4554
rect 11704 4490 11756 4496
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11624 3534 11652 4422
rect 11716 4078 11744 4490
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11612 3052 11664 3058
rect 11716 3040 11744 4014
rect 11808 3058 11836 5034
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 4146 12388 4966
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12544 3942 12572 5782
rect 12636 5710 12664 12038
rect 13188 11558 13216 12786
rect 13372 11898 13400 12786
rect 13556 12442 13584 12786
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13740 12102 13768 12786
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 12238 13952 12582
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 14016 12170 14044 14010
rect 14568 14006 14596 16186
rect 14738 15464 14794 15473
rect 14738 15399 14740 15408
rect 14792 15399 14794 15408
rect 14740 15370 14792 15376
rect 14738 15056 14794 15065
rect 14738 14991 14740 15000
rect 14792 14991 14794 15000
rect 14740 14962 14792 14968
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14646 14376 14702 14385
rect 14646 14311 14702 14320
rect 14464 14000 14516 14006
rect 14462 13968 14464 13977
rect 14556 14000 14608 14006
rect 14516 13968 14518 13977
rect 14556 13942 14608 13948
rect 14462 13903 14518 13912
rect 14660 13326 14688 14311
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14200 12850 14228 12922
rect 14752 12850 14780 14418
rect 14844 13190 14872 16458
rect 14936 14278 14964 25706
rect 15120 24410 15148 27950
rect 15108 24404 15160 24410
rect 15108 24346 15160 24352
rect 15120 24206 15148 24346
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 17236 22778 17264 31726
rect 17880 30802 17908 34478
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 20824 31346 20852 35430
rect 21178 35320 21234 35329
rect 21178 35255 21234 35264
rect 21192 35154 21220 35255
rect 21180 35148 21232 35154
rect 21180 35090 21232 35096
rect 21192 35057 21220 35090
rect 21732 35080 21784 35086
rect 21178 35048 21234 35057
rect 21178 34983 21234 34992
rect 21730 35048 21732 35057
rect 21784 35048 21786 35057
rect 21730 34983 21786 34992
rect 20812 31340 20864 31346
rect 20812 31282 20864 31288
rect 17868 30796 17920 30802
rect 17868 30738 17920 30744
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 21928 29102 21956 38354
rect 22008 37868 22060 37874
rect 22008 37810 22060 37816
rect 22020 34202 22048 37810
rect 22376 37324 22428 37330
rect 22376 37266 22428 37272
rect 22388 37233 22416 37266
rect 22374 37224 22430 37233
rect 22374 37159 22430 37168
rect 22284 36304 22336 36310
rect 22284 36246 22336 36252
rect 22296 35834 22324 36246
rect 22284 35828 22336 35834
rect 22284 35770 22336 35776
rect 22008 34196 22060 34202
rect 22008 34138 22060 34144
rect 22388 30258 22416 37159
rect 22558 36680 22614 36689
rect 22558 36615 22560 36624
rect 22612 36615 22614 36624
rect 22560 36586 22612 36592
rect 22652 36576 22704 36582
rect 22652 36518 22704 36524
rect 22560 35556 22612 35562
rect 22560 35498 22612 35504
rect 22572 34678 22600 35498
rect 22560 34672 22612 34678
rect 22560 34614 22612 34620
rect 22664 34066 22692 36518
rect 22652 34060 22704 34066
rect 22652 34002 22704 34008
rect 22756 31754 22784 38966
rect 22848 38654 22876 52430
rect 22928 44804 22980 44810
rect 22928 44746 22980 44752
rect 22940 39370 22968 44746
rect 23848 42696 23900 42702
rect 23848 42638 23900 42644
rect 23388 42628 23440 42634
rect 23388 42570 23440 42576
rect 23400 40730 23428 42570
rect 23860 42022 23888 42638
rect 23848 42016 23900 42022
rect 23848 41958 23900 41964
rect 23388 40724 23440 40730
rect 23388 40666 23440 40672
rect 23572 40384 23624 40390
rect 23386 40352 23442 40361
rect 23572 40326 23624 40332
rect 23386 40287 23442 40296
rect 23400 40050 23428 40287
rect 23388 40044 23440 40050
rect 23388 39986 23440 39992
rect 22928 39364 22980 39370
rect 22928 39306 22980 39312
rect 22940 39098 22968 39306
rect 23480 39296 23532 39302
rect 23480 39238 23532 39244
rect 22928 39092 22980 39098
rect 22928 39034 22980 39040
rect 23020 38888 23072 38894
rect 23020 38830 23072 38836
rect 23032 38654 23060 38830
rect 22848 38626 22968 38654
rect 23032 38626 23152 38654
rect 22940 36038 22968 38626
rect 23124 37942 23152 38626
rect 23492 38593 23520 39238
rect 23584 39098 23612 40326
rect 23860 40050 23888 41958
rect 24044 41138 24072 52906
rect 24504 52154 24532 53110
rect 24596 53106 24624 55270
rect 25594 55270 25728 55298
rect 25594 55200 25650 55270
rect 25596 53236 25648 53242
rect 25596 53178 25648 53184
rect 24584 53100 24636 53106
rect 24584 53042 24636 53048
rect 25412 52896 25464 52902
rect 25412 52838 25464 52844
rect 24492 52148 24544 52154
rect 24492 52090 24544 52096
rect 25424 52086 25452 52838
rect 25504 52352 25556 52358
rect 25504 52294 25556 52300
rect 25412 52080 25464 52086
rect 25412 52022 25464 52028
rect 25516 52018 25544 52294
rect 25504 52012 25556 52018
rect 25504 51954 25556 51960
rect 25516 51610 25544 51954
rect 25504 51604 25556 51610
rect 25504 51546 25556 51552
rect 25136 50448 25188 50454
rect 25136 50390 25188 50396
rect 24768 44260 24820 44266
rect 24768 44202 24820 44208
rect 24216 42152 24268 42158
rect 24216 42094 24268 42100
rect 24032 41132 24084 41138
rect 24032 41074 24084 41080
rect 23848 40044 23900 40050
rect 23848 39986 23900 39992
rect 23940 39296 23992 39302
rect 23940 39238 23992 39244
rect 23572 39092 23624 39098
rect 23572 39034 23624 39040
rect 23952 38826 23980 39238
rect 23940 38820 23992 38826
rect 23940 38762 23992 38768
rect 23478 38584 23534 38593
rect 23478 38519 23534 38528
rect 23112 37936 23164 37942
rect 23112 37878 23164 37884
rect 23124 37738 23152 37878
rect 23112 37732 23164 37738
rect 23112 37674 23164 37680
rect 23020 37120 23072 37126
rect 23020 37062 23072 37068
rect 22928 36032 22980 36038
rect 22926 36000 22928 36009
rect 22980 36000 22982 36009
rect 22926 35935 22982 35944
rect 23032 35601 23060 37062
rect 23018 35592 23074 35601
rect 23018 35527 23074 35536
rect 23032 35494 23060 35527
rect 23020 35488 23072 35494
rect 23020 35430 23072 35436
rect 23032 34474 23060 35430
rect 23124 35086 23152 37674
rect 23492 36378 23520 38519
rect 23572 37664 23624 37670
rect 23572 37606 23624 37612
rect 23480 36372 23532 36378
rect 23480 36314 23532 36320
rect 23584 36038 23612 37606
rect 23952 37262 23980 38762
rect 24032 38208 24084 38214
rect 24030 38176 24032 38185
rect 24084 38176 24086 38185
rect 24030 38111 24086 38120
rect 24030 37496 24086 37505
rect 24030 37431 24032 37440
rect 24084 37431 24086 37440
rect 24032 37402 24084 37408
rect 23940 37256 23992 37262
rect 23940 37198 23992 37204
rect 23664 36916 23716 36922
rect 23664 36858 23716 36864
rect 23676 36582 23704 36858
rect 23664 36576 23716 36582
rect 23664 36518 23716 36524
rect 23572 36032 23624 36038
rect 23572 35974 23624 35980
rect 24228 35834 24256 42094
rect 24492 41676 24544 41682
rect 24492 41618 24544 41624
rect 24400 41472 24452 41478
rect 24400 41414 24452 41420
rect 24412 41206 24440 41414
rect 24504 41274 24532 41618
rect 24676 41540 24728 41546
rect 24676 41482 24728 41488
rect 24492 41268 24544 41274
rect 24492 41210 24544 41216
rect 24400 41200 24452 41206
rect 24400 41142 24452 41148
rect 24412 40186 24440 41142
rect 24504 40458 24532 41210
rect 24688 40526 24716 41482
rect 24676 40520 24728 40526
rect 24676 40462 24728 40468
rect 24492 40452 24544 40458
rect 24492 40394 24544 40400
rect 24400 40180 24452 40186
rect 24400 40122 24452 40128
rect 24308 39296 24360 39302
rect 24308 39238 24360 39244
rect 24320 39098 24348 39238
rect 24308 39092 24360 39098
rect 24308 39034 24360 39040
rect 24412 38758 24440 40122
rect 24584 39568 24636 39574
rect 24584 39510 24636 39516
rect 24596 39030 24624 39510
rect 24584 39024 24636 39030
rect 24584 38966 24636 38972
rect 24400 38752 24452 38758
rect 24400 38694 24452 38700
rect 24780 38654 24808 44202
rect 24860 42220 24912 42226
rect 24860 42162 24912 42168
rect 24872 41818 24900 42162
rect 24950 41984 25006 41993
rect 24950 41919 25006 41928
rect 24860 41812 24912 41818
rect 24860 41754 24912 41760
rect 24964 41478 24992 41919
rect 25044 41744 25096 41750
rect 25044 41686 25096 41692
rect 24952 41472 25004 41478
rect 24952 41414 25004 41420
rect 24964 39098 24992 41414
rect 25056 40186 25084 41686
rect 25044 40180 25096 40186
rect 25044 40122 25096 40128
rect 25044 40044 25096 40050
rect 25044 39986 25096 39992
rect 25056 39438 25084 39986
rect 25044 39432 25096 39438
rect 25044 39374 25096 39380
rect 24952 39092 25004 39098
rect 24952 39034 25004 39040
rect 24858 38992 24914 39001
rect 24858 38927 24914 38936
rect 24872 38758 24900 38927
rect 24860 38752 24912 38758
rect 24860 38694 24912 38700
rect 24596 38626 24808 38654
rect 24308 37800 24360 37806
rect 24308 37742 24360 37748
rect 23296 35828 23348 35834
rect 23296 35770 23348 35776
rect 23664 35828 23716 35834
rect 23664 35770 23716 35776
rect 24032 35828 24084 35834
rect 24032 35770 24084 35776
rect 24216 35828 24268 35834
rect 24216 35770 24268 35776
rect 23308 35494 23336 35770
rect 23480 35760 23532 35766
rect 23478 35728 23480 35737
rect 23532 35728 23534 35737
rect 23478 35663 23534 35672
rect 23572 35692 23624 35698
rect 23572 35634 23624 35640
rect 23296 35488 23348 35494
rect 23296 35430 23348 35436
rect 23112 35080 23164 35086
rect 23112 35022 23164 35028
rect 23296 35080 23348 35086
rect 23480 35080 23532 35086
rect 23296 35022 23348 35028
rect 23478 35048 23480 35057
rect 23532 35048 23534 35057
rect 23020 34468 23072 34474
rect 23020 34410 23072 34416
rect 22836 34400 22888 34406
rect 22836 34342 22888 34348
rect 22848 34202 22876 34342
rect 22836 34196 22888 34202
rect 22836 34138 22888 34144
rect 23032 32230 23060 34410
rect 23124 33658 23152 35022
rect 23112 33652 23164 33658
rect 23112 33594 23164 33600
rect 23020 32224 23072 32230
rect 23020 32166 23072 32172
rect 22572 31726 22784 31754
rect 22376 30252 22428 30258
rect 22376 30194 22428 30200
rect 21916 29096 21968 29102
rect 21916 29038 21968 29044
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 18788 22704 18840 22710
rect 18788 22646 18840 22652
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15304 22098 15332 22374
rect 15292 22092 15344 22098
rect 18800 22094 18828 22646
rect 15292 22034 15344 22040
rect 18708 22066 18828 22094
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15396 16250 15424 17614
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15108 16176 15160 16182
rect 15106 16144 15108 16153
rect 15160 16144 15162 16153
rect 15106 16079 15162 16088
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 13938 14964 14214
rect 15028 14074 15056 15302
rect 15120 14618 15148 15370
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15396 14822 15424 14962
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15106 14512 15162 14521
rect 15106 14447 15108 14456
rect 15160 14447 15162 14456
rect 15108 14418 15160 14424
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14922 13560 14978 13569
rect 14922 13495 14924 13504
rect 14976 13495 14978 13504
rect 14924 13466 14976 13472
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11014 13768 11494
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13832 10606 13860 11018
rect 14016 10742 14044 11018
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12728 3738 12756 6122
rect 12820 4826 12848 6122
rect 12912 5914 12940 7822
rect 13004 7342 13032 7890
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13004 6458 13032 6734
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 13096 6458 13124 6666
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 13004 5846 13032 6190
rect 13096 5914 13124 6258
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12912 4826 12940 5170
rect 13004 5098 13032 5782
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 11664 3012 11744 3040
rect 11796 3052 11848 3058
rect 11612 2994 11664 3000
rect 11796 2994 11848 3000
rect 11808 2666 11836 2994
rect 11520 2644 11572 2650
rect 11808 2638 12020 2666
rect 11520 2586 11572 2592
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 11612 2440 11664 2446
rect 10928 2400 11284 2428
rect 10876 2382 10928 2388
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10888 800 10916 2042
rect 11256 800 11284 2400
rect 11612 2382 11664 2388
rect 11624 2038 11652 2382
rect 11612 2032 11664 2038
rect 11612 1974 11664 1980
rect 11624 800 11652 1974
rect 11992 800 12020 2638
rect 12360 800 12388 3470
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12530 2816 12586 2825
rect 12530 2751 12586 2760
rect 12544 2650 12572 2751
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12728 800 12756 2926
rect 12820 2446 12848 4558
rect 13004 4486 13032 5034
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12912 3194 12940 3878
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 12912 2825 12940 2994
rect 13004 2922 13032 4150
rect 13096 3670 13124 4694
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 12992 2916 13044 2922
rect 12992 2858 13044 2864
rect 12898 2816 12954 2825
rect 13188 2774 13216 10134
rect 14016 10130 14044 10678
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14016 9654 14044 10066
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 12898 2751 12954 2760
rect 13096 2746 13216 2774
rect 13096 2650 13124 2746
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 12820 762 12848 2382
rect 13280 2310 13308 9046
rect 13372 3738 13400 9386
rect 14108 8974 14136 9454
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13464 6798 13492 7278
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13464 5914 13492 6734
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13556 5846 13584 6734
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13464 4554 13492 5102
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13556 4078 13584 5646
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 13004 870 13124 898
rect 13004 762 13032 870
rect 13096 800 13124 870
rect 13464 800 13492 3470
rect 13648 3194 13676 8298
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13740 7546 13768 7890
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 14200 6458 14228 12786
rect 14844 12434 14872 13126
rect 15120 12918 15148 13942
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 13326 15332 13670
rect 15396 13394 15424 14758
rect 15488 14482 15516 18838
rect 15566 16008 15622 16017
rect 15566 15943 15622 15952
rect 15580 15910 15608 15943
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15580 14618 15608 15438
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 15488 12434 15516 14214
rect 15580 13530 15608 14282
rect 15672 13734 15700 14350
rect 15856 13938 15884 19858
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15948 15094 15976 15506
rect 15936 15088 15988 15094
rect 15936 15030 15988 15036
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15948 14278 15976 14758
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15948 13870 15976 14214
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15948 13326 15976 13806
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15948 12782 15976 13262
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 15856 12442 15884 12650
rect 14844 12406 14964 12434
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 13820 5160 13872 5166
rect 13818 5128 13820 5137
rect 13872 5128 13874 5137
rect 13728 5092 13780 5098
rect 13818 5063 13874 5072
rect 13728 5034 13780 5040
rect 13740 4214 13768 5034
rect 13912 4548 13964 4554
rect 13912 4490 13964 4496
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13740 3534 13768 3878
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13648 2938 13676 2994
rect 13648 2910 13860 2938
rect 13832 800 13860 2910
rect 13924 2446 13952 4490
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14108 3058 14136 3878
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 13924 2106 13952 2382
rect 14200 2378 14228 5170
rect 14292 3194 14320 10474
rect 14384 10266 14412 10474
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14476 9602 14504 11222
rect 14384 9574 14504 9602
rect 14556 9580 14608 9586
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14384 2774 14412 9574
rect 14556 9522 14608 9528
rect 14568 9178 14596 9522
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14660 8974 14688 9454
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14476 8566 14504 8774
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14568 8480 14596 8842
rect 14648 8492 14700 8498
rect 14568 8452 14648 8480
rect 14648 8434 14700 8440
rect 14660 8401 14688 8434
rect 14646 8392 14702 8401
rect 14646 8327 14702 8336
rect 14660 8090 14688 8327
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14752 5098 14780 8910
rect 14844 5302 14872 12038
rect 14936 11694 14964 12406
rect 15396 12406 15516 12434
rect 15844 12436 15896 12442
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14936 10606 14964 11630
rect 15028 11150 15056 12038
rect 15212 11778 15240 12106
rect 15120 11750 15240 11778
rect 15120 11694 15148 11750
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14832 5296 14884 5302
rect 14832 5238 14884 5244
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14462 3632 14518 3641
rect 14462 3567 14464 3576
rect 14516 3567 14518 3576
rect 14464 3538 14516 3544
rect 14568 3534 14596 4422
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14660 3602 14688 4014
rect 14936 3942 14964 10542
rect 15028 10266 15056 10610
rect 15212 10470 15240 11630
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15304 11354 15332 11562
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15304 10606 15332 11154
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15304 10198 15332 10542
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15028 9382 15056 9998
rect 15212 9722 15240 9998
rect 15396 9722 15424 12406
rect 15844 12378 15896 12384
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15764 11898 15792 12242
rect 15948 12238 15976 12718
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15856 11762 15884 12038
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15948 11694 15976 12174
rect 15936 11688 15988 11694
rect 15856 11636 15936 11642
rect 15856 11630 15988 11636
rect 15856 11614 15976 11630
rect 15856 11014 15884 11614
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15120 9450 15148 9522
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15120 4010 15148 8366
rect 15212 8090 15240 9658
rect 15488 8634 15516 9998
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15304 7970 15332 8298
rect 15212 7942 15332 7970
rect 15212 4622 15240 7942
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14292 2746 14412 2774
rect 14292 2650 14320 2746
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 13912 2100 13964 2106
rect 13912 2042 13964 2048
rect 14200 800 14228 2314
rect 14568 800 14596 2994
rect 14660 2922 14688 3334
rect 14648 2916 14700 2922
rect 14648 2858 14700 2864
rect 14844 2446 14872 3878
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14936 3194 14964 3470
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 15212 2990 15240 4558
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15396 3058 15424 3878
rect 15580 3194 15608 10474
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15672 9450 15700 10066
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15660 9444 15712 9450
rect 15660 9386 15712 9392
rect 15764 9217 15792 9454
rect 15750 9208 15806 9217
rect 15750 9143 15806 9152
rect 15764 7546 15792 9143
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15856 3738 15884 10950
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15396 2774 15424 2994
rect 15304 2746 15424 2774
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 14924 2100 14976 2106
rect 14924 2042 14976 2048
rect 14936 800 14964 2042
rect 15304 800 15332 2746
rect 15948 2582 15976 11222
rect 16040 10266 16068 14350
rect 16132 13530 16160 16594
rect 16500 15706 16528 17138
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16500 14482 16528 14758
rect 16592 14618 16620 16526
rect 16684 15026 16712 16934
rect 16762 16688 16818 16697
rect 16762 16623 16764 16632
rect 16816 16623 16818 16632
rect 16948 16652 17000 16658
rect 16764 16594 16816 16600
rect 16948 16594 17000 16600
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16592 13938 16620 14282
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16132 12986 16160 13466
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16316 12850 16344 13126
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16132 12170 16160 12786
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 16132 11694 16160 12106
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16132 11218 16160 11630
rect 16224 11354 16252 12718
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16212 9648 16264 9654
rect 16210 9616 16212 9625
rect 16264 9616 16266 9625
rect 16210 9551 16266 9560
rect 16408 9518 16436 13806
rect 16684 13326 16712 14962
rect 16776 13734 16804 15982
rect 16868 15706 16896 16050
rect 16960 16046 16988 16594
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16960 15502 16988 15982
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16500 9178 16528 13262
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16684 12238 16712 12310
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16592 10810 16620 12174
rect 16868 11082 16896 13874
rect 16960 11830 16988 15438
rect 17052 13852 17080 19450
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 17236 18086 17264 18634
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17144 17202 17172 17478
rect 17236 17338 17264 18022
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17696 16998 17724 17478
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17236 16232 17264 16526
rect 17972 16522 18000 18158
rect 18156 17270 18184 21286
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 18426 18368 18566
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18234 17776 18290 17785
rect 18234 17711 18236 17720
rect 18288 17711 18290 17720
rect 18236 17682 18288 17688
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 17316 16244 17368 16250
rect 17236 16204 17316 16232
rect 17316 16186 17368 16192
rect 17500 16176 17552 16182
rect 17500 16118 17552 16124
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17224 16040 17276 16046
rect 17144 16000 17224 16028
rect 17144 15502 17172 16000
rect 17420 16017 17448 16050
rect 17224 15982 17276 15988
rect 17406 16008 17462 16017
rect 17406 15943 17462 15952
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17144 14890 17172 15438
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17144 14346 17172 14826
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 17132 13864 17184 13870
rect 17052 13824 17132 13852
rect 17132 13806 17184 13812
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17052 12986 17080 13194
rect 17144 12986 17172 13398
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 16040 5030 16068 5306
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 15936 2576 15988 2582
rect 15936 2518 15988 2524
rect 16132 2446 16160 3334
rect 16224 2650 16252 9046
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16408 3058 16436 3334
rect 16592 3194 16620 9386
rect 16684 8362 16712 11018
rect 16856 10192 16908 10198
rect 16776 10140 16856 10146
rect 16776 10134 16908 10140
rect 16776 10118 16896 10134
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16776 3194 16804 10118
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16960 8906 16988 9114
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 12820 734 13032 762
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15396 762 15424 2382
rect 15580 870 15700 898
rect 15580 762 15608 870
rect 15672 800 15700 870
rect 16040 800 16068 2382
rect 16408 800 16436 2994
rect 17052 2650 17080 12310
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17144 10062 17172 12174
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 17144 9722 17172 9998
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17144 8566 17172 9658
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17144 8090 17172 8502
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17144 7750 17172 8026
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17144 7410 17172 7686
rect 17236 7546 17264 15438
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17328 12442 17356 14894
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17420 14482 17448 14758
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17328 10606 17356 10950
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17328 9654 17356 10542
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17328 9178 17356 9590
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17314 8936 17370 8945
rect 17314 8871 17316 8880
rect 17368 8871 17370 8880
rect 17316 8842 17368 8848
rect 17420 8634 17448 13806
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17512 8090 17540 16118
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17604 15434 17632 15982
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17604 14074 17632 14894
rect 17696 14770 17724 15030
rect 17788 14890 17816 15642
rect 17776 14884 17828 14890
rect 17776 14826 17828 14832
rect 17696 14742 17816 14770
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17604 13569 17632 13874
rect 17590 13560 17646 13569
rect 17590 13495 17646 13504
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17604 12918 17632 13262
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17604 11762 17632 12378
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17512 6866 17540 7346
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17236 5710 17264 6054
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16776 800 16804 2382
rect 17144 2310 17172 2994
rect 17420 2650 17448 6802
rect 17512 6458 17540 6802
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17604 3194 17632 8298
rect 17696 6662 17724 14350
rect 17788 11558 17816 14742
rect 17880 14414 17908 15846
rect 17972 15570 18000 15846
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 18156 15450 18184 17206
rect 18248 16794 18276 17546
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18248 16590 18276 16730
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18340 16182 18368 17070
rect 18328 16176 18380 16182
rect 18328 16118 18380 16124
rect 18156 15422 18276 15450
rect 18248 15366 18276 15422
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 17868 14408 17920 14414
rect 18156 14385 18184 15302
rect 18340 15094 18368 16118
rect 18432 16114 18460 18022
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18420 15088 18472 15094
rect 18420 15030 18472 15036
rect 18432 14618 18460 15030
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 17868 14350 17920 14356
rect 18142 14376 18198 14385
rect 17960 14340 18012 14346
rect 18142 14311 18198 14320
rect 17960 14282 18012 14288
rect 17972 13190 18000 14282
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17972 12714 18000 13126
rect 18156 12782 18184 14214
rect 18616 14074 18644 15302
rect 18708 15162 18736 22066
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 21192 21418 21220 21966
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21180 21412 21232 21418
rect 21180 21354 21232 21360
rect 21376 21146 21404 21422
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 19984 21072 20036 21078
rect 19984 21014 20036 21020
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18708 14278 18736 15098
rect 18800 14482 18828 15506
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18236 14000 18288 14006
rect 18236 13942 18288 13948
rect 18248 12986 18276 13942
rect 18340 13326 18368 14010
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17880 12238 17908 12310
rect 18248 12306 18276 12922
rect 18432 12434 18460 13670
rect 18800 12434 18828 14418
rect 18984 13734 19012 20334
rect 19248 20256 19300 20262
rect 19248 20198 19300 20204
rect 19260 19378 19288 20198
rect 19628 20058 19656 20402
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19996 19854 20024 21014
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21468 20398 21496 20742
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 20088 19514 20116 19654
rect 20180 19514 20208 19858
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19352 18358 19380 19382
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19062 17776 19118 17785
rect 19352 17746 19380 18294
rect 19062 17711 19118 17720
rect 19340 17740 19392 17746
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18432 12406 18552 12434
rect 18800 12406 18920 12434
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17776 11552 17828 11558
rect 17828 11500 17908 11506
rect 17776 11494 17908 11500
rect 17788 11478 17908 11494
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17788 10266 17816 11018
rect 17880 10554 17908 11478
rect 17972 10742 18000 11698
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 18064 10674 18092 12038
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17880 10526 18000 10554
rect 17972 10418 18000 10526
rect 18052 10532 18104 10538
rect 18156 10520 18184 12174
rect 18524 12102 18552 12406
rect 18892 12306 18920 12406
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11898 18552 12038
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18696 11280 18748 11286
rect 18696 11222 18748 11228
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18104 10492 18184 10520
rect 18052 10474 18104 10480
rect 17972 10390 18184 10418
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17880 10062 17908 10202
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17788 8945 17816 9522
rect 17972 9042 18000 9998
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17774 8936 17830 8945
rect 17774 8871 17830 8880
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17788 3058 17816 3334
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 17144 800 17172 2246
rect 17512 800 17540 2994
rect 17880 2446 17908 3878
rect 17972 3194 18000 7210
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18064 2650 18092 7958
rect 18156 5098 18184 10390
rect 18248 9178 18276 10610
rect 18616 9926 18644 10950
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 18616 9625 18644 9862
rect 18602 9616 18658 9625
rect 18708 9586 18736 11222
rect 18602 9551 18658 9560
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18800 9450 18828 11834
rect 18892 10130 18920 12242
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 19076 9994 19104 17711
rect 19340 17682 19392 17688
rect 19444 17610 19472 18566
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20364 18426 20392 18702
rect 20548 18698 20576 20266
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20640 19378 20668 20198
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 20812 19984 20864 19990
rect 20812 19926 20864 19932
rect 20824 19718 20852 19926
rect 21284 19922 21312 19994
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 18766 20760 19110
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19248 17536 19300 17542
rect 19300 17484 19472 17490
rect 19248 17478 19472 17484
rect 19260 17462 19472 17478
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19352 15162 19380 17274
rect 19444 15586 19472 17462
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20076 17060 20128 17066
rect 20076 17002 20128 17008
rect 20088 16454 20116 17002
rect 20258 16688 20314 16697
rect 20258 16623 20314 16632
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19444 15558 19564 15586
rect 19536 15502 19564 15558
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19444 14414 19472 15438
rect 19996 15366 20024 15982
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20088 15026 20116 16390
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19614 13968 19670 13977
rect 19614 13903 19616 13912
rect 19668 13903 19670 13912
rect 19616 13874 19668 13880
rect 20088 13870 20116 14350
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 19892 13796 19944 13802
rect 19892 13738 19944 13744
rect 19904 13326 19932 13738
rect 20088 13462 20116 13806
rect 20076 13456 20128 13462
rect 20076 13398 20128 13404
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19996 12986 20024 13262
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 20088 12850 20116 13398
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20180 12986 20208 13126
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19260 11558 19288 12174
rect 19352 11694 19380 12582
rect 19800 12368 19852 12374
rect 19798 12336 19800 12345
rect 19852 12336 19854 12345
rect 19798 12271 19854 12280
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19352 11150 19380 11630
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19248 10532 19300 10538
rect 19248 10474 19300 10480
rect 19260 10062 19288 10474
rect 19352 10470 19380 11086
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19064 9988 19116 9994
rect 19064 9930 19116 9936
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18418 9208 18474 9217
rect 18236 9172 18288 9178
rect 18418 9143 18474 9152
rect 18236 9114 18288 9120
rect 18432 9110 18460 9143
rect 18328 9104 18380 9110
rect 18328 9046 18380 9052
rect 18420 9104 18472 9110
rect 18420 9046 18472 9052
rect 18340 7410 18368 9046
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18892 8634 18920 8774
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18524 6458 18552 8434
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18616 7546 18644 7686
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18616 7002 18644 7482
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18800 6798 18828 8434
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18984 6322 19012 9318
rect 19352 8566 19380 10406
rect 19444 10266 19472 11698
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10266 20024 12786
rect 20074 12200 20130 12209
rect 20074 12135 20130 12144
rect 20088 12102 20116 12135
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20180 11286 20208 12038
rect 20168 11280 20220 11286
rect 20168 11222 20220 11228
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 20088 10606 20116 10950
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19444 9042 19472 9862
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9674 20024 9862
rect 19904 9646 20024 9674
rect 19904 9602 19932 9646
rect 19536 9574 19932 9602
rect 19984 9580 20036 9586
rect 19536 9518 19564 9574
rect 19984 9522 20036 9528
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19628 9058 19656 9454
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19536 9042 19656 9058
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19524 9036 19656 9042
rect 19576 9030 19656 9036
rect 19524 8978 19576 8984
rect 19536 8922 19564 8978
rect 19444 8894 19564 8922
rect 19812 8906 19840 9318
rect 19800 8900 19852 8906
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19352 8430 19380 8502
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19444 7954 19472 8894
rect 19800 8842 19852 8848
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19996 8616 20024 9522
rect 20088 9450 20116 10542
rect 20272 9926 20300 16623
rect 20640 16250 20668 18022
rect 20732 17542 20760 18158
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20628 16244 20680 16250
rect 20548 16204 20628 16232
rect 20548 15978 20576 16204
rect 20628 16186 20680 16192
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20640 15978 20668 16050
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20352 15428 20404 15434
rect 20352 15370 20404 15376
rect 20364 12850 20392 15370
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20548 9722 20576 14894
rect 20640 13734 20668 15642
rect 20732 14822 20760 17478
rect 20824 16776 20852 19654
rect 21284 19310 21312 19858
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21560 19378 21588 19654
rect 21548 19372 21600 19378
rect 21548 19314 21600 19320
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21192 18902 21220 19246
rect 21180 18896 21232 18902
rect 21180 18838 21232 18844
rect 21284 18222 21312 19246
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21364 17264 21416 17270
rect 21364 17206 21416 17212
rect 20904 17128 20956 17134
rect 20956 17088 21128 17116
rect 20904 17070 20956 17076
rect 20824 16748 21036 16776
rect 20902 16144 20958 16153
rect 20902 16079 20904 16088
rect 20956 16079 20958 16088
rect 20904 16050 20956 16056
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20824 15638 20852 15846
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20810 15464 20866 15473
rect 20810 15399 20866 15408
rect 20824 15162 20852 15399
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20812 14884 20864 14890
rect 20812 14826 20864 14832
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20732 14521 20760 14554
rect 20718 14512 20774 14521
rect 20718 14447 20774 14456
rect 20720 14340 20772 14346
rect 20720 14282 20772 14288
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20732 13190 20760 14282
rect 20824 14278 20852 14826
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20732 12730 20760 12786
rect 20640 12702 20760 12730
rect 20640 12306 20668 12702
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20732 12238 20760 12582
rect 20824 12442 20852 14214
rect 20916 13802 20944 14758
rect 21008 13938 21036 16748
rect 21100 16046 21128 17088
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 21192 14482 21220 14894
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 21192 13802 21220 14418
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 21180 13796 21232 13802
rect 21180 13738 21232 13744
rect 21192 12646 21220 13738
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 21192 12306 21220 12582
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 20916 11898 20944 12038
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20916 11558 20944 11834
rect 21008 11762 21036 12038
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 19904 8588 20024 8616
rect 19904 8362 19932 8588
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19616 8356 19668 8362
rect 19616 8298 19668 8304
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19628 7886 19656 8298
rect 19996 7886 20024 8366
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19248 7812 19300 7818
rect 19248 7754 19300 7760
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18602 3904 18658 3913
rect 18602 3839 18658 3848
rect 18616 3398 18644 3839
rect 19076 3602 19104 7346
rect 19260 6662 19288 7754
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19260 5642 19288 6598
rect 19352 6322 19380 7686
rect 19444 6798 19472 7754
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19996 7478 20024 7822
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 20088 7324 20116 8774
rect 19996 7296 20116 7324
rect 19996 7206 20024 7296
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6458 20024 6666
rect 20180 6458 20208 9658
rect 20640 9586 20668 10406
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20824 9450 20852 11018
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21008 10674 21036 10746
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 21008 10198 21036 10610
rect 21192 10606 21220 12242
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 20996 10192 21048 10198
rect 20996 10134 21048 10140
rect 21192 10130 21220 10542
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 21284 10062 21312 14214
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20732 6458 20760 9318
rect 21376 9178 21404 17206
rect 21468 15473 21496 19178
rect 21652 18154 21680 25774
rect 22572 22030 22600 31726
rect 23308 29714 23336 35022
rect 23478 34983 23534 34992
rect 23584 34746 23612 35634
rect 23676 35018 23704 35770
rect 23756 35692 23808 35698
rect 23756 35634 23808 35640
rect 23768 35601 23796 35634
rect 23754 35592 23810 35601
rect 23754 35527 23810 35536
rect 23848 35080 23900 35086
rect 23848 35022 23900 35028
rect 23664 35012 23716 35018
rect 23664 34954 23716 34960
rect 23480 34740 23532 34746
rect 23480 34682 23532 34688
rect 23572 34740 23624 34746
rect 23572 34682 23624 34688
rect 23492 34610 23520 34682
rect 23480 34604 23532 34610
rect 23480 34546 23532 34552
rect 23492 34202 23520 34546
rect 23676 34406 23704 34954
rect 23664 34400 23716 34406
rect 23664 34342 23716 34348
rect 23480 34196 23532 34202
rect 23480 34138 23532 34144
rect 23860 34134 23888 35022
rect 24044 34762 24072 35770
rect 24216 35488 24268 35494
rect 24216 35430 24268 35436
rect 23952 34734 24072 34762
rect 23952 34678 23980 34734
rect 24228 34678 24256 35430
rect 24320 34762 24348 37742
rect 24400 35760 24452 35766
rect 24400 35702 24452 35708
rect 24412 35329 24440 35702
rect 24596 35698 24624 38626
rect 24872 38554 24900 38694
rect 24860 38548 24912 38554
rect 24860 38490 24912 38496
rect 24674 38448 24730 38457
rect 24674 38383 24730 38392
rect 24688 37466 24716 38383
rect 24768 37868 24820 37874
rect 24768 37810 24820 37816
rect 24780 37466 24808 37810
rect 24676 37460 24728 37466
rect 24676 37402 24728 37408
rect 24768 37460 24820 37466
rect 24768 37402 24820 37408
rect 25056 37074 25084 39374
rect 25148 37754 25176 50390
rect 25412 50380 25464 50386
rect 25412 50322 25464 50328
rect 25320 43648 25372 43654
rect 25320 43590 25372 43596
rect 25228 39840 25280 39846
rect 25228 39782 25280 39788
rect 25240 39438 25268 39782
rect 25332 39506 25360 43590
rect 25424 43382 25452 50322
rect 25412 43376 25464 43382
rect 25412 43318 25464 43324
rect 25424 42362 25452 43318
rect 25412 42356 25464 42362
rect 25412 42298 25464 42304
rect 25608 42294 25636 53178
rect 25700 53106 25728 55270
rect 26620 55270 26846 55298
rect 26620 53242 26648 55270
rect 26790 55200 26846 55270
rect 27986 55298 28042 56000
rect 27986 55270 28304 55298
rect 27986 55200 28042 55270
rect 26608 53236 26660 53242
rect 26608 53178 26660 53184
rect 28276 53106 28304 55270
rect 29182 55200 29238 56000
rect 30378 55298 30434 56000
rect 31574 55298 31630 56000
rect 30378 55270 30696 55298
rect 30378 55200 30434 55270
rect 29196 53242 29224 55200
rect 29184 53236 29236 53242
rect 29184 53178 29236 53184
rect 30668 53106 30696 55270
rect 31574 55270 31708 55298
rect 31574 55200 31630 55270
rect 31680 53802 31708 55270
rect 32770 55200 32826 56000
rect 33966 55298 34022 56000
rect 35162 55298 35218 56000
rect 36358 55298 36414 56000
rect 37554 55298 37610 56000
rect 38750 55298 38806 56000
rect 33966 55270 34284 55298
rect 33966 55200 34022 55270
rect 31680 53774 31800 53802
rect 31772 53242 31800 53774
rect 31760 53236 31812 53242
rect 31760 53178 31812 53184
rect 32220 53168 32272 53174
rect 32220 53110 32272 53116
rect 25688 53100 25740 53106
rect 25688 53042 25740 53048
rect 28264 53100 28316 53106
rect 28264 53042 28316 53048
rect 30656 53100 30708 53106
rect 30656 53042 30708 53048
rect 25700 52698 25728 53042
rect 26700 52964 26752 52970
rect 26700 52906 26752 52912
rect 25964 52896 26016 52902
rect 25964 52838 26016 52844
rect 25688 52692 25740 52698
rect 25688 52634 25740 52640
rect 25780 42832 25832 42838
rect 25780 42774 25832 42780
rect 25596 42288 25648 42294
rect 25596 42230 25648 42236
rect 25412 41540 25464 41546
rect 25412 41482 25464 41488
rect 25424 39846 25452 41482
rect 25792 41002 25820 42774
rect 25872 42764 25924 42770
rect 25872 42706 25924 42712
rect 25884 41682 25912 42706
rect 25872 41676 25924 41682
rect 25872 41618 25924 41624
rect 25780 40996 25832 41002
rect 25780 40938 25832 40944
rect 25792 40497 25820 40938
rect 25872 40928 25924 40934
rect 25872 40870 25924 40876
rect 25778 40488 25834 40497
rect 25778 40423 25834 40432
rect 25504 40384 25556 40390
rect 25504 40326 25556 40332
rect 25596 40384 25648 40390
rect 25596 40326 25648 40332
rect 25516 40186 25544 40326
rect 25504 40180 25556 40186
rect 25504 40122 25556 40128
rect 25412 39840 25464 39846
rect 25412 39782 25464 39788
rect 25320 39500 25372 39506
rect 25320 39442 25372 39448
rect 25228 39432 25280 39438
rect 25228 39374 25280 39380
rect 25332 39370 25360 39442
rect 25320 39364 25372 39370
rect 25320 39306 25372 39312
rect 25228 39296 25280 39302
rect 25228 39238 25280 39244
rect 25240 38214 25268 39238
rect 25332 38758 25360 39306
rect 25320 38752 25372 38758
rect 25320 38694 25372 38700
rect 25228 38208 25280 38214
rect 25228 38150 25280 38156
rect 25424 37874 25452 39782
rect 25504 38752 25556 38758
rect 25504 38694 25556 38700
rect 25412 37868 25464 37874
rect 25412 37810 25464 37816
rect 25148 37726 25360 37754
rect 25228 37664 25280 37670
rect 25228 37606 25280 37612
rect 25240 37262 25268 37606
rect 25228 37256 25280 37262
rect 25228 37198 25280 37204
rect 25056 37046 25268 37074
rect 24676 36576 24728 36582
rect 24676 36518 24728 36524
rect 24584 35692 24636 35698
rect 24584 35634 24636 35640
rect 24398 35320 24454 35329
rect 24398 35255 24454 35264
rect 24320 34734 24624 34762
rect 23940 34672 23992 34678
rect 23940 34614 23992 34620
rect 24216 34672 24268 34678
rect 24216 34614 24268 34620
rect 24228 34406 24256 34614
rect 24308 34604 24360 34610
rect 24308 34546 24360 34552
rect 24216 34400 24268 34406
rect 24216 34342 24268 34348
rect 24228 34202 24256 34342
rect 24216 34196 24268 34202
rect 24216 34138 24268 34144
rect 23848 34128 23900 34134
rect 23848 34070 23900 34076
rect 24214 34096 24270 34105
rect 24214 34031 24270 34040
rect 24228 33658 24256 34031
rect 24032 33652 24084 33658
rect 24032 33594 24084 33600
rect 24216 33652 24268 33658
rect 24216 33594 24268 33600
rect 23480 33516 23532 33522
rect 23480 33458 23532 33464
rect 23492 33114 23520 33458
rect 23480 33108 23532 33114
rect 23480 33050 23532 33056
rect 24044 32774 24072 33594
rect 24032 32768 24084 32774
rect 24032 32710 24084 32716
rect 24044 32570 24072 32710
rect 24032 32564 24084 32570
rect 24032 32506 24084 32512
rect 23296 29708 23348 29714
rect 23296 29650 23348 29656
rect 22744 29504 22796 29510
rect 22744 29446 22796 29452
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22284 21956 22336 21962
rect 22284 21898 22336 21904
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22112 21350 22140 21830
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 22204 20466 22232 21830
rect 22296 21622 22324 21898
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22296 20890 22324 21558
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22388 21010 22416 21286
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22296 20862 22416 20890
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 21916 19984 21968 19990
rect 21916 19926 21968 19932
rect 21928 19802 21956 19926
rect 21928 19774 22140 19802
rect 22112 19718 22140 19774
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22296 19514 22324 19722
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22008 18216 22060 18222
rect 22008 18158 22060 18164
rect 21640 18148 21692 18154
rect 21640 18090 21692 18096
rect 21652 17678 21680 18090
rect 22020 17746 22048 18158
rect 22388 17762 22416 20862
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 22468 19440 22520 19446
rect 22468 19382 22520 19388
rect 22480 18834 22508 19382
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22480 17882 22508 18226
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22008 17740 22060 17746
rect 22388 17734 22508 17762
rect 22008 17682 22060 17688
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21640 16516 21692 16522
rect 21640 16458 21692 16464
rect 21652 15706 21680 16458
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21744 15638 21772 17478
rect 21836 17202 21864 17478
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21836 15502 21864 16934
rect 22020 16046 22048 17682
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22204 16794 22232 17070
rect 22388 16794 22416 17138
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 22204 16538 22232 16730
rect 22112 16250 22140 16526
rect 22204 16510 22324 16538
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22008 16040 22060 16046
rect 22008 15982 22060 15988
rect 21824 15496 21876 15502
rect 21454 15464 21510 15473
rect 21824 15438 21876 15444
rect 21454 15399 21510 15408
rect 22020 15178 22048 15982
rect 22204 15434 22232 16390
rect 22296 15570 22324 16510
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 22020 15150 22140 15178
rect 21914 15056 21970 15065
rect 21914 14991 21970 15000
rect 21640 14884 21692 14890
rect 21640 14826 21692 14832
rect 21652 14414 21680 14826
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21744 14006 21772 14214
rect 21836 14074 21864 14214
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21732 14000 21784 14006
rect 21732 13942 21784 13948
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21468 12850 21496 13874
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21468 12714 21496 12786
rect 21456 12708 21508 12714
rect 21456 12650 21508 12656
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 21468 9450 21496 11018
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21456 9444 21508 9450
rect 21456 9386 21508 9392
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21560 9042 21588 9862
rect 21548 9036 21600 9042
rect 21548 8978 21600 8984
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21284 7750 21312 8366
rect 21376 8362 21404 8774
rect 21364 8356 21416 8362
rect 21364 8298 21416 8304
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 21284 4690 21312 7686
rect 21364 7404 21416 7410
rect 21364 7346 21416 7352
rect 21376 7002 21404 7346
rect 21364 6996 21416 7002
rect 21364 6938 21416 6944
rect 21468 6458 21496 8910
rect 21560 8362 21588 8978
rect 21652 8974 21680 10202
rect 21928 9382 21956 14991
rect 22112 14006 22140 15150
rect 22296 14482 22324 15506
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 22112 12850 22140 13942
rect 22296 13530 22324 14418
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22296 12918 22324 13466
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22112 10130 22140 12786
rect 22480 12730 22508 17734
rect 22572 17678 22600 19450
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22664 17270 22692 18022
rect 22652 17264 22704 17270
rect 22652 17206 22704 17212
rect 22756 17218 22784 29446
rect 23940 27532 23992 27538
rect 23940 27474 23992 27480
rect 23952 26858 23980 27474
rect 23940 26852 23992 26858
rect 23940 26794 23992 26800
rect 23664 26580 23716 26586
rect 23664 26522 23716 26528
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23400 23526 23428 24210
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23388 23520 23440 23526
rect 23388 23462 23440 23468
rect 23400 23322 23428 23462
rect 22928 23316 22980 23322
rect 22928 23258 22980 23264
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 22940 22778 22968 23258
rect 23584 23118 23612 24006
rect 23676 23730 23704 26522
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 23020 22976 23072 22982
rect 23020 22918 23072 22924
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23756 22976 23808 22982
rect 23756 22918 23808 22924
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 22940 22234 22968 22714
rect 22928 22228 22980 22234
rect 22928 22170 22980 22176
rect 22940 22094 22968 22170
rect 23032 22166 23060 22918
rect 23492 22642 23520 22918
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23492 22166 23520 22374
rect 23020 22160 23072 22166
rect 23020 22102 23072 22108
rect 23480 22160 23532 22166
rect 23480 22102 23532 22108
rect 22848 22066 22968 22094
rect 22848 21350 22876 22066
rect 23110 21856 23166 21865
rect 23110 21791 23166 21800
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 22848 19922 22876 20266
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 23124 17660 23152 21791
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 23308 21146 23336 21286
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 23204 18284 23256 18290
rect 23204 18226 23256 18232
rect 23216 17814 23244 18226
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 23124 17632 23244 17660
rect 22756 17190 22876 17218
rect 22652 17060 22704 17066
rect 22652 17002 22704 17008
rect 22664 16522 22692 17002
rect 22652 16516 22704 16522
rect 22652 16458 22704 16464
rect 22848 16182 22876 17190
rect 23110 16824 23166 16833
rect 23110 16759 23112 16768
rect 23164 16759 23166 16768
rect 23112 16730 23164 16736
rect 22836 16176 22888 16182
rect 22836 16118 22888 16124
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 22756 15162 22784 16050
rect 22836 15972 22888 15978
rect 22836 15914 22888 15920
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22572 14822 22600 14962
rect 22848 14958 22876 15914
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22560 14816 22612 14822
rect 22560 14758 22612 14764
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22296 12702 22508 12730
rect 22190 12336 22246 12345
rect 22190 12271 22246 12280
rect 22204 12170 22232 12271
rect 22192 12164 22244 12170
rect 22192 12106 22244 12112
rect 22204 12073 22232 12106
rect 22190 12064 22246 12073
rect 22190 11999 22246 12008
rect 22296 11830 22324 12702
rect 22572 12442 22600 12854
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22664 12288 22692 13670
rect 22744 12708 22796 12714
rect 22744 12650 22796 12656
rect 22572 12260 22692 12288
rect 22468 12164 22520 12170
rect 22468 12106 22520 12112
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22100 10124 22152 10130
rect 22100 10066 22152 10072
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22112 9586 22140 9862
rect 22204 9586 22232 11494
rect 22296 11150 22324 11630
rect 22388 11626 22416 12038
rect 22376 11620 22428 11626
rect 22376 11562 22428 11568
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22296 10062 22324 11086
rect 22480 10656 22508 12106
rect 22388 10628 22508 10656
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 21916 9376 21968 9382
rect 21916 9318 21968 9324
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 22296 8498 22324 9998
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 21548 8356 21600 8362
rect 21548 8298 21600 8304
rect 22008 8356 22060 8362
rect 22008 8298 22060 8304
rect 22020 7410 22048 8298
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 21640 7200 21692 7206
rect 21640 7142 21692 7148
rect 21652 6798 21680 7142
rect 22204 7002 22232 7482
rect 22296 7478 22324 8434
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22296 7342 22324 7414
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22192 6996 22244 7002
rect 22192 6938 22244 6944
rect 22296 6866 22324 7278
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 22388 6662 22416 10628
rect 22468 10532 22520 10538
rect 22468 10474 22520 10480
rect 22480 10062 22508 10474
rect 22572 10470 22600 12260
rect 22652 11824 22704 11830
rect 22652 11766 22704 11772
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22572 9994 22600 10406
rect 22560 9988 22612 9994
rect 22560 9930 22612 9936
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22572 7886 22600 8774
rect 22664 8650 22692 11766
rect 22756 10674 22784 12650
rect 22848 12102 22876 14894
rect 23216 14890 23244 17632
rect 23204 14884 23256 14890
rect 23204 14826 23256 14832
rect 23020 12912 23072 12918
rect 23018 12880 23020 12889
rect 23072 12880 23074 12889
rect 23018 12815 23074 12824
rect 23204 12368 23256 12374
rect 23204 12310 23256 12316
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 22836 11688 22888 11694
rect 22836 11630 22888 11636
rect 22848 11082 22876 11630
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 22836 10736 22888 10742
rect 22836 10678 22888 10684
rect 22744 10668 22796 10674
rect 22744 10610 22796 10616
rect 22848 9722 22876 10678
rect 23032 10606 23060 12038
rect 23020 10600 23072 10606
rect 23020 10542 23072 10548
rect 22836 9716 22888 9722
rect 22836 9658 22888 9664
rect 23112 9512 23164 9518
rect 23112 9454 23164 9460
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22664 8622 22784 8650
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22664 7954 22692 8434
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22468 7880 22520 7886
rect 22468 7822 22520 7828
rect 22560 7880 22612 7886
rect 22560 7822 22612 7828
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21468 5846 21496 6394
rect 21456 5840 21508 5846
rect 21456 5782 21508 5788
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18524 3058 18552 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17880 800 17908 2382
rect 18248 800 18276 2994
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18616 800 18644 2382
rect 18984 800 19012 2790
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19352 800 19380 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19720 870 19840 898
rect 19720 800 19748 870
rect 15396 734 15608 762
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 19812 762 19840 870
rect 19996 762 20024 3470
rect 22112 3466 22140 4082
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 20088 800 20116 2790
rect 20456 800 20484 2790
rect 20812 2576 20864 2582
rect 20812 2518 20864 2524
rect 20824 800 20852 2518
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 21192 800 21220 2382
rect 21560 800 21588 2790
rect 22204 2514 22232 6598
rect 22480 6186 22508 7822
rect 22468 6180 22520 6186
rect 22468 6122 22520 6128
rect 22560 4548 22612 4554
rect 22560 4490 22612 4496
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 21928 800 21956 2382
rect 22296 800 22324 2790
rect 22572 2446 22600 4490
rect 22756 3466 22784 8622
rect 22848 6662 22876 8978
rect 23124 8838 23152 9454
rect 23216 8974 23244 12310
rect 23308 9568 23336 21082
rect 23492 20398 23520 22102
rect 23768 22030 23796 22918
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23584 21690 23612 21830
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 23676 21554 23704 21830
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23570 21040 23626 21049
rect 23570 20975 23626 20984
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23480 19440 23532 19446
rect 23480 19382 23532 19388
rect 23492 18358 23520 19382
rect 23584 19174 23612 20975
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23860 20602 23888 20878
rect 23848 20596 23900 20602
rect 23848 20538 23900 20544
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23676 18766 23704 19110
rect 23940 18828 23992 18834
rect 23940 18770 23992 18776
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23400 16046 23428 17614
rect 23492 16182 23520 18294
rect 23848 17808 23900 17814
rect 23848 17750 23900 17756
rect 23860 17542 23888 17750
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23952 17202 23980 18770
rect 24044 17746 24072 32506
rect 24320 29646 24348 34546
rect 24596 34542 24624 34734
rect 24584 34536 24636 34542
rect 24584 34478 24636 34484
rect 24688 34202 24716 36518
rect 25240 36378 25268 37046
rect 25332 36768 25360 37726
rect 25516 37126 25544 38694
rect 25608 37874 25636 40326
rect 25688 40112 25740 40118
rect 25688 40054 25740 40060
rect 25700 39642 25728 40054
rect 25780 39976 25832 39982
rect 25780 39918 25832 39924
rect 25688 39636 25740 39642
rect 25688 39578 25740 39584
rect 25688 38004 25740 38010
rect 25688 37946 25740 37952
rect 25596 37868 25648 37874
rect 25596 37810 25648 37816
rect 25596 37664 25648 37670
rect 25596 37606 25648 37612
rect 25608 37126 25636 37606
rect 25504 37120 25556 37126
rect 25504 37062 25556 37068
rect 25596 37120 25648 37126
rect 25596 37062 25648 37068
rect 25412 36780 25464 36786
rect 25332 36740 25412 36768
rect 25412 36722 25464 36728
rect 25424 36553 25452 36722
rect 25410 36544 25466 36553
rect 25410 36479 25466 36488
rect 25516 36417 25544 37062
rect 25502 36408 25558 36417
rect 25136 36372 25188 36378
rect 25136 36314 25188 36320
rect 25228 36372 25280 36378
rect 25502 36343 25558 36352
rect 25228 36314 25280 36320
rect 25044 35760 25096 35766
rect 25042 35728 25044 35737
rect 25096 35728 25098 35737
rect 24860 35692 24912 35698
rect 25042 35663 25098 35672
rect 24860 35634 24912 35640
rect 24676 34196 24728 34202
rect 24676 34138 24728 34144
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 24584 33380 24636 33386
rect 24584 33322 24636 33328
rect 24596 32502 24624 33322
rect 24584 32496 24636 32502
rect 24584 32438 24636 32444
rect 24308 29640 24360 29646
rect 24308 29582 24360 29588
rect 24400 29164 24452 29170
rect 24400 29106 24452 29112
rect 24412 27606 24440 29106
rect 24584 28552 24636 28558
rect 24584 28494 24636 28500
rect 24400 27600 24452 27606
rect 24400 27542 24452 27548
rect 24412 27130 24440 27542
rect 24400 27124 24452 27130
rect 24400 27066 24452 27072
rect 24596 26382 24624 28494
rect 24676 28484 24728 28490
rect 24676 28426 24728 28432
rect 24688 28218 24716 28426
rect 24676 28212 24728 28218
rect 24676 28154 24728 28160
rect 24584 26376 24636 26382
rect 24584 26318 24636 26324
rect 24308 24608 24360 24614
rect 24308 24550 24360 24556
rect 24320 23662 24348 24550
rect 24584 24404 24636 24410
rect 24584 24346 24636 24352
rect 24596 23798 24624 24346
rect 24584 23792 24636 23798
rect 24584 23734 24636 23740
rect 24308 23656 24360 23662
rect 24308 23598 24360 23604
rect 24320 22778 24348 23598
rect 24400 23588 24452 23594
rect 24452 23548 24532 23576
rect 24400 23530 24452 23536
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 24308 22228 24360 22234
rect 24308 22170 24360 22176
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24228 19378 24256 20334
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24136 17882 24164 19314
rect 24124 17876 24176 17882
rect 24124 17818 24176 17824
rect 24032 17740 24084 17746
rect 24032 17682 24084 17688
rect 24032 17536 24084 17542
rect 24030 17504 24032 17513
rect 24124 17536 24176 17542
rect 24084 17504 24086 17513
rect 24124 17478 24176 17484
rect 24030 17439 24086 17448
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23756 17060 23808 17066
rect 23756 17002 23808 17008
rect 23768 16794 23796 17002
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23768 16590 23796 16730
rect 23756 16584 23808 16590
rect 23756 16526 23808 16532
rect 23480 16176 23532 16182
rect 23480 16118 23532 16124
rect 23388 16040 23440 16046
rect 23388 15982 23440 15988
rect 24044 15434 24072 16934
rect 24136 16794 24164 17478
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 24216 16584 24268 16590
rect 24216 16526 24268 16532
rect 24228 15910 24256 16526
rect 24124 15904 24176 15910
rect 24124 15846 24176 15852
rect 24216 15904 24268 15910
rect 24216 15846 24268 15852
rect 24032 15428 24084 15434
rect 24032 15370 24084 15376
rect 24136 15366 24164 15846
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 23676 15026 23704 15302
rect 23756 15088 23808 15094
rect 23754 15056 23756 15065
rect 23808 15056 23810 15065
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23664 15020 23716 15026
rect 23754 14991 23810 15000
rect 23664 14962 23716 14968
rect 23400 14074 23428 14962
rect 23848 14952 23900 14958
rect 23848 14894 23900 14900
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23768 14074 23796 14554
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23400 10674 23428 13262
rect 23676 12238 23704 13466
rect 23768 13394 23796 14010
rect 23860 13954 23888 14894
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23952 14074 23980 14758
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 23860 13926 23980 13954
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23860 12782 23888 13926
rect 23952 13870 23980 13926
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 24032 13456 24084 13462
rect 24032 13398 24084 13404
rect 24044 12850 24072 13398
rect 24136 13190 24164 14418
rect 24228 14414 24256 15846
rect 24320 14482 24348 22170
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24412 20602 24440 20878
rect 24400 20596 24452 20602
rect 24400 20538 24452 20544
rect 24412 20505 24440 20538
rect 24398 20496 24454 20505
rect 24398 20431 24454 20440
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24412 16250 24440 17274
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24308 14476 24360 14482
rect 24308 14418 24360 14424
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24228 13938 24256 14350
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24504 13870 24532 23548
rect 24596 23186 24624 23734
rect 24584 23180 24636 23186
rect 24584 23122 24636 23128
rect 24780 22234 24808 33594
rect 24872 32570 24900 35634
rect 25044 34944 25096 34950
rect 25044 34886 25096 34892
rect 24952 33856 25004 33862
rect 24952 33798 25004 33804
rect 24964 33522 24992 33798
rect 24952 33516 25004 33522
rect 24952 33458 25004 33464
rect 24860 32564 24912 32570
rect 24860 32506 24912 32512
rect 24952 32292 25004 32298
rect 24952 32234 25004 32240
rect 24860 32224 24912 32230
rect 24860 32166 24912 32172
rect 24872 31686 24900 32166
rect 24964 32026 24992 32234
rect 24952 32020 25004 32026
rect 24952 31962 25004 31968
rect 24964 31929 24992 31962
rect 24950 31920 25006 31929
rect 24950 31855 25006 31864
rect 25056 31754 25084 34886
rect 25148 33454 25176 36314
rect 25240 36174 25268 36314
rect 25228 36168 25280 36174
rect 25228 36110 25280 36116
rect 25412 36100 25464 36106
rect 25516 36088 25544 36343
rect 25596 36168 25648 36174
rect 25464 36060 25544 36088
rect 25594 36136 25596 36145
rect 25648 36136 25650 36145
rect 25594 36071 25650 36080
rect 25412 36042 25464 36048
rect 25596 36032 25648 36038
rect 25596 35974 25648 35980
rect 25320 35828 25372 35834
rect 25320 35770 25372 35776
rect 25332 34678 25360 35770
rect 25608 35630 25636 35974
rect 25596 35624 25648 35630
rect 25596 35566 25648 35572
rect 25596 35148 25648 35154
rect 25700 35136 25728 37946
rect 25648 35108 25728 35136
rect 25596 35090 25648 35096
rect 25700 34746 25728 35108
rect 25792 34746 25820 39918
rect 25884 38758 25912 40870
rect 25976 39506 26004 52838
rect 26056 52488 26108 52494
rect 26056 52430 26108 52436
rect 26068 52154 26096 52430
rect 26056 52148 26108 52154
rect 26056 52090 26108 52096
rect 26068 51270 26096 52090
rect 26056 51264 26108 51270
rect 26056 51206 26108 51212
rect 26068 43382 26096 51206
rect 26424 45552 26476 45558
rect 26424 45494 26476 45500
rect 26436 44402 26464 45494
rect 26424 44396 26476 44402
rect 26424 44338 26476 44344
rect 26056 43376 26108 43382
rect 26056 43318 26108 43324
rect 26068 42906 26096 43318
rect 26056 42900 26108 42906
rect 26056 42842 26108 42848
rect 26068 42294 26096 42842
rect 26436 42770 26464 44338
rect 26608 43648 26660 43654
rect 26608 43590 26660 43596
rect 26424 42764 26476 42770
rect 26424 42706 26476 42712
rect 26240 42696 26292 42702
rect 26240 42638 26292 42644
rect 26056 42288 26108 42294
rect 26056 42230 26108 42236
rect 26068 41721 26096 42230
rect 26054 41712 26110 41721
rect 26054 41647 26110 41656
rect 26148 41676 26200 41682
rect 25964 39500 26016 39506
rect 25964 39442 26016 39448
rect 26068 39386 26096 41647
rect 26148 41618 26200 41624
rect 26160 40769 26188 41618
rect 26252 41313 26280 42638
rect 26332 42628 26384 42634
rect 26332 42570 26384 42576
rect 26344 42226 26372 42570
rect 26332 42220 26384 42226
rect 26332 42162 26384 42168
rect 26238 41304 26294 41313
rect 26344 41274 26372 42162
rect 26238 41239 26294 41248
rect 26332 41268 26384 41274
rect 26332 41210 26384 41216
rect 26436 41138 26464 42706
rect 26516 42016 26568 42022
rect 26516 41958 26568 41964
rect 26528 41585 26556 41958
rect 26514 41576 26570 41585
rect 26514 41511 26570 41520
rect 26516 41268 26568 41274
rect 26516 41210 26568 41216
rect 26424 41132 26476 41138
rect 26424 41074 26476 41080
rect 26528 41018 26556 41210
rect 26344 40990 26556 41018
rect 26146 40760 26202 40769
rect 26146 40695 26202 40704
rect 26146 40624 26202 40633
rect 26146 40559 26202 40568
rect 26160 40526 26188 40559
rect 26148 40520 26200 40526
rect 26148 40462 26200 40468
rect 26148 40384 26200 40390
rect 26148 40326 26200 40332
rect 26160 40050 26188 40326
rect 26240 40180 26292 40186
rect 26240 40122 26292 40128
rect 26148 40044 26200 40050
rect 26148 39986 26200 39992
rect 26252 39574 26280 40122
rect 26344 40050 26372 40990
rect 26516 40928 26568 40934
rect 26516 40870 26568 40876
rect 26528 40526 26556 40870
rect 26424 40520 26476 40526
rect 26424 40462 26476 40468
rect 26516 40520 26568 40526
rect 26516 40462 26568 40468
rect 26436 40089 26464 40462
rect 26422 40080 26478 40089
rect 26332 40044 26384 40050
rect 26422 40015 26478 40024
rect 26516 40044 26568 40050
rect 26332 39986 26384 39992
rect 26516 39986 26568 39992
rect 26240 39568 26292 39574
rect 26240 39510 26292 39516
rect 25976 39358 26096 39386
rect 26148 39432 26200 39438
rect 26148 39374 26200 39380
rect 25872 38752 25924 38758
rect 25872 38694 25924 38700
rect 25872 38208 25924 38214
rect 25872 38150 25924 38156
rect 25884 37652 25912 38150
rect 25976 37806 26004 39358
rect 26056 39296 26108 39302
rect 26056 39238 26108 39244
rect 26068 39098 26096 39238
rect 26160 39098 26188 39374
rect 26056 39092 26108 39098
rect 26056 39034 26108 39040
rect 26148 39092 26200 39098
rect 26148 39034 26200 39040
rect 26054 38856 26110 38865
rect 26054 38791 26110 38800
rect 26068 38758 26096 38791
rect 26056 38752 26108 38758
rect 26056 38694 26108 38700
rect 26240 38752 26292 38758
rect 26240 38694 26292 38700
rect 26252 38486 26280 38694
rect 26240 38480 26292 38486
rect 26240 38422 26292 38428
rect 26056 38276 26108 38282
rect 26056 38218 26108 38224
rect 26068 37874 26096 38218
rect 26056 37868 26108 37874
rect 26056 37810 26108 37816
rect 25964 37800 26016 37806
rect 25964 37742 26016 37748
rect 26240 37732 26292 37738
rect 26240 37674 26292 37680
rect 26148 37664 26200 37670
rect 25884 37624 26004 37652
rect 25872 36780 25924 36786
rect 25872 36722 25924 36728
rect 25884 36689 25912 36722
rect 25870 36680 25926 36689
rect 25870 36615 25926 36624
rect 25976 36174 26004 37624
rect 26252 37641 26280 37674
rect 26148 37606 26200 37612
rect 26238 37632 26294 37641
rect 26054 37360 26110 37369
rect 26054 37295 26110 37304
rect 26068 37194 26096 37295
rect 26056 37188 26108 37194
rect 26056 37130 26108 37136
rect 26056 36780 26108 36786
rect 26056 36722 26108 36728
rect 25964 36168 26016 36174
rect 25964 36110 26016 36116
rect 25964 36032 26016 36038
rect 25964 35974 26016 35980
rect 25976 35494 26004 35974
rect 25872 35488 25924 35494
rect 25872 35430 25924 35436
rect 25964 35488 26016 35494
rect 25964 35430 26016 35436
rect 25884 35086 25912 35430
rect 25872 35080 25924 35086
rect 25872 35022 25924 35028
rect 25964 35012 26016 35018
rect 25964 34954 26016 34960
rect 25976 34762 26004 34954
rect 25688 34740 25740 34746
rect 25688 34682 25740 34688
rect 25780 34740 25832 34746
rect 25780 34682 25832 34688
rect 25884 34734 26004 34762
rect 25320 34672 25372 34678
rect 25792 34626 25820 34682
rect 25320 34614 25372 34620
rect 25504 34604 25556 34610
rect 25504 34546 25556 34552
rect 25608 34598 25820 34626
rect 25410 34504 25466 34513
rect 25410 34439 25466 34448
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 25136 33448 25188 33454
rect 25136 33390 25188 33396
rect 25332 33386 25360 33934
rect 25424 33522 25452 34439
rect 25412 33516 25464 33522
rect 25412 33458 25464 33464
rect 25320 33380 25372 33386
rect 25320 33322 25372 33328
rect 25332 32978 25360 33322
rect 25320 32972 25372 32978
rect 25320 32914 25372 32920
rect 25056 31726 25176 31754
rect 24860 31680 24912 31686
rect 24860 31622 24912 31628
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 24872 22778 24900 25230
rect 25044 25152 25096 25158
rect 25044 25094 25096 25100
rect 25056 24886 25084 25094
rect 25044 24880 25096 24886
rect 25044 24822 25096 24828
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 25056 24206 25084 24686
rect 25044 24200 25096 24206
rect 25044 24142 25096 24148
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 24768 22228 24820 22234
rect 24768 22170 24820 22176
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24584 21616 24636 21622
rect 24584 21558 24636 21564
rect 24596 20942 24624 21558
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 24596 19446 24624 20878
rect 24584 19440 24636 19446
rect 24584 19382 24636 19388
rect 24688 18766 24716 21830
rect 24780 20058 24808 21966
rect 25056 21622 25084 22170
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 25148 21350 25176 31726
rect 25424 28762 25452 33458
rect 25516 31346 25544 34546
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 25412 28756 25464 28762
rect 25412 28698 25464 28704
rect 25228 28416 25280 28422
rect 25228 28358 25280 28364
rect 25240 28150 25268 28358
rect 25228 28144 25280 28150
rect 25228 28086 25280 28092
rect 25240 28014 25268 28086
rect 25228 28008 25280 28014
rect 25228 27950 25280 27956
rect 25240 27470 25268 27950
rect 25228 27464 25280 27470
rect 25228 27406 25280 27412
rect 25424 27418 25452 28698
rect 25240 27130 25268 27406
rect 25424 27390 25544 27418
rect 25412 27328 25464 27334
rect 25412 27270 25464 27276
rect 25228 27124 25280 27130
rect 25228 27066 25280 27072
rect 25424 27062 25452 27270
rect 25412 27056 25464 27062
rect 25412 26998 25464 27004
rect 25412 25900 25464 25906
rect 25412 25842 25464 25848
rect 25228 25696 25280 25702
rect 25228 25638 25280 25644
rect 25240 24138 25268 25638
rect 25228 24132 25280 24138
rect 25228 24074 25280 24080
rect 25320 24132 25372 24138
rect 25320 24074 25372 24080
rect 25332 23730 25360 24074
rect 25424 23866 25452 25842
rect 25412 23860 25464 23866
rect 25412 23802 25464 23808
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 25516 23662 25544 27390
rect 25412 23656 25464 23662
rect 25412 23598 25464 23604
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 24860 20528 24912 20534
rect 24860 20470 24912 20476
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24872 19922 24900 20470
rect 25148 20466 25176 20742
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 25320 20460 25372 20466
rect 25320 20402 25372 20408
rect 25044 20392 25096 20398
rect 25096 20340 25176 20346
rect 25044 20334 25176 20340
rect 25056 20318 25176 20334
rect 25148 19922 25176 20318
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 25136 19916 25188 19922
rect 25136 19858 25188 19864
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24872 18290 24900 19858
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 25056 19446 25084 19654
rect 25044 19440 25096 19446
rect 25044 19382 25096 19388
rect 24952 19304 25004 19310
rect 24952 19246 25004 19252
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24964 18086 24992 19246
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24584 17604 24636 17610
rect 24584 17546 24636 17552
rect 24596 16794 24624 17546
rect 24688 17338 24716 17614
rect 24964 17542 24992 18022
rect 25044 17876 25096 17882
rect 25044 17818 25096 17824
rect 25056 17785 25084 17818
rect 25042 17776 25098 17785
rect 25148 17746 25176 19858
rect 25332 18970 25360 20402
rect 25320 18964 25372 18970
rect 25320 18906 25372 18912
rect 25320 18624 25372 18630
rect 25320 18566 25372 18572
rect 25228 18284 25280 18290
rect 25332 18272 25360 18566
rect 25280 18244 25360 18272
rect 25228 18226 25280 18232
rect 25042 17711 25098 17720
rect 25136 17740 25188 17746
rect 25056 17542 25084 17711
rect 25136 17682 25188 17688
rect 25148 17649 25176 17682
rect 25134 17640 25190 17649
rect 25134 17575 25190 17584
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 25044 17536 25096 17542
rect 25044 17478 25096 17484
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24674 17232 24730 17241
rect 24674 17167 24676 17176
rect 24728 17167 24730 17176
rect 24676 17138 24728 17144
rect 24676 17060 24728 17066
rect 24676 17002 24728 17008
rect 24688 16794 24716 17002
rect 24584 16788 24636 16794
rect 24584 16730 24636 16736
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 25042 16688 25098 16697
rect 25148 16658 25176 17575
rect 25424 17270 25452 23598
rect 25516 23186 25544 23598
rect 25504 23180 25556 23186
rect 25504 23122 25556 23128
rect 25608 22094 25636 34598
rect 25884 33946 25912 34734
rect 25964 34672 26016 34678
rect 25964 34614 26016 34620
rect 25792 33918 25912 33946
rect 25792 33114 25820 33918
rect 25872 33856 25924 33862
rect 25872 33798 25924 33804
rect 25884 33454 25912 33798
rect 25872 33448 25924 33454
rect 25872 33390 25924 33396
rect 25780 33108 25832 33114
rect 25780 33050 25832 33056
rect 25884 32434 25912 33390
rect 25872 32428 25924 32434
rect 25872 32370 25924 32376
rect 25884 31754 25912 32370
rect 25976 32026 26004 34614
rect 26068 34134 26096 36722
rect 26160 36650 26188 37606
rect 26238 37567 26294 37576
rect 26240 36780 26292 36786
rect 26240 36722 26292 36728
rect 26148 36644 26200 36650
rect 26148 36586 26200 36592
rect 26160 35698 26188 36586
rect 26148 35692 26200 35698
rect 26148 35634 26200 35640
rect 26148 35556 26200 35562
rect 26148 35498 26200 35504
rect 26160 35465 26188 35498
rect 26146 35456 26202 35465
rect 26146 35391 26202 35400
rect 26252 34678 26280 36722
rect 26344 35018 26372 39986
rect 26424 38344 26476 38350
rect 26424 38286 26476 38292
rect 26436 37398 26464 38286
rect 26424 37392 26476 37398
rect 26424 37334 26476 37340
rect 26528 36961 26556 39986
rect 26620 38962 26648 43590
rect 26712 40186 26740 52906
rect 26976 52896 27028 52902
rect 26976 52838 27028 52844
rect 28080 52896 28132 52902
rect 28080 52838 28132 52844
rect 26792 45892 26844 45898
rect 26792 45834 26844 45840
rect 26804 43382 26832 45834
rect 26884 44736 26936 44742
rect 26884 44678 26936 44684
rect 26896 44402 26924 44678
rect 26884 44396 26936 44402
rect 26884 44338 26936 44344
rect 26792 43376 26844 43382
rect 26792 43318 26844 43324
rect 26792 42560 26844 42566
rect 26792 42502 26844 42508
rect 26804 41750 26832 42502
rect 26792 41744 26844 41750
rect 26792 41686 26844 41692
rect 26884 41608 26936 41614
rect 26884 41550 26936 41556
rect 26896 41414 26924 41550
rect 26804 41386 26924 41414
rect 26700 40180 26752 40186
rect 26700 40122 26752 40128
rect 26804 39386 26832 41386
rect 26884 40520 26936 40526
rect 26884 40462 26936 40468
rect 26896 40390 26924 40462
rect 26884 40384 26936 40390
rect 26884 40326 26936 40332
rect 26896 39545 26924 40326
rect 26882 39536 26938 39545
rect 26882 39471 26938 39480
rect 26712 39358 26832 39386
rect 26988 39370 27016 52838
rect 27160 52488 27212 52494
rect 27160 52430 27212 52436
rect 27172 52086 27200 52430
rect 28092 52086 28120 52838
rect 28276 52698 28304 53042
rect 32128 52964 32180 52970
rect 32128 52906 32180 52912
rect 28724 52896 28776 52902
rect 28724 52838 28776 52844
rect 30104 52896 30156 52902
rect 30104 52838 30156 52844
rect 31208 52896 31260 52902
rect 31208 52838 31260 52844
rect 28264 52692 28316 52698
rect 28264 52634 28316 52640
rect 27160 52080 27212 52086
rect 27160 52022 27212 52028
rect 28080 52080 28132 52086
rect 28080 52022 28132 52028
rect 27896 52012 27948 52018
rect 27896 51954 27948 51960
rect 27620 51808 27672 51814
rect 27620 51750 27672 51756
rect 27436 45076 27488 45082
rect 27436 45018 27488 45024
rect 27448 44470 27476 45018
rect 27068 44464 27120 44470
rect 27068 44406 27120 44412
rect 27436 44464 27488 44470
rect 27436 44406 27488 44412
rect 27080 41414 27108 44406
rect 27448 43790 27476 44406
rect 27436 43784 27488 43790
rect 27436 43726 27488 43732
rect 27252 43376 27304 43382
rect 27252 43318 27304 43324
rect 27264 41614 27292 43318
rect 27436 42084 27488 42090
rect 27436 42026 27488 42032
rect 27252 41608 27304 41614
rect 27252 41550 27304 41556
rect 27252 41472 27304 41478
rect 27252 41414 27304 41420
rect 27080 41386 27200 41414
rect 27068 41132 27120 41138
rect 27068 41074 27120 41080
rect 27080 39438 27108 41074
rect 27068 39432 27120 39438
rect 27068 39374 27120 39380
rect 26976 39364 27028 39370
rect 26608 38956 26660 38962
rect 26608 38898 26660 38904
rect 26608 38344 26660 38350
rect 26606 38312 26608 38321
rect 26660 38312 26662 38321
rect 26606 38247 26662 38256
rect 26608 38004 26660 38010
rect 26608 37946 26660 37952
rect 26514 36952 26570 36961
rect 26514 36887 26570 36896
rect 26424 36372 26476 36378
rect 26424 36314 26476 36320
rect 26436 36174 26464 36314
rect 26424 36168 26476 36174
rect 26424 36110 26476 36116
rect 26436 35698 26464 36110
rect 26424 35692 26476 35698
rect 26424 35634 26476 35640
rect 26332 35012 26384 35018
rect 26332 34954 26384 34960
rect 26240 34672 26292 34678
rect 26160 34620 26240 34626
rect 26160 34614 26292 34620
rect 26160 34598 26280 34614
rect 26056 34128 26108 34134
rect 26056 34070 26108 34076
rect 26160 33114 26188 34598
rect 26436 34406 26464 35634
rect 26516 35556 26568 35562
rect 26516 35498 26568 35504
rect 26528 35222 26556 35498
rect 26516 35216 26568 35222
rect 26516 35158 26568 35164
rect 26516 35080 26568 35086
rect 26516 35022 26568 35028
rect 26424 34400 26476 34406
rect 26424 34342 26476 34348
rect 26332 34060 26384 34066
rect 26332 34002 26384 34008
rect 26344 33538 26372 34002
rect 26528 33998 26556 35022
rect 26516 33992 26568 33998
rect 26516 33934 26568 33940
rect 26516 33584 26568 33590
rect 26344 33522 26464 33538
rect 26516 33526 26568 33532
rect 26240 33516 26292 33522
rect 26240 33458 26292 33464
rect 26344 33516 26476 33522
rect 26344 33510 26424 33516
rect 26148 33108 26200 33114
rect 26148 33050 26200 33056
rect 26252 32910 26280 33458
rect 26240 32904 26292 32910
rect 26240 32846 26292 32852
rect 26252 32434 26280 32846
rect 26344 32774 26372 33510
rect 26424 33458 26476 33464
rect 26424 32972 26476 32978
rect 26424 32914 26476 32920
rect 26332 32768 26384 32774
rect 26332 32710 26384 32716
rect 26240 32428 26292 32434
rect 26240 32370 26292 32376
rect 25964 32020 26016 32026
rect 25964 31962 26016 31968
rect 25976 31754 26004 31962
rect 25688 31748 25740 31754
rect 25688 31690 25740 31696
rect 25792 31726 25912 31754
rect 25964 31748 26016 31754
rect 25700 26926 25728 31690
rect 25792 31278 25820 31726
rect 25964 31690 26016 31696
rect 26148 31680 26200 31686
rect 26148 31622 26200 31628
rect 25872 31408 25924 31414
rect 25872 31350 25924 31356
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 25792 28014 25820 31214
rect 25884 28150 25912 31350
rect 26056 31272 26108 31278
rect 26056 31214 26108 31220
rect 26068 30802 26096 31214
rect 26160 30870 26188 31622
rect 26344 31414 26372 32710
rect 26436 32366 26464 32914
rect 26528 32502 26556 33526
rect 26516 32496 26568 32502
rect 26516 32438 26568 32444
rect 26424 32360 26476 32366
rect 26424 32302 26476 32308
rect 26436 31482 26464 32302
rect 26620 31822 26648 37946
rect 26712 37913 26740 39358
rect 26976 39306 27028 39312
rect 26792 39296 26844 39302
rect 26792 39238 26844 39244
rect 26884 39296 26936 39302
rect 26884 39238 26936 39244
rect 26804 38729 26832 39238
rect 26896 38758 26924 39238
rect 27066 38992 27122 39001
rect 27066 38927 27122 38936
rect 26976 38820 27028 38826
rect 26976 38762 27028 38768
rect 26884 38752 26936 38758
rect 26790 38720 26846 38729
rect 26884 38694 26936 38700
rect 26790 38655 26846 38664
rect 26792 38344 26844 38350
rect 26792 38286 26844 38292
rect 26804 38214 26832 38286
rect 26988 38282 27016 38762
rect 26976 38276 27028 38282
rect 26976 38218 27028 38224
rect 26792 38208 26844 38214
rect 27080 38162 27108 38927
rect 27172 38457 27200 41386
rect 27264 40934 27292 41414
rect 27448 41313 27476 42026
rect 27528 42016 27580 42022
rect 27526 41984 27528 41993
rect 27580 41984 27582 41993
rect 27526 41919 27582 41928
rect 27434 41304 27490 41313
rect 27434 41239 27490 41248
rect 27448 41002 27476 41239
rect 27436 40996 27488 41002
rect 27436 40938 27488 40944
rect 27252 40928 27304 40934
rect 27252 40870 27304 40876
rect 27448 40338 27476 40938
rect 27526 40624 27582 40633
rect 27526 40559 27582 40568
rect 27540 40458 27568 40559
rect 27528 40452 27580 40458
rect 27528 40394 27580 40400
rect 27264 40310 27476 40338
rect 27264 39506 27292 40310
rect 27342 40216 27398 40225
rect 27342 40151 27398 40160
rect 27356 40050 27384 40151
rect 27344 40044 27396 40050
rect 27344 39986 27396 39992
rect 27436 40044 27488 40050
rect 27436 39986 27488 39992
rect 27252 39500 27304 39506
rect 27252 39442 27304 39448
rect 27344 39432 27396 39438
rect 27344 39374 27396 39380
rect 27356 38842 27384 39374
rect 27448 39001 27476 39986
rect 27528 39840 27580 39846
rect 27528 39782 27580 39788
rect 27540 39302 27568 39782
rect 27632 39642 27660 51750
rect 27908 51610 27936 51954
rect 27896 51604 27948 51610
rect 27896 51546 27948 51552
rect 28264 47456 28316 47462
rect 28264 47398 28316 47404
rect 27804 44328 27856 44334
rect 27804 44270 27856 44276
rect 27712 43104 27764 43110
rect 27712 43046 27764 43052
rect 27724 42226 27752 43046
rect 27712 42220 27764 42226
rect 27712 42162 27764 42168
rect 27816 41614 27844 44270
rect 27988 44192 28040 44198
rect 27988 44134 28040 44140
rect 27896 42832 27948 42838
rect 27896 42774 27948 42780
rect 27908 42566 27936 42774
rect 27896 42560 27948 42566
rect 27896 42502 27948 42508
rect 28000 42226 28028 44134
rect 28080 43784 28132 43790
rect 28080 43726 28132 43732
rect 27988 42220 28040 42226
rect 27988 42162 28040 42168
rect 28000 42022 28028 42162
rect 27988 42016 28040 42022
rect 27988 41958 28040 41964
rect 27986 41848 28042 41857
rect 27986 41783 27988 41792
rect 28040 41783 28042 41792
rect 27988 41754 28040 41760
rect 27986 41712 28042 41721
rect 27986 41647 28042 41656
rect 27804 41608 27856 41614
rect 27804 41550 27856 41556
rect 28000 41546 28028 41647
rect 28092 41614 28120 43726
rect 28276 43382 28304 47398
rect 28540 45416 28592 45422
rect 28540 45358 28592 45364
rect 28356 44872 28408 44878
rect 28356 44814 28408 44820
rect 28264 43376 28316 43382
rect 28264 43318 28316 43324
rect 28276 42634 28304 43318
rect 28368 42770 28396 44814
rect 28448 43104 28500 43110
rect 28448 43046 28500 43052
rect 28356 42764 28408 42770
rect 28356 42706 28408 42712
rect 28264 42628 28316 42634
rect 28264 42570 28316 42576
rect 28172 42220 28224 42226
rect 28172 42162 28224 42168
rect 28080 41608 28132 41614
rect 28080 41550 28132 41556
rect 27988 41540 28040 41546
rect 27988 41482 28040 41488
rect 27986 41440 28042 41449
rect 27986 41375 28042 41384
rect 27710 41304 27766 41313
rect 27710 41239 27766 41248
rect 27724 41138 27752 41239
rect 27712 41132 27764 41138
rect 27712 41074 27764 41080
rect 27712 40928 27764 40934
rect 27712 40870 27764 40876
rect 27620 39636 27672 39642
rect 27620 39578 27672 39584
rect 27724 39438 27752 40870
rect 27802 40760 27858 40769
rect 27802 40695 27858 40704
rect 27816 40118 27844 40695
rect 27896 40656 27948 40662
rect 27896 40598 27948 40604
rect 27804 40112 27856 40118
rect 27804 40054 27856 40060
rect 27804 39840 27856 39846
rect 27804 39782 27856 39788
rect 27712 39432 27764 39438
rect 27712 39374 27764 39380
rect 27528 39296 27580 39302
rect 27528 39238 27580 39244
rect 27434 38992 27490 39001
rect 27540 38962 27568 39238
rect 27618 38992 27674 39001
rect 27434 38927 27490 38936
rect 27528 38956 27580 38962
rect 27618 38927 27620 38936
rect 27528 38898 27580 38904
rect 27672 38927 27674 38936
rect 27620 38898 27672 38904
rect 27356 38814 27568 38842
rect 27252 38752 27304 38758
rect 27252 38694 27304 38700
rect 27264 38554 27292 38694
rect 27540 38593 27568 38814
rect 27724 38654 27752 39374
rect 27632 38626 27752 38654
rect 27526 38584 27582 38593
rect 27252 38548 27304 38554
rect 27526 38519 27582 38528
rect 27252 38490 27304 38496
rect 27158 38448 27214 38457
rect 27158 38383 27214 38392
rect 27436 38276 27488 38282
rect 27436 38218 27488 38224
rect 26792 38150 26844 38156
rect 26896 38134 27108 38162
rect 27158 38176 27214 38185
rect 26698 37904 26754 37913
rect 26698 37839 26754 37848
rect 26712 37806 26740 37839
rect 26700 37800 26752 37806
rect 26700 37742 26752 37748
rect 26700 37664 26752 37670
rect 26698 37632 26700 37641
rect 26752 37632 26754 37641
rect 26698 37567 26754 37576
rect 26896 37262 26924 38134
rect 27158 38111 27214 38120
rect 27172 37806 27200 38111
rect 27344 37868 27396 37874
rect 27344 37810 27396 37816
rect 27160 37800 27212 37806
rect 27160 37742 27212 37748
rect 27356 37505 27384 37810
rect 27342 37496 27398 37505
rect 27448 37466 27476 38218
rect 27342 37431 27344 37440
rect 27396 37431 27398 37440
rect 27436 37460 27488 37466
rect 27344 37402 27396 37408
rect 27436 37402 27488 37408
rect 27356 37371 27384 37402
rect 27436 37324 27488 37330
rect 27436 37266 27488 37272
rect 26884 37256 26936 37262
rect 26790 37224 26846 37233
rect 27068 37256 27120 37262
rect 26884 37198 26936 37204
rect 27066 37224 27068 37233
rect 27160 37256 27212 37262
rect 27120 37224 27122 37233
rect 26790 37159 26792 37168
rect 26844 37159 26846 37168
rect 27160 37198 27212 37204
rect 27344 37256 27396 37262
rect 27344 37198 27396 37204
rect 27066 37159 27122 37168
rect 26792 37130 26844 37136
rect 26700 37120 26752 37126
rect 26700 37062 26752 37068
rect 26712 36922 26740 37062
rect 27066 36952 27122 36961
rect 26700 36916 26752 36922
rect 27066 36887 27122 36896
rect 26700 36858 26752 36864
rect 26700 36576 26752 36582
rect 26700 36518 26752 36524
rect 26712 36242 26740 36518
rect 26700 36236 26752 36242
rect 26700 36178 26752 36184
rect 26712 35737 26740 36178
rect 26884 36100 26936 36106
rect 26884 36042 26936 36048
rect 26698 35728 26754 35737
rect 26698 35663 26754 35672
rect 26712 35442 26740 35663
rect 26712 35414 26832 35442
rect 26804 35086 26832 35414
rect 26700 35080 26752 35086
rect 26700 35022 26752 35028
rect 26792 35080 26844 35086
rect 26792 35022 26844 35028
rect 26712 34202 26740 35022
rect 26896 34218 26924 36042
rect 27080 35222 27108 36887
rect 27172 35834 27200 37198
rect 27356 36786 27384 37198
rect 27344 36780 27396 36786
rect 27344 36722 27396 36728
rect 27356 36174 27384 36722
rect 27448 36650 27476 37266
rect 27436 36644 27488 36650
rect 27436 36586 27488 36592
rect 27540 36281 27568 38519
rect 27632 38321 27660 38626
rect 27712 38344 27764 38350
rect 27618 38312 27674 38321
rect 27712 38286 27764 38292
rect 27618 38247 27674 38256
rect 27632 37262 27660 38247
rect 27620 37256 27672 37262
rect 27620 37198 27672 37204
rect 27620 36780 27672 36786
rect 27620 36722 27672 36728
rect 27632 36378 27660 36722
rect 27620 36372 27672 36378
rect 27620 36314 27672 36320
rect 27526 36272 27582 36281
rect 27526 36207 27582 36216
rect 27540 36174 27568 36207
rect 27344 36168 27396 36174
rect 27344 36110 27396 36116
rect 27528 36168 27580 36174
rect 27528 36110 27580 36116
rect 27160 35828 27212 35834
rect 27160 35770 27212 35776
rect 27160 35488 27212 35494
rect 27160 35430 27212 35436
rect 27068 35216 27120 35222
rect 27068 35158 27120 35164
rect 27172 35154 27200 35430
rect 27356 35329 27384 36110
rect 27436 36100 27488 36106
rect 27436 36042 27488 36048
rect 27448 36009 27476 36042
rect 27434 36000 27490 36009
rect 27434 35935 27490 35944
rect 27526 35864 27582 35873
rect 27526 35799 27582 35808
rect 27540 35766 27568 35799
rect 27528 35760 27580 35766
rect 27528 35702 27580 35708
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 27448 35601 27476 35634
rect 27434 35592 27490 35601
rect 27434 35527 27490 35536
rect 27618 35592 27674 35601
rect 27618 35527 27674 35536
rect 27342 35320 27398 35329
rect 27632 35290 27660 35527
rect 27342 35255 27398 35264
rect 27620 35284 27672 35290
rect 27620 35226 27672 35232
rect 27160 35148 27212 35154
rect 27160 35090 27212 35096
rect 27068 35012 27120 35018
rect 27068 34954 27120 34960
rect 27160 35012 27212 35018
rect 27160 34954 27212 34960
rect 27080 34610 27108 34954
rect 27068 34604 27120 34610
rect 27068 34546 27120 34552
rect 27172 34218 27200 34954
rect 27620 34672 27672 34678
rect 27620 34614 27672 34620
rect 26700 34196 26752 34202
rect 26896 34190 27200 34218
rect 26700 34138 26752 34144
rect 26976 34060 27028 34066
rect 26976 34002 27028 34008
rect 26700 33924 26752 33930
rect 26700 33866 26752 33872
rect 26712 33590 26740 33866
rect 26884 33856 26936 33862
rect 26884 33798 26936 33804
rect 26700 33584 26752 33590
rect 26700 33526 26752 33532
rect 26712 33046 26740 33526
rect 26896 33386 26924 33798
rect 26988 33658 27016 34002
rect 27068 33992 27120 33998
rect 27068 33934 27120 33940
rect 27080 33658 27108 33934
rect 26976 33652 27028 33658
rect 26976 33594 27028 33600
rect 27068 33652 27120 33658
rect 27068 33594 27120 33600
rect 26884 33380 26936 33386
rect 26884 33322 26936 33328
rect 26700 33040 26752 33046
rect 26700 32982 26752 32988
rect 26608 31816 26660 31822
rect 26608 31758 26660 31764
rect 26424 31476 26476 31482
rect 26424 31418 26476 31424
rect 26332 31408 26384 31414
rect 26332 31350 26384 31356
rect 26148 30864 26200 30870
rect 26148 30806 26200 30812
rect 26056 30796 26108 30802
rect 26056 30738 26108 30744
rect 25964 29572 26016 29578
rect 25964 29514 26016 29520
rect 25976 29306 26004 29514
rect 25964 29300 26016 29306
rect 25964 29242 26016 29248
rect 25872 28144 25924 28150
rect 25872 28086 25924 28092
rect 25780 28008 25832 28014
rect 25780 27950 25832 27956
rect 25688 26920 25740 26926
rect 25688 26862 25740 26868
rect 25792 26858 25820 27950
rect 25884 27554 25912 28086
rect 25884 27526 26004 27554
rect 25872 27464 25924 27470
rect 25872 27406 25924 27412
rect 25884 27130 25912 27406
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25976 26994 26004 27526
rect 26068 27402 26096 30738
rect 26160 30598 26188 30806
rect 26148 30592 26200 30598
rect 26148 30534 26200 30540
rect 26160 29170 26188 30534
rect 26148 29164 26200 29170
rect 26148 29106 26200 29112
rect 26436 28082 26464 31418
rect 26608 31408 26660 31414
rect 26608 31350 26660 31356
rect 26516 28484 26568 28490
rect 26516 28426 26568 28432
rect 26528 28218 26556 28426
rect 26516 28212 26568 28218
rect 26516 28154 26568 28160
rect 26424 28076 26476 28082
rect 26424 28018 26476 28024
rect 26436 27690 26464 28018
rect 26344 27662 26464 27690
rect 26056 27396 26108 27402
rect 26056 27338 26108 27344
rect 26148 27396 26200 27402
rect 26148 27338 26200 27344
rect 25964 26988 26016 26994
rect 25964 26930 26016 26936
rect 25780 26852 25832 26858
rect 25780 26794 25832 26800
rect 25792 25362 25820 26794
rect 25976 26314 26004 26930
rect 26160 26450 26188 27338
rect 26148 26444 26200 26450
rect 26148 26386 26200 26392
rect 25964 26308 26016 26314
rect 25964 26250 26016 26256
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26252 25498 26280 26250
rect 26344 26042 26372 27662
rect 26424 27600 26476 27606
rect 26422 27568 26424 27577
rect 26476 27568 26478 27577
rect 26422 27503 26478 27512
rect 26528 27470 26556 28154
rect 26620 27946 26648 31350
rect 26712 28626 26740 32982
rect 26896 32910 26924 33322
rect 26884 32904 26936 32910
rect 26884 32846 26936 32852
rect 27080 32842 27108 33594
rect 27068 32836 27120 32842
rect 27068 32778 27120 32784
rect 26884 32496 26936 32502
rect 26884 32438 26936 32444
rect 26790 31784 26846 31793
rect 26790 31719 26846 31728
rect 26700 28620 26752 28626
rect 26700 28562 26752 28568
rect 26608 27940 26660 27946
rect 26608 27882 26660 27888
rect 26516 27464 26568 27470
rect 26516 27406 26568 27412
rect 26516 26920 26568 26926
rect 26516 26862 26568 26868
rect 26424 26784 26476 26790
rect 26424 26726 26476 26732
rect 26436 26382 26464 26726
rect 26424 26376 26476 26382
rect 26424 26318 26476 26324
rect 26332 26036 26384 26042
rect 26332 25978 26384 25984
rect 26240 25492 26292 25498
rect 26240 25434 26292 25440
rect 25780 25356 25832 25362
rect 25780 25298 25832 25304
rect 25792 25242 25820 25298
rect 25700 25214 25820 25242
rect 25700 24410 25728 25214
rect 25872 25152 25924 25158
rect 25872 25094 25924 25100
rect 25780 24608 25832 24614
rect 25780 24550 25832 24556
rect 25688 24404 25740 24410
rect 25688 24346 25740 24352
rect 25700 22778 25728 24346
rect 25792 23322 25820 24550
rect 25884 23730 25912 25094
rect 25872 23724 25924 23730
rect 25872 23666 25924 23672
rect 25780 23316 25832 23322
rect 25780 23258 25832 23264
rect 25884 23118 25912 23666
rect 26252 23118 26280 25434
rect 26344 23798 26372 25978
rect 26436 25362 26464 26318
rect 26424 25356 26476 25362
rect 26424 25298 26476 25304
rect 26436 24614 26464 25298
rect 26424 24608 26476 24614
rect 26424 24550 26476 24556
rect 26436 23866 26464 24550
rect 26528 24070 26556 26862
rect 26620 26790 26648 27882
rect 26608 26784 26660 26790
rect 26608 26726 26660 26732
rect 26712 26518 26740 28562
rect 26700 26512 26752 26518
rect 26700 26454 26752 26460
rect 26608 26444 26660 26450
rect 26608 26386 26660 26392
rect 26620 25294 26648 26386
rect 26712 25906 26740 26454
rect 26700 25900 26752 25906
rect 26700 25842 26752 25848
rect 26712 25294 26740 25842
rect 26608 25288 26660 25294
rect 26608 25230 26660 25236
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 26620 24954 26648 25230
rect 26608 24948 26660 24954
rect 26608 24890 26660 24896
rect 26712 24410 26740 25230
rect 26804 25158 26832 31719
rect 26896 26926 26924 32438
rect 26976 32428 27028 32434
rect 26976 32370 27028 32376
rect 26988 32230 27016 32370
rect 26976 32224 27028 32230
rect 26976 32166 27028 32172
rect 26974 31920 27030 31929
rect 26974 31855 27030 31864
rect 26988 31822 27016 31855
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 27080 31414 27108 32778
rect 27068 31408 27120 31414
rect 27068 31350 27120 31356
rect 26976 30660 27028 30666
rect 26976 30602 27028 30608
rect 26988 30394 27016 30602
rect 26976 30388 27028 30394
rect 26976 30330 27028 30336
rect 27068 28416 27120 28422
rect 27068 28358 27120 28364
rect 27080 27470 27108 28358
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 27068 27328 27120 27334
rect 27068 27270 27120 27276
rect 27080 26994 27108 27270
rect 27068 26988 27120 26994
rect 27068 26930 27120 26936
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 26792 25152 26844 25158
rect 26792 25094 26844 25100
rect 26884 24744 26936 24750
rect 26884 24686 26936 24692
rect 26700 24404 26752 24410
rect 26700 24346 26752 24352
rect 26896 24206 26924 24686
rect 26884 24200 26936 24206
rect 26884 24142 26936 24148
rect 26516 24064 26568 24070
rect 26516 24006 26568 24012
rect 26424 23860 26476 23866
rect 26424 23802 26476 23808
rect 26332 23792 26384 23798
rect 26332 23734 26384 23740
rect 26332 23180 26384 23186
rect 26332 23122 26384 23128
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 25688 22772 25740 22778
rect 25688 22714 25740 22720
rect 26344 22710 26372 23122
rect 26424 22976 26476 22982
rect 26424 22918 26476 22924
rect 26332 22704 26384 22710
rect 26332 22646 26384 22652
rect 25688 22500 25740 22506
rect 25688 22442 25740 22448
rect 25516 22066 25636 22094
rect 25516 21962 25544 22066
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25412 17264 25464 17270
rect 25412 17206 25464 17212
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25042 16623 25044 16632
rect 25096 16623 25098 16632
rect 25136 16652 25188 16658
rect 25044 16594 25096 16600
rect 25136 16594 25188 16600
rect 25240 16590 25268 16934
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 24584 16516 24636 16522
rect 24584 16458 24636 16464
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23572 11824 23624 11830
rect 23572 11766 23624 11772
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23584 10266 23612 11766
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23676 11014 23704 11630
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23584 9654 23612 10202
rect 23676 10062 23704 10950
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23480 9580 23532 9586
rect 23308 9540 23480 9568
rect 23480 9522 23532 9528
rect 23572 9512 23624 9518
rect 23570 9480 23572 9489
rect 23624 9480 23626 9489
rect 23768 9450 23796 11766
rect 23860 11354 23888 12718
rect 23940 12300 23992 12306
rect 23940 12242 23992 12248
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23952 11286 23980 12242
rect 24032 12164 24084 12170
rect 24032 12106 24084 12112
rect 23940 11280 23992 11286
rect 23940 11222 23992 11228
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23570 9415 23626 9424
rect 23756 9444 23808 9450
rect 23756 9386 23808 9392
rect 23860 8974 23888 10406
rect 23940 9988 23992 9994
rect 23940 9930 23992 9936
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 23756 8900 23808 8906
rect 23756 8842 23808 8848
rect 23112 8832 23164 8838
rect 23112 8774 23164 8780
rect 23124 8634 23152 8774
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22848 5370 22876 6598
rect 23124 6458 23152 8570
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23584 8090 23612 8434
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23768 8022 23796 8842
rect 23756 8016 23808 8022
rect 23756 7958 23808 7964
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23216 7546 23244 7822
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23124 5710 23152 6394
rect 23216 5914 23244 7482
rect 23754 7440 23810 7449
rect 23754 7375 23810 7384
rect 23572 7200 23624 7206
rect 23572 7142 23624 7148
rect 23584 6730 23612 7142
rect 23572 6724 23624 6730
rect 23572 6666 23624 6672
rect 23664 6724 23716 6730
rect 23664 6666 23716 6672
rect 23676 6458 23704 6666
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23768 6338 23796 7375
rect 23676 6310 23796 6338
rect 23204 5908 23256 5914
rect 23204 5850 23256 5856
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 22836 5364 22888 5370
rect 22836 5306 22888 5312
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 23308 4486 23336 4626
rect 23676 4486 23704 6310
rect 23296 4480 23348 4486
rect 23296 4422 23348 4428
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 23112 4072 23164 4078
rect 23112 4014 23164 4020
rect 23124 3670 23152 4014
rect 23112 3664 23164 3670
rect 23112 3606 23164 3612
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 22664 800 22692 2790
rect 23308 2446 23336 4422
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 23492 3466 23520 3878
rect 23480 3460 23532 3466
rect 23480 3402 23532 3408
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 23032 800 23060 2246
rect 23400 800 23428 2790
rect 23492 2446 23520 3402
rect 23676 3058 23704 4422
rect 23952 4078 23980 9930
rect 24044 9178 24072 12106
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 24228 11694 24256 12038
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 24136 5914 24164 9318
rect 24228 6118 24256 11630
rect 24320 7818 24348 13806
rect 24596 13530 24624 16458
rect 25516 15978 25544 21286
rect 25504 15972 25556 15978
rect 25504 15914 25556 15920
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24688 14006 24716 15438
rect 24780 15026 24808 15642
rect 25136 15088 25188 15094
rect 25136 15030 25188 15036
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24768 14884 24820 14890
rect 24768 14826 24820 14832
rect 24676 14000 24728 14006
rect 24676 13942 24728 13948
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24308 7812 24360 7818
rect 24308 7754 24360 7760
rect 24216 6112 24268 6118
rect 24216 6054 24268 6060
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23768 3058 23796 3878
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 24136 2990 24164 5850
rect 24308 5704 24360 5710
rect 24308 5646 24360 5652
rect 24124 2984 24176 2990
rect 24124 2926 24176 2932
rect 24124 2848 24176 2854
rect 24124 2790 24176 2796
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23756 2304 23808 2310
rect 23756 2246 23808 2252
rect 23768 800 23796 2246
rect 24136 800 24164 2790
rect 24320 2650 24348 5646
rect 24412 3194 24440 13126
rect 24584 8832 24636 8838
rect 24584 8774 24636 8780
rect 24492 8356 24544 8362
rect 24492 8298 24544 8304
rect 24504 6254 24532 8298
rect 24596 6322 24624 8774
rect 24688 8090 24716 13942
rect 24780 13802 24808 14826
rect 24768 13796 24820 13802
rect 24768 13738 24820 13744
rect 25148 13326 25176 15030
rect 25320 14952 25372 14958
rect 25318 14920 25320 14929
rect 25372 14920 25374 14929
rect 25318 14855 25374 14864
rect 25332 13394 25360 14855
rect 25516 14278 25544 15914
rect 25504 14272 25556 14278
rect 25504 14214 25556 14220
rect 25320 13388 25372 13394
rect 25320 13330 25372 13336
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25412 13320 25464 13326
rect 25412 13262 25464 13268
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 24952 12640 25004 12646
rect 24872 12588 24952 12594
rect 24872 12582 25004 12588
rect 24872 12566 24992 12582
rect 24872 11762 24900 12566
rect 25056 12170 25084 13194
rect 25320 12844 25372 12850
rect 25320 12786 25372 12792
rect 25044 12164 25096 12170
rect 25044 12106 25096 12112
rect 24860 11756 24912 11762
rect 24860 11698 24912 11704
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24780 11082 24808 11630
rect 25056 11354 25084 12106
rect 25044 11348 25096 11354
rect 25044 11290 25096 11296
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24768 11076 24820 11082
rect 24768 11018 24820 11024
rect 24780 10810 24808 11018
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24768 9580 24820 9586
rect 24768 9522 24820 9528
rect 24780 9178 24808 9522
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24676 8084 24728 8090
rect 24676 8026 24728 8032
rect 24688 6730 24716 8026
rect 24768 7812 24820 7818
rect 24768 7754 24820 7760
rect 24780 7206 24808 7754
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24872 6882 24900 7686
rect 24964 7562 24992 11086
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 25056 9722 25084 9862
rect 25044 9716 25096 9722
rect 25044 9658 25096 9664
rect 25240 9489 25268 10066
rect 25332 9625 25360 12786
rect 25424 12238 25452 13262
rect 25412 12232 25464 12238
rect 25412 12174 25464 12180
rect 25318 9616 25374 9625
rect 25318 9551 25374 9560
rect 25226 9480 25282 9489
rect 25226 9415 25282 9424
rect 25136 9036 25188 9042
rect 25136 8978 25188 8984
rect 25148 8634 25176 8978
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25148 7954 25176 8570
rect 25240 8090 25268 9415
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 24964 7534 25084 7562
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 24964 7002 24992 7346
rect 24952 6996 25004 7002
rect 24952 6938 25004 6944
rect 24872 6854 24992 6882
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24492 6248 24544 6254
rect 24492 6190 24544 6196
rect 24676 6180 24728 6186
rect 24676 6122 24728 6128
rect 24688 5914 24716 6122
rect 24676 5908 24728 5914
rect 24676 5850 24728 5856
rect 24964 5030 24992 6854
rect 25056 6458 25084 7534
rect 25148 6866 25176 7890
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 25056 5370 25084 6394
rect 25148 6254 25176 6802
rect 25332 6798 25360 9551
rect 25412 8424 25464 8430
rect 25412 8366 25464 8372
rect 25320 6792 25372 6798
rect 25320 6734 25372 6740
rect 25332 6458 25360 6734
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25044 5364 25096 5370
rect 25044 5306 25096 5312
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24964 3534 24992 4966
rect 25424 4486 25452 8366
rect 25412 4480 25464 4486
rect 25412 4422 25464 4428
rect 25320 4276 25372 4282
rect 25320 4218 25372 4224
rect 25136 4072 25188 4078
rect 25136 4014 25188 4020
rect 25044 3936 25096 3942
rect 25044 3878 25096 3884
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24400 3188 24452 3194
rect 24400 3130 24452 3136
rect 24308 2644 24360 2650
rect 24308 2586 24360 2592
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 24504 800 24532 2246
rect 24872 800 24900 3334
rect 25056 3058 25084 3878
rect 25044 3052 25096 3058
rect 25044 2994 25096 3000
rect 25148 2774 25176 4014
rect 25332 3534 25360 4218
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 25424 3126 25452 4422
rect 25516 4078 25544 14214
rect 25700 8634 25728 22442
rect 26332 21888 26384 21894
rect 26332 21830 26384 21836
rect 26148 21616 26200 21622
rect 26148 21558 26200 21564
rect 25780 20528 25832 20534
rect 25780 20470 25832 20476
rect 25792 19922 25820 20470
rect 26160 20058 26188 21558
rect 26344 21146 26372 21830
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 26148 20052 26200 20058
rect 26148 19994 26200 20000
rect 25780 19916 25832 19922
rect 25780 19858 25832 19864
rect 26056 19780 26108 19786
rect 26056 19722 26108 19728
rect 26068 19514 26096 19722
rect 26160 19718 26188 19994
rect 26148 19712 26200 19718
rect 26148 19654 26200 19660
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26160 17270 26188 17478
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 26148 17264 26200 17270
rect 26148 17206 26200 17212
rect 25872 16176 25924 16182
rect 25872 16118 25924 16124
rect 25780 14952 25832 14958
rect 25780 14894 25832 14900
rect 25792 13938 25820 14894
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 25884 10470 25912 16118
rect 25872 10464 25924 10470
rect 25872 10406 25924 10412
rect 25884 10062 25912 10406
rect 25872 10056 25924 10062
rect 25872 9998 25924 10004
rect 25872 9580 25924 9586
rect 25872 9522 25924 9528
rect 25780 9376 25832 9382
rect 25780 9318 25832 9324
rect 25792 9110 25820 9318
rect 25780 9104 25832 9110
rect 25780 9046 25832 9052
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 25792 5574 25820 6394
rect 25780 5568 25832 5574
rect 25780 5510 25832 5516
rect 25792 4826 25820 5510
rect 25884 5370 25912 9522
rect 25976 9450 26004 17206
rect 26238 16824 26294 16833
rect 26238 16759 26294 16768
rect 26252 16590 26280 16759
rect 26240 16584 26292 16590
rect 26240 16526 26292 16532
rect 26240 16040 26292 16046
rect 26240 15982 26292 15988
rect 26332 16040 26384 16046
rect 26332 15982 26384 15988
rect 26252 15570 26280 15982
rect 26344 15706 26372 15982
rect 26332 15700 26384 15706
rect 26332 15642 26384 15648
rect 26240 15564 26292 15570
rect 26240 15506 26292 15512
rect 26054 15192 26110 15201
rect 26054 15127 26056 15136
rect 26108 15127 26110 15136
rect 26056 15098 26108 15104
rect 26068 13938 26096 15098
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 26240 14340 26292 14346
rect 26240 14282 26292 14288
rect 26056 13932 26108 13938
rect 26056 13874 26108 13880
rect 26252 13530 26280 14282
rect 26240 13524 26292 13530
rect 26240 13466 26292 13472
rect 26240 12912 26292 12918
rect 26240 12854 26292 12860
rect 26148 12708 26200 12714
rect 26148 12650 26200 12656
rect 26160 11082 26188 12650
rect 26252 11898 26280 12854
rect 26344 12209 26372 14894
rect 26330 12200 26386 12209
rect 26330 12135 26386 12144
rect 26332 12096 26384 12102
rect 26332 12038 26384 12044
rect 26240 11892 26292 11898
rect 26240 11834 26292 11840
rect 26344 11150 26372 12038
rect 26332 11144 26384 11150
rect 26332 11086 26384 11092
rect 26148 11076 26200 11082
rect 26148 11018 26200 11024
rect 26436 10810 26464 22918
rect 26516 22432 26568 22438
rect 26516 22374 26568 22380
rect 26528 21486 26556 22374
rect 26896 22234 26924 24142
rect 26976 23656 27028 23662
rect 26976 23598 27028 23604
rect 26884 22228 26936 22234
rect 26884 22170 26936 22176
rect 26608 21956 26660 21962
rect 26608 21898 26660 21904
rect 26792 21956 26844 21962
rect 26792 21898 26844 21904
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 26528 21049 26556 21422
rect 26620 21146 26648 21898
rect 26608 21140 26660 21146
rect 26608 21082 26660 21088
rect 26514 21040 26570 21049
rect 26514 20975 26570 20984
rect 26516 20800 26568 20806
rect 26516 20742 26568 20748
rect 26528 20602 26556 20742
rect 26516 20596 26568 20602
rect 26516 20538 26568 20544
rect 26528 19514 26556 20538
rect 26620 20466 26648 21082
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 26804 20398 26832 21898
rect 26884 21412 26936 21418
rect 26884 21354 26936 21360
rect 26896 21146 26924 21354
rect 26884 21140 26936 21146
rect 26884 21082 26936 21088
rect 26792 20392 26844 20398
rect 26792 20334 26844 20340
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 26516 19304 26568 19310
rect 26516 19246 26568 19252
rect 26528 18970 26556 19246
rect 26516 18964 26568 18970
rect 26516 18906 26568 18912
rect 26516 18352 26568 18358
rect 26516 18294 26568 18300
rect 26528 17270 26556 18294
rect 26884 17808 26936 17814
rect 26884 17750 26936 17756
rect 26516 17264 26568 17270
rect 26516 17206 26568 17212
rect 26896 17066 26924 17750
rect 26884 17060 26936 17066
rect 26884 17002 26936 17008
rect 26516 15496 26568 15502
rect 26516 15438 26568 15444
rect 26528 15162 26556 15438
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26516 15156 26568 15162
rect 26516 15098 26568 15104
rect 26608 14340 26660 14346
rect 26608 14282 26660 14288
rect 26620 13802 26648 14282
rect 26700 13932 26752 13938
rect 26700 13874 26752 13880
rect 26608 13796 26660 13802
rect 26608 13738 26660 13744
rect 26620 12986 26648 13738
rect 26608 12980 26660 12986
rect 26608 12922 26660 12928
rect 26516 12640 26568 12646
rect 26516 12582 26568 12588
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 25964 9444 26016 9450
rect 25964 9386 26016 9392
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 25976 5370 26004 8774
rect 26068 5914 26096 9998
rect 26148 9580 26200 9586
rect 26148 9522 26200 9528
rect 26160 9353 26188 9522
rect 26146 9344 26202 9353
rect 26146 9279 26202 9288
rect 26056 5908 26108 5914
rect 26056 5850 26108 5856
rect 26148 5704 26200 5710
rect 26252 5658 26280 10610
rect 26332 10600 26384 10606
rect 26332 10542 26384 10548
rect 26344 9994 26372 10542
rect 26332 9988 26384 9994
rect 26332 9930 26384 9936
rect 26344 9654 26372 9930
rect 26332 9648 26384 9654
rect 26332 9590 26384 9596
rect 26344 9518 26372 9590
rect 26332 9512 26384 9518
rect 26332 9454 26384 9460
rect 26344 8838 26372 9454
rect 26422 9072 26478 9081
rect 26422 9007 26424 9016
rect 26476 9007 26478 9016
rect 26424 8978 26476 8984
rect 26332 8832 26384 8838
rect 26332 8774 26384 8780
rect 26424 8832 26476 8838
rect 26424 8774 26476 8780
rect 26344 8412 26372 8774
rect 26436 8566 26464 8774
rect 26424 8560 26476 8566
rect 26424 8502 26476 8508
rect 26424 8424 26476 8430
rect 26344 8384 26424 8412
rect 26424 8366 26476 8372
rect 26436 7954 26464 8366
rect 26424 7948 26476 7954
rect 26424 7890 26476 7896
rect 26424 7744 26476 7750
rect 26424 7686 26476 7692
rect 26436 7206 26464 7686
rect 26424 7200 26476 7206
rect 26424 7142 26476 7148
rect 26528 6866 26556 12582
rect 26620 12442 26648 12922
rect 26608 12436 26660 12442
rect 26608 12378 26660 12384
rect 26620 11218 26648 12378
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 26200 5652 26280 5658
rect 26148 5646 26280 5652
rect 26160 5630 26280 5646
rect 26332 5636 26384 5642
rect 26332 5578 26384 5584
rect 25872 5364 25924 5370
rect 25872 5306 25924 5312
rect 25964 5364 26016 5370
rect 25964 5306 26016 5312
rect 25884 5166 25912 5306
rect 25872 5160 25924 5166
rect 25872 5102 25924 5108
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 26344 4214 26372 5578
rect 26332 4208 26384 4214
rect 26332 4150 26384 4156
rect 26712 4146 26740 13874
rect 26804 13530 26832 15302
rect 26884 14952 26936 14958
rect 26884 14894 26936 14900
rect 26792 13524 26844 13530
rect 26792 13466 26844 13472
rect 26896 12102 26924 14894
rect 26884 12096 26936 12102
rect 26884 12038 26936 12044
rect 26988 9450 27016 23598
rect 27080 21010 27108 26930
rect 27172 26586 27200 34190
rect 27344 33992 27396 33998
rect 27344 33934 27396 33940
rect 27252 33924 27304 33930
rect 27252 33866 27304 33872
rect 27264 32230 27292 33866
rect 27356 33454 27384 33934
rect 27344 33448 27396 33454
rect 27344 33390 27396 33396
rect 27632 32978 27660 34614
rect 27620 32972 27672 32978
rect 27620 32914 27672 32920
rect 27344 32904 27396 32910
rect 27344 32846 27396 32852
rect 27252 32224 27304 32230
rect 27252 32166 27304 32172
rect 27160 26580 27212 26586
rect 27160 26522 27212 26528
rect 27264 26042 27292 32166
rect 27356 31754 27384 32846
rect 27632 32502 27660 32914
rect 27620 32496 27672 32502
rect 27620 32438 27672 32444
rect 27436 32292 27488 32298
rect 27436 32234 27488 32240
rect 27448 32026 27476 32234
rect 27436 32020 27488 32026
rect 27436 31962 27488 31968
rect 27356 31726 27476 31754
rect 27344 29844 27396 29850
rect 27344 29786 27396 29792
rect 27356 29170 27384 29786
rect 27344 29164 27396 29170
rect 27344 29106 27396 29112
rect 27344 29028 27396 29034
rect 27344 28970 27396 28976
rect 27356 28082 27384 28970
rect 27344 28076 27396 28082
rect 27344 28018 27396 28024
rect 27356 27946 27384 28018
rect 27344 27940 27396 27946
rect 27344 27882 27396 27888
rect 27448 26994 27476 31726
rect 27724 30938 27752 38286
rect 27816 31754 27844 39782
rect 27908 37777 27936 40598
rect 28000 39098 28028 41375
rect 28078 40488 28134 40497
rect 28078 40423 28080 40432
rect 28132 40423 28134 40432
rect 28080 40394 28132 40400
rect 28184 40050 28212 42162
rect 28264 42016 28316 42022
rect 28264 41958 28316 41964
rect 28276 41721 28304 41958
rect 28262 41712 28318 41721
rect 28262 41647 28318 41656
rect 28368 41290 28396 42706
rect 28460 42702 28488 43046
rect 28448 42696 28500 42702
rect 28448 42638 28500 42644
rect 28460 41614 28488 42638
rect 28552 41818 28580 45358
rect 28632 45008 28684 45014
rect 28632 44950 28684 44956
rect 28644 44538 28672 44950
rect 28632 44532 28684 44538
rect 28632 44474 28684 44480
rect 28644 43858 28672 44474
rect 28632 43852 28684 43858
rect 28632 43794 28684 43800
rect 28632 42220 28684 42226
rect 28632 42162 28684 42168
rect 28540 41812 28592 41818
rect 28540 41754 28592 41760
rect 28448 41608 28500 41614
rect 28448 41550 28500 41556
rect 28552 41449 28580 41754
rect 28538 41440 28594 41449
rect 28538 41375 28594 41384
rect 28368 41262 28580 41290
rect 28644 41274 28672 42162
rect 28736 41857 28764 52838
rect 29828 51808 29880 51814
rect 29828 51750 29880 51756
rect 29644 51604 29696 51610
rect 29644 51546 29696 51552
rect 29656 47802 29684 51546
rect 29644 47796 29696 47802
rect 29644 47738 29696 47744
rect 29092 47660 29144 47666
rect 29092 47602 29144 47608
rect 29104 47258 29132 47602
rect 29092 47252 29144 47258
rect 29092 47194 29144 47200
rect 29656 47122 29684 47738
rect 29644 47116 29696 47122
rect 29644 47058 29696 47064
rect 29656 45558 29684 47058
rect 29644 45552 29696 45558
rect 29644 45494 29696 45500
rect 28908 43716 28960 43722
rect 28908 43658 28960 43664
rect 28816 42220 28868 42226
rect 28816 42162 28868 42168
rect 28828 41993 28856 42162
rect 28920 42158 28948 43658
rect 29000 43648 29052 43654
rect 29000 43590 29052 43596
rect 29012 43314 29040 43590
rect 29184 43376 29236 43382
rect 29184 43318 29236 43324
rect 29000 43308 29052 43314
rect 29000 43250 29052 43256
rect 29012 42294 29040 43250
rect 29092 43104 29144 43110
rect 29092 43046 29144 43052
rect 29000 42288 29052 42294
rect 29000 42230 29052 42236
rect 28908 42152 28960 42158
rect 28908 42094 28960 42100
rect 28814 41984 28870 41993
rect 28814 41919 28870 41928
rect 28722 41848 28778 41857
rect 28722 41783 28778 41792
rect 28816 41676 28868 41682
rect 28816 41618 28868 41624
rect 28722 41576 28778 41585
rect 28722 41511 28778 41520
rect 28264 40520 28316 40526
rect 28264 40462 28316 40468
rect 28080 40044 28132 40050
rect 28080 39986 28132 39992
rect 28172 40044 28224 40050
rect 28172 39986 28224 39992
rect 27988 39092 28040 39098
rect 27988 39034 28040 39040
rect 28092 38865 28120 39986
rect 28172 39636 28224 39642
rect 28172 39578 28224 39584
rect 28078 38856 28134 38865
rect 28078 38791 28134 38800
rect 27988 38752 28040 38758
rect 27988 38694 28040 38700
rect 27894 37768 27950 37777
rect 27894 37703 27950 37712
rect 27894 37224 27950 37233
rect 27894 37159 27896 37168
rect 27948 37159 27950 37168
rect 27896 37130 27948 37136
rect 27896 36712 27948 36718
rect 27894 36680 27896 36689
rect 27948 36680 27950 36689
rect 27894 36615 27950 36624
rect 27894 36544 27950 36553
rect 27894 36479 27950 36488
rect 27908 36242 27936 36479
rect 27896 36236 27948 36242
rect 27896 36178 27948 36184
rect 27896 36032 27948 36038
rect 27896 35974 27948 35980
rect 27804 31748 27856 31754
rect 27804 31690 27856 31696
rect 27712 30932 27764 30938
rect 27712 30874 27764 30880
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 27816 29578 27844 29786
rect 27804 29572 27856 29578
rect 27804 29514 27856 29520
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27540 29034 27568 29106
rect 27528 29028 27580 29034
rect 27528 28970 27580 28976
rect 27528 28484 27580 28490
rect 27528 28426 27580 28432
rect 27804 28484 27856 28490
rect 27804 28426 27856 28432
rect 27540 28150 27568 28426
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 27528 28144 27580 28150
rect 27528 28086 27580 28092
rect 27632 28082 27660 28358
rect 27816 28218 27844 28426
rect 27804 28212 27856 28218
rect 27804 28154 27856 28160
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 27908 27470 27936 35974
rect 28000 34105 28028 38694
rect 28092 37874 28120 38791
rect 28184 38418 28212 39578
rect 28276 39545 28304 40462
rect 28552 40225 28580 41262
rect 28632 41268 28684 41274
rect 28632 41210 28684 41216
rect 28736 41206 28764 41511
rect 28724 41200 28776 41206
rect 28724 41142 28776 41148
rect 28632 41132 28684 41138
rect 28632 41074 28684 41080
rect 28644 41002 28672 41074
rect 28632 40996 28684 41002
rect 28632 40938 28684 40944
rect 28538 40216 28594 40225
rect 28448 40180 28500 40186
rect 28538 40151 28594 40160
rect 28448 40122 28500 40128
rect 28460 39982 28488 40122
rect 28448 39976 28500 39982
rect 28448 39918 28500 39924
rect 28356 39908 28408 39914
rect 28356 39850 28408 39856
rect 28262 39536 28318 39545
rect 28262 39471 28318 39480
rect 28276 39438 28304 39471
rect 28264 39432 28316 39438
rect 28264 39374 28316 39380
rect 28368 38962 28396 39850
rect 28264 38956 28316 38962
rect 28264 38898 28316 38904
rect 28356 38956 28408 38962
rect 28356 38898 28408 38904
rect 28172 38412 28224 38418
rect 28172 38354 28224 38360
rect 28276 38049 28304 38898
rect 28540 38480 28592 38486
rect 28460 38457 28540 38468
rect 28446 38448 28540 38457
rect 28502 38440 28540 38448
rect 28540 38422 28592 38428
rect 28446 38383 28502 38392
rect 28356 38208 28408 38214
rect 28356 38150 28408 38156
rect 28262 38040 28318 38049
rect 28172 38004 28224 38010
rect 28262 37975 28318 37984
rect 28172 37946 28224 37952
rect 28080 37868 28132 37874
rect 28080 37810 28132 37816
rect 28092 36174 28120 37810
rect 28184 37466 28212 37946
rect 28264 37664 28316 37670
rect 28262 37632 28264 37641
rect 28316 37632 28318 37641
rect 28262 37567 28318 37576
rect 28172 37460 28224 37466
rect 28172 37402 28224 37408
rect 28172 37256 28224 37262
rect 28172 37198 28224 37204
rect 28184 37097 28212 37198
rect 28170 37088 28226 37097
rect 28170 37023 28226 37032
rect 28262 36952 28318 36961
rect 28262 36887 28318 36896
rect 28276 36786 28304 36887
rect 28368 36854 28396 38150
rect 28460 37330 28488 38383
rect 28540 38208 28592 38214
rect 28540 38150 28592 38156
rect 28448 37324 28500 37330
rect 28448 37266 28500 37272
rect 28356 36848 28408 36854
rect 28356 36790 28408 36796
rect 28264 36780 28316 36786
rect 28264 36722 28316 36728
rect 28080 36168 28132 36174
rect 28080 36110 28132 36116
rect 28172 36032 28224 36038
rect 28172 35974 28224 35980
rect 28080 34604 28132 34610
rect 28080 34546 28132 34552
rect 28092 34513 28120 34546
rect 28078 34504 28134 34513
rect 28078 34439 28134 34448
rect 28080 34128 28132 34134
rect 27986 34096 28042 34105
rect 28080 34070 28132 34076
rect 27986 34031 28042 34040
rect 27988 33992 28040 33998
rect 27988 33934 28040 33940
rect 28000 33114 28028 33934
rect 27988 33108 28040 33114
rect 27988 33050 28040 33056
rect 28092 32910 28120 34070
rect 28080 32904 28132 32910
rect 28080 32846 28132 32852
rect 27988 31272 28040 31278
rect 27988 31214 28040 31220
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27896 27464 27948 27470
rect 27896 27406 27948 27412
rect 27436 26988 27488 26994
rect 27436 26930 27488 26936
rect 27448 26450 27476 26930
rect 27436 26444 27488 26450
rect 27436 26386 27488 26392
rect 27724 26382 27752 27406
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 27528 26308 27580 26314
rect 27528 26250 27580 26256
rect 27252 26036 27304 26042
rect 27252 25978 27304 25984
rect 27160 24132 27212 24138
rect 27160 24074 27212 24080
rect 27172 23322 27200 24074
rect 27264 23730 27292 25978
rect 27540 25294 27568 26250
rect 27528 25288 27580 25294
rect 27528 25230 27580 25236
rect 27252 23724 27304 23730
rect 27252 23666 27304 23672
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27436 23588 27488 23594
rect 27436 23530 27488 23536
rect 27252 23520 27304 23526
rect 27252 23462 27304 23468
rect 27160 23316 27212 23322
rect 27160 23258 27212 23264
rect 27264 23118 27292 23462
rect 27252 23112 27304 23118
rect 27252 23054 27304 23060
rect 27344 22976 27396 22982
rect 27344 22918 27396 22924
rect 27356 22574 27384 22918
rect 27344 22568 27396 22574
rect 27344 22510 27396 22516
rect 27356 22166 27384 22510
rect 27448 22506 27476 23530
rect 27724 23186 27752 23598
rect 27712 23180 27764 23186
rect 27712 23122 27764 23128
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 27436 22500 27488 22506
rect 27436 22442 27488 22448
rect 27436 22228 27488 22234
rect 27436 22170 27488 22176
rect 27344 22160 27396 22166
rect 27344 22102 27396 22108
rect 27448 22098 27476 22170
rect 27436 22092 27488 22098
rect 27436 22034 27488 22040
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 27172 20602 27200 21966
rect 27540 21690 27568 22578
rect 28000 22094 28028 31214
rect 28080 28960 28132 28966
rect 28080 28902 28132 28908
rect 28092 27878 28120 28902
rect 28184 28014 28212 35974
rect 28356 35692 28408 35698
rect 28356 35634 28408 35640
rect 28264 35012 28316 35018
rect 28264 34954 28316 34960
rect 28276 34202 28304 34954
rect 28264 34196 28316 34202
rect 28264 34138 28316 34144
rect 28276 33658 28304 34138
rect 28368 34134 28396 35634
rect 28460 35290 28488 37266
rect 28552 36786 28580 38150
rect 28540 36780 28592 36786
rect 28540 36722 28592 36728
rect 28644 36174 28672 40938
rect 28828 40746 28856 41618
rect 28736 40718 28856 40746
rect 28736 40633 28764 40718
rect 28816 40656 28868 40662
rect 28722 40624 28778 40633
rect 28816 40598 28868 40604
rect 28722 40559 28724 40568
rect 28776 40559 28778 40568
rect 28724 40530 28776 40536
rect 28736 38826 28764 40530
rect 28828 40361 28856 40598
rect 28814 40352 28870 40361
rect 28814 40287 28870 40296
rect 28920 40186 28948 42094
rect 29104 41138 29132 43046
rect 29196 42362 29224 43318
rect 29644 43240 29696 43246
rect 29366 43208 29422 43217
rect 29366 43143 29422 43152
rect 29642 43208 29644 43217
rect 29696 43208 29698 43217
rect 29642 43143 29698 43152
rect 29184 42356 29236 42362
rect 29184 42298 29236 42304
rect 29276 41608 29328 41614
rect 29276 41550 29328 41556
rect 29092 41132 29144 41138
rect 29092 41074 29144 41080
rect 29184 41132 29236 41138
rect 29184 41074 29236 41080
rect 29104 40905 29132 41074
rect 29090 40896 29146 40905
rect 29090 40831 29146 40840
rect 29092 40520 29144 40526
rect 29092 40462 29144 40468
rect 29104 40390 29132 40462
rect 29092 40384 29144 40390
rect 29092 40326 29144 40332
rect 28908 40180 28960 40186
rect 28908 40122 28960 40128
rect 28908 39908 28960 39914
rect 28908 39850 28960 39856
rect 28920 39098 28948 39850
rect 29000 39840 29052 39846
rect 29000 39782 29052 39788
rect 28908 39092 28960 39098
rect 28908 39034 28960 39040
rect 28816 38956 28868 38962
rect 28816 38898 28868 38904
rect 28724 38820 28776 38826
rect 28724 38762 28776 38768
rect 28736 38214 28764 38762
rect 28828 38418 28856 38898
rect 29012 38593 29040 39782
rect 29104 39438 29132 40326
rect 29092 39432 29144 39438
rect 29092 39374 29144 39380
rect 28998 38584 29054 38593
rect 28998 38519 29054 38528
rect 28954 38480 29006 38486
rect 29006 38448 29054 38457
rect 28954 38422 28998 38428
rect 28816 38412 28868 38418
rect 28966 38406 28998 38422
rect 28998 38383 29054 38392
rect 28816 38354 28868 38360
rect 29000 38344 29052 38350
rect 29000 38286 29052 38292
rect 28816 38276 28868 38282
rect 28816 38218 28868 38224
rect 28724 38208 28776 38214
rect 28724 38150 28776 38156
rect 28828 37913 28856 38218
rect 29012 38214 29040 38286
rect 29000 38208 29052 38214
rect 29000 38150 29052 38156
rect 28908 37936 28960 37942
rect 28814 37904 28870 37913
rect 28724 37868 28776 37874
rect 28908 37878 28960 37884
rect 28814 37839 28870 37848
rect 28724 37810 28776 37816
rect 28736 37482 28764 37810
rect 28736 37454 28856 37482
rect 28828 37330 28856 37454
rect 28920 37330 28948 37878
rect 29104 37874 29132 39374
rect 29196 38706 29224 41074
rect 29288 41002 29316 41550
rect 29380 41274 29408 43143
rect 29644 42764 29696 42770
rect 29644 42706 29696 42712
rect 29460 42628 29512 42634
rect 29460 42570 29512 42576
rect 29472 42362 29500 42570
rect 29552 42560 29604 42566
rect 29552 42502 29604 42508
rect 29460 42356 29512 42362
rect 29460 42298 29512 42304
rect 29472 41682 29500 42298
rect 29460 41676 29512 41682
rect 29460 41618 29512 41624
rect 29368 41268 29420 41274
rect 29368 41210 29420 41216
rect 29276 40996 29328 41002
rect 29276 40938 29328 40944
rect 29460 40928 29512 40934
rect 29458 40896 29460 40905
rect 29512 40896 29514 40905
rect 29458 40831 29514 40840
rect 29460 39976 29512 39982
rect 29460 39918 29512 39924
rect 29276 39432 29328 39438
rect 29276 39374 29328 39380
rect 29288 38962 29316 39374
rect 29472 39302 29500 39918
rect 29460 39296 29512 39302
rect 29460 39238 29512 39244
rect 29472 38962 29500 39238
rect 29276 38956 29328 38962
rect 29276 38898 29328 38904
rect 29460 38956 29512 38962
rect 29460 38898 29512 38904
rect 29191 38678 29224 38706
rect 29368 38752 29420 38758
rect 29368 38694 29420 38700
rect 29191 38536 29219 38678
rect 29380 38654 29408 38694
rect 29380 38626 29409 38654
rect 29191 38508 29224 38536
rect 29092 37868 29144 37874
rect 29092 37810 29144 37816
rect 28816 37324 28868 37330
rect 28816 37266 28868 37272
rect 28908 37324 28960 37330
rect 28908 37266 28960 37272
rect 28724 37256 28776 37262
rect 28724 37198 28776 37204
rect 28736 36922 28764 37198
rect 29092 37120 29144 37126
rect 29092 37062 29144 37068
rect 28724 36916 28776 36922
rect 28724 36858 28776 36864
rect 28724 36712 28776 36718
rect 28722 36680 28724 36689
rect 28776 36680 28778 36689
rect 28722 36615 28778 36624
rect 28908 36644 28960 36650
rect 28908 36586 28960 36592
rect 28722 36408 28778 36417
rect 28920 36378 28948 36586
rect 28998 36544 29054 36553
rect 28998 36479 29054 36488
rect 28722 36343 28778 36352
rect 28908 36372 28960 36378
rect 28632 36168 28684 36174
rect 28632 36110 28684 36116
rect 28644 35873 28672 36110
rect 28736 36038 28764 36343
rect 28908 36314 28960 36320
rect 28814 36272 28870 36281
rect 28814 36207 28816 36216
rect 28868 36207 28870 36216
rect 28816 36178 28868 36184
rect 28724 36032 28776 36038
rect 28724 35974 28776 35980
rect 28630 35864 28686 35873
rect 28630 35799 28686 35808
rect 28538 35728 28594 35737
rect 28538 35663 28540 35672
rect 28592 35663 28594 35672
rect 28540 35634 28592 35640
rect 28644 35630 28672 35799
rect 28736 35766 28764 35974
rect 28724 35760 28776 35766
rect 28724 35702 28776 35708
rect 28632 35624 28684 35630
rect 28632 35566 28684 35572
rect 28814 35592 28870 35601
rect 28814 35527 28870 35536
rect 28632 35488 28684 35494
rect 28632 35430 28684 35436
rect 28448 35284 28500 35290
rect 28448 35226 28500 35232
rect 28540 34740 28592 34746
rect 28540 34682 28592 34688
rect 28552 34610 28580 34682
rect 28644 34610 28672 35430
rect 28722 35320 28778 35329
rect 28722 35255 28778 35264
rect 28736 35018 28764 35255
rect 28828 35204 28856 35527
rect 28920 35494 28948 36314
rect 29012 36242 29040 36479
rect 29000 36236 29052 36242
rect 29000 36178 29052 36184
rect 28998 36136 29054 36145
rect 28998 36071 29000 36080
rect 29052 36071 29054 36080
rect 29000 36042 29052 36048
rect 29104 35766 29132 37062
rect 29092 35760 29144 35766
rect 29092 35702 29144 35708
rect 28908 35488 28960 35494
rect 29092 35488 29144 35494
rect 28908 35430 28960 35436
rect 29090 35456 29092 35465
rect 29144 35456 29146 35465
rect 29090 35391 29146 35400
rect 29196 35290 29224 38508
rect 29381 38434 29409 38626
rect 29472 38554 29500 38898
rect 29564 38654 29592 42502
rect 29656 42090 29684 42706
rect 29644 42084 29696 42090
rect 29644 42026 29696 42032
rect 29840 41750 29868 51750
rect 29920 50380 29972 50386
rect 29920 50322 29972 50328
rect 29828 41744 29880 41750
rect 29828 41686 29880 41692
rect 29736 41472 29788 41478
rect 29736 41414 29788 41420
rect 29932 41414 29960 50322
rect 30116 47054 30144 52838
rect 31116 48272 31168 48278
rect 31116 48214 31168 48220
rect 30472 48068 30524 48074
rect 30472 48010 30524 48016
rect 30104 47048 30156 47054
rect 30104 46990 30156 46996
rect 30484 46986 30512 48010
rect 31128 47462 31156 48214
rect 31116 47456 31168 47462
rect 31116 47398 31168 47404
rect 31128 46986 31156 47398
rect 31220 47054 31248 52838
rect 31852 48000 31904 48006
rect 31852 47942 31904 47948
rect 31668 47456 31720 47462
rect 31668 47398 31720 47404
rect 31300 47184 31352 47190
rect 31300 47126 31352 47132
rect 31208 47048 31260 47054
rect 31208 46990 31260 46996
rect 30012 46980 30064 46986
rect 30012 46922 30064 46928
rect 30472 46980 30524 46986
rect 30472 46922 30524 46928
rect 31116 46980 31168 46986
rect 31116 46922 31168 46928
rect 30024 46646 30052 46922
rect 30484 46714 30512 46922
rect 30932 46912 30984 46918
rect 30932 46854 30984 46860
rect 30472 46708 30524 46714
rect 30472 46650 30524 46656
rect 30012 46640 30064 46646
rect 30012 46582 30064 46588
rect 30840 44192 30892 44198
rect 30840 44134 30892 44140
rect 30012 43920 30064 43926
rect 30012 43862 30064 43868
rect 30024 42702 30052 43862
rect 30472 43716 30524 43722
rect 30472 43658 30524 43664
rect 30196 43104 30248 43110
rect 30196 43046 30248 43052
rect 30012 42696 30064 42702
rect 30012 42638 30064 42644
rect 30208 42548 30236 43046
rect 30286 42800 30342 42809
rect 30286 42735 30342 42744
rect 30300 42702 30328 42735
rect 30288 42696 30340 42702
rect 30288 42638 30340 42644
rect 30288 42560 30340 42566
rect 30208 42520 30288 42548
rect 30288 42502 30340 42508
rect 30300 42362 30328 42502
rect 30288 42356 30340 42362
rect 30288 42298 30340 42304
rect 30196 42084 30248 42090
rect 30196 42026 30248 42032
rect 30012 42016 30064 42022
rect 30012 41958 30064 41964
rect 29644 40384 29696 40390
rect 29644 40326 29696 40332
rect 29656 39030 29684 40326
rect 29748 40118 29776 41414
rect 29840 41386 29960 41414
rect 29840 40390 29868 41386
rect 29920 40928 29972 40934
rect 29920 40870 29972 40876
rect 29828 40384 29880 40390
rect 29828 40326 29880 40332
rect 29736 40112 29788 40118
rect 29736 40054 29788 40060
rect 29736 39296 29788 39302
rect 29736 39238 29788 39244
rect 29748 39030 29776 39238
rect 29644 39024 29696 39030
rect 29644 38966 29696 38972
rect 29736 39024 29788 39030
rect 29736 38966 29788 38972
rect 29748 38894 29776 38966
rect 29736 38888 29788 38894
rect 29736 38830 29788 38836
rect 29736 38752 29788 38758
rect 29828 38752 29880 38758
rect 29736 38694 29788 38700
rect 29826 38720 29828 38729
rect 29880 38720 29882 38729
rect 29564 38626 29684 38654
rect 29460 38548 29512 38554
rect 29460 38490 29512 38496
rect 29381 38406 29500 38434
rect 29472 38332 29500 38406
rect 29472 38304 29592 38332
rect 29564 38196 29592 38304
rect 29380 38168 29592 38196
rect 29276 37936 29328 37942
rect 29276 37878 29328 37884
rect 29288 37777 29316 37878
rect 29274 37768 29330 37777
rect 29274 37703 29330 37712
rect 29276 36576 29328 36582
rect 29276 36518 29328 36524
rect 29288 36009 29316 36518
rect 29274 36000 29330 36009
rect 29274 35935 29330 35944
rect 29380 35850 29408 38168
rect 29458 38040 29514 38049
rect 29656 37992 29684 38626
rect 29748 38486 29776 38694
rect 29826 38655 29882 38664
rect 29828 38548 29880 38554
rect 29828 38490 29880 38496
rect 29736 38480 29788 38486
rect 29736 38422 29788 38428
rect 29458 37975 29514 37984
rect 29472 37942 29500 37975
rect 29564 37964 29684 37992
rect 29734 38040 29790 38049
rect 29840 38010 29868 38490
rect 29932 38350 29960 40870
rect 29920 38344 29972 38350
rect 29920 38286 29972 38292
rect 29920 38208 29972 38214
rect 29920 38150 29972 38156
rect 29734 37975 29790 37984
rect 29828 38004 29880 38010
rect 29460 37936 29512 37942
rect 29460 37878 29512 37884
rect 29458 36408 29514 36417
rect 29458 36343 29514 36352
rect 29472 36174 29500 36343
rect 29460 36168 29512 36174
rect 29460 36110 29512 36116
rect 29288 35822 29408 35850
rect 29184 35284 29236 35290
rect 29184 35226 29236 35232
rect 29092 35216 29144 35222
rect 28828 35176 29092 35204
rect 29092 35158 29144 35164
rect 28998 35048 29054 35057
rect 28724 35012 28776 35018
rect 28998 34983 29054 34992
rect 28724 34954 28776 34960
rect 29012 34950 29040 34983
rect 29000 34944 29052 34950
rect 29000 34886 29052 34892
rect 29012 34626 29040 34886
rect 28540 34604 28592 34610
rect 28540 34546 28592 34552
rect 28632 34604 28684 34610
rect 28632 34546 28684 34552
rect 28920 34598 29040 34626
rect 29288 34610 29316 35822
rect 29460 35624 29512 35630
rect 29460 35566 29512 35572
rect 29366 35456 29422 35465
rect 29366 35391 29422 35400
rect 29276 34604 29328 34610
rect 28356 34128 28408 34134
rect 28356 34070 28408 34076
rect 28448 33856 28500 33862
rect 28448 33798 28500 33804
rect 28264 33652 28316 33658
rect 28264 33594 28316 33600
rect 28262 33144 28318 33153
rect 28262 33079 28318 33088
rect 28276 28082 28304 33079
rect 28460 32910 28488 33798
rect 28448 32904 28500 32910
rect 28448 32846 28500 32852
rect 28356 31680 28408 31686
rect 28356 31622 28408 31628
rect 28368 31346 28396 31622
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28356 29572 28408 29578
rect 28356 29514 28408 29520
rect 28368 28558 28396 29514
rect 28356 28552 28408 28558
rect 28356 28494 28408 28500
rect 28264 28076 28316 28082
rect 28264 28018 28316 28024
rect 28172 28008 28224 28014
rect 28172 27950 28224 27956
rect 28356 28008 28408 28014
rect 28356 27950 28408 27956
rect 28080 27872 28132 27878
rect 28080 27814 28132 27820
rect 28368 27606 28396 27950
rect 28632 27872 28684 27878
rect 28632 27814 28684 27820
rect 28356 27600 28408 27606
rect 28356 27542 28408 27548
rect 28644 27538 28672 27814
rect 28632 27532 28684 27538
rect 28632 27474 28684 27480
rect 28264 26784 28316 26790
rect 28264 26726 28316 26732
rect 28276 26518 28304 26726
rect 28264 26512 28316 26518
rect 28264 26454 28316 26460
rect 28276 25770 28304 26454
rect 28264 25764 28316 25770
rect 28264 25706 28316 25712
rect 28172 25288 28224 25294
rect 28172 25230 28224 25236
rect 28184 24818 28212 25230
rect 28540 25220 28592 25226
rect 28540 25162 28592 25168
rect 28552 24954 28580 25162
rect 28540 24948 28592 24954
rect 28540 24890 28592 24896
rect 28172 24812 28224 24818
rect 28172 24754 28224 24760
rect 28184 24410 28212 24754
rect 28172 24404 28224 24410
rect 28172 24346 28224 24352
rect 28920 23526 28948 34598
rect 29276 34546 29328 34552
rect 29092 34400 29144 34406
rect 29092 34342 29144 34348
rect 29104 33522 29132 34342
rect 29092 33516 29144 33522
rect 29092 33458 29144 33464
rect 29090 33416 29146 33425
rect 29000 33380 29052 33386
rect 29090 33351 29146 33360
rect 29000 33322 29052 33328
rect 29012 33114 29040 33322
rect 29000 33108 29052 33114
rect 29000 33050 29052 33056
rect 29000 25900 29052 25906
rect 29000 25842 29052 25848
rect 29012 25498 29040 25842
rect 29000 25492 29052 25498
rect 29000 25434 29052 25440
rect 29000 25356 29052 25362
rect 29000 25298 29052 25304
rect 28908 23520 28960 23526
rect 28908 23462 28960 23468
rect 28908 23316 28960 23322
rect 28908 23258 28960 23264
rect 28724 23180 28776 23186
rect 28724 23122 28776 23128
rect 28172 22432 28224 22438
rect 28172 22374 28224 22380
rect 27908 22066 28028 22094
rect 27804 21888 27856 21894
rect 27804 21830 27856 21836
rect 27528 21684 27580 21690
rect 27528 21626 27580 21632
rect 27434 21584 27490 21593
rect 27816 21554 27844 21830
rect 27434 21519 27490 21528
rect 27804 21548 27856 21554
rect 27448 21486 27476 21519
rect 27804 21490 27856 21496
rect 27436 21480 27488 21486
rect 27436 21422 27488 21428
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27160 20596 27212 20602
rect 27160 20538 27212 20544
rect 27172 18834 27200 20538
rect 27528 20392 27580 20398
rect 27526 20360 27528 20369
rect 27580 20360 27582 20369
rect 27526 20295 27582 20304
rect 27540 19378 27568 20295
rect 27632 20058 27660 21286
rect 27816 20602 27844 21490
rect 27804 20596 27856 20602
rect 27804 20538 27856 20544
rect 27620 20052 27672 20058
rect 27620 19994 27672 20000
rect 27632 19378 27660 19994
rect 27804 19848 27856 19854
rect 27804 19790 27856 19796
rect 27528 19372 27580 19378
rect 27528 19314 27580 19320
rect 27620 19372 27672 19378
rect 27620 19314 27672 19320
rect 27160 18828 27212 18834
rect 27160 18770 27212 18776
rect 27436 18352 27488 18358
rect 27436 18294 27488 18300
rect 27448 17241 27476 18294
rect 27540 18154 27568 19314
rect 27632 18834 27660 19314
rect 27816 19310 27844 19790
rect 27804 19304 27856 19310
rect 27804 19246 27856 19252
rect 27816 18834 27844 19246
rect 27620 18828 27672 18834
rect 27620 18770 27672 18776
rect 27804 18828 27856 18834
rect 27804 18770 27856 18776
rect 27620 18692 27672 18698
rect 27620 18634 27672 18640
rect 27528 18148 27580 18154
rect 27528 18090 27580 18096
rect 27632 17762 27660 18634
rect 27710 17776 27766 17785
rect 27528 17740 27580 17746
rect 27632 17734 27710 17762
rect 27710 17711 27712 17720
rect 27528 17682 27580 17688
rect 27764 17711 27766 17720
rect 27712 17682 27764 17688
rect 27434 17232 27490 17241
rect 27434 17167 27490 17176
rect 27448 16726 27476 17167
rect 27436 16720 27488 16726
rect 27436 16662 27488 16668
rect 27540 16640 27568 17682
rect 27908 17626 27936 22066
rect 28184 22030 28212 22374
rect 28540 22092 28592 22098
rect 28540 22034 28592 22040
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28552 21486 28580 22034
rect 28540 21480 28592 21486
rect 28632 21480 28684 21486
rect 28540 21422 28592 21428
rect 28630 21448 28632 21457
rect 28684 21448 28686 21457
rect 28552 21010 28580 21422
rect 28736 21418 28764 23122
rect 28816 21888 28868 21894
rect 28816 21830 28868 21836
rect 28828 21486 28856 21830
rect 28816 21480 28868 21486
rect 28816 21422 28868 21428
rect 28630 21383 28686 21392
rect 28724 21412 28776 21418
rect 28644 21078 28672 21383
rect 28724 21354 28776 21360
rect 28632 21072 28684 21078
rect 28632 21014 28684 21020
rect 28540 21004 28592 21010
rect 28540 20946 28592 20952
rect 28920 20890 28948 23258
rect 28644 20874 28948 20890
rect 28632 20868 28948 20874
rect 28684 20862 28948 20868
rect 28632 20810 28684 20816
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28354 19544 28410 19553
rect 28080 19508 28132 19514
rect 28354 19479 28410 19488
rect 28080 19450 28132 19456
rect 28092 18358 28120 19450
rect 28368 19446 28396 19479
rect 28356 19440 28408 19446
rect 28356 19382 28408 19388
rect 28460 19378 28488 19790
rect 28448 19372 28500 19378
rect 28644 19357 28672 20810
rect 28816 20596 28868 20602
rect 28816 20538 28868 20544
rect 28828 20369 28856 20538
rect 28814 20360 28870 20369
rect 28814 20295 28870 20304
rect 28448 19314 28500 19320
rect 28630 19348 28686 19357
rect 28630 19283 28686 19292
rect 28264 19236 28316 19242
rect 28264 19178 28316 19184
rect 28172 18760 28224 18766
rect 28172 18702 28224 18708
rect 28276 18714 28304 19178
rect 28448 19168 28500 19174
rect 28368 19128 28448 19156
rect 28368 18834 28396 19128
rect 28448 19110 28500 19116
rect 28632 18964 28684 18970
rect 28632 18906 28684 18912
rect 28448 18896 28500 18902
rect 28448 18838 28500 18844
rect 28356 18828 28408 18834
rect 28356 18770 28408 18776
rect 28080 18352 28132 18358
rect 28080 18294 28132 18300
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 28000 17882 28028 18226
rect 27988 17876 28040 17882
rect 27988 17818 28040 17824
rect 27816 17598 27936 17626
rect 27712 17128 27764 17134
rect 27712 17070 27764 17076
rect 27724 16998 27752 17070
rect 27712 16992 27764 16998
rect 27712 16934 27764 16940
rect 27540 16612 27660 16640
rect 27068 16584 27120 16590
rect 27068 16526 27120 16532
rect 27080 14958 27108 16526
rect 27528 16516 27580 16522
rect 27528 16458 27580 16464
rect 27436 16448 27488 16454
rect 27436 16390 27488 16396
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 27068 14952 27120 14958
rect 27068 14894 27120 14900
rect 27172 14890 27200 16050
rect 27356 15978 27384 16050
rect 27344 15972 27396 15978
rect 27344 15914 27396 15920
rect 27448 15162 27476 16390
rect 27436 15156 27488 15162
rect 27436 15098 27488 15104
rect 27448 14958 27476 15098
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27160 14884 27212 14890
rect 27160 14826 27212 14832
rect 27252 14408 27304 14414
rect 27252 14350 27304 14356
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 27068 13320 27120 13326
rect 27068 13262 27120 13268
rect 27080 11642 27108 13262
rect 27172 12918 27200 13670
rect 27264 13190 27292 14350
rect 27540 13818 27568 16458
rect 27632 16454 27660 16612
rect 27816 16590 27844 17598
rect 27896 17536 27948 17542
rect 27988 17536 28040 17542
rect 27896 17478 27948 17484
rect 27986 17504 27988 17513
rect 28040 17504 28042 17513
rect 27908 17338 27936 17478
rect 27986 17439 28042 17448
rect 27896 17332 27948 17338
rect 27896 17274 27948 17280
rect 27804 16584 27856 16590
rect 27804 16526 27856 16532
rect 27620 16448 27672 16454
rect 27620 16390 27672 16396
rect 27632 15366 27660 16390
rect 27896 15496 27948 15502
rect 27896 15438 27948 15444
rect 27620 15360 27672 15366
rect 27620 15302 27672 15308
rect 27710 15328 27766 15337
rect 27710 15263 27766 15272
rect 27620 14952 27672 14958
rect 27618 14920 27620 14929
rect 27672 14920 27674 14929
rect 27618 14855 27674 14864
rect 27724 14414 27752 15263
rect 27804 14952 27856 14958
rect 27804 14894 27856 14900
rect 27816 14618 27844 14894
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 27724 13938 27752 14350
rect 27712 13932 27764 13938
rect 27712 13874 27764 13880
rect 27540 13790 27752 13818
rect 27344 13728 27396 13734
rect 27344 13670 27396 13676
rect 27356 13530 27384 13670
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27160 12912 27212 12918
rect 27160 12854 27212 12860
rect 27436 12912 27488 12918
rect 27724 12889 27752 13790
rect 27436 12854 27488 12860
rect 27710 12880 27766 12889
rect 27172 12306 27200 12854
rect 27344 12640 27396 12646
rect 27344 12582 27396 12588
rect 27160 12300 27212 12306
rect 27160 12242 27212 12248
rect 27356 11898 27384 12582
rect 27344 11892 27396 11898
rect 27344 11834 27396 11840
rect 27080 11614 27292 11642
rect 27160 11552 27212 11558
rect 27160 11494 27212 11500
rect 27172 11354 27200 11494
rect 27160 11348 27212 11354
rect 27160 11290 27212 11296
rect 27068 11144 27120 11150
rect 27068 11086 27120 11092
rect 26976 9444 27028 9450
rect 26976 9386 27028 9392
rect 26884 7744 26936 7750
rect 26884 7686 26936 7692
rect 26896 7478 26924 7686
rect 26884 7472 26936 7478
rect 26884 7414 26936 7420
rect 27080 6730 27108 11086
rect 27172 10742 27200 11290
rect 27160 10736 27212 10742
rect 27160 10678 27212 10684
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 27068 6724 27120 6730
rect 27068 6666 27120 6672
rect 27080 6458 27108 6666
rect 27068 6452 27120 6458
rect 27068 6394 27120 6400
rect 27172 5778 27200 9522
rect 27264 9058 27292 11614
rect 27448 11150 27476 12854
rect 27710 12815 27766 12824
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27436 11144 27488 11150
rect 27436 11086 27488 11092
rect 27344 11008 27396 11014
rect 27344 10950 27396 10956
rect 27356 10674 27384 10950
rect 27344 10668 27396 10674
rect 27344 10610 27396 10616
rect 27528 10464 27580 10470
rect 27528 10406 27580 10412
rect 27540 10130 27568 10406
rect 27528 10124 27580 10130
rect 27528 10066 27580 10072
rect 27632 9926 27660 11494
rect 27620 9920 27672 9926
rect 27620 9862 27672 9868
rect 27434 9480 27490 9489
rect 27434 9415 27490 9424
rect 27264 9030 27384 9058
rect 27252 8900 27304 8906
rect 27252 8842 27304 8848
rect 27264 7546 27292 8842
rect 27252 7540 27304 7546
rect 27252 7482 27304 7488
rect 27356 6866 27384 9030
rect 27448 8974 27476 9415
rect 27632 8974 27660 9862
rect 27436 8968 27488 8974
rect 27436 8910 27488 8916
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 27632 8566 27660 8910
rect 27620 8560 27672 8566
rect 27620 8502 27672 8508
rect 27620 8016 27672 8022
rect 27620 7958 27672 7964
rect 27344 6860 27396 6866
rect 27344 6802 27396 6808
rect 27436 6316 27488 6322
rect 27436 6258 27488 6264
rect 27160 5772 27212 5778
rect 27160 5714 27212 5720
rect 26884 5092 26936 5098
rect 26884 5034 26936 5040
rect 26896 4758 26924 5034
rect 26884 4752 26936 4758
rect 26884 4694 26936 4700
rect 27448 4690 27476 6258
rect 27632 5370 27660 7958
rect 27620 5364 27672 5370
rect 27620 5306 27672 5312
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 26700 4140 26752 4146
rect 26700 4082 26752 4088
rect 25504 4072 25556 4078
rect 25504 4014 25556 4020
rect 25872 4072 25924 4078
rect 25872 4014 25924 4020
rect 25412 3120 25464 3126
rect 25412 3062 25464 3068
rect 25228 2848 25280 2854
rect 25228 2790 25280 2796
rect 25056 2746 25176 2774
rect 25056 2446 25084 2746
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 25240 800 25268 2790
rect 25884 2446 25912 4014
rect 26252 3058 26280 4082
rect 26790 3768 26846 3777
rect 26790 3703 26792 3712
rect 26844 3703 26846 3712
rect 26792 3674 26844 3680
rect 26332 3460 26384 3466
rect 26332 3402 26384 3408
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 25964 2848 26016 2854
rect 25964 2790 26016 2796
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 25596 2304 25648 2310
rect 25596 2246 25648 2252
rect 25608 800 25636 2246
rect 25976 800 26004 2790
rect 26344 2446 26372 3402
rect 26804 3058 26832 3674
rect 27724 3466 27752 12815
rect 27908 12481 27936 15438
rect 28000 15348 28028 17439
rect 28184 16250 28212 18702
rect 28276 18698 28396 18714
rect 28276 18692 28408 18698
rect 28276 18686 28356 18692
rect 28356 18634 28408 18640
rect 28264 18624 28316 18630
rect 28264 18566 28316 18572
rect 28172 16244 28224 16250
rect 28172 16186 28224 16192
rect 28276 15978 28304 18566
rect 28356 18352 28408 18358
rect 28354 18320 28356 18329
rect 28408 18320 28410 18329
rect 28354 18255 28410 18264
rect 28356 17740 28408 17746
rect 28356 17682 28408 17688
rect 28368 16522 28396 17682
rect 28460 17202 28488 18838
rect 28540 18692 28592 18698
rect 28540 18634 28592 18640
rect 28552 18290 28580 18634
rect 28644 18358 28672 18906
rect 28722 18864 28778 18873
rect 28722 18799 28778 18808
rect 28632 18352 28684 18358
rect 28632 18294 28684 18300
rect 28540 18284 28592 18290
rect 28540 18226 28592 18232
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 28356 16516 28408 16522
rect 28356 16458 28408 16464
rect 28552 16250 28580 18226
rect 28632 18148 28684 18154
rect 28632 18090 28684 18096
rect 28644 17377 28672 18090
rect 28630 17368 28686 17377
rect 28630 17303 28686 17312
rect 28632 16584 28684 16590
rect 28632 16526 28684 16532
rect 28540 16244 28592 16250
rect 28540 16186 28592 16192
rect 28264 15972 28316 15978
rect 28264 15914 28316 15920
rect 28448 15904 28500 15910
rect 28448 15846 28500 15852
rect 28078 15600 28134 15609
rect 28078 15535 28134 15544
rect 28092 15502 28120 15535
rect 28080 15496 28132 15502
rect 28080 15438 28132 15444
rect 28000 15320 28120 15348
rect 27988 13932 28040 13938
rect 27988 13874 28040 13880
rect 28000 12986 28028 13874
rect 27988 12980 28040 12986
rect 27988 12922 28040 12928
rect 27894 12472 27950 12481
rect 27816 12416 27894 12434
rect 27816 12407 27950 12416
rect 27816 12406 27936 12407
rect 27816 3738 27844 12406
rect 27986 12064 28042 12073
rect 27986 11999 28042 12008
rect 28000 11218 28028 11999
rect 27988 11212 28040 11218
rect 27988 11154 28040 11160
rect 27988 10464 28040 10470
rect 27988 10406 28040 10412
rect 27896 9988 27948 9994
rect 27896 9930 27948 9936
rect 27908 9586 27936 9930
rect 27896 9580 27948 9586
rect 27896 9522 27948 9528
rect 28000 8634 28028 10406
rect 27988 8628 28040 8634
rect 27988 8570 28040 8576
rect 27988 7268 28040 7274
rect 27988 7210 28040 7216
rect 27896 6860 27948 6866
rect 27896 6802 27948 6808
rect 27908 3942 27936 6802
rect 28000 4078 28028 7210
rect 27988 4072 28040 4078
rect 27988 4014 28040 4020
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 28092 3738 28120 15320
rect 28262 15192 28318 15201
rect 28262 15127 28318 15136
rect 28356 15156 28408 15162
rect 28276 15026 28304 15127
rect 28356 15098 28408 15104
rect 28264 15020 28316 15026
rect 28264 14962 28316 14968
rect 28172 14816 28224 14822
rect 28172 14758 28224 14764
rect 28184 14618 28212 14758
rect 28172 14612 28224 14618
rect 28172 14554 28224 14560
rect 28368 13410 28396 15098
rect 28460 14346 28488 15846
rect 28644 15706 28672 16526
rect 28632 15700 28684 15706
rect 28632 15642 28684 15648
rect 28540 15496 28592 15502
rect 28540 15438 28592 15444
rect 28552 15026 28580 15438
rect 28632 15360 28684 15366
rect 28632 15302 28684 15308
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28552 14414 28580 14962
rect 28540 14408 28592 14414
rect 28540 14350 28592 14356
rect 28448 14340 28500 14346
rect 28448 14282 28500 14288
rect 28552 14278 28580 14350
rect 28540 14272 28592 14278
rect 28540 14214 28592 14220
rect 28368 13382 28488 13410
rect 28356 13320 28408 13326
rect 28356 13262 28408 13268
rect 28264 12096 28316 12102
rect 28264 12038 28316 12044
rect 28172 10668 28224 10674
rect 28172 10610 28224 10616
rect 28184 9178 28212 10610
rect 28276 10062 28304 12038
rect 28368 10266 28396 13262
rect 28460 12918 28488 13382
rect 28448 12912 28500 12918
rect 28448 12854 28500 12860
rect 28540 12300 28592 12306
rect 28540 12242 28592 12248
rect 28552 11694 28580 12242
rect 28540 11688 28592 11694
rect 28540 11630 28592 11636
rect 28644 11150 28672 15302
rect 28736 12730 28764 18799
rect 28816 18080 28868 18086
rect 28816 18022 28868 18028
rect 28828 17678 28856 18022
rect 28908 17740 28960 17746
rect 29012 17728 29040 25298
rect 29104 23322 29132 33351
rect 29184 23520 29236 23526
rect 29184 23462 29236 23468
rect 29092 23316 29144 23322
rect 29092 23258 29144 23264
rect 29092 21344 29144 21350
rect 29092 21286 29144 21292
rect 29104 21078 29132 21286
rect 29092 21072 29144 21078
rect 29092 21014 29144 21020
rect 29196 20466 29224 23462
rect 29380 22094 29408 35391
rect 29472 34610 29500 35566
rect 29460 34604 29512 34610
rect 29460 34546 29512 34552
rect 29564 34134 29592 37964
rect 29748 37942 29776 37975
rect 29828 37946 29880 37952
rect 29736 37936 29788 37942
rect 29642 37904 29698 37913
rect 29736 37878 29788 37884
rect 29642 37839 29644 37848
rect 29696 37839 29698 37848
rect 29828 37868 29880 37874
rect 29644 37810 29696 37816
rect 29828 37810 29880 37816
rect 29840 37670 29868 37810
rect 29828 37664 29880 37670
rect 29828 37606 29880 37612
rect 29840 37330 29868 37606
rect 29828 37324 29880 37330
rect 29828 37266 29880 37272
rect 29828 37120 29880 37126
rect 29828 37062 29880 37068
rect 29736 36780 29788 36786
rect 29736 36722 29788 36728
rect 29748 36122 29776 36722
rect 29656 36094 29776 36122
rect 29656 36038 29684 36094
rect 29644 36032 29696 36038
rect 29644 35974 29696 35980
rect 29736 36032 29788 36038
rect 29736 35974 29788 35980
rect 29644 35692 29696 35698
rect 29644 35634 29696 35640
rect 29656 35494 29684 35634
rect 29644 35488 29696 35494
rect 29644 35430 29696 35436
rect 29644 35216 29696 35222
rect 29644 35158 29696 35164
rect 29656 35086 29684 35158
rect 29644 35080 29696 35086
rect 29644 35022 29696 35028
rect 29748 35018 29776 35974
rect 29736 35012 29788 35018
rect 29736 34954 29788 34960
rect 29748 34746 29776 34954
rect 29736 34740 29788 34746
rect 29736 34682 29788 34688
rect 29642 34640 29698 34649
rect 29642 34575 29644 34584
rect 29696 34575 29698 34584
rect 29644 34546 29696 34552
rect 29552 34128 29604 34134
rect 29552 34070 29604 34076
rect 29460 34060 29512 34066
rect 29460 34002 29512 34008
rect 29472 33454 29500 34002
rect 29736 33516 29788 33522
rect 29736 33458 29788 33464
rect 29460 33448 29512 33454
rect 29460 33390 29512 33396
rect 29748 32570 29776 33458
rect 29736 32564 29788 32570
rect 29736 32506 29788 32512
rect 29552 28688 29604 28694
rect 29552 28630 29604 28636
rect 29288 22066 29408 22094
rect 29092 20460 29144 20466
rect 29092 20402 29144 20408
rect 29184 20460 29236 20466
rect 29184 20402 29236 20408
rect 29104 19514 29132 20402
rect 29196 19922 29224 20402
rect 29184 19916 29236 19922
rect 29184 19858 29236 19864
rect 29092 19508 29144 19514
rect 29092 19450 29144 19456
rect 29092 19372 29144 19378
rect 29092 19314 29144 19320
rect 29104 18329 29132 19314
rect 29184 19304 29236 19310
rect 29184 19246 29236 19252
rect 29196 18970 29224 19246
rect 29184 18964 29236 18970
rect 29184 18906 29236 18912
rect 29090 18320 29146 18329
rect 29288 18272 29316 22066
rect 29368 21548 29420 21554
rect 29368 21490 29420 21496
rect 29090 18255 29146 18264
rect 29196 18244 29316 18272
rect 29012 17700 29132 17728
rect 28908 17682 28960 17688
rect 28816 17672 28868 17678
rect 28920 17649 28948 17682
rect 28816 17614 28868 17620
rect 28906 17640 28962 17649
rect 28828 17490 28856 17614
rect 28906 17575 28962 17584
rect 29104 17542 29132 17700
rect 29092 17536 29144 17542
rect 28828 17462 28948 17490
rect 29092 17478 29144 17484
rect 28814 17368 28870 17377
rect 28814 17303 28870 17312
rect 28828 16114 28856 17303
rect 28920 17202 28948 17462
rect 28908 17196 28960 17202
rect 28908 17138 28960 17144
rect 29092 16720 29144 16726
rect 29092 16662 29144 16668
rect 28998 16280 29054 16289
rect 28998 16215 29054 16224
rect 29012 16182 29040 16215
rect 29000 16176 29052 16182
rect 29000 16118 29052 16124
rect 29104 16114 29132 16662
rect 28816 16108 28868 16114
rect 28816 16050 28868 16056
rect 29092 16108 29144 16114
rect 29092 16050 29144 16056
rect 28816 15972 28868 15978
rect 28816 15914 28868 15920
rect 28828 15366 28856 15914
rect 29196 15722 29224 18244
rect 29276 18148 29328 18154
rect 29276 18090 29328 18096
rect 29104 15694 29224 15722
rect 28908 15564 28960 15570
rect 28908 15506 28960 15512
rect 28920 15450 28948 15506
rect 28920 15422 29040 15450
rect 28816 15360 28868 15366
rect 28816 15302 28868 15308
rect 29012 15162 29040 15422
rect 29000 15156 29052 15162
rect 29000 15098 29052 15104
rect 28908 15088 28960 15094
rect 28908 15030 28960 15036
rect 28920 14550 28948 15030
rect 29104 14906 29132 15694
rect 29288 15434 29316 18090
rect 29380 17746 29408 21490
rect 29460 20256 29512 20262
rect 29460 20198 29512 20204
rect 29472 19961 29500 20198
rect 29458 19952 29514 19961
rect 29458 19887 29514 19896
rect 29564 19802 29592 28630
rect 29840 28558 29868 37062
rect 29932 35578 29960 38150
rect 30024 35698 30052 41958
rect 30102 41712 30158 41721
rect 30102 41647 30104 41656
rect 30156 41647 30158 41656
rect 30104 41618 30156 41624
rect 30104 41540 30156 41546
rect 30104 41482 30156 41488
rect 30116 41070 30144 41482
rect 30208 41138 30236 42026
rect 30196 41132 30248 41138
rect 30196 41074 30248 41080
rect 30104 41064 30156 41070
rect 30300 41018 30328 42298
rect 30380 42288 30432 42294
rect 30378 42256 30380 42265
rect 30432 42256 30434 42265
rect 30378 42191 30434 42200
rect 30484 41546 30512 43658
rect 30564 43648 30616 43654
rect 30564 43590 30616 43596
rect 30576 42838 30604 43590
rect 30748 43104 30800 43110
rect 30748 43046 30800 43052
rect 30760 42906 30788 43046
rect 30748 42900 30800 42906
rect 30748 42842 30800 42848
rect 30564 42832 30616 42838
rect 30564 42774 30616 42780
rect 30576 42226 30604 42774
rect 30564 42220 30616 42226
rect 30564 42162 30616 42168
rect 30576 41614 30604 42162
rect 30564 41608 30616 41614
rect 30564 41550 30616 41556
rect 30472 41540 30524 41546
rect 30472 41482 30524 41488
rect 30576 41274 30604 41550
rect 30564 41268 30616 41274
rect 30564 41210 30616 41216
rect 30156 41012 30420 41018
rect 30104 41006 30420 41012
rect 30116 40990 30420 41006
rect 30116 40941 30144 40990
rect 30196 40928 30248 40934
rect 30196 40870 30248 40876
rect 30104 40588 30156 40594
rect 30104 40530 30156 40536
rect 30116 40186 30144 40530
rect 30104 40180 30156 40186
rect 30104 40122 30156 40128
rect 30208 39982 30236 40870
rect 30288 40656 30340 40662
rect 30288 40598 30340 40604
rect 30196 39976 30248 39982
rect 30196 39918 30248 39924
rect 30104 38276 30156 38282
rect 30104 38218 30156 38224
rect 30116 38010 30144 38218
rect 30196 38208 30248 38214
rect 30196 38150 30248 38156
rect 30104 38004 30156 38010
rect 30104 37946 30156 37952
rect 30104 37460 30156 37466
rect 30104 37402 30156 37408
rect 30116 37194 30144 37402
rect 30208 37330 30236 38150
rect 30300 37346 30328 40598
rect 30392 37466 30420 40990
rect 30576 40662 30604 41210
rect 30760 41002 30788 42842
rect 30852 42770 30880 44134
rect 30840 42764 30892 42770
rect 30840 42706 30892 42712
rect 30852 42566 30880 42706
rect 30840 42560 30892 42566
rect 30840 42502 30892 42508
rect 30748 40996 30800 41002
rect 30748 40938 30800 40944
rect 30564 40656 30616 40662
rect 30564 40598 30616 40604
rect 30576 40050 30604 40598
rect 30564 40044 30616 40050
rect 30616 40004 30696 40032
rect 30564 39986 30616 39992
rect 30472 39840 30524 39846
rect 30472 39782 30524 39788
rect 30380 37460 30432 37466
rect 30380 37402 30432 37408
rect 30196 37324 30248 37330
rect 30300 37318 30420 37346
rect 30196 37266 30248 37272
rect 30392 37262 30420 37318
rect 30380 37256 30432 37262
rect 30286 37224 30342 37233
rect 30104 37188 30156 37194
rect 30380 37198 30432 37204
rect 30286 37159 30342 37168
rect 30104 37130 30156 37136
rect 30012 35692 30064 35698
rect 30012 35634 30064 35640
rect 29932 35550 30052 35578
rect 29920 34740 29972 34746
rect 29920 34682 29972 34688
rect 29932 34610 29960 34682
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 29932 32774 29960 34546
rect 29920 32768 29972 32774
rect 29920 32710 29972 32716
rect 29932 28762 29960 32710
rect 29920 28756 29972 28762
rect 29920 28698 29972 28704
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 29828 27464 29880 27470
rect 29828 27406 29880 27412
rect 29644 24268 29696 24274
rect 29644 24210 29696 24216
rect 29656 22642 29684 24210
rect 29644 22636 29696 22642
rect 29644 22578 29696 22584
rect 29656 22438 29684 22578
rect 29644 22432 29696 22438
rect 29644 22374 29696 22380
rect 29840 22094 29868 27406
rect 30024 25362 30052 35550
rect 30116 34950 30144 37130
rect 30300 37126 30328 37159
rect 30288 37120 30340 37126
rect 30288 37062 30340 37068
rect 30288 35692 30340 35698
rect 30288 35634 30340 35640
rect 30300 35562 30328 35634
rect 30288 35556 30340 35562
rect 30288 35498 30340 35504
rect 30380 35216 30432 35222
rect 30380 35158 30432 35164
rect 30392 35018 30420 35158
rect 30380 35012 30432 35018
rect 30380 34954 30432 34960
rect 30104 34944 30156 34950
rect 30104 34886 30156 34892
rect 30116 29578 30144 34886
rect 30378 34776 30434 34785
rect 30378 34711 30434 34720
rect 30392 34610 30420 34711
rect 30484 34610 30512 39782
rect 30564 39432 30616 39438
rect 30668 39420 30696 40004
rect 30944 39914 30972 46854
rect 31208 46368 31260 46374
rect 31208 46310 31260 46316
rect 31220 45082 31248 46310
rect 31208 45076 31260 45082
rect 31208 45018 31260 45024
rect 31024 44192 31076 44198
rect 31024 44134 31076 44140
rect 31036 42809 31064 44134
rect 31022 42800 31078 42809
rect 31022 42735 31078 42744
rect 31208 42152 31260 42158
rect 31208 42094 31260 42100
rect 31220 41682 31248 42094
rect 31208 41676 31260 41682
rect 31208 41618 31260 41624
rect 31312 40118 31340 47126
rect 31680 47054 31708 47398
rect 31864 47258 31892 47942
rect 32036 47524 32088 47530
rect 32036 47466 32088 47472
rect 31852 47252 31904 47258
rect 31852 47194 31904 47200
rect 32048 47054 32076 47466
rect 31668 47048 31720 47054
rect 31668 46990 31720 46996
rect 32036 47048 32088 47054
rect 32036 46990 32088 46996
rect 31392 46096 31444 46102
rect 31392 46038 31444 46044
rect 31404 45898 31432 46038
rect 31392 45892 31444 45898
rect 31392 45834 31444 45840
rect 31852 45280 31904 45286
rect 31852 45222 31904 45228
rect 31484 43104 31536 43110
rect 31484 43046 31536 43052
rect 31392 42356 31444 42362
rect 31392 42298 31444 42304
rect 31404 41614 31432 42298
rect 31496 41721 31524 43046
rect 31576 42560 31628 42566
rect 31576 42502 31628 42508
rect 31588 42158 31616 42502
rect 31576 42152 31628 42158
rect 31576 42094 31628 42100
rect 31482 41712 31538 41721
rect 31482 41647 31538 41656
rect 31392 41608 31444 41614
rect 31392 41550 31444 41556
rect 31300 40112 31352 40118
rect 31300 40054 31352 40060
rect 30932 39908 30984 39914
rect 30932 39850 30984 39856
rect 31404 39642 31432 41550
rect 31482 40080 31538 40089
rect 31482 40015 31484 40024
rect 31536 40015 31538 40024
rect 31484 39986 31536 39992
rect 31392 39636 31444 39642
rect 31392 39578 31444 39584
rect 30616 39392 30696 39420
rect 30564 39374 30616 39380
rect 30668 39098 30696 39392
rect 30748 39296 30800 39302
rect 30748 39238 30800 39244
rect 31208 39296 31260 39302
rect 31208 39238 31260 39244
rect 30656 39092 30708 39098
rect 30656 39034 30708 39040
rect 30564 39024 30616 39030
rect 30564 38966 30616 38972
rect 30576 37874 30604 38966
rect 30564 37868 30616 37874
rect 30564 37810 30616 37816
rect 30656 35080 30708 35086
rect 30656 35022 30708 35028
rect 30564 34944 30616 34950
rect 30562 34912 30564 34921
rect 30616 34912 30618 34921
rect 30562 34847 30618 34856
rect 30380 34604 30432 34610
rect 30380 34546 30432 34552
rect 30472 34604 30524 34610
rect 30472 34546 30524 34552
rect 30380 34468 30432 34474
rect 30380 34410 30432 34416
rect 30288 34128 30340 34134
rect 30288 34070 30340 34076
rect 30300 33998 30328 34070
rect 30392 33998 30420 34410
rect 30668 34066 30696 35022
rect 30656 34060 30708 34066
rect 30656 34002 30708 34008
rect 30288 33992 30340 33998
rect 30288 33934 30340 33940
rect 30380 33992 30432 33998
rect 30380 33934 30432 33940
rect 30564 33856 30616 33862
rect 30564 33798 30616 33804
rect 30380 31136 30432 31142
rect 30380 31078 30432 31084
rect 30104 29572 30156 29578
rect 30104 29514 30156 29520
rect 30392 29306 30420 31078
rect 30472 29504 30524 29510
rect 30472 29446 30524 29452
rect 30484 29306 30512 29446
rect 30380 29300 30432 29306
rect 30380 29242 30432 29248
rect 30472 29300 30524 29306
rect 30472 29242 30524 29248
rect 30104 28416 30156 28422
rect 30104 28358 30156 28364
rect 30116 27470 30144 28358
rect 30104 27464 30156 27470
rect 30104 27406 30156 27412
rect 30012 25356 30064 25362
rect 30012 25298 30064 25304
rect 30012 23724 30064 23730
rect 30012 23666 30064 23672
rect 30024 22778 30052 23666
rect 30196 23520 30248 23526
rect 30196 23462 30248 23468
rect 30208 23050 30236 23462
rect 30380 23112 30432 23118
rect 30380 23054 30432 23060
rect 30196 23044 30248 23050
rect 30196 22986 30248 22992
rect 30012 22772 30064 22778
rect 30012 22714 30064 22720
rect 30392 22642 30420 23054
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 30288 22160 30340 22166
rect 30288 22102 30340 22108
rect 29840 22066 29960 22094
rect 29828 21888 29880 21894
rect 29828 21830 29880 21836
rect 29840 21690 29868 21830
rect 29828 21684 29880 21690
rect 29828 21626 29880 21632
rect 29736 20800 29788 20806
rect 29736 20742 29788 20748
rect 29644 20596 29696 20602
rect 29644 20538 29696 20544
rect 29656 20466 29684 20538
rect 29644 20460 29696 20466
rect 29644 20402 29696 20408
rect 29644 20256 29696 20262
rect 29644 20198 29696 20204
rect 29472 19774 29592 19802
rect 29368 17740 29420 17746
rect 29368 17682 29420 17688
rect 29472 17678 29500 19774
rect 29552 19712 29604 19718
rect 29552 19654 29604 19660
rect 29564 19378 29592 19654
rect 29552 19372 29604 19378
rect 29552 19314 29604 19320
rect 29460 17672 29512 17678
rect 29460 17614 29512 17620
rect 29472 16658 29500 17614
rect 29552 16788 29604 16794
rect 29552 16730 29604 16736
rect 29460 16652 29512 16658
rect 29460 16594 29512 16600
rect 29368 15564 29420 15570
rect 29368 15506 29420 15512
rect 29184 15428 29236 15434
rect 29184 15370 29236 15376
rect 29276 15428 29328 15434
rect 29276 15370 29328 15376
rect 29012 14878 29132 14906
rect 29196 14890 29224 15370
rect 29184 14884 29236 14890
rect 28908 14544 28960 14550
rect 28908 14486 28960 14492
rect 28908 13728 28960 13734
rect 28908 13670 28960 13676
rect 28920 13190 28948 13670
rect 29012 13258 29040 14878
rect 29184 14826 29236 14832
rect 29276 14476 29328 14482
rect 29276 14418 29328 14424
rect 29092 14408 29144 14414
rect 29092 14350 29144 14356
rect 29104 13938 29132 14350
rect 29184 14340 29236 14346
rect 29184 14282 29236 14288
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 29104 13530 29132 13874
rect 29092 13524 29144 13530
rect 29092 13466 29144 13472
rect 29000 13252 29052 13258
rect 29000 13194 29052 13200
rect 28816 13184 28868 13190
rect 28816 13126 28868 13132
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 28828 12850 28856 13126
rect 28816 12844 28868 12850
rect 28816 12786 28868 12792
rect 28736 12702 28856 12730
rect 28632 11144 28684 11150
rect 28632 11086 28684 11092
rect 28724 11076 28776 11082
rect 28724 11018 28776 11024
rect 28356 10260 28408 10266
rect 28356 10202 28408 10208
rect 28264 10056 28316 10062
rect 28264 9998 28316 10004
rect 28356 9648 28408 9654
rect 28356 9590 28408 9596
rect 28446 9616 28502 9625
rect 28368 9178 28396 9590
rect 28446 9551 28502 9560
rect 28460 9518 28488 9551
rect 28448 9512 28500 9518
rect 28448 9454 28500 9460
rect 28736 9382 28764 11018
rect 28724 9376 28776 9382
rect 28724 9318 28776 9324
rect 28172 9172 28224 9178
rect 28172 9114 28224 9120
rect 28356 9172 28408 9178
rect 28356 9114 28408 9120
rect 28540 9172 28592 9178
rect 28540 9114 28592 9120
rect 28448 9036 28500 9042
rect 28448 8978 28500 8984
rect 28460 8634 28488 8978
rect 28448 8628 28500 8634
rect 28448 8570 28500 8576
rect 28356 7744 28408 7750
rect 28356 7686 28408 7692
rect 28368 7410 28396 7686
rect 28552 7410 28580 9114
rect 28736 8838 28764 9318
rect 28632 8832 28684 8838
rect 28630 8800 28632 8809
rect 28724 8832 28776 8838
rect 28684 8800 28686 8809
rect 28724 8774 28776 8780
rect 28630 8735 28686 8744
rect 28644 8378 28672 8735
rect 28644 8350 28764 8378
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 28644 7886 28672 8230
rect 28632 7880 28684 7886
rect 28632 7822 28684 7828
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 28540 7404 28592 7410
rect 28540 7346 28592 7352
rect 28644 5370 28672 7822
rect 28736 7818 28764 8350
rect 28724 7812 28776 7818
rect 28724 7754 28776 7760
rect 28736 5914 28764 7754
rect 28724 5908 28776 5914
rect 28724 5850 28776 5856
rect 28632 5364 28684 5370
rect 28632 5306 28684 5312
rect 28736 4826 28764 5850
rect 28724 4820 28776 4826
rect 28724 4762 28776 4768
rect 28630 3768 28686 3777
rect 27804 3732 27856 3738
rect 27804 3674 27856 3680
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 28080 3732 28132 3738
rect 28630 3703 28632 3712
rect 28080 3674 28132 3680
rect 28684 3703 28686 3712
rect 28632 3674 28684 3680
rect 27712 3460 27764 3466
rect 27712 3402 27764 3408
rect 27816 3058 27844 3674
rect 26792 3052 26844 3058
rect 26792 2994 26844 3000
rect 27804 3052 27856 3058
rect 27804 2994 27856 3000
rect 26700 2848 26752 2854
rect 26700 2790 26752 2796
rect 27436 2848 27488 2854
rect 27436 2790 27488 2796
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 26332 2304 26384 2310
rect 26332 2246 26384 2252
rect 26344 800 26372 2246
rect 26712 800 26740 2790
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 27080 800 27108 2246
rect 27448 800 27476 2790
rect 27908 2446 27936 3674
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 27804 2304 27856 2310
rect 27804 2246 27856 2252
rect 27816 800 27844 2246
rect 28184 800 28212 2790
rect 28644 2774 28672 3674
rect 28828 3194 28856 12702
rect 29092 12436 29144 12442
rect 29092 12378 29144 12384
rect 29000 12368 29052 12374
rect 29000 12310 29052 12316
rect 28908 12164 28960 12170
rect 28908 12106 28960 12112
rect 28920 11830 28948 12106
rect 28908 11824 28960 11830
rect 28908 11766 28960 11772
rect 29012 10062 29040 12310
rect 29104 11830 29132 12378
rect 29092 11824 29144 11830
rect 29092 11766 29144 11772
rect 29092 11688 29144 11694
rect 29090 11656 29092 11665
rect 29144 11656 29146 11665
rect 29090 11591 29146 11600
rect 29090 11384 29146 11393
rect 29090 11319 29146 11328
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 29104 9674 29132 11319
rect 29196 10810 29224 14282
rect 29288 14006 29316 14418
rect 29276 14000 29328 14006
rect 29276 13942 29328 13948
rect 29276 12164 29328 12170
rect 29276 12106 29328 12112
rect 29184 10804 29236 10810
rect 29184 10746 29236 10752
rect 29184 10600 29236 10606
rect 29184 10542 29236 10548
rect 29012 9646 29132 9674
rect 28908 9580 28960 9586
rect 28908 9522 28960 9528
rect 28920 9353 28948 9522
rect 28906 9344 28962 9353
rect 28906 9279 28962 9288
rect 29012 7970 29040 9646
rect 29092 9036 29144 9042
rect 29092 8978 29144 8984
rect 28920 7942 29040 7970
rect 29104 7954 29132 8978
rect 29196 7954 29224 10542
rect 29288 10266 29316 12106
rect 29276 10260 29328 10266
rect 29276 10202 29328 10208
rect 29380 8401 29408 15506
rect 29472 15502 29500 16594
rect 29460 15496 29512 15502
rect 29460 15438 29512 15444
rect 29564 15094 29592 16730
rect 29656 16590 29684 20198
rect 29748 19990 29776 20742
rect 29840 20641 29868 21626
rect 29826 20632 29882 20641
rect 29826 20567 29882 20576
rect 29828 20528 29880 20534
rect 29828 20470 29880 20476
rect 29736 19984 29788 19990
rect 29736 19926 29788 19932
rect 29840 19854 29868 20470
rect 29828 19848 29880 19854
rect 29828 19790 29880 19796
rect 29932 19530 29960 22066
rect 30300 21554 30328 22102
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 30288 21548 30340 21554
rect 30288 21490 30340 21496
rect 30484 21457 30512 21830
rect 30470 21448 30526 21457
rect 30470 21383 30526 21392
rect 30104 21344 30156 21350
rect 30104 21286 30156 21292
rect 30012 20936 30064 20942
rect 30012 20878 30064 20884
rect 30024 20466 30052 20878
rect 30116 20534 30144 21286
rect 30288 20936 30340 20942
rect 30288 20878 30340 20884
rect 30196 20800 30248 20806
rect 30196 20742 30248 20748
rect 30104 20528 30156 20534
rect 30104 20470 30156 20476
rect 30012 20460 30064 20466
rect 30012 20402 30064 20408
rect 30012 20324 30064 20330
rect 30012 20266 30064 20272
rect 30024 20058 30052 20266
rect 30012 20052 30064 20058
rect 30012 19994 30064 20000
rect 29748 19502 29960 19530
rect 29644 16584 29696 16590
rect 29644 16526 29696 16532
rect 29552 15088 29604 15094
rect 29552 15030 29604 15036
rect 29550 13560 29606 13569
rect 29550 13495 29606 13504
rect 29564 13326 29592 13495
rect 29552 13320 29604 13326
rect 29552 13262 29604 13268
rect 29460 11620 29512 11626
rect 29460 11562 29512 11568
rect 29472 11393 29500 11562
rect 29458 11384 29514 11393
rect 29458 11319 29514 11328
rect 29460 11280 29512 11286
rect 29460 11222 29512 11228
rect 29472 9654 29500 11222
rect 29460 9648 29512 9654
rect 29460 9590 29512 9596
rect 29472 9518 29500 9590
rect 29460 9512 29512 9518
rect 29460 9454 29512 9460
rect 29472 9042 29500 9454
rect 29460 9036 29512 9042
rect 29460 8978 29512 8984
rect 29460 8492 29512 8498
rect 29460 8434 29512 8440
rect 29366 8392 29422 8401
rect 29366 8327 29422 8336
rect 29092 7948 29144 7954
rect 28920 7426 28948 7942
rect 29092 7890 29144 7896
rect 29184 7948 29236 7954
rect 29184 7890 29236 7896
rect 29000 7880 29052 7886
rect 29000 7822 29052 7828
rect 29012 7546 29040 7822
rect 29000 7540 29052 7546
rect 29000 7482 29052 7488
rect 28920 7398 29040 7426
rect 29012 6662 29040 7398
rect 29104 7342 29132 7890
rect 29196 7410 29224 7890
rect 29184 7404 29236 7410
rect 29184 7346 29236 7352
rect 29368 7404 29420 7410
rect 29368 7346 29420 7352
rect 29092 7336 29144 7342
rect 29092 7278 29144 7284
rect 29000 6656 29052 6662
rect 29000 6598 29052 6604
rect 29012 5710 29040 6598
rect 29196 6458 29224 7346
rect 29380 6934 29408 7346
rect 29472 7274 29500 8434
rect 29460 7268 29512 7274
rect 29460 7210 29512 7216
rect 29368 6928 29420 6934
rect 29368 6870 29420 6876
rect 29380 6730 29408 6870
rect 29564 6866 29592 13262
rect 29748 12986 29776 19502
rect 29920 19440 29972 19446
rect 29920 19382 29972 19388
rect 29828 17536 29880 17542
rect 29828 17478 29880 17484
rect 29840 17134 29868 17478
rect 29828 17128 29880 17134
rect 29828 17070 29880 17076
rect 29932 16454 29960 19382
rect 30208 19242 30236 20742
rect 30300 20602 30328 20878
rect 30288 20596 30340 20602
rect 30288 20538 30340 20544
rect 30472 20324 30524 20330
rect 30472 20266 30524 20272
rect 30288 19916 30340 19922
rect 30288 19858 30340 19864
rect 30300 19825 30328 19858
rect 30286 19816 30342 19825
rect 30286 19751 30342 19760
rect 30288 19712 30340 19718
rect 30286 19680 30288 19689
rect 30340 19680 30342 19689
rect 30286 19615 30342 19624
rect 30484 19514 30512 20266
rect 30472 19508 30524 19514
rect 30472 19450 30524 19456
rect 30196 19236 30248 19242
rect 30196 19178 30248 19184
rect 30104 18760 30156 18766
rect 30104 18702 30156 18708
rect 30288 18760 30340 18766
rect 30288 18702 30340 18708
rect 30116 18358 30144 18702
rect 30104 18352 30156 18358
rect 30010 18320 30066 18329
rect 30104 18294 30156 18300
rect 30010 18255 30066 18264
rect 30024 16454 30052 18255
rect 30300 18086 30328 18702
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 30300 17746 30328 18022
rect 30104 17740 30156 17746
rect 30104 17682 30156 17688
rect 30288 17740 30340 17746
rect 30288 17682 30340 17688
rect 30380 17740 30432 17746
rect 30380 17682 30432 17688
rect 30116 17626 30144 17682
rect 30392 17626 30420 17682
rect 30116 17598 30420 17626
rect 30380 17536 30432 17542
rect 30380 17478 30432 17484
rect 30392 16794 30420 17478
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 29920 16448 29972 16454
rect 29920 16390 29972 16396
rect 30012 16448 30064 16454
rect 30012 16390 30064 16396
rect 30024 16114 30052 16390
rect 30300 16250 30328 16594
rect 30288 16244 30340 16250
rect 30288 16186 30340 16192
rect 30012 16108 30064 16114
rect 30012 16050 30064 16056
rect 29920 15496 29972 15502
rect 29920 15438 29972 15444
rect 29826 14512 29882 14521
rect 29826 14447 29828 14456
rect 29880 14447 29882 14456
rect 29828 14418 29880 14424
rect 29932 14414 29960 15438
rect 30380 15360 30432 15366
rect 30380 15302 30432 15308
rect 30470 15328 30526 15337
rect 30104 14816 30156 14822
rect 30104 14758 30156 14764
rect 29920 14408 29972 14414
rect 29920 14350 29972 14356
rect 30012 13932 30064 13938
rect 30012 13874 30064 13880
rect 30024 13841 30052 13874
rect 30010 13832 30066 13841
rect 30010 13767 30066 13776
rect 29920 13728 29972 13734
rect 29920 13670 29972 13676
rect 29932 13258 29960 13670
rect 29920 13252 29972 13258
rect 29840 13212 29920 13240
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 29840 12918 29868 13212
rect 29920 13194 29972 13200
rect 29828 12912 29880 12918
rect 29828 12854 29880 12860
rect 29736 12844 29788 12850
rect 29736 12786 29788 12792
rect 30012 12844 30064 12850
rect 30012 12786 30064 12792
rect 29748 12442 29776 12786
rect 30024 12442 30052 12786
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 30012 12436 30064 12442
rect 30012 12378 30064 12384
rect 29644 12232 29696 12238
rect 29644 12174 29696 12180
rect 29828 12232 29880 12238
rect 29828 12174 29880 12180
rect 29656 11898 29684 12174
rect 29644 11892 29696 11898
rect 29644 11834 29696 11840
rect 29840 11665 29868 12174
rect 30024 11898 30052 12378
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 29920 11824 29972 11830
rect 29918 11792 29920 11801
rect 29972 11792 29974 11801
rect 29918 11727 29974 11736
rect 29826 11656 29882 11665
rect 29826 11591 29882 11600
rect 29644 11552 29696 11558
rect 29932 11540 29960 11727
rect 29932 11512 30052 11540
rect 29644 11494 29696 11500
rect 29656 11082 29684 11494
rect 29644 11076 29696 11082
rect 29644 11018 29696 11024
rect 29918 10840 29974 10849
rect 29918 10775 29974 10784
rect 29932 10742 29960 10775
rect 29644 10736 29696 10742
rect 29644 10678 29696 10684
rect 29920 10736 29972 10742
rect 29920 10678 29972 10684
rect 29656 7834 29684 10678
rect 29828 10668 29880 10674
rect 29828 10610 29880 10616
rect 29736 10600 29788 10606
rect 29736 10542 29788 10548
rect 29748 10266 29776 10542
rect 29736 10260 29788 10266
rect 29736 10202 29788 10208
rect 29840 10198 29868 10610
rect 29920 10600 29972 10606
rect 29920 10542 29972 10548
rect 29828 10192 29880 10198
rect 29828 10134 29880 10140
rect 29932 9994 29960 10542
rect 29920 9988 29972 9994
rect 29920 9930 29972 9936
rect 29918 9752 29974 9761
rect 29918 9687 29974 9696
rect 29736 9580 29788 9586
rect 29736 9522 29788 9528
rect 29748 9489 29776 9522
rect 29734 9480 29790 9489
rect 29734 9415 29790 9424
rect 29828 9376 29880 9382
rect 29828 9318 29880 9324
rect 29840 8974 29868 9318
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 29748 8566 29776 8910
rect 29736 8560 29788 8566
rect 29736 8502 29788 8508
rect 29748 7954 29776 8502
rect 29736 7948 29788 7954
rect 29736 7890 29788 7896
rect 29656 7806 29776 7834
rect 29642 7032 29698 7041
rect 29642 6967 29698 6976
rect 29552 6860 29604 6866
rect 29552 6802 29604 6808
rect 29368 6724 29420 6730
rect 29368 6666 29420 6672
rect 29184 6452 29236 6458
rect 29184 6394 29236 6400
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 29012 3466 29040 5646
rect 29196 5234 29224 6394
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 29000 3460 29052 3466
rect 29000 3402 29052 3408
rect 29656 3194 29684 6967
rect 29748 6322 29776 7806
rect 29736 6316 29788 6322
rect 29736 6258 29788 6264
rect 29932 3194 29960 9687
rect 30024 6730 30052 11512
rect 30116 10810 30144 14758
rect 30194 13832 30250 13841
rect 30194 13767 30250 13776
rect 30208 11082 30236 13767
rect 30392 13326 30420 15302
rect 30470 15263 30526 15272
rect 30484 14958 30512 15263
rect 30576 15201 30604 33798
rect 30656 33380 30708 33386
rect 30656 33322 30708 33328
rect 30668 15552 30696 33322
rect 30760 30938 30788 39238
rect 30932 38412 30984 38418
rect 30932 38354 30984 38360
rect 30840 37936 30892 37942
rect 30838 37904 30840 37913
rect 30892 37904 30894 37913
rect 30944 37874 30972 38354
rect 31220 38350 31248 39238
rect 31496 38418 31524 39986
rect 31588 38418 31616 42094
rect 31864 41138 31892 45222
rect 31944 43648 31996 43654
rect 31944 43590 31996 43596
rect 31956 42362 31984 43590
rect 32036 43308 32088 43314
rect 32036 43250 32088 43256
rect 31944 42356 31996 42362
rect 31944 42298 31996 42304
rect 31944 42016 31996 42022
rect 31944 41958 31996 41964
rect 31852 41132 31904 41138
rect 31852 41074 31904 41080
rect 31956 41018 31984 41958
rect 32048 41818 32076 43250
rect 32036 41812 32088 41818
rect 32036 41754 32088 41760
rect 31772 40990 31984 41018
rect 31772 40934 31800 40990
rect 31760 40928 31812 40934
rect 31760 40870 31812 40876
rect 31944 40928 31996 40934
rect 31944 40870 31996 40876
rect 31668 39840 31720 39846
rect 31668 39782 31720 39788
rect 31680 39030 31708 39782
rect 31668 39024 31720 39030
rect 31668 38966 31720 38972
rect 31484 38412 31536 38418
rect 31484 38354 31536 38360
rect 31576 38412 31628 38418
rect 31576 38354 31628 38360
rect 31208 38344 31260 38350
rect 31208 38286 31260 38292
rect 31482 38312 31538 38321
rect 31482 38247 31484 38256
rect 31536 38247 31538 38256
rect 31484 38218 31536 38224
rect 31668 38208 31720 38214
rect 31668 38150 31720 38156
rect 31022 38040 31078 38049
rect 31022 37975 31078 37984
rect 31206 38040 31262 38049
rect 31206 37975 31262 37984
rect 31036 37942 31064 37975
rect 31024 37936 31076 37942
rect 31024 37878 31076 37884
rect 31220 37874 31248 37975
rect 30838 37839 30894 37848
rect 30932 37868 30984 37874
rect 30932 37810 30984 37816
rect 31208 37868 31260 37874
rect 31208 37810 31260 37816
rect 30840 37188 30892 37194
rect 30840 37130 30892 37136
rect 30852 36854 30880 37130
rect 31220 37097 31248 37810
rect 31576 37324 31628 37330
rect 31576 37266 31628 37272
rect 31206 37088 31262 37097
rect 31206 37023 31262 37032
rect 30840 36848 30892 36854
rect 30840 36790 30892 36796
rect 31208 36644 31260 36650
rect 31208 36586 31260 36592
rect 31220 36417 31248 36586
rect 31206 36408 31262 36417
rect 31206 36343 31262 36352
rect 31208 36032 31260 36038
rect 31208 35974 31260 35980
rect 30840 35488 30892 35494
rect 30840 35430 30892 35436
rect 31024 35488 31076 35494
rect 31024 35430 31076 35436
rect 30852 34950 30880 35430
rect 31036 35290 31064 35430
rect 31024 35284 31076 35290
rect 31024 35226 31076 35232
rect 30932 35080 30984 35086
rect 30932 35022 30984 35028
rect 31116 35080 31168 35086
rect 31116 35022 31168 35028
rect 30840 34944 30892 34950
rect 30840 34886 30892 34892
rect 30852 34524 30880 34886
rect 30944 34785 30972 35022
rect 30930 34776 30986 34785
rect 30930 34711 30986 34720
rect 30932 34536 30984 34542
rect 30852 34496 30932 34524
rect 31128 34513 31156 35022
rect 30932 34478 30984 34484
rect 31114 34504 31170 34513
rect 31114 34439 31116 34448
rect 31168 34439 31170 34448
rect 31116 34410 31168 34416
rect 30932 34400 30984 34406
rect 31128 34379 31156 34410
rect 30932 34342 30984 34348
rect 30748 30932 30800 30938
rect 30748 30874 30800 30880
rect 30944 27713 30972 34342
rect 31220 34202 31248 35974
rect 31392 35624 31444 35630
rect 31392 35566 31444 35572
rect 31298 34640 31354 34649
rect 31298 34575 31354 34584
rect 31312 34202 31340 34575
rect 31208 34196 31260 34202
rect 31208 34138 31260 34144
rect 31300 34196 31352 34202
rect 31300 34138 31352 34144
rect 31220 33998 31248 34138
rect 31208 33992 31260 33998
rect 31208 33934 31260 33940
rect 31312 31754 31340 34138
rect 31220 31726 31340 31754
rect 31404 31754 31432 35566
rect 31484 35488 31536 35494
rect 31484 35430 31536 35436
rect 31496 35057 31524 35430
rect 31482 35048 31538 35057
rect 31482 34983 31538 34992
rect 31484 34740 31536 34746
rect 31484 34682 31536 34688
rect 31496 34542 31524 34682
rect 31484 34536 31536 34542
rect 31484 34478 31536 34484
rect 31588 31793 31616 37266
rect 31574 31784 31630 31793
rect 31404 31726 31524 31754
rect 30930 27704 30986 27713
rect 30930 27639 30986 27648
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30944 24410 30972 24754
rect 30932 24404 30984 24410
rect 30932 24346 30984 24352
rect 31220 24342 31248 31726
rect 31300 24608 31352 24614
rect 31300 24550 31352 24556
rect 31208 24336 31260 24342
rect 31208 24278 31260 24284
rect 31208 23860 31260 23866
rect 31208 23802 31260 23808
rect 31220 23730 31248 23802
rect 31208 23724 31260 23730
rect 31208 23666 31260 23672
rect 30840 23520 30892 23526
rect 30840 23462 30892 23468
rect 30852 23322 30880 23462
rect 30840 23316 30892 23322
rect 30840 23258 30892 23264
rect 30852 22098 30880 23258
rect 31312 23050 31340 24550
rect 31392 24064 31444 24070
rect 31392 24006 31444 24012
rect 31300 23044 31352 23050
rect 31300 22986 31352 22992
rect 31208 22976 31260 22982
rect 31208 22918 31260 22924
rect 30932 22704 30984 22710
rect 30932 22646 30984 22652
rect 30944 22234 30972 22646
rect 30932 22228 30984 22234
rect 30932 22170 30984 22176
rect 30840 22092 30892 22098
rect 30840 22034 30892 22040
rect 31220 22030 31248 22918
rect 31300 22432 31352 22438
rect 31300 22374 31352 22380
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31220 21554 31248 21966
rect 31208 21548 31260 21554
rect 31208 21490 31260 21496
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30840 19916 30892 19922
rect 30840 19858 30892 19864
rect 30748 19848 30800 19854
rect 30748 19790 30800 19796
rect 30760 19446 30788 19790
rect 30748 19440 30800 19446
rect 30748 19382 30800 19388
rect 30852 18834 30880 19858
rect 30840 18828 30892 18834
rect 30840 18770 30892 18776
rect 30840 18624 30892 18630
rect 30838 18592 30840 18601
rect 30892 18592 30894 18601
rect 30838 18527 30894 18536
rect 30944 18358 30972 21286
rect 31312 21128 31340 22374
rect 31404 21894 31432 24006
rect 31392 21888 31444 21894
rect 31390 21856 31392 21865
rect 31444 21856 31446 21865
rect 31390 21791 31446 21800
rect 31312 21100 31432 21128
rect 31300 21004 31352 21010
rect 31300 20946 31352 20952
rect 31116 19848 31168 19854
rect 31022 19816 31078 19825
rect 31168 19808 31248 19836
rect 31116 19790 31168 19796
rect 31022 19751 31078 19760
rect 31036 19310 31064 19751
rect 31220 19514 31248 19808
rect 31208 19508 31260 19514
rect 31208 19450 31260 19456
rect 31116 19372 31168 19378
rect 31116 19314 31168 19320
rect 31024 19304 31076 19310
rect 31024 19246 31076 19252
rect 31036 18358 31064 19246
rect 30748 18352 30800 18358
rect 30746 18320 30748 18329
rect 30932 18352 30984 18358
rect 30800 18320 30802 18329
rect 30932 18294 30984 18300
rect 31024 18352 31076 18358
rect 31024 18294 31076 18300
rect 30746 18255 30802 18264
rect 31128 17785 31156 19314
rect 31114 17776 31170 17785
rect 31114 17711 31170 17720
rect 30748 17604 30800 17610
rect 30748 17546 30800 17552
rect 30760 17270 30788 17546
rect 30748 17264 30800 17270
rect 30748 17206 30800 17212
rect 31024 17196 31076 17202
rect 31024 17138 31076 17144
rect 31036 16794 31064 17138
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 31128 16114 31156 17711
rect 31312 16153 31340 20946
rect 31404 19378 31432 21100
rect 31392 19372 31444 19378
rect 31392 19314 31444 19320
rect 31390 18456 31446 18465
rect 31390 18391 31392 18400
rect 31444 18391 31446 18400
rect 31392 18362 31444 18368
rect 31390 17776 31446 17785
rect 31390 17711 31446 17720
rect 31404 17678 31432 17711
rect 31392 17672 31444 17678
rect 31392 17614 31444 17620
rect 31298 16144 31354 16153
rect 31116 16108 31168 16114
rect 31298 16079 31354 16088
rect 31116 16050 31168 16056
rect 30668 15524 31064 15552
rect 30932 15428 30984 15434
rect 30932 15370 30984 15376
rect 30840 15360 30892 15366
rect 30840 15302 30892 15308
rect 30562 15192 30618 15201
rect 30562 15127 30618 15136
rect 30472 14952 30524 14958
rect 30472 14894 30524 14900
rect 30748 14272 30800 14278
rect 30748 14214 30800 14220
rect 30472 14000 30524 14006
rect 30472 13942 30524 13948
rect 30484 13394 30512 13942
rect 30472 13388 30524 13394
rect 30472 13330 30524 13336
rect 30760 13326 30788 14214
rect 30852 13326 30880 15302
rect 30944 14414 30972 15370
rect 30932 14408 30984 14414
rect 30932 14350 30984 14356
rect 30944 13938 30972 14350
rect 30932 13932 30984 13938
rect 30932 13874 30984 13880
rect 30932 13796 30984 13802
rect 30932 13738 30984 13744
rect 30380 13320 30432 13326
rect 30380 13262 30432 13268
rect 30748 13320 30800 13326
rect 30748 13262 30800 13268
rect 30840 13320 30892 13326
rect 30840 13262 30892 13268
rect 30380 13184 30432 13190
rect 30380 13126 30432 13132
rect 30656 13184 30708 13190
rect 30656 13126 30708 13132
rect 30288 12640 30340 12646
rect 30288 12582 30340 12588
rect 30300 11762 30328 12582
rect 30288 11756 30340 11762
rect 30288 11698 30340 11704
rect 30286 11384 30342 11393
rect 30286 11319 30342 11328
rect 30196 11076 30248 11082
rect 30196 11018 30248 11024
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 30104 9376 30156 9382
rect 30104 9318 30156 9324
rect 30116 8498 30144 9318
rect 30104 8492 30156 8498
rect 30104 8434 30156 8440
rect 30208 7750 30236 11018
rect 30300 9994 30328 11319
rect 30392 10198 30420 13126
rect 30564 12980 30616 12986
rect 30564 12922 30616 12928
rect 30576 11150 30604 12922
rect 30668 12918 30696 13126
rect 30656 12912 30708 12918
rect 30656 12854 30708 12860
rect 30760 12850 30788 13262
rect 30748 12844 30800 12850
rect 30748 12786 30800 12792
rect 30654 12472 30710 12481
rect 30654 12407 30710 12416
rect 30668 12170 30696 12407
rect 30760 12238 30788 12786
rect 30852 12306 30880 13262
rect 30840 12300 30892 12306
rect 30840 12242 30892 12248
rect 30748 12232 30800 12238
rect 30748 12174 30800 12180
rect 30656 12164 30708 12170
rect 30656 12106 30708 12112
rect 30748 11824 30800 11830
rect 30800 11784 30880 11812
rect 30748 11766 30800 11772
rect 30656 11620 30708 11626
rect 30656 11562 30708 11568
rect 30564 11144 30616 11150
rect 30564 11086 30616 11092
rect 30668 10198 30696 11562
rect 30852 11150 30880 11784
rect 30944 11234 30972 13738
rect 31036 12889 31064 15524
rect 31300 15496 31352 15502
rect 31300 15438 31352 15444
rect 31116 15428 31168 15434
rect 31116 15370 31168 15376
rect 31128 13530 31156 15370
rect 31312 14482 31340 15438
rect 31300 14476 31352 14482
rect 31300 14418 31352 14424
rect 31208 14272 31260 14278
rect 31208 14214 31260 14220
rect 31116 13524 31168 13530
rect 31116 13466 31168 13472
rect 31220 13394 31248 14214
rect 31312 14074 31340 14418
rect 31300 14068 31352 14074
rect 31300 14010 31352 14016
rect 31496 13954 31524 31726
rect 31574 31719 31630 31728
rect 31576 24200 31628 24206
rect 31576 24142 31628 24148
rect 31588 21894 31616 24142
rect 31576 21888 31628 21894
rect 31576 21830 31628 21836
rect 31680 21690 31708 38150
rect 31772 37913 31800 40870
rect 31852 39976 31904 39982
rect 31852 39918 31904 39924
rect 31864 38554 31892 39918
rect 31852 38548 31904 38554
rect 31852 38490 31904 38496
rect 31758 37904 31814 37913
rect 31758 37839 31814 37848
rect 31864 36922 31892 38490
rect 31852 36916 31904 36922
rect 31852 36858 31904 36864
rect 31956 36786 31984 40870
rect 32140 40458 32168 52906
rect 32232 41274 32260 53110
rect 32784 53106 32812 55200
rect 34256 53106 34284 55270
rect 35162 55270 35480 55298
rect 35162 55200 35218 55270
rect 35452 53106 35480 55270
rect 36358 55270 36676 55298
rect 36358 55200 36414 55270
rect 36648 53106 36676 55270
rect 37554 55270 37872 55298
rect 37554 55200 37610 55270
rect 37844 53106 37872 55270
rect 38750 55270 39068 55298
rect 38750 55200 38806 55270
rect 39040 53106 39068 55270
rect 39946 55200 40002 56000
rect 41142 55298 41198 56000
rect 41142 55270 41368 55298
rect 41142 55200 41198 55270
rect 32772 53100 32824 53106
rect 32772 53042 32824 53048
rect 34244 53100 34296 53106
rect 34244 53042 34296 53048
rect 35440 53100 35492 53106
rect 35440 53042 35492 53048
rect 36636 53100 36688 53106
rect 36636 53042 36688 53048
rect 37832 53100 37884 53106
rect 37832 53042 37884 53048
rect 39028 53100 39080 53106
rect 39960 53088 39988 55200
rect 40040 53100 40092 53106
rect 39960 53060 40040 53088
rect 39028 53042 39080 53048
rect 41340 53088 41368 55270
rect 42338 55200 42394 56000
rect 43534 55298 43590 56000
rect 43534 55270 43668 55298
rect 43534 55200 43590 55270
rect 42352 53106 42380 55200
rect 43640 53106 43668 55270
rect 44730 55200 44786 56000
rect 45926 55298 45982 56000
rect 45926 55270 46060 55298
rect 45926 55200 45982 55270
rect 44744 53106 44772 55200
rect 41420 53100 41472 53106
rect 41340 53060 41420 53088
rect 40040 53042 40092 53048
rect 41420 53042 41472 53048
rect 42340 53100 42392 53106
rect 42340 53042 42392 53048
rect 43628 53100 43680 53106
rect 43628 53042 43680 53048
rect 44732 53100 44784 53106
rect 44732 53042 44784 53048
rect 45192 53100 45244 53106
rect 45192 53042 45244 53048
rect 32588 52896 32640 52902
rect 32588 52838 32640 52844
rect 32404 47456 32456 47462
rect 32404 47398 32456 47404
rect 32416 47054 32444 47398
rect 32600 47122 32628 52838
rect 32784 52698 32812 53042
rect 34256 52698 34284 53042
rect 34796 53032 34848 53038
rect 34796 52974 34848 52980
rect 34704 52964 34756 52970
rect 34704 52906 34756 52912
rect 34336 52896 34388 52902
rect 34336 52838 34388 52844
rect 32772 52692 32824 52698
rect 32772 52634 32824 52640
rect 34244 52692 34296 52698
rect 34244 52634 34296 52640
rect 33048 52556 33100 52562
rect 33048 52498 33100 52504
rect 32680 51876 32732 51882
rect 32680 51818 32732 51824
rect 32588 47116 32640 47122
rect 32588 47058 32640 47064
rect 32404 47048 32456 47054
rect 32404 46990 32456 46996
rect 32404 45960 32456 45966
rect 32404 45902 32456 45908
rect 32416 45830 32444 45902
rect 32404 45824 32456 45830
rect 32404 45766 32456 45772
rect 32310 44296 32366 44305
rect 32310 44231 32312 44240
rect 32364 44231 32366 44240
rect 32312 44202 32364 44208
rect 32324 42770 32352 44202
rect 32692 43738 32720 51818
rect 33060 51074 33088 52498
rect 32968 51046 33088 51074
rect 32864 49088 32916 49094
rect 32864 49030 32916 49036
rect 32876 48618 32904 49030
rect 32864 48612 32916 48618
rect 32864 48554 32916 48560
rect 32772 47728 32824 47734
rect 32772 47670 32824 47676
rect 32784 46646 32812 47670
rect 32772 46640 32824 46646
rect 32772 46582 32824 46588
rect 32784 45966 32812 46582
rect 32772 45960 32824 45966
rect 32772 45902 32824 45908
rect 32784 45286 32812 45902
rect 32772 45280 32824 45286
rect 32772 45222 32824 45228
rect 32772 44192 32824 44198
rect 32772 44134 32824 44140
rect 32600 43710 32720 43738
rect 32600 43314 32628 43710
rect 32784 43654 32812 44134
rect 32968 43994 32996 51046
rect 33508 49088 33560 49094
rect 33508 49030 33560 49036
rect 33140 48544 33192 48550
rect 33140 48486 33192 48492
rect 33232 48544 33284 48550
rect 33232 48486 33284 48492
rect 33152 47666 33180 48486
rect 33244 48074 33272 48486
rect 33416 48272 33468 48278
rect 33416 48214 33468 48220
rect 33428 48142 33456 48214
rect 33520 48142 33548 49030
rect 34060 48544 34112 48550
rect 34060 48486 34112 48492
rect 33416 48136 33468 48142
rect 33416 48078 33468 48084
rect 33508 48136 33560 48142
rect 33508 48078 33560 48084
rect 33968 48136 34020 48142
rect 33968 48078 34020 48084
rect 33232 48068 33284 48074
rect 33232 48010 33284 48016
rect 33244 47734 33272 48010
rect 33520 47818 33548 48078
rect 33336 47802 33548 47818
rect 33324 47796 33548 47802
rect 33376 47790 33548 47796
rect 33324 47738 33376 47744
rect 33232 47728 33284 47734
rect 33232 47670 33284 47676
rect 33140 47660 33192 47666
rect 33140 47602 33192 47608
rect 33508 47660 33560 47666
rect 33508 47602 33560 47608
rect 33520 47122 33548 47602
rect 33876 47524 33928 47530
rect 33876 47466 33928 47472
rect 33692 47456 33744 47462
rect 33692 47398 33744 47404
rect 33508 47116 33560 47122
rect 33508 47058 33560 47064
rect 33140 47048 33192 47054
rect 33324 47048 33376 47054
rect 33140 46990 33192 46996
rect 33322 47016 33324 47025
rect 33376 47016 33378 47025
rect 33048 46368 33100 46374
rect 33048 46310 33100 46316
rect 32956 43988 33008 43994
rect 32956 43930 33008 43936
rect 32968 43874 32996 43930
rect 32876 43846 32996 43874
rect 32680 43648 32732 43654
rect 32680 43590 32732 43596
rect 32772 43648 32824 43654
rect 32772 43590 32824 43596
rect 32692 43450 32720 43590
rect 32680 43444 32732 43450
rect 32680 43386 32732 43392
rect 32588 43308 32640 43314
rect 32588 43250 32640 43256
rect 32404 43240 32456 43246
rect 32404 43182 32456 43188
rect 32312 42764 32364 42770
rect 32312 42706 32364 42712
rect 32416 42294 32444 43182
rect 32588 43172 32640 43178
rect 32588 43114 32640 43120
rect 32496 42696 32548 42702
rect 32496 42638 32548 42644
rect 32404 42288 32456 42294
rect 32404 42230 32456 42236
rect 32508 41818 32536 42638
rect 32600 42226 32628 43114
rect 32588 42220 32640 42226
rect 32588 42162 32640 42168
rect 32588 42016 32640 42022
rect 32588 41958 32640 41964
rect 32496 41812 32548 41818
rect 32496 41754 32548 41760
rect 32600 41614 32628 41958
rect 32692 41614 32720 43386
rect 32784 42634 32812 43590
rect 32876 42702 32904 43846
rect 32864 42696 32916 42702
rect 32864 42638 32916 42644
rect 32772 42628 32824 42634
rect 32772 42570 32824 42576
rect 32784 42226 32812 42570
rect 32864 42288 32916 42294
rect 32864 42230 32916 42236
rect 32772 42220 32824 42226
rect 32772 42162 32824 42168
rect 32784 42022 32812 42162
rect 32876 42022 32904 42230
rect 32772 42016 32824 42022
rect 32772 41958 32824 41964
rect 32864 42016 32916 42022
rect 32864 41958 32916 41964
rect 32588 41608 32640 41614
rect 32586 41576 32588 41585
rect 32680 41608 32732 41614
rect 32640 41576 32642 41585
rect 32680 41550 32732 41556
rect 32586 41511 32642 41520
rect 32220 41268 32272 41274
rect 32220 41210 32272 41216
rect 32680 41268 32732 41274
rect 32680 41210 32732 41216
rect 32232 40526 32260 41210
rect 32692 40905 32720 41210
rect 32772 41200 32824 41206
rect 32770 41168 32772 41177
rect 32824 41168 32826 41177
rect 32770 41103 32826 41112
rect 32772 40928 32824 40934
rect 32678 40896 32734 40905
rect 32772 40870 32824 40876
rect 32678 40831 32734 40840
rect 32692 40594 32720 40831
rect 32680 40588 32732 40594
rect 32680 40530 32732 40536
rect 32220 40520 32272 40526
rect 32588 40520 32640 40526
rect 32220 40462 32272 40468
rect 32586 40488 32588 40497
rect 32640 40488 32642 40497
rect 32128 40452 32180 40458
rect 32586 40423 32642 40432
rect 32128 40394 32180 40400
rect 32220 40384 32272 40390
rect 32220 40326 32272 40332
rect 32404 40384 32456 40390
rect 32404 40326 32456 40332
rect 32496 40384 32548 40390
rect 32496 40326 32548 40332
rect 32036 38752 32088 38758
rect 32036 38694 32088 38700
rect 32128 38752 32180 38758
rect 32128 38694 32180 38700
rect 31944 36780 31996 36786
rect 31944 36722 31996 36728
rect 31944 36372 31996 36378
rect 31944 36314 31996 36320
rect 31760 36304 31812 36310
rect 31956 36281 31984 36314
rect 31760 36246 31812 36252
rect 31942 36272 31998 36281
rect 31772 34134 31800 36246
rect 31942 36207 31998 36216
rect 31760 34128 31812 34134
rect 31760 34070 31812 34076
rect 31760 33924 31812 33930
rect 31760 33866 31812 33872
rect 31772 33318 31800 33866
rect 31760 33312 31812 33318
rect 31760 33254 31812 33260
rect 31772 26926 31800 33254
rect 31760 26920 31812 26926
rect 31760 26862 31812 26868
rect 31944 26240 31996 26246
rect 31944 26182 31996 26188
rect 31956 25498 31984 26182
rect 31944 25492 31996 25498
rect 31944 25434 31996 25440
rect 31956 24954 31984 25434
rect 31944 24948 31996 24954
rect 31944 24890 31996 24896
rect 31956 24274 31984 24890
rect 31944 24268 31996 24274
rect 31944 24210 31996 24216
rect 31758 23896 31814 23905
rect 31758 23831 31760 23840
rect 31812 23831 31814 23840
rect 31944 23860 31996 23866
rect 31760 23802 31812 23808
rect 31944 23802 31996 23808
rect 31760 23724 31812 23730
rect 31760 23666 31812 23672
rect 31772 22778 31800 23666
rect 31760 22772 31812 22778
rect 31760 22714 31812 22720
rect 31772 22030 31800 22714
rect 31760 22024 31812 22030
rect 31760 21966 31812 21972
rect 31668 21684 31720 21690
rect 31668 21626 31720 21632
rect 31852 21412 31904 21418
rect 31852 21354 31904 21360
rect 31668 19372 31720 19378
rect 31668 19314 31720 19320
rect 31680 18766 31708 19314
rect 31668 18760 31720 18766
rect 31668 18702 31720 18708
rect 31864 18630 31892 21354
rect 31852 18624 31904 18630
rect 31852 18566 31904 18572
rect 31758 18320 31814 18329
rect 31758 18255 31760 18264
rect 31812 18255 31814 18264
rect 31760 18226 31812 18232
rect 31852 17536 31904 17542
rect 31852 17478 31904 17484
rect 31576 16720 31628 16726
rect 31576 16662 31628 16668
rect 31404 13926 31524 13954
rect 31208 13388 31260 13394
rect 31128 13348 31208 13376
rect 31022 12880 31078 12889
rect 31022 12815 31024 12824
rect 31076 12815 31078 12824
rect 31024 12786 31076 12792
rect 31036 11393 31064 12786
rect 31128 12442 31156 13348
rect 31208 13330 31260 13336
rect 31208 13184 31260 13190
rect 31208 13126 31260 13132
rect 31220 12850 31248 13126
rect 31404 12918 31432 13926
rect 31484 13796 31536 13802
rect 31484 13738 31536 13744
rect 31496 13326 31524 13738
rect 31484 13320 31536 13326
rect 31484 13262 31536 13268
rect 31392 12912 31444 12918
rect 31392 12854 31444 12860
rect 31208 12844 31260 12850
rect 31208 12786 31260 12792
rect 31404 12714 31432 12854
rect 31208 12708 31260 12714
rect 31208 12650 31260 12656
rect 31392 12708 31444 12714
rect 31392 12650 31444 12656
rect 31116 12436 31168 12442
rect 31116 12378 31168 12384
rect 31220 12220 31248 12650
rect 31484 12436 31536 12442
rect 31484 12378 31536 12384
rect 31220 12192 31340 12220
rect 31208 11756 31260 11762
rect 31208 11698 31260 11704
rect 31022 11384 31078 11393
rect 31022 11319 31078 11328
rect 30944 11206 31156 11234
rect 30748 11144 30800 11150
rect 30748 11086 30800 11092
rect 30840 11144 30892 11150
rect 30840 11086 30892 11092
rect 31024 11144 31076 11150
rect 31024 11086 31076 11092
rect 30760 10713 30788 11086
rect 30746 10704 30802 10713
rect 30746 10639 30748 10648
rect 30800 10639 30802 10648
rect 30852 10656 30880 11086
rect 30932 10668 30984 10674
rect 30748 10610 30800 10616
rect 30852 10628 30932 10656
rect 30748 10464 30800 10470
rect 30748 10406 30800 10412
rect 30380 10192 30432 10198
rect 30380 10134 30432 10140
rect 30564 10192 30616 10198
rect 30564 10134 30616 10140
rect 30656 10192 30708 10198
rect 30656 10134 30708 10140
rect 30288 9988 30340 9994
rect 30288 9930 30340 9936
rect 30472 9988 30524 9994
rect 30472 9930 30524 9936
rect 30380 9920 30432 9926
rect 30378 9888 30380 9897
rect 30432 9888 30434 9897
rect 30378 9823 30434 9832
rect 30380 9580 30432 9586
rect 30380 9522 30432 9528
rect 30392 8430 30420 9522
rect 30380 8424 30432 8430
rect 30380 8366 30432 8372
rect 30380 7812 30432 7818
rect 30380 7754 30432 7760
rect 30196 7744 30248 7750
rect 30196 7686 30248 7692
rect 30392 7546 30420 7754
rect 30380 7540 30432 7546
rect 30380 7482 30432 7488
rect 30288 7268 30340 7274
rect 30288 7210 30340 7216
rect 30012 6724 30064 6730
rect 30012 6666 30064 6672
rect 30024 5370 30052 6666
rect 30300 6322 30328 7210
rect 30484 6866 30512 9930
rect 30576 9674 30604 10134
rect 30760 9994 30788 10406
rect 30852 10062 30880 10628
rect 30932 10610 30984 10616
rect 30840 10056 30892 10062
rect 30840 9998 30892 10004
rect 30748 9988 30800 9994
rect 30748 9930 30800 9936
rect 30576 9646 30880 9674
rect 30656 9580 30708 9586
rect 30656 9522 30708 9528
rect 30564 7744 30616 7750
rect 30564 7686 30616 7692
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30380 6792 30432 6798
rect 30380 6734 30432 6740
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30012 5364 30064 5370
rect 30012 5306 30064 5312
rect 30392 4146 30420 6734
rect 30484 6458 30512 6802
rect 30472 6452 30524 6458
rect 30472 6394 30524 6400
rect 30484 5914 30512 6394
rect 30576 6322 30604 7686
rect 30668 7478 30696 9522
rect 30656 7472 30708 7478
rect 30748 7472 30800 7478
rect 30656 7414 30708 7420
rect 30746 7440 30748 7449
rect 30800 7440 30802 7449
rect 30746 7375 30802 7384
rect 30852 7206 30880 9646
rect 30932 9648 30984 9654
rect 30932 9590 30984 9596
rect 30944 8294 30972 9590
rect 31036 8906 31064 11086
rect 31128 9654 31156 11206
rect 31116 9648 31168 9654
rect 31116 9590 31168 9596
rect 31116 9512 31168 9518
rect 31116 9454 31168 9460
rect 31024 8900 31076 8906
rect 31024 8842 31076 8848
rect 31036 8362 31064 8842
rect 31024 8356 31076 8362
rect 31024 8298 31076 8304
rect 30932 8288 30984 8294
rect 30932 8230 30984 8236
rect 30944 7546 30972 8230
rect 30932 7540 30984 7546
rect 30932 7482 30984 7488
rect 31036 7342 31064 8298
rect 31128 8090 31156 9454
rect 31220 9178 31248 11698
rect 31208 9172 31260 9178
rect 31208 9114 31260 9120
rect 31208 8288 31260 8294
rect 31208 8230 31260 8236
rect 31116 8084 31168 8090
rect 31116 8026 31168 8032
rect 31220 7410 31248 8230
rect 31208 7404 31260 7410
rect 31208 7346 31260 7352
rect 31024 7336 31076 7342
rect 31024 7278 31076 7284
rect 30840 7200 30892 7206
rect 30840 7142 30892 7148
rect 31312 6798 31340 12192
rect 31496 11898 31524 12378
rect 31588 12102 31616 16662
rect 31864 16114 31892 17478
rect 31852 16108 31904 16114
rect 31852 16050 31904 16056
rect 31668 14952 31720 14958
rect 31668 14894 31720 14900
rect 31680 14618 31708 14894
rect 31668 14612 31720 14618
rect 31668 14554 31720 14560
rect 31760 14476 31812 14482
rect 31760 14418 31812 14424
rect 31668 12164 31720 12170
rect 31668 12106 31720 12112
rect 31576 12096 31628 12102
rect 31576 12038 31628 12044
rect 31680 11898 31708 12106
rect 31772 12102 31800 14418
rect 31852 13320 31904 13326
rect 31852 13262 31904 13268
rect 31760 12096 31812 12102
rect 31760 12038 31812 12044
rect 31484 11892 31536 11898
rect 31484 11834 31536 11840
rect 31668 11892 31720 11898
rect 31668 11834 31720 11840
rect 31760 11824 31812 11830
rect 31760 11766 31812 11772
rect 31772 11370 31800 11766
rect 31864 11558 31892 13262
rect 31852 11552 31904 11558
rect 31852 11494 31904 11500
rect 31772 11342 31892 11370
rect 31864 11150 31892 11342
rect 31484 11144 31536 11150
rect 31484 11086 31536 11092
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 31852 11144 31904 11150
rect 31852 11086 31904 11092
rect 31390 10840 31446 10849
rect 31390 10775 31446 10784
rect 31404 10742 31432 10775
rect 31392 10736 31444 10742
rect 31392 10678 31444 10684
rect 31496 10674 31524 11086
rect 31680 10810 31708 11086
rect 31668 10804 31720 10810
rect 31668 10746 31720 10752
rect 31864 10742 31892 11086
rect 31852 10736 31904 10742
rect 31850 10704 31852 10713
rect 31904 10704 31906 10713
rect 31484 10668 31536 10674
rect 31850 10639 31906 10648
rect 31484 10610 31536 10616
rect 31496 10282 31524 10610
rect 31404 10254 31524 10282
rect 31404 6866 31432 10254
rect 31852 10124 31904 10130
rect 31852 10066 31904 10072
rect 31588 9676 31800 9704
rect 31588 9450 31616 9676
rect 31772 9586 31800 9676
rect 31864 9654 31892 10066
rect 31852 9648 31904 9654
rect 31852 9590 31904 9596
rect 31668 9580 31720 9586
rect 31668 9522 31720 9528
rect 31760 9580 31812 9586
rect 31760 9522 31812 9528
rect 31576 9444 31628 9450
rect 31576 9386 31628 9392
rect 31680 9178 31708 9522
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 31668 9172 31720 9178
rect 31668 9114 31720 9120
rect 31772 8498 31800 9318
rect 31850 9072 31906 9081
rect 31850 9007 31852 9016
rect 31904 9007 31906 9016
rect 31852 8978 31904 8984
rect 31852 8832 31904 8838
rect 31852 8774 31904 8780
rect 31864 8673 31892 8774
rect 31850 8664 31906 8673
rect 31850 8599 31906 8608
rect 31760 8492 31812 8498
rect 31760 8434 31812 8440
rect 31576 8424 31628 8430
rect 31576 8366 31628 8372
rect 31484 8356 31536 8362
rect 31484 8298 31536 8304
rect 31392 6860 31444 6866
rect 31392 6802 31444 6808
rect 31300 6792 31352 6798
rect 31300 6734 31352 6740
rect 31496 6458 31524 8298
rect 31588 7886 31616 8366
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 31576 7200 31628 7206
rect 31576 7142 31628 7148
rect 31588 6730 31616 7142
rect 31576 6724 31628 6730
rect 31576 6666 31628 6672
rect 31484 6452 31536 6458
rect 31484 6394 31536 6400
rect 31588 6390 31616 6666
rect 31576 6384 31628 6390
rect 31576 6326 31628 6332
rect 30564 6316 30616 6322
rect 30564 6258 30616 6264
rect 30472 5908 30524 5914
rect 30472 5850 30524 5856
rect 30484 5710 30512 5850
rect 30472 5704 30524 5710
rect 30472 5646 30524 5652
rect 30484 5370 30512 5646
rect 30472 5364 30524 5370
rect 30472 5306 30524 5312
rect 31956 4162 31984 23802
rect 32048 21418 32076 38694
rect 32140 37670 32168 38694
rect 32128 37664 32180 37670
rect 32128 37606 32180 37612
rect 32140 37466 32168 37606
rect 32128 37460 32180 37466
rect 32128 37402 32180 37408
rect 32232 26081 32260 40326
rect 32312 39840 32364 39846
rect 32312 39782 32364 39788
rect 32324 39438 32352 39782
rect 32416 39438 32444 40326
rect 32508 40186 32536 40326
rect 32496 40180 32548 40186
rect 32496 40122 32548 40128
rect 32496 40044 32548 40050
rect 32692 40032 32720 40530
rect 32548 40004 32720 40032
rect 32496 39986 32548 39992
rect 32680 39840 32732 39846
rect 32680 39782 32732 39788
rect 32692 39506 32720 39782
rect 32680 39500 32732 39506
rect 32680 39442 32732 39448
rect 32312 39432 32364 39438
rect 32312 39374 32364 39380
rect 32404 39432 32456 39438
rect 32404 39374 32456 39380
rect 32784 39030 32812 40870
rect 33060 40526 33088 46310
rect 33152 46170 33180 46990
rect 33322 46951 33378 46960
rect 33232 46912 33284 46918
rect 33232 46854 33284 46860
rect 33600 46912 33652 46918
rect 33600 46854 33652 46860
rect 33140 46164 33192 46170
rect 33140 46106 33192 46112
rect 33140 42696 33192 42702
rect 33140 42638 33192 42644
rect 33152 40662 33180 42638
rect 33244 42344 33272 46854
rect 33324 46572 33376 46578
rect 33324 46514 33376 46520
rect 33336 45558 33364 46514
rect 33416 46368 33468 46374
rect 33416 46310 33468 46316
rect 33324 45552 33376 45558
rect 33324 45494 33376 45500
rect 33244 42316 33364 42344
rect 33232 42220 33284 42226
rect 33232 42162 33284 42168
rect 33244 41546 33272 42162
rect 33336 42090 33364 42316
rect 33324 42084 33376 42090
rect 33324 42026 33376 42032
rect 33322 41848 33378 41857
rect 33322 41783 33378 41792
rect 33336 41682 33364 41783
rect 33324 41676 33376 41682
rect 33324 41618 33376 41624
rect 33232 41540 33284 41546
rect 33232 41482 33284 41488
rect 33324 41472 33376 41478
rect 33324 41414 33376 41420
rect 33232 41268 33284 41274
rect 33232 41210 33284 41216
rect 33244 41138 33272 41210
rect 33232 41132 33284 41138
rect 33232 41074 33284 41080
rect 33140 40656 33192 40662
rect 33140 40598 33192 40604
rect 33232 40656 33284 40662
rect 33232 40598 33284 40604
rect 33048 40520 33100 40526
rect 33048 40462 33100 40468
rect 33244 40118 33272 40598
rect 33336 40526 33364 41414
rect 33428 41002 33456 46310
rect 33508 45824 33560 45830
rect 33508 45766 33560 45772
rect 33520 45626 33548 45766
rect 33508 45620 33560 45626
rect 33508 45562 33560 45568
rect 33612 43654 33640 46854
rect 33600 43648 33652 43654
rect 33600 43590 33652 43596
rect 33600 42628 33652 42634
rect 33600 42570 33652 42576
rect 33508 42560 33560 42566
rect 33508 42502 33560 42508
rect 33520 42294 33548 42502
rect 33612 42362 33640 42570
rect 33600 42356 33652 42362
rect 33600 42298 33652 42304
rect 33508 42288 33560 42294
rect 33508 42230 33560 42236
rect 33508 42084 33560 42090
rect 33508 42026 33560 42032
rect 33416 40996 33468 41002
rect 33416 40938 33468 40944
rect 33324 40520 33376 40526
rect 33324 40462 33376 40468
rect 33520 40118 33548 42026
rect 33600 41608 33652 41614
rect 33600 41550 33652 41556
rect 33612 40905 33640 41550
rect 33704 41206 33732 47398
rect 33784 47184 33836 47190
rect 33784 47126 33836 47132
rect 33692 41200 33744 41206
rect 33692 41142 33744 41148
rect 33598 40896 33654 40905
rect 33598 40831 33654 40840
rect 33692 40452 33744 40458
rect 33692 40394 33744 40400
rect 33600 40384 33652 40390
rect 33600 40326 33652 40332
rect 33232 40112 33284 40118
rect 33232 40054 33284 40060
rect 33508 40112 33560 40118
rect 33508 40054 33560 40060
rect 32864 40044 32916 40050
rect 32864 39986 32916 39992
rect 32876 39438 32904 39986
rect 33612 39506 33640 40326
rect 33600 39500 33652 39506
rect 33600 39442 33652 39448
rect 32864 39432 32916 39438
rect 32864 39374 32916 39380
rect 32864 39296 32916 39302
rect 32864 39238 32916 39244
rect 33324 39296 33376 39302
rect 33324 39238 33376 39244
rect 32772 39024 32824 39030
rect 32772 38966 32824 38972
rect 32680 38412 32732 38418
rect 32680 38354 32732 38360
rect 32692 38010 32720 38354
rect 32876 38350 32904 39238
rect 33336 38350 33364 39238
rect 33704 39030 33732 40394
rect 33796 39438 33824 47126
rect 33888 41750 33916 47466
rect 33980 46578 34008 48078
rect 34072 47666 34100 48486
rect 34152 48000 34204 48006
rect 34152 47942 34204 47948
rect 34060 47660 34112 47666
rect 34060 47602 34112 47608
rect 34072 47462 34100 47602
rect 34060 47456 34112 47462
rect 34060 47398 34112 47404
rect 34072 47054 34100 47398
rect 34060 47048 34112 47054
rect 34060 46990 34112 46996
rect 33968 46572 34020 46578
rect 33968 46514 34020 46520
rect 33980 46442 34008 46514
rect 33968 46436 34020 46442
rect 33968 46378 34020 46384
rect 33968 43648 34020 43654
rect 33968 43590 34020 43596
rect 33980 42566 34008 43590
rect 34060 42628 34112 42634
rect 34060 42570 34112 42576
rect 33968 42560 34020 42566
rect 33968 42502 34020 42508
rect 33980 42226 34008 42502
rect 33968 42220 34020 42226
rect 33968 42162 34020 42168
rect 33876 41744 33928 41750
rect 33876 41686 33928 41692
rect 33876 41540 33928 41546
rect 33980 41528 34008 42162
rect 33928 41500 34008 41528
rect 33876 41482 33928 41488
rect 33888 41070 33916 41482
rect 34072 41478 34100 42570
rect 34060 41472 34112 41478
rect 34060 41414 34112 41420
rect 33968 41132 34020 41138
rect 34072 41120 34100 41414
rect 34020 41092 34100 41120
rect 33968 41074 34020 41080
rect 33876 41064 33928 41070
rect 33876 41006 33928 41012
rect 33888 40662 33916 41006
rect 33876 40656 33928 40662
rect 33876 40598 33928 40604
rect 33876 40384 33928 40390
rect 33876 40326 33928 40332
rect 33784 39432 33836 39438
rect 33784 39374 33836 39380
rect 33888 39030 33916 40326
rect 33980 40118 34008 41074
rect 34164 40118 34192 47942
rect 34244 47524 34296 47530
rect 34244 47466 34296 47472
rect 34256 46714 34284 47466
rect 34348 46714 34376 52838
rect 34520 52624 34572 52630
rect 34520 52566 34572 52572
rect 34532 51074 34560 52566
rect 34532 51046 34652 51074
rect 34428 48544 34480 48550
rect 34428 48486 34480 48492
rect 34440 48314 34468 48486
rect 34440 48286 34560 48314
rect 34532 47666 34560 48286
rect 34520 47660 34572 47666
rect 34520 47602 34572 47608
rect 34428 47048 34480 47054
rect 34428 46990 34480 46996
rect 34244 46708 34296 46714
rect 34244 46650 34296 46656
rect 34336 46708 34388 46714
rect 34336 46650 34388 46656
rect 34244 46572 34296 46578
rect 34244 46514 34296 46520
rect 34256 46102 34284 46514
rect 34244 46096 34296 46102
rect 34244 46038 34296 46044
rect 34336 43104 34388 43110
rect 34336 43046 34388 43052
rect 34244 42628 34296 42634
rect 34244 42570 34296 42576
rect 34256 41018 34284 42570
rect 34348 41857 34376 43046
rect 34334 41848 34390 41857
rect 34334 41783 34390 41792
rect 34348 41750 34376 41783
rect 34336 41744 34388 41750
rect 34336 41686 34388 41692
rect 34256 40990 34376 41018
rect 34244 40928 34296 40934
rect 34244 40870 34296 40876
rect 33968 40112 34020 40118
rect 33966 40080 33968 40089
rect 34152 40112 34204 40118
rect 34020 40080 34022 40089
rect 34152 40054 34204 40060
rect 33966 40015 34022 40024
rect 34256 39438 34284 40870
rect 34244 39432 34296 39438
rect 34244 39374 34296 39380
rect 33692 39024 33744 39030
rect 33692 38966 33744 38972
rect 33876 39024 33928 39030
rect 33876 38966 33928 38972
rect 32864 38344 32916 38350
rect 32864 38286 32916 38292
rect 33324 38344 33376 38350
rect 33324 38286 33376 38292
rect 32864 38208 32916 38214
rect 32864 38150 32916 38156
rect 33416 38208 33468 38214
rect 33416 38150 33468 38156
rect 32588 38004 32640 38010
rect 32588 37946 32640 37952
rect 32680 38004 32732 38010
rect 32680 37946 32732 37952
rect 32312 37460 32364 37466
rect 32312 37402 32364 37408
rect 32324 36310 32352 37402
rect 32312 36304 32364 36310
rect 32312 36246 32364 36252
rect 32312 36100 32364 36106
rect 32312 36042 32364 36048
rect 32324 34678 32352 36042
rect 32600 36038 32628 37946
rect 32588 36032 32640 36038
rect 32588 35974 32640 35980
rect 32312 34672 32364 34678
rect 32312 34614 32364 34620
rect 32324 34202 32352 34614
rect 32312 34196 32364 34202
rect 32312 34138 32364 34144
rect 32600 32434 32628 35974
rect 32588 32428 32640 32434
rect 32588 32370 32640 32376
rect 32404 30932 32456 30938
rect 32404 30874 32456 30880
rect 32218 26072 32274 26081
rect 32218 26007 32274 26016
rect 32416 25498 32444 30874
rect 32876 26042 32904 38150
rect 33230 37904 33286 37913
rect 33048 37868 33100 37874
rect 33230 37839 33232 37848
rect 33048 37810 33100 37816
rect 33284 37839 33286 37848
rect 33232 37810 33284 37816
rect 33060 37670 33088 37810
rect 33048 37664 33100 37670
rect 33048 37606 33100 37612
rect 33060 37126 33088 37606
rect 33232 37188 33284 37194
rect 33232 37130 33284 37136
rect 33048 37120 33100 37126
rect 33048 37062 33100 37068
rect 33060 36378 33088 37062
rect 33244 36582 33272 37130
rect 33232 36576 33284 36582
rect 33230 36544 33232 36553
rect 33284 36544 33286 36553
rect 33230 36479 33286 36488
rect 33048 36372 33100 36378
rect 33048 36314 33100 36320
rect 33048 28212 33100 28218
rect 33048 28154 33100 28160
rect 32864 26036 32916 26042
rect 32864 25978 32916 25984
rect 33060 25838 33088 28154
rect 33428 26194 33456 38150
rect 34348 38010 34376 40990
rect 34440 40497 34468 46990
rect 34532 46918 34560 47602
rect 34520 46912 34572 46918
rect 34520 46854 34572 46860
rect 34624 43450 34652 51046
rect 34716 46986 34744 52906
rect 34704 46980 34756 46986
rect 34704 46922 34756 46928
rect 34612 43444 34664 43450
rect 34612 43386 34664 43392
rect 34624 42022 34652 43386
rect 34808 42634 34836 52974
rect 35348 52896 35400 52902
rect 35348 52838 35400 52844
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34888 48000 34940 48006
rect 34888 47942 34940 47948
rect 34900 47462 34928 47942
rect 35360 47802 35388 52838
rect 36648 52698 36676 53042
rect 38844 52896 38896 52902
rect 38844 52838 38896 52844
rect 38936 52896 38988 52902
rect 38936 52838 38988 52844
rect 36636 52692 36688 52698
rect 36636 52634 36688 52640
rect 38660 49224 38712 49230
rect 38660 49166 38712 49172
rect 35624 48544 35676 48550
rect 35624 48486 35676 48492
rect 35348 47796 35400 47802
rect 35348 47738 35400 47744
rect 35440 47796 35492 47802
rect 35440 47738 35492 47744
rect 35452 47530 35480 47738
rect 35440 47524 35492 47530
rect 35440 47466 35492 47472
rect 34888 47456 34940 47462
rect 34888 47398 34940 47404
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 35636 47025 35664 48486
rect 35808 47456 35860 47462
rect 35808 47398 35860 47404
rect 35820 47190 35848 47398
rect 35808 47184 35860 47190
rect 35808 47126 35860 47132
rect 35622 47016 35678 47025
rect 35622 46951 35678 46960
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 35636 46170 35664 46951
rect 35624 46164 35676 46170
rect 35624 46106 35676 46112
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 35440 43104 35492 43110
rect 35440 43046 35492 43052
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34796 42628 34848 42634
rect 34796 42570 34848 42576
rect 34796 42356 34848 42362
rect 34796 42298 34848 42304
rect 34702 42256 34758 42265
rect 34702 42191 34758 42200
rect 34716 42090 34744 42191
rect 34704 42084 34756 42090
rect 34704 42026 34756 42032
rect 34612 42016 34664 42022
rect 34612 41958 34664 41964
rect 34808 41614 34836 42298
rect 35452 42294 35480 43046
rect 35532 42764 35584 42770
rect 35532 42706 35584 42712
rect 35544 42566 35572 42706
rect 35532 42560 35584 42566
rect 35532 42502 35584 42508
rect 35544 42362 35572 42502
rect 38672 42362 38700 49166
rect 38752 48680 38804 48686
rect 38752 48622 38804 48628
rect 35532 42356 35584 42362
rect 35532 42298 35584 42304
rect 38660 42356 38712 42362
rect 38660 42298 38712 42304
rect 35440 42288 35492 42294
rect 35440 42230 35492 42236
rect 35348 42016 35400 42022
rect 35348 41958 35400 41964
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 35360 41818 35388 41958
rect 35348 41812 35400 41818
rect 35268 41772 35348 41800
rect 34796 41608 34848 41614
rect 34796 41550 34848 41556
rect 35268 41274 35296 41772
rect 35348 41754 35400 41760
rect 35452 41546 35480 42230
rect 35530 41712 35586 41721
rect 38764 41682 38792 48622
rect 38856 48278 38884 52838
rect 38844 48272 38896 48278
rect 38844 48214 38896 48220
rect 38948 47734 38976 52838
rect 39040 52698 39068 53042
rect 41236 52896 41288 52902
rect 41236 52838 41288 52844
rect 39028 52692 39080 52698
rect 39028 52634 39080 52640
rect 41248 52630 41276 52838
rect 42352 52698 42380 53042
rect 42616 52896 42668 52902
rect 42616 52838 42668 52844
rect 42340 52692 42392 52698
rect 42340 52634 42392 52640
rect 41236 52624 41288 52630
rect 41236 52566 41288 52572
rect 42628 52562 42656 52838
rect 43640 52698 43668 53042
rect 43904 53032 43956 53038
rect 43904 52974 43956 52980
rect 43628 52692 43680 52698
rect 43628 52634 43680 52640
rect 42616 52556 42668 52562
rect 42616 52498 42668 52504
rect 38936 47728 38988 47734
rect 38936 47670 38988 47676
rect 35530 41647 35586 41656
rect 36820 41676 36872 41682
rect 35440 41540 35492 41546
rect 35440 41482 35492 41488
rect 35348 41472 35400 41478
rect 35348 41414 35400 41420
rect 35256 41268 35308 41274
rect 35256 41210 35308 41216
rect 35254 41168 35310 41177
rect 35254 41103 35256 41112
rect 35308 41103 35310 41112
rect 35256 41074 35308 41080
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35360 40526 35388 41414
rect 35348 40520 35400 40526
rect 34426 40488 34482 40497
rect 34426 40423 34482 40432
rect 34610 40488 34666 40497
rect 35348 40462 35400 40468
rect 34610 40423 34666 40432
rect 34796 40452 34848 40458
rect 34624 40390 34652 40423
rect 34796 40394 34848 40400
rect 34612 40384 34664 40390
rect 34612 40326 34664 40332
rect 34428 39568 34480 39574
rect 34428 39510 34480 39516
rect 34440 38418 34468 39510
rect 34520 38752 34572 38758
rect 34520 38694 34572 38700
rect 34428 38412 34480 38418
rect 34428 38354 34480 38360
rect 34336 38004 34388 38010
rect 34336 37946 34388 37952
rect 34348 37777 34376 37946
rect 34334 37768 34390 37777
rect 34334 37703 34390 37712
rect 33784 37324 33836 37330
rect 33784 37266 33836 37272
rect 33796 37233 33824 37266
rect 33782 37224 33838 37233
rect 33782 37159 33838 37168
rect 33692 35828 33744 35834
rect 33692 35770 33744 35776
rect 33704 35630 33732 35770
rect 33692 35624 33744 35630
rect 33692 35566 33744 35572
rect 33508 34944 33560 34950
rect 33506 34912 33508 34921
rect 33560 34912 33562 34921
rect 33506 34847 33562 34856
rect 33520 28490 33548 34847
rect 33796 31210 33824 37159
rect 33784 31204 33836 31210
rect 33784 31146 33836 31152
rect 33508 28484 33560 28490
rect 33508 28426 33560 28432
rect 33784 27328 33836 27334
rect 33784 27270 33836 27276
rect 33428 26166 33548 26194
rect 33416 26036 33468 26042
rect 33416 25978 33468 25984
rect 33048 25832 33100 25838
rect 33048 25774 33100 25780
rect 32864 25764 32916 25770
rect 32864 25706 32916 25712
rect 32404 25492 32456 25498
rect 32404 25434 32456 25440
rect 32312 24132 32364 24138
rect 32312 24074 32364 24080
rect 32220 24064 32272 24070
rect 32220 24006 32272 24012
rect 32128 23656 32180 23662
rect 32128 23598 32180 23604
rect 32140 22574 32168 23598
rect 32232 22642 32260 24006
rect 32324 22778 32352 24074
rect 32416 23866 32444 25434
rect 32588 25220 32640 25226
rect 32588 25162 32640 25168
rect 32404 23860 32456 23866
rect 32404 23802 32456 23808
rect 32404 23656 32456 23662
rect 32404 23598 32456 23604
rect 32416 23322 32444 23598
rect 32404 23316 32456 23322
rect 32404 23258 32456 23264
rect 32312 22772 32364 22778
rect 32312 22714 32364 22720
rect 32416 22642 32444 23258
rect 32220 22636 32272 22642
rect 32220 22578 32272 22584
rect 32404 22636 32456 22642
rect 32404 22578 32456 22584
rect 32128 22568 32180 22574
rect 32128 22510 32180 22516
rect 32312 22024 32364 22030
rect 32312 21966 32364 21972
rect 32036 21412 32088 21418
rect 32036 21354 32088 21360
rect 32324 21010 32352 21966
rect 32416 21486 32444 22578
rect 32600 22506 32628 25162
rect 32876 24818 32904 25706
rect 33140 25288 33192 25294
rect 33140 25230 33192 25236
rect 33152 24954 33180 25230
rect 33324 25152 33376 25158
rect 33324 25094 33376 25100
rect 33140 24948 33192 24954
rect 33140 24890 33192 24896
rect 33336 24886 33364 25094
rect 33324 24880 33376 24886
rect 33324 24822 33376 24828
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 33232 24064 33284 24070
rect 33232 24006 33284 24012
rect 33140 22976 33192 22982
rect 33140 22918 33192 22924
rect 33152 22778 33180 22918
rect 33140 22772 33192 22778
rect 33140 22714 33192 22720
rect 32772 22568 32824 22574
rect 32772 22510 32824 22516
rect 32864 22568 32916 22574
rect 32864 22510 32916 22516
rect 32588 22500 32640 22506
rect 32588 22442 32640 22448
rect 32600 21894 32628 22442
rect 32784 22234 32812 22510
rect 32772 22228 32824 22234
rect 32772 22170 32824 22176
rect 32876 22166 32904 22510
rect 32864 22160 32916 22166
rect 33244 22137 33272 24006
rect 33324 22772 33376 22778
rect 33324 22714 33376 22720
rect 32864 22102 32916 22108
rect 33230 22128 33286 22137
rect 33230 22063 33286 22072
rect 33336 22030 33364 22714
rect 33428 22710 33456 25978
rect 33520 24041 33548 26166
rect 33598 26072 33654 26081
rect 33598 26007 33600 26016
rect 33652 26007 33654 26016
rect 33600 25978 33652 25984
rect 33612 25294 33640 25978
rect 33600 25288 33652 25294
rect 33598 25256 33600 25265
rect 33652 25256 33654 25265
rect 33598 25191 33654 25200
rect 33692 24812 33744 24818
rect 33692 24754 33744 24760
rect 33600 24744 33652 24750
rect 33600 24686 33652 24692
rect 33612 24614 33640 24686
rect 33600 24608 33652 24614
rect 33600 24550 33652 24556
rect 33612 24274 33640 24550
rect 33704 24410 33732 24754
rect 33692 24404 33744 24410
rect 33692 24346 33744 24352
rect 33600 24268 33652 24274
rect 33600 24210 33652 24216
rect 33506 24032 33562 24041
rect 33506 23967 33562 23976
rect 33506 23896 33562 23905
rect 33506 23831 33562 23840
rect 33416 22704 33468 22710
rect 33416 22646 33468 22652
rect 33140 22024 33192 22030
rect 33140 21966 33192 21972
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 32588 21888 32640 21894
rect 32588 21830 32640 21836
rect 32496 21548 32548 21554
rect 32496 21490 32548 21496
rect 32404 21480 32456 21486
rect 32404 21422 32456 21428
rect 32312 21004 32364 21010
rect 32312 20946 32364 20952
rect 32036 20936 32088 20942
rect 32036 20878 32088 20884
rect 32048 18970 32076 20878
rect 32220 20392 32272 20398
rect 32220 20334 32272 20340
rect 32126 19680 32182 19689
rect 32126 19615 32182 19624
rect 32140 19310 32168 19615
rect 32232 19514 32260 20334
rect 32324 20058 32352 20946
rect 32312 20052 32364 20058
rect 32312 19994 32364 20000
rect 32508 19990 32536 21490
rect 32600 21146 32628 21830
rect 32864 21344 32916 21350
rect 32864 21286 32916 21292
rect 32588 21140 32640 21146
rect 32588 21082 32640 21088
rect 32876 20942 32904 21286
rect 32864 20936 32916 20942
rect 32864 20878 32916 20884
rect 32864 20800 32916 20806
rect 32864 20742 32916 20748
rect 32496 19984 32548 19990
rect 32496 19926 32548 19932
rect 32220 19508 32272 19514
rect 32220 19450 32272 19456
rect 32128 19304 32180 19310
rect 32128 19246 32180 19252
rect 32312 19168 32364 19174
rect 32312 19110 32364 19116
rect 32036 18964 32088 18970
rect 32036 18906 32088 18912
rect 32034 18728 32090 18737
rect 32034 18663 32090 18672
rect 32048 16046 32076 18663
rect 32324 18086 32352 19110
rect 32876 18834 32904 20742
rect 33152 19496 33180 21966
rect 33060 19468 33180 19496
rect 33060 18902 33088 19468
rect 33140 19372 33192 19378
rect 33520 19334 33548 23831
rect 33612 23118 33640 24210
rect 33796 23322 33824 27270
rect 34532 27130 34560 38694
rect 34624 37670 34652 40326
rect 34612 37664 34664 37670
rect 34612 37606 34664 37612
rect 34520 27124 34572 27130
rect 34520 27066 34572 27072
rect 34336 26784 34388 26790
rect 34336 26726 34388 26732
rect 34348 26586 34376 26726
rect 34336 26580 34388 26586
rect 34336 26522 34388 26528
rect 34348 25294 34376 26522
rect 34428 26240 34480 26246
rect 34428 26182 34480 26188
rect 34440 25838 34468 26182
rect 34532 26058 34560 27066
rect 34532 26030 34652 26058
rect 34520 25900 34572 25906
rect 34520 25842 34572 25848
rect 34428 25832 34480 25838
rect 34428 25774 34480 25780
rect 34440 25294 34468 25774
rect 34336 25288 34388 25294
rect 34336 25230 34388 25236
rect 34428 25288 34480 25294
rect 34428 25230 34480 25236
rect 33968 25220 34020 25226
rect 33968 25162 34020 25168
rect 33876 25152 33928 25158
rect 33876 25094 33928 25100
rect 33888 24410 33916 25094
rect 33876 24404 33928 24410
rect 33876 24346 33928 24352
rect 33888 24206 33916 24346
rect 33876 24200 33928 24206
rect 33876 24142 33928 24148
rect 33980 24154 34008 25162
rect 34152 24812 34204 24818
rect 34152 24754 34204 24760
rect 34164 24206 34192 24754
rect 34244 24404 34296 24410
rect 34244 24346 34296 24352
rect 34152 24200 34204 24206
rect 33980 24138 34100 24154
rect 34152 24142 34204 24148
rect 33980 24132 34112 24138
rect 33980 24126 34060 24132
rect 34060 24074 34112 24080
rect 33876 24064 33928 24070
rect 33876 24006 33928 24012
rect 33784 23316 33836 23322
rect 33784 23258 33836 23264
rect 33784 23180 33836 23186
rect 33784 23122 33836 23128
rect 33600 23112 33652 23118
rect 33600 23054 33652 23060
rect 33692 21888 33744 21894
rect 33692 21830 33744 21836
rect 33600 20392 33652 20398
rect 33600 20334 33652 20340
rect 33140 19314 33192 19320
rect 33048 18896 33100 18902
rect 33048 18838 33100 18844
rect 32864 18828 32916 18834
rect 32864 18770 32916 18776
rect 32496 18760 32548 18766
rect 32496 18702 32548 18708
rect 32508 18290 32536 18702
rect 32680 18624 32732 18630
rect 32680 18566 32732 18572
rect 32692 18290 32720 18566
rect 32876 18290 32904 18770
rect 32496 18284 32548 18290
rect 32496 18226 32548 18232
rect 32680 18284 32732 18290
rect 32680 18226 32732 18232
rect 32864 18284 32916 18290
rect 32864 18226 32916 18232
rect 33152 18154 33180 19314
rect 33336 19306 33548 19334
rect 33232 18216 33284 18222
rect 33232 18158 33284 18164
rect 33140 18148 33192 18154
rect 33140 18090 33192 18096
rect 32312 18080 32364 18086
rect 32312 18022 32364 18028
rect 33140 17740 33192 17746
rect 33140 17682 33192 17688
rect 32312 17672 32364 17678
rect 32312 17614 32364 17620
rect 32402 17640 32458 17649
rect 32324 16998 32352 17614
rect 32402 17575 32458 17584
rect 32416 17542 32444 17575
rect 32404 17536 32456 17542
rect 32404 17478 32456 17484
rect 32312 16992 32364 16998
rect 32312 16934 32364 16940
rect 32324 16658 32352 16934
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 32036 16040 32088 16046
rect 32324 16017 32352 16050
rect 32036 15982 32088 15988
rect 32310 16008 32366 16017
rect 32416 15994 32444 17478
rect 33152 16794 33180 17682
rect 33244 17270 33272 18158
rect 33232 17264 33284 17270
rect 33232 17206 33284 17212
rect 33140 16788 33192 16794
rect 33140 16730 33192 16736
rect 32956 16720 33008 16726
rect 32956 16662 33008 16668
rect 32494 16144 32550 16153
rect 32968 16114 32996 16662
rect 33048 16652 33100 16658
rect 33048 16594 33100 16600
rect 33060 16114 33088 16594
rect 33336 16538 33364 19306
rect 33416 19168 33468 19174
rect 33416 19110 33468 19116
rect 33428 16658 33456 19110
rect 33508 18828 33560 18834
rect 33508 18770 33560 18776
rect 33520 18358 33548 18770
rect 33508 18352 33560 18358
rect 33508 18294 33560 18300
rect 33612 18222 33640 20334
rect 33704 19242 33732 21830
rect 33796 21010 33824 23122
rect 33888 22094 33916 24006
rect 34072 23730 34100 24074
rect 34256 23730 34284 24346
rect 34336 24064 34388 24070
rect 34336 24006 34388 24012
rect 34060 23724 34112 23730
rect 34060 23666 34112 23672
rect 34244 23724 34296 23730
rect 34244 23666 34296 23672
rect 34072 23610 34100 23666
rect 34072 23582 34192 23610
rect 34348 23594 34376 24006
rect 34532 23866 34560 25842
rect 34624 24206 34652 26030
rect 34704 25696 34756 25702
rect 34704 25638 34756 25644
rect 34716 25362 34744 25638
rect 34704 25356 34756 25362
rect 34704 25298 34756 25304
rect 34704 24336 34756 24342
rect 34704 24278 34756 24284
rect 34612 24200 34664 24206
rect 34612 24142 34664 24148
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 34060 23316 34112 23322
rect 34060 23258 34112 23264
rect 33888 22066 34008 22094
rect 33784 21004 33836 21010
rect 33784 20946 33836 20952
rect 33692 19236 33744 19242
rect 33692 19178 33744 19184
rect 33704 18748 33732 19178
rect 33876 18828 33928 18834
rect 33876 18770 33928 18776
rect 33784 18760 33836 18766
rect 33704 18720 33784 18748
rect 33704 18630 33732 18720
rect 33784 18702 33836 18708
rect 33692 18624 33744 18630
rect 33692 18566 33744 18572
rect 33888 18290 33916 18770
rect 33876 18284 33928 18290
rect 33876 18226 33928 18232
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 33506 17096 33562 17105
rect 33506 17031 33562 17040
rect 33520 16658 33548 17031
rect 33416 16652 33468 16658
rect 33416 16594 33468 16600
rect 33508 16652 33560 16658
rect 33508 16594 33560 16600
rect 33600 16584 33652 16590
rect 33336 16532 33600 16538
rect 33336 16526 33652 16532
rect 33336 16510 33640 16526
rect 33692 16516 33744 16522
rect 32956 16108 33008 16114
rect 32494 16079 32496 16088
rect 32548 16079 32550 16088
rect 32496 16050 32548 16056
rect 32784 16068 32956 16096
rect 32416 15966 32536 15994
rect 32310 15943 32366 15952
rect 32220 15496 32272 15502
rect 32324 15484 32352 15943
rect 32272 15456 32352 15484
rect 32220 15438 32272 15444
rect 32036 14476 32088 14482
rect 32036 14418 32088 14424
rect 32048 14074 32076 14418
rect 32128 14408 32180 14414
rect 32128 14350 32180 14356
rect 32036 14068 32088 14074
rect 32036 14010 32088 14016
rect 32140 13938 32168 14350
rect 32128 13932 32180 13938
rect 32128 13874 32180 13880
rect 32140 13530 32168 13874
rect 32402 13696 32458 13705
rect 32402 13631 32458 13640
rect 32128 13524 32180 13530
rect 32128 13466 32180 13472
rect 32128 12980 32180 12986
rect 32128 12922 32180 12928
rect 32140 12646 32168 12922
rect 32416 12782 32444 13631
rect 32404 12776 32456 12782
rect 32402 12744 32404 12753
rect 32456 12744 32458 12753
rect 32220 12708 32272 12714
rect 32402 12679 32458 12688
rect 32220 12650 32272 12656
rect 32128 12640 32180 12646
rect 32128 12582 32180 12588
rect 32128 12300 32180 12306
rect 32128 12242 32180 12248
rect 32036 11280 32088 11286
rect 32034 11248 32036 11257
rect 32088 11248 32090 11257
rect 32034 11183 32090 11192
rect 32036 11144 32088 11150
rect 32036 11086 32088 11092
rect 32048 9586 32076 11086
rect 32036 9580 32088 9586
rect 32036 9522 32088 9528
rect 32140 9450 32168 12242
rect 32128 9444 32180 9450
rect 32128 9386 32180 9392
rect 32036 9376 32088 9382
rect 32036 9318 32088 9324
rect 32048 8634 32076 9318
rect 32140 8838 32168 9386
rect 32128 8832 32180 8838
rect 32128 8774 32180 8780
rect 32036 8628 32088 8634
rect 32036 8570 32088 8576
rect 32232 8090 32260 12650
rect 32312 12640 32364 12646
rect 32312 12582 32364 12588
rect 32324 10606 32352 12582
rect 32312 10600 32364 10606
rect 32312 10542 32364 10548
rect 32310 9072 32366 9081
rect 32310 9007 32312 9016
rect 32364 9007 32366 9016
rect 32312 8978 32364 8984
rect 32324 8090 32352 8978
rect 32220 8084 32272 8090
rect 32220 8026 32272 8032
rect 32312 8084 32364 8090
rect 32312 8026 32364 8032
rect 30380 4140 30432 4146
rect 30380 4082 30432 4088
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 31680 4134 31984 4162
rect 30944 3942 30972 4082
rect 30932 3936 30984 3942
rect 30932 3878 30984 3884
rect 30288 3664 30340 3670
rect 30288 3606 30340 3612
rect 30380 3664 30432 3670
rect 30380 3606 30432 3612
rect 28816 3188 28868 3194
rect 28816 3130 28868 3136
rect 29644 3188 29696 3194
rect 29644 3130 29696 3136
rect 29920 3188 29972 3194
rect 29920 3130 29972 3136
rect 28828 3058 28856 3130
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 28552 2746 28672 2774
rect 28552 2446 28580 2746
rect 28908 2576 28960 2582
rect 28908 2518 28960 2524
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 28540 2304 28592 2310
rect 28540 2246 28592 2252
rect 28552 800 28580 2246
rect 28920 800 28948 2518
rect 29656 2446 29684 3130
rect 29932 2446 29960 3130
rect 30012 2848 30064 2854
rect 30012 2790 30064 2796
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 29920 2440 29972 2446
rect 29920 2382 29972 2388
rect 29276 2304 29328 2310
rect 29276 2246 29328 2252
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 29288 800 29316 2246
rect 29656 800 29684 2246
rect 30024 800 30052 2790
rect 30300 2650 30328 3606
rect 30392 3058 30420 3606
rect 30380 3052 30432 3058
rect 30380 2994 30432 3000
rect 30748 2848 30800 2854
rect 30748 2790 30800 2796
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 30380 2576 30432 2582
rect 30380 2518 30432 2524
rect 30392 800 30420 2518
rect 30760 800 30788 2790
rect 30944 2446 30972 3878
rect 31680 3670 31708 4134
rect 31760 3732 31812 3738
rect 31760 3674 31812 3680
rect 31668 3664 31720 3670
rect 31668 3606 31720 3612
rect 31772 3058 31800 3674
rect 31852 3664 31904 3670
rect 31852 3606 31904 3612
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 31484 2916 31536 2922
rect 31484 2858 31536 2864
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 31116 2304 31168 2310
rect 31116 2246 31168 2252
rect 31128 800 31156 2246
rect 31496 800 31524 2858
rect 31864 2774 31892 3606
rect 32232 2990 32260 8026
rect 32416 4554 32444 12679
rect 32508 10538 32536 15966
rect 32680 14884 32732 14890
rect 32680 14826 32732 14832
rect 32692 14278 32720 14826
rect 32680 14272 32732 14278
rect 32680 14214 32732 14220
rect 32680 13252 32732 13258
rect 32680 13194 32732 13200
rect 32586 12880 32642 12889
rect 32586 12815 32588 12824
rect 32640 12815 32642 12824
rect 32588 12786 32640 12792
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 32600 11121 32628 11630
rect 32586 11112 32642 11121
rect 32586 11047 32588 11056
rect 32640 11047 32642 11056
rect 32588 11018 32640 11024
rect 32692 11014 32720 13194
rect 32784 12918 32812 16068
rect 32956 16050 33008 16056
rect 33048 16108 33100 16114
rect 33048 16050 33100 16056
rect 33140 15904 33192 15910
rect 33140 15846 33192 15852
rect 33324 15904 33376 15910
rect 33324 15846 33376 15852
rect 33152 15570 33180 15846
rect 33140 15564 33192 15570
rect 33140 15506 33192 15512
rect 32956 14476 33008 14482
rect 32956 14418 33008 14424
rect 32864 14408 32916 14414
rect 32864 14350 32916 14356
rect 32876 13530 32904 14350
rect 32968 13870 32996 14418
rect 32956 13864 33008 13870
rect 32956 13806 33008 13812
rect 32864 13524 32916 13530
rect 32864 13466 32916 13472
rect 32772 12912 32824 12918
rect 32772 12854 32824 12860
rect 32772 12776 32824 12782
rect 32772 12718 32824 12724
rect 32680 11008 32732 11014
rect 32680 10950 32732 10956
rect 32692 10690 32720 10950
rect 32784 10810 32812 12718
rect 32864 11620 32916 11626
rect 32864 11562 32916 11568
rect 32876 11218 32904 11562
rect 32864 11212 32916 11218
rect 32864 11154 32916 11160
rect 32968 11082 32996 13806
rect 33140 13388 33192 13394
rect 33140 13330 33192 13336
rect 33048 13184 33100 13190
rect 33048 13126 33100 13132
rect 32956 11076 33008 11082
rect 32956 11018 33008 11024
rect 32772 10804 32824 10810
rect 32772 10746 32824 10752
rect 32770 10704 32826 10713
rect 32692 10662 32770 10690
rect 32770 10639 32772 10648
rect 32824 10639 32826 10648
rect 32772 10610 32824 10616
rect 32496 10532 32548 10538
rect 32496 10474 32548 10480
rect 32784 10062 32812 10610
rect 33060 10198 33088 13126
rect 33152 12850 33180 13330
rect 33140 12844 33192 12850
rect 33140 12786 33192 12792
rect 33336 12434 33364 15846
rect 33428 13569 33456 16510
rect 33692 16458 33744 16464
rect 33704 15706 33732 16458
rect 33692 15700 33744 15706
rect 33692 15642 33744 15648
rect 33600 15632 33652 15638
rect 33652 15580 33732 15586
rect 33600 15574 33732 15580
rect 33612 15558 33732 15574
rect 33704 14958 33732 15558
rect 33692 14952 33744 14958
rect 33692 14894 33744 14900
rect 33508 14816 33560 14822
rect 33508 14758 33560 14764
rect 33414 13560 33470 13569
rect 33414 13495 33470 13504
rect 33520 13394 33548 14758
rect 33704 14521 33732 14894
rect 33876 14884 33928 14890
rect 33876 14826 33928 14832
rect 33784 14816 33836 14822
rect 33784 14758 33836 14764
rect 33690 14512 33746 14521
rect 33796 14482 33824 14758
rect 33690 14447 33746 14456
rect 33784 14476 33836 14482
rect 33600 14408 33652 14414
rect 33600 14350 33652 14356
rect 33612 14278 33640 14350
rect 33600 14272 33652 14278
rect 33600 14214 33652 14220
rect 33612 13870 33640 14214
rect 33704 14006 33732 14447
rect 33784 14418 33836 14424
rect 33692 14000 33744 14006
rect 33692 13942 33744 13948
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33692 13728 33744 13734
rect 33692 13670 33744 13676
rect 33508 13388 33560 13394
rect 33508 13330 33560 13336
rect 33244 12406 33364 12434
rect 33140 12232 33192 12238
rect 33140 12174 33192 12180
rect 33152 10674 33180 12174
rect 33244 11626 33272 12406
rect 33520 12170 33548 13330
rect 33704 12782 33732 13670
rect 33784 12844 33836 12850
rect 33888 12832 33916 14826
rect 33836 12804 33916 12832
rect 33784 12786 33836 12792
rect 33692 12776 33744 12782
rect 33692 12718 33744 12724
rect 33508 12164 33560 12170
rect 33508 12106 33560 12112
rect 33520 11898 33548 12106
rect 33600 12096 33652 12102
rect 33600 12038 33652 12044
rect 33508 11892 33560 11898
rect 33508 11834 33560 11840
rect 33232 11620 33284 11626
rect 33232 11562 33284 11568
rect 33244 11098 33272 11562
rect 33416 11280 33468 11286
rect 33416 11222 33468 11228
rect 33244 11070 33364 11098
rect 33232 11008 33284 11014
rect 33232 10950 33284 10956
rect 33140 10668 33192 10674
rect 33140 10610 33192 10616
rect 33048 10192 33100 10198
rect 33048 10134 33100 10140
rect 32772 10056 32824 10062
rect 33060 10033 33088 10134
rect 33152 10062 33180 10610
rect 33140 10056 33192 10062
rect 32772 9998 32824 10004
rect 33046 10024 33102 10033
rect 33140 9998 33192 10004
rect 33046 9959 33102 9968
rect 32956 9920 33008 9926
rect 32956 9862 33008 9868
rect 32496 9580 32548 9586
rect 32496 9522 32548 9528
rect 32508 8634 32536 9522
rect 32968 9042 32996 9862
rect 32956 9036 33008 9042
rect 32956 8978 33008 8984
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 33060 6866 33088 9959
rect 33152 9722 33180 9998
rect 33140 9716 33192 9722
rect 33140 9658 33192 9664
rect 33244 8362 33272 10950
rect 33336 10062 33364 11070
rect 33428 10282 33456 11222
rect 33520 11150 33548 11834
rect 33612 11150 33640 12038
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 33600 11144 33652 11150
rect 33600 11086 33652 11092
rect 33704 11014 33732 12718
rect 33876 11552 33928 11558
rect 33876 11494 33928 11500
rect 33888 11286 33916 11494
rect 33876 11280 33928 11286
rect 33876 11222 33928 11228
rect 33692 11008 33744 11014
rect 33692 10950 33744 10956
rect 33428 10266 33732 10282
rect 33428 10260 33744 10266
rect 33428 10254 33692 10260
rect 33692 10202 33744 10208
rect 33324 10056 33376 10062
rect 33324 9998 33376 10004
rect 33784 10056 33836 10062
rect 33784 9998 33836 10004
rect 33692 9512 33744 9518
rect 33692 9454 33744 9460
rect 33598 9072 33654 9081
rect 33598 9007 33600 9016
rect 33652 9007 33654 9016
rect 33600 8978 33652 8984
rect 33324 8968 33376 8974
rect 33324 8910 33376 8916
rect 33232 8356 33284 8362
rect 33232 8298 33284 8304
rect 33336 8090 33364 8910
rect 33508 8832 33560 8838
rect 33508 8774 33560 8780
rect 33520 8498 33548 8774
rect 33704 8634 33732 9454
rect 33796 9042 33824 9998
rect 33784 9036 33836 9042
rect 33784 8978 33836 8984
rect 33692 8628 33744 8634
rect 33692 8570 33744 8576
rect 33508 8492 33560 8498
rect 33508 8434 33560 8440
rect 33324 8084 33376 8090
rect 33324 8026 33376 8032
rect 33796 7546 33824 8978
rect 33876 8832 33928 8838
rect 33874 8800 33876 8809
rect 33928 8800 33930 8809
rect 33874 8735 33930 8744
rect 33876 7880 33928 7886
rect 33876 7822 33928 7828
rect 33784 7540 33836 7546
rect 33784 7482 33836 7488
rect 33888 7002 33916 7822
rect 33876 6996 33928 7002
rect 33876 6938 33928 6944
rect 33048 6860 33100 6866
rect 33048 6802 33100 6808
rect 33060 6458 33088 6802
rect 33048 6452 33100 6458
rect 33048 6394 33100 6400
rect 32772 5568 32824 5574
rect 32772 5510 32824 5516
rect 32404 4548 32456 4554
rect 32404 4490 32456 4496
rect 32404 4276 32456 4282
rect 32404 4218 32456 4224
rect 32416 3738 32444 4218
rect 32784 4214 32812 5510
rect 32772 4208 32824 4214
rect 32772 4150 32824 4156
rect 32864 4208 32916 4214
rect 32864 4150 32916 4156
rect 32496 4140 32548 4146
rect 32496 4082 32548 4088
rect 32508 4026 32536 4082
rect 32508 3998 32720 4026
rect 32692 3942 32720 3998
rect 32680 3936 32732 3942
rect 32680 3878 32732 3884
rect 32404 3732 32456 3738
rect 32404 3674 32456 3680
rect 32220 2984 32272 2990
rect 32220 2926 32272 2932
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 31772 2746 31892 2774
rect 31772 2446 31800 2746
rect 31852 2576 31904 2582
rect 31852 2518 31904 2524
rect 31760 2440 31812 2446
rect 31760 2382 31812 2388
rect 31864 800 31892 2518
rect 32232 800 32260 2790
rect 32784 2774 32812 4150
rect 32876 3738 32904 4150
rect 33322 3768 33378 3777
rect 32864 3732 32916 3738
rect 33980 3738 34008 22066
rect 34072 12374 34100 23258
rect 34164 20466 34192 23582
rect 34336 23588 34388 23594
rect 34336 23530 34388 23536
rect 34348 23497 34376 23530
rect 34428 23520 34480 23526
rect 34334 23488 34390 23497
rect 34428 23462 34480 23468
rect 34334 23423 34390 23432
rect 34440 23322 34468 23462
rect 34428 23316 34480 23322
rect 34428 23258 34480 23264
rect 34716 23100 34744 24278
rect 34808 24070 34836 40394
rect 35544 39982 35572 41647
rect 36820 41618 36872 41624
rect 38752 41676 38804 41682
rect 38752 41618 38804 41624
rect 36268 41608 36320 41614
rect 35622 41576 35678 41585
rect 36268 41550 36320 41556
rect 35622 41511 35678 41520
rect 35636 41478 35664 41511
rect 36280 41478 36308 41550
rect 36832 41478 36860 41618
rect 35624 41472 35676 41478
rect 35624 41414 35676 41420
rect 36268 41472 36320 41478
rect 36268 41414 36320 41420
rect 36820 41472 36872 41478
rect 36820 41414 36872 41420
rect 36544 41268 36596 41274
rect 36544 41210 36596 41216
rect 35900 40996 35952 41002
rect 35900 40938 35952 40944
rect 35808 40656 35860 40662
rect 35808 40598 35860 40604
rect 35532 39976 35584 39982
rect 35532 39918 35584 39924
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35820 35222 35848 40598
rect 35912 36922 35940 40938
rect 36556 40730 36584 41210
rect 36544 40724 36596 40730
rect 36544 40666 36596 40672
rect 36084 39908 36136 39914
rect 36084 39850 36136 39856
rect 35992 38820 36044 38826
rect 35992 38762 36044 38768
rect 35900 36916 35952 36922
rect 35900 36858 35952 36864
rect 35808 35216 35860 35222
rect 35808 35158 35860 35164
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35900 29028 35952 29034
rect 35900 28970 35952 28976
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35716 26784 35768 26790
rect 35716 26726 35768 26732
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35728 26042 35756 26726
rect 35912 26518 35940 28970
rect 36004 26586 36032 38762
rect 36096 27130 36124 39850
rect 36544 39364 36596 39370
rect 36544 39306 36596 39312
rect 36084 27124 36136 27130
rect 36084 27066 36136 27072
rect 35992 26580 36044 26586
rect 35992 26522 36044 26528
rect 35900 26512 35952 26518
rect 35900 26454 35952 26460
rect 35912 26330 35940 26454
rect 35820 26302 35940 26330
rect 35716 26036 35768 26042
rect 35716 25978 35768 25984
rect 35440 25900 35492 25906
rect 35440 25842 35492 25848
rect 35348 25696 35400 25702
rect 35348 25638 35400 25644
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34980 25288 35032 25294
rect 34980 25230 35032 25236
rect 34992 24614 35020 25230
rect 34980 24608 35032 24614
rect 34980 24550 35032 24556
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24138 35388 25638
rect 35452 25498 35480 25842
rect 35532 25764 35584 25770
rect 35532 25706 35584 25712
rect 35440 25492 35492 25498
rect 35440 25434 35492 25440
rect 35544 24954 35572 25706
rect 35820 25430 35848 26302
rect 35808 25424 35860 25430
rect 35808 25366 35860 25372
rect 35820 25276 35848 25366
rect 35820 25248 35940 25276
rect 35716 25152 35768 25158
rect 35716 25094 35768 25100
rect 35808 25152 35860 25158
rect 35808 25094 35860 25100
rect 35532 24948 35584 24954
rect 35532 24890 35584 24896
rect 35728 24886 35756 25094
rect 35716 24880 35768 24886
rect 35716 24822 35768 24828
rect 35624 24608 35676 24614
rect 35624 24550 35676 24556
rect 35716 24608 35768 24614
rect 35716 24550 35768 24556
rect 35348 24132 35400 24138
rect 35348 24074 35400 24080
rect 34796 24064 34848 24070
rect 34796 24006 34848 24012
rect 35438 24032 35494 24041
rect 35438 23967 35494 23976
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34980 23180 35032 23186
rect 34980 23122 35032 23128
rect 34624 23072 34744 23100
rect 34244 22704 34296 22710
rect 34244 22646 34296 22652
rect 34520 22704 34572 22710
rect 34520 22646 34572 22652
rect 34152 20460 34204 20466
rect 34152 20402 34204 20408
rect 34256 20346 34284 22646
rect 34428 20460 34480 20466
rect 34428 20402 34480 20408
rect 34164 20318 34284 20346
rect 34336 20392 34388 20398
rect 34336 20334 34388 20340
rect 34060 12368 34112 12374
rect 34060 12310 34112 12316
rect 34060 10804 34112 10810
rect 34060 10746 34112 10752
rect 34072 10062 34100 10746
rect 34060 10056 34112 10062
rect 34060 9998 34112 10004
rect 34060 9920 34112 9926
rect 34060 9862 34112 9868
rect 34072 9654 34100 9862
rect 34060 9648 34112 9654
rect 34060 9590 34112 9596
rect 34060 7744 34112 7750
rect 34060 7686 34112 7692
rect 33322 3703 33324 3712
rect 32864 3674 32916 3680
rect 33376 3703 33378 3712
rect 33784 3732 33836 3738
rect 33324 3674 33376 3680
rect 33784 3674 33836 3680
rect 33968 3732 34020 3738
rect 33968 3674 34020 3680
rect 32876 3058 32904 3674
rect 33336 3058 33364 3674
rect 32864 3052 32916 3058
rect 32864 2994 32916 3000
rect 33324 3052 33376 3058
rect 33324 2994 33376 3000
rect 32956 2984 33008 2990
rect 32956 2926 33008 2932
rect 32784 2746 32904 2774
rect 32876 2446 32904 2746
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32588 2304 32640 2310
rect 32588 2246 32640 2252
rect 32600 800 32628 2246
rect 32968 800 32996 2926
rect 33692 2916 33744 2922
rect 33692 2858 33744 2864
rect 33416 2508 33468 2514
rect 33416 2450 33468 2456
rect 33428 1170 33456 2450
rect 33336 1142 33456 1170
rect 33336 800 33364 1142
rect 33704 800 33732 2858
rect 33796 2446 33824 3674
rect 34072 3534 34100 7686
rect 34164 3942 34192 20318
rect 34244 20256 34296 20262
rect 34244 20198 34296 20204
rect 34256 19446 34284 20198
rect 34348 19854 34376 20334
rect 34336 19848 34388 19854
rect 34336 19790 34388 19796
rect 34244 19440 34296 19446
rect 34244 19382 34296 19388
rect 34348 19310 34376 19790
rect 34336 19304 34388 19310
rect 34336 19246 34388 19252
rect 34348 18970 34376 19246
rect 34336 18964 34388 18970
rect 34336 18906 34388 18912
rect 34348 18290 34376 18906
rect 34336 18284 34388 18290
rect 34336 18226 34388 18232
rect 34440 18170 34468 20402
rect 34532 19334 34560 22646
rect 34624 21146 34652 23072
rect 34704 22636 34756 22642
rect 34704 22578 34756 22584
rect 34716 21894 34744 22578
rect 34992 22574 35020 23122
rect 35164 22976 35216 22982
rect 35216 22936 35296 22964
rect 35164 22918 35216 22924
rect 35268 22642 35296 22936
rect 35256 22636 35308 22642
rect 35256 22578 35308 22584
rect 34796 22568 34848 22574
rect 34796 22510 34848 22516
rect 34980 22568 35032 22574
rect 34980 22510 35032 22516
rect 34704 21888 34756 21894
rect 34704 21830 34756 21836
rect 34716 21486 34744 21830
rect 34808 21486 34836 22510
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35452 21894 35480 23967
rect 35532 23724 35584 23730
rect 35532 23666 35584 23672
rect 35544 23594 35572 23666
rect 35636 23662 35664 24550
rect 35624 23656 35676 23662
rect 35624 23598 35676 23604
rect 35532 23588 35584 23594
rect 35532 23530 35584 23536
rect 35728 23338 35756 24550
rect 35820 23866 35848 25094
rect 35912 24410 35940 25248
rect 35900 24404 35952 24410
rect 35900 24346 35952 24352
rect 35808 23860 35860 23866
rect 35808 23802 35860 23808
rect 35636 23310 35756 23338
rect 35530 22808 35586 22817
rect 35530 22743 35532 22752
rect 35584 22743 35586 22752
rect 35532 22714 35584 22720
rect 35532 22636 35584 22642
rect 35532 22578 35584 22584
rect 35544 22094 35572 22578
rect 35636 22506 35664 23310
rect 36004 23202 36032 26522
rect 35728 23174 36032 23202
rect 35728 22710 35756 23174
rect 35992 23044 36044 23050
rect 35992 22986 36044 22992
rect 35808 22976 35860 22982
rect 35808 22918 35860 22924
rect 35716 22704 35768 22710
rect 35716 22646 35768 22652
rect 35624 22500 35676 22506
rect 35624 22442 35676 22448
rect 35544 22066 35664 22094
rect 35440 21888 35492 21894
rect 35440 21830 35492 21836
rect 35452 21690 35480 21830
rect 35440 21684 35492 21690
rect 35440 21626 35492 21632
rect 34704 21480 34756 21486
rect 34704 21422 34756 21428
rect 34796 21480 34848 21486
rect 34796 21422 34848 21428
rect 34612 21140 34664 21146
rect 34612 21082 34664 21088
rect 34716 20874 34744 21422
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35348 21004 35400 21010
rect 35348 20946 35400 20952
rect 34704 20868 34756 20874
rect 34704 20810 34756 20816
rect 34612 20800 34664 20806
rect 34612 20742 34664 20748
rect 34796 20800 34848 20806
rect 34796 20742 34848 20748
rect 34624 20466 34652 20742
rect 34612 20460 34664 20466
rect 34612 20402 34664 20408
rect 34808 19718 34836 20742
rect 35360 20466 35388 20946
rect 35348 20460 35400 20466
rect 35348 20402 35400 20408
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34796 19712 34848 19718
rect 34796 19654 34848 19660
rect 34532 19306 34652 19334
rect 34520 18760 34572 18766
rect 34520 18702 34572 18708
rect 34348 18142 34468 18170
rect 34244 14340 34296 14346
rect 34244 14282 34296 14288
rect 34256 12646 34284 14282
rect 34348 12730 34376 18142
rect 34428 18080 34480 18086
rect 34428 18022 34480 18028
rect 34440 17678 34468 18022
rect 34532 17814 34560 18702
rect 34520 17808 34572 17814
rect 34520 17750 34572 17756
rect 34428 17672 34480 17678
rect 34428 17614 34480 17620
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 34426 17096 34482 17105
rect 34532 17066 34560 17614
rect 34426 17031 34482 17040
rect 34520 17060 34572 17066
rect 34440 15910 34468 17031
rect 34520 17002 34572 17008
rect 34428 15904 34480 15910
rect 34428 15846 34480 15852
rect 34520 15904 34572 15910
rect 34520 15846 34572 15852
rect 34532 15502 34560 15846
rect 34520 15496 34572 15502
rect 34520 15438 34572 15444
rect 34428 14272 34480 14278
rect 34428 14214 34480 14220
rect 34440 13938 34468 14214
rect 34428 13932 34480 13938
rect 34428 13874 34480 13880
rect 34532 13818 34560 15438
rect 34624 14498 34652 19306
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34888 18896 34940 18902
rect 34888 18838 34940 18844
rect 35348 18896 35400 18902
rect 35348 18838 35400 18844
rect 34900 18358 34928 18838
rect 34978 18456 35034 18465
rect 34978 18391 35034 18400
rect 34992 18358 35020 18391
rect 34888 18352 34940 18358
rect 34702 18320 34758 18329
rect 34888 18294 34940 18300
rect 34980 18352 35032 18358
rect 34980 18294 35032 18300
rect 34702 18255 34758 18264
rect 34716 17134 34744 18255
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17542 35388 18838
rect 34796 17536 34848 17542
rect 34796 17478 34848 17484
rect 35164 17536 35216 17542
rect 35164 17478 35216 17484
rect 35348 17536 35400 17542
rect 35348 17478 35400 17484
rect 34704 17128 34756 17134
rect 34704 17070 34756 17076
rect 34808 16590 34836 17478
rect 35176 16998 35204 17478
rect 35164 16992 35216 16998
rect 35164 16934 35216 16940
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35348 16720 35400 16726
rect 35348 16662 35400 16668
rect 34888 16652 34940 16658
rect 35164 16652 35216 16658
rect 34940 16612 35164 16640
rect 34888 16594 34940 16600
rect 35164 16594 35216 16600
rect 34796 16584 34848 16590
rect 34796 16526 34848 16532
rect 35162 16280 35218 16289
rect 35162 16215 35218 16224
rect 35176 16182 35204 16215
rect 35164 16176 35216 16182
rect 35164 16118 35216 16124
rect 34704 16040 34756 16046
rect 34704 15982 34756 15988
rect 34716 15706 34744 15982
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34704 15700 34756 15706
rect 34704 15642 34756 15648
rect 35164 15496 35216 15502
rect 35164 15438 35216 15444
rect 34796 15360 34848 15366
rect 34796 15302 34848 15308
rect 34704 14952 34756 14958
rect 34704 14894 34756 14900
rect 34716 14618 34744 14894
rect 34704 14612 34756 14618
rect 34704 14554 34756 14560
rect 34624 14470 34744 14498
rect 34612 14340 34664 14346
rect 34612 14282 34664 14288
rect 34440 13790 34560 13818
rect 34440 13258 34468 13790
rect 34428 13252 34480 13258
rect 34428 13194 34480 13200
rect 34348 12702 34560 12730
rect 34532 12646 34560 12702
rect 34244 12640 34296 12646
rect 34520 12640 34572 12646
rect 34296 12600 34376 12628
rect 34244 12582 34296 12588
rect 34244 12368 34296 12374
rect 34244 12310 34296 12316
rect 34256 7750 34284 12310
rect 34348 12209 34376 12600
rect 34520 12582 34572 12588
rect 34520 12368 34572 12374
rect 34520 12310 34572 12316
rect 34334 12200 34390 12209
rect 34334 12135 34390 12144
rect 34348 11150 34376 12135
rect 34336 11144 34388 11150
rect 34336 11086 34388 11092
rect 34532 10198 34560 12310
rect 34520 10192 34572 10198
rect 34520 10134 34572 10140
rect 34520 9988 34572 9994
rect 34520 9930 34572 9936
rect 34532 9178 34560 9930
rect 34520 9172 34572 9178
rect 34520 9114 34572 9120
rect 34428 8832 34480 8838
rect 34428 8774 34480 8780
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34440 8566 34468 8774
rect 34428 8560 34480 8566
rect 34428 8502 34480 8508
rect 34532 7954 34560 8774
rect 34520 7948 34572 7954
rect 34520 7890 34572 7896
rect 34244 7744 34296 7750
rect 34244 7686 34296 7692
rect 34624 5574 34652 14282
rect 34716 12374 34744 14470
rect 34808 12374 34836 15302
rect 35176 15026 35204 15438
rect 35360 15366 35388 16662
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 35452 15144 35480 21626
rect 35532 21548 35584 21554
rect 35532 21490 35584 21496
rect 35544 20097 35572 21490
rect 35530 20088 35586 20097
rect 35530 20023 35532 20032
rect 35584 20023 35586 20032
rect 35532 19994 35584 20000
rect 35544 19963 35572 19994
rect 35532 17740 35584 17746
rect 35532 17682 35584 17688
rect 35544 17105 35572 17682
rect 35530 17096 35586 17105
rect 35530 17031 35586 17040
rect 35532 15564 35584 15570
rect 35532 15506 35584 15512
rect 35360 15116 35480 15144
rect 35164 15020 35216 15026
rect 35164 14962 35216 14968
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14362 35388 15116
rect 35440 15020 35492 15026
rect 35440 14962 35492 14968
rect 35268 14346 35388 14362
rect 35256 14340 35388 14346
rect 35308 14334 35388 14340
rect 35256 14282 35308 14288
rect 35348 14272 35400 14278
rect 35348 14214 35400 14220
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35360 12850 35388 14214
rect 35452 13734 35480 14962
rect 35544 13802 35572 15506
rect 35532 13796 35584 13802
rect 35532 13738 35584 13744
rect 35440 13728 35492 13734
rect 35440 13670 35492 13676
rect 35532 13184 35584 13190
rect 35530 13152 35532 13161
rect 35584 13152 35586 13161
rect 35530 13087 35586 13096
rect 35348 12844 35400 12850
rect 35400 12804 35572 12832
rect 35348 12786 35400 12792
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34704 12368 34756 12374
rect 34704 12310 34756 12316
rect 34796 12368 34848 12374
rect 34796 12310 34848 12316
rect 35346 12200 35402 12209
rect 35346 12135 35348 12144
rect 35400 12135 35402 12144
rect 35348 12106 35400 12112
rect 34704 12096 34756 12102
rect 34704 12038 34756 12044
rect 34796 12096 34848 12102
rect 34796 12038 34848 12044
rect 34716 11082 34744 12038
rect 34808 11762 34836 12038
rect 34796 11756 34848 11762
rect 34796 11698 34848 11704
rect 35348 11688 35400 11694
rect 35348 11630 35400 11636
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 34704 11076 34756 11082
rect 34704 11018 34756 11024
rect 34808 10674 34836 11086
rect 34796 10668 34848 10674
rect 34796 10610 34848 10616
rect 34704 9580 34756 9586
rect 34704 9522 34756 9528
rect 34716 8634 34744 9522
rect 34808 8922 34836 10610
rect 35360 10606 35388 11630
rect 35544 10810 35572 12804
rect 35636 12434 35664 22066
rect 35716 20868 35768 20874
rect 35716 20810 35768 20816
rect 35728 19514 35756 20810
rect 35716 19508 35768 19514
rect 35716 19450 35768 19456
rect 35820 18154 35848 22918
rect 36004 22094 36032 22986
rect 36096 22642 36124 27066
rect 36556 26586 36584 39306
rect 43916 34610 43944 52974
rect 45204 52698 45232 53042
rect 45468 53032 45520 53038
rect 45468 52974 45520 52980
rect 45192 52692 45244 52698
rect 45192 52634 45244 52640
rect 45480 50386 45508 52974
rect 46032 52562 46060 55270
rect 47122 55200 47178 56000
rect 48318 55298 48374 56000
rect 49514 55298 49570 56000
rect 50710 55298 50766 56000
rect 48318 55270 48452 55298
rect 48318 55200 48374 55270
rect 47136 53242 47164 55200
rect 47124 53236 47176 53242
rect 47124 53178 47176 53184
rect 47032 53168 47084 53174
rect 47032 53110 47084 53116
rect 47044 52630 47072 53110
rect 48044 53032 48096 53038
rect 48044 52974 48096 52980
rect 47032 52624 47084 52630
rect 47032 52566 47084 52572
rect 46020 52556 46072 52562
rect 46020 52498 46072 52504
rect 46032 52154 46060 52498
rect 46296 52488 46348 52494
rect 46296 52430 46348 52436
rect 46020 52148 46072 52154
rect 46020 52090 46072 52096
rect 45468 50380 45520 50386
rect 45468 50322 45520 50328
rect 46112 40044 46164 40050
rect 46112 39986 46164 39992
rect 46124 39642 46152 39986
rect 46112 39636 46164 39642
rect 46112 39578 46164 39584
rect 46308 39506 46336 52430
rect 47032 46640 47084 46646
rect 47032 46582 47084 46588
rect 47044 44878 47072 46582
rect 47032 44872 47084 44878
rect 47032 44814 47084 44820
rect 48056 42090 48084 52974
rect 48424 52562 48452 55270
rect 49514 55270 49648 55298
rect 49514 55200 49570 55270
rect 49620 53666 49648 55270
rect 50710 55270 51028 55298
rect 50710 55200 50766 55270
rect 49620 53638 49740 53666
rect 49712 53242 49740 53638
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 51000 53258 51028 55270
rect 51906 55200 51962 56000
rect 53102 55298 53158 56000
rect 53102 55270 53236 55298
rect 53102 55200 53158 55270
rect 49700 53236 49752 53242
rect 51000 53230 51120 53258
rect 49700 53178 49752 53184
rect 51092 53174 51120 53230
rect 51080 53168 51132 53174
rect 51080 53110 51132 53116
rect 51448 53168 51500 53174
rect 51448 53110 51500 53116
rect 50160 53032 50212 53038
rect 50160 52974 50212 52980
rect 49516 52896 49568 52902
rect 49516 52838 49568 52844
rect 48412 52556 48464 52562
rect 48412 52498 48464 52504
rect 49528 51882 49556 52838
rect 49516 51876 49568 51882
rect 49516 51818 49568 51824
rect 48136 49904 48188 49910
rect 48136 49846 48188 49852
rect 48148 46374 48176 49846
rect 48228 47048 48280 47054
rect 48228 46990 48280 46996
rect 48136 46368 48188 46374
rect 48136 46310 48188 46316
rect 48240 45966 48268 46990
rect 48228 45960 48280 45966
rect 48228 45902 48280 45908
rect 48044 42084 48096 42090
rect 48044 42026 48096 42032
rect 50172 41274 50200 52974
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 51460 52154 51488 53110
rect 51920 52698 51948 55200
rect 53208 53106 53236 55270
rect 54298 55200 54354 56000
rect 53196 53100 53248 53106
rect 53196 53042 53248 53048
rect 53208 52698 53236 53042
rect 51908 52692 51960 52698
rect 51908 52634 51960 52640
rect 53196 52692 53248 52698
rect 53196 52634 53248 52640
rect 51920 52494 51948 52634
rect 51998 52592 52054 52601
rect 51998 52527 52000 52536
rect 52052 52527 52054 52536
rect 52000 52498 52052 52504
rect 51908 52488 51960 52494
rect 51908 52430 51960 52436
rect 54024 52488 54076 52494
rect 54024 52430 54076 52436
rect 51448 52148 51500 52154
rect 51448 52090 51500 52096
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 53564 50720 53616 50726
rect 53564 50662 53616 50668
rect 53932 50720 53984 50726
rect 53932 50662 53984 50668
rect 52276 50448 52328 50454
rect 52276 50390 52328 50396
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 51172 49768 51224 49774
rect 51172 49710 51224 49716
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 51184 47530 51212 49710
rect 52184 48884 52236 48890
rect 52184 48826 52236 48832
rect 51264 48544 51316 48550
rect 51264 48486 51316 48492
rect 51276 48278 51304 48486
rect 51264 48272 51316 48278
rect 51264 48214 51316 48220
rect 51276 48006 51304 48214
rect 52196 48142 52224 48826
rect 51816 48136 51868 48142
rect 51816 48078 51868 48084
rect 52184 48136 52236 48142
rect 52184 48078 52236 48084
rect 51356 48068 51408 48074
rect 51356 48010 51408 48016
rect 51264 48000 51316 48006
rect 51264 47942 51316 47948
rect 51276 47598 51304 47942
rect 51264 47592 51316 47598
rect 51264 47534 51316 47540
rect 51172 47524 51224 47530
rect 51172 47466 51224 47472
rect 50896 47048 50948 47054
rect 50894 47016 50896 47025
rect 50948 47016 50950 47025
rect 50894 46951 50950 46960
rect 51276 46918 51304 47534
rect 51368 47530 51396 48010
rect 51632 48000 51684 48006
rect 51632 47942 51684 47948
rect 51448 47660 51500 47666
rect 51448 47602 51500 47608
rect 51356 47524 51408 47530
rect 51356 47466 51408 47472
rect 51460 47161 51488 47602
rect 51540 47184 51592 47190
rect 51446 47152 51502 47161
rect 51540 47126 51592 47132
rect 51446 47087 51502 47096
rect 51552 47002 51580 47126
rect 51644 47025 51672 47942
rect 51724 47728 51776 47734
rect 51724 47670 51776 47676
rect 51736 47462 51764 47670
rect 51828 47530 51856 48078
rect 52000 48000 52052 48006
rect 52000 47942 52052 47948
rect 52012 47802 52040 47942
rect 52000 47796 52052 47802
rect 52000 47738 52052 47744
rect 52092 47796 52144 47802
rect 52092 47738 52144 47744
rect 51816 47524 51868 47530
rect 51816 47466 51868 47472
rect 51724 47456 51776 47462
rect 51724 47398 51776 47404
rect 51908 47048 51960 47054
rect 51460 46986 51580 47002
rect 51448 46980 51580 46986
rect 51500 46974 51580 46980
rect 51630 47016 51686 47025
rect 51630 46951 51686 46960
rect 51814 47016 51870 47025
rect 51908 46990 51960 46996
rect 51814 46951 51816 46960
rect 51448 46922 51500 46928
rect 51868 46951 51870 46960
rect 51816 46922 51868 46928
rect 51264 46912 51316 46918
rect 51264 46854 51316 46860
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 51080 46504 51132 46510
rect 51080 46446 51132 46452
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50160 41268 50212 41274
rect 50160 41210 50212 41216
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 46296 39500 46348 39506
rect 46296 39442 46348 39448
rect 51092 39302 51120 46446
rect 51276 46374 51304 46854
rect 51264 46368 51316 46374
rect 51264 46310 51316 46316
rect 51276 45830 51304 46310
rect 51264 45824 51316 45830
rect 51264 45766 51316 45772
rect 51172 45620 51224 45626
rect 51172 45562 51224 45568
rect 51184 41206 51212 45562
rect 51172 41200 51224 41206
rect 51172 41142 51224 41148
rect 51080 39296 51132 39302
rect 51080 39238 51132 39244
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 44180 37256 44232 37262
rect 44180 37198 44232 37204
rect 44192 35698 44220 37198
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 49608 36644 49660 36650
rect 49608 36586 49660 36592
rect 49620 36242 49648 36586
rect 49608 36236 49660 36242
rect 49608 36178 49660 36184
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 44180 35692 44232 35698
rect 44180 35634 44232 35640
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 43904 34604 43956 34610
rect 43904 34546 43956 34552
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 51276 33658 51304 45766
rect 51356 43920 51408 43926
rect 51356 43862 51408 43868
rect 51368 38010 51396 43862
rect 51920 40730 51948 46990
rect 52104 46986 52132 47738
rect 52092 46980 52144 46986
rect 52092 46922 52144 46928
rect 52196 46889 52224 48078
rect 52288 47666 52316 50390
rect 53104 50176 53156 50182
rect 53104 50118 53156 50124
rect 52920 49632 52972 49638
rect 52920 49574 52972 49580
rect 52644 49224 52696 49230
rect 52644 49166 52696 49172
rect 52368 49156 52420 49162
rect 52368 49098 52420 49104
rect 52380 48754 52408 49098
rect 52460 49088 52512 49094
rect 52460 49030 52512 49036
rect 52368 48748 52420 48754
rect 52368 48690 52420 48696
rect 52380 47977 52408 48690
rect 52366 47968 52422 47977
rect 52366 47903 52422 47912
rect 52276 47660 52328 47666
rect 52276 47602 52328 47608
rect 52472 47054 52500 49030
rect 52656 48142 52684 49166
rect 52932 48314 52960 49574
rect 53116 49230 53144 50118
rect 53576 49230 53604 50662
rect 53656 49836 53708 49842
rect 53656 49778 53708 49784
rect 53104 49224 53156 49230
rect 53104 49166 53156 49172
rect 53564 49224 53616 49230
rect 53564 49166 53616 49172
rect 52840 48286 52960 48314
rect 52840 48210 52868 48286
rect 52828 48204 52880 48210
rect 52828 48146 52880 48152
rect 52644 48136 52696 48142
rect 52644 48078 52696 48084
rect 52460 47048 52512 47054
rect 52460 46990 52512 46996
rect 52182 46880 52238 46889
rect 52182 46815 52238 46824
rect 52656 46617 52684 48078
rect 52840 47734 52868 48146
rect 53012 48000 53064 48006
rect 53012 47942 53064 47948
rect 52828 47728 52880 47734
rect 52828 47670 52880 47676
rect 52736 47524 52788 47530
rect 52736 47466 52788 47472
rect 52642 46608 52698 46617
rect 52642 46543 52698 46552
rect 52644 46028 52696 46034
rect 52644 45970 52696 45976
rect 52184 45960 52236 45966
rect 52184 45902 52236 45908
rect 52552 45960 52604 45966
rect 52552 45902 52604 45908
rect 52196 45801 52224 45902
rect 52182 45792 52238 45801
rect 52182 45727 52238 45736
rect 52458 44976 52514 44985
rect 52458 44911 52460 44920
rect 52512 44911 52514 44920
rect 52460 44882 52512 44888
rect 52184 44872 52236 44878
rect 52184 44814 52236 44820
rect 52196 44713 52224 44814
rect 52182 44704 52238 44713
rect 52182 44639 52238 44648
rect 52092 44328 52144 44334
rect 52092 44270 52144 44276
rect 52104 43450 52132 44270
rect 52564 43654 52592 45902
rect 52656 44470 52684 45970
rect 52644 44464 52696 44470
rect 52644 44406 52696 44412
rect 52748 43858 52776 47466
rect 52840 47054 52868 47670
rect 53024 47054 53052 47942
rect 53116 47705 53144 49166
rect 53470 49056 53526 49065
rect 53470 48991 53526 49000
rect 53484 48822 53512 48991
rect 53472 48816 53524 48822
rect 53576 48793 53604 49166
rect 53472 48758 53524 48764
rect 53562 48784 53618 48793
rect 53484 48686 53512 48758
rect 53562 48719 53618 48728
rect 53472 48680 53524 48686
rect 53472 48622 53524 48628
rect 53668 48521 53696 49778
rect 53654 48512 53710 48521
rect 53654 48447 53710 48456
rect 53196 48000 53248 48006
rect 53196 47942 53248 47948
rect 53840 48000 53892 48006
rect 53840 47942 53892 47948
rect 53102 47696 53158 47705
rect 53102 47631 53158 47640
rect 52828 47048 52880 47054
rect 52828 46990 52880 46996
rect 53012 47048 53064 47054
rect 53012 46990 53064 46996
rect 52920 46980 52972 46986
rect 52920 46922 52972 46928
rect 52932 45014 52960 46922
rect 53012 46368 53064 46374
rect 53010 46336 53012 46345
rect 53064 46336 53066 46345
rect 53010 46271 53066 46280
rect 53012 45280 53064 45286
rect 53010 45248 53012 45257
rect 53064 45248 53066 45257
rect 53010 45183 53066 45192
rect 52920 45008 52972 45014
rect 52920 44950 52972 44956
rect 53104 44396 53156 44402
rect 53104 44338 53156 44344
rect 53012 44192 53064 44198
rect 53010 44160 53012 44169
rect 53064 44160 53066 44169
rect 53010 44095 53066 44104
rect 52736 43852 52788 43858
rect 52736 43794 52788 43800
rect 52920 43716 52972 43722
rect 52920 43658 52972 43664
rect 52552 43648 52604 43654
rect 52552 43590 52604 43596
rect 52828 43648 52880 43654
rect 52828 43590 52880 43596
rect 52092 43444 52144 43450
rect 52092 43386 52144 43392
rect 52644 43172 52696 43178
rect 52644 43114 52696 43120
rect 52552 42900 52604 42906
rect 52552 42842 52604 42848
rect 52368 42696 52420 42702
rect 52368 42638 52420 42644
rect 52380 42566 52408 42638
rect 52368 42560 52420 42566
rect 52368 42502 52420 42508
rect 52460 42560 52512 42566
rect 52460 42502 52512 42508
rect 52276 42016 52328 42022
rect 52276 41958 52328 41964
rect 52288 41478 52316 41958
rect 52380 41721 52408 42502
rect 52366 41712 52422 41721
rect 52472 41682 52500 42502
rect 52564 42226 52592 42842
rect 52552 42220 52604 42226
rect 52552 42162 52604 42168
rect 52366 41647 52422 41656
rect 52460 41676 52512 41682
rect 52460 41618 52512 41624
rect 52368 41608 52420 41614
rect 52368 41550 52420 41556
rect 52276 41472 52328 41478
rect 52380 41449 52408 41550
rect 52276 41414 52328 41420
rect 52366 41440 52422 41449
rect 52366 41375 52422 41384
rect 51908 40724 51960 40730
rect 51908 40666 51960 40672
rect 52656 40662 52684 43114
rect 52644 40656 52696 40662
rect 52644 40598 52696 40604
rect 52368 40520 52420 40526
rect 52368 40462 52420 40468
rect 52380 40361 52408 40462
rect 52366 40352 52422 40361
rect 52366 40287 52422 40296
rect 52090 38992 52146 39001
rect 52090 38927 52092 38936
rect 52144 38927 52146 38936
rect 52092 38898 52144 38904
rect 52184 38344 52236 38350
rect 52184 38286 52236 38292
rect 52196 38185 52224 38286
rect 52182 38176 52238 38185
rect 52182 38111 52238 38120
rect 51356 38004 51408 38010
rect 51356 37946 51408 37952
rect 52368 36168 52420 36174
rect 52368 36110 52420 36116
rect 52380 35193 52408 36110
rect 52366 35184 52422 35193
rect 52366 35119 52422 35128
rect 51264 33652 51316 33658
rect 51264 33594 51316 33600
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50066 32464 50122 32473
rect 47860 32428 47912 32434
rect 50066 32399 50122 32408
rect 47860 32370 47912 32376
rect 44824 30592 44876 30598
rect 44824 30534 44876 30540
rect 37648 30048 37700 30054
rect 37648 29990 37700 29996
rect 37464 27872 37516 27878
rect 37464 27814 37516 27820
rect 37476 26586 37504 27814
rect 36176 26580 36228 26586
rect 36176 26522 36228 26528
rect 36544 26580 36596 26586
rect 36544 26522 36596 26528
rect 37464 26580 37516 26586
rect 37464 26522 37516 26528
rect 36188 22710 36216 26522
rect 36820 25152 36872 25158
rect 36820 25094 36872 25100
rect 36268 24880 36320 24886
rect 36268 24822 36320 24828
rect 36280 23905 36308 24822
rect 36832 24206 36860 25094
rect 37280 24676 37332 24682
rect 37280 24618 37332 24624
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 36820 24200 36872 24206
rect 36820 24142 36872 24148
rect 36266 23896 36322 23905
rect 36266 23831 36322 23840
rect 36176 22704 36228 22710
rect 36176 22646 36228 22652
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 36084 22500 36136 22506
rect 36084 22442 36136 22448
rect 35912 22066 36032 22094
rect 35912 21350 35940 22066
rect 36096 21690 36124 22442
rect 36372 22166 36400 24142
rect 36728 23724 36780 23730
rect 36728 23666 36780 23672
rect 36740 22778 36768 23666
rect 37292 23526 37320 24618
rect 37476 24410 37504 26522
rect 37660 25498 37688 29990
rect 39580 26852 39632 26858
rect 39580 26794 39632 26800
rect 38200 26036 38252 26042
rect 38200 25978 38252 25984
rect 37648 25492 37700 25498
rect 37648 25434 37700 25440
rect 37660 24682 37688 25434
rect 38212 25226 38240 25978
rect 39028 25696 39080 25702
rect 39028 25638 39080 25644
rect 39040 25498 39068 25638
rect 39028 25492 39080 25498
rect 39028 25434 39080 25440
rect 38384 25288 38436 25294
rect 38384 25230 38436 25236
rect 38200 25220 38252 25226
rect 38200 25162 38252 25168
rect 37832 25152 37884 25158
rect 37832 25094 37884 25100
rect 37740 24812 37792 24818
rect 37740 24754 37792 24760
rect 37648 24676 37700 24682
rect 37648 24618 37700 24624
rect 37752 24410 37780 24754
rect 37464 24404 37516 24410
rect 37464 24346 37516 24352
rect 37740 24404 37792 24410
rect 37740 24346 37792 24352
rect 37476 23866 37504 24346
rect 37844 24274 37872 25094
rect 37924 24608 37976 24614
rect 37924 24550 37976 24556
rect 37832 24268 37884 24274
rect 37832 24210 37884 24216
rect 37464 23860 37516 23866
rect 37464 23802 37516 23808
rect 37740 23792 37792 23798
rect 37740 23734 37792 23740
rect 37648 23724 37700 23730
rect 37648 23666 37700 23672
rect 37280 23520 37332 23526
rect 37280 23462 37332 23468
rect 37660 23322 37688 23666
rect 37648 23316 37700 23322
rect 37648 23258 37700 23264
rect 37752 23118 37780 23734
rect 37844 23594 37872 24210
rect 37936 23798 37964 24550
rect 37924 23792 37976 23798
rect 37924 23734 37976 23740
rect 37832 23588 37884 23594
rect 37832 23530 37884 23536
rect 37464 23112 37516 23118
rect 37464 23054 37516 23060
rect 37740 23112 37792 23118
rect 37740 23054 37792 23060
rect 37476 22778 37504 23054
rect 37752 22778 37780 23054
rect 36728 22772 36780 22778
rect 36728 22714 36780 22720
rect 37464 22772 37516 22778
rect 37464 22714 37516 22720
rect 37740 22772 37792 22778
rect 37740 22714 37792 22720
rect 36452 22636 36504 22642
rect 36452 22578 36504 22584
rect 36360 22160 36412 22166
rect 36360 22102 36412 22108
rect 36084 21684 36136 21690
rect 36084 21626 36136 21632
rect 36372 21622 36400 22102
rect 36360 21616 36412 21622
rect 36360 21558 36412 21564
rect 36176 21548 36228 21554
rect 36176 21490 36228 21496
rect 35900 21344 35952 21350
rect 35900 21286 35952 21292
rect 35900 21140 35952 21146
rect 35900 21082 35952 21088
rect 35912 21010 35940 21082
rect 35900 21004 35952 21010
rect 35900 20946 35952 20952
rect 35992 19304 36044 19310
rect 35992 19246 36044 19252
rect 36004 18970 36032 19246
rect 35992 18964 36044 18970
rect 35992 18906 36044 18912
rect 36188 18766 36216 21490
rect 36372 21010 36400 21558
rect 36360 21004 36412 21010
rect 36360 20946 36412 20952
rect 36268 19848 36320 19854
rect 36266 19816 36268 19825
rect 36320 19816 36322 19825
rect 36266 19751 36322 19760
rect 36268 19304 36320 19310
rect 36268 19246 36320 19252
rect 36280 18834 36308 19246
rect 36268 18828 36320 18834
rect 36268 18770 36320 18776
rect 36176 18760 36228 18766
rect 36176 18702 36228 18708
rect 36360 18760 36412 18766
rect 36360 18702 36412 18708
rect 36188 18290 36216 18702
rect 36176 18284 36228 18290
rect 36176 18226 36228 18232
rect 35808 18148 35860 18154
rect 35808 18090 35860 18096
rect 35820 17678 35848 18090
rect 36372 18086 36400 18702
rect 36360 18080 36412 18086
rect 36360 18022 36412 18028
rect 35808 17672 35860 17678
rect 35808 17614 35860 17620
rect 36084 17536 36136 17542
rect 36082 17504 36084 17513
rect 36136 17504 36138 17513
rect 36082 17439 36138 17448
rect 36096 17270 36124 17439
rect 36084 17264 36136 17270
rect 36464 17218 36492 22578
rect 36636 22160 36688 22166
rect 36820 22160 36872 22166
rect 36688 22120 36820 22148
rect 36636 22102 36688 22108
rect 36820 22102 36872 22108
rect 36910 22128 36966 22137
rect 36910 22063 36966 22072
rect 36924 22030 36952 22063
rect 36912 22024 36964 22030
rect 36912 21966 36964 21972
rect 37096 22024 37148 22030
rect 37096 21966 37148 21972
rect 36728 21548 36780 21554
rect 36648 21508 36728 21536
rect 36544 21344 36596 21350
rect 36544 21286 36596 21292
rect 36556 20806 36584 21286
rect 36544 20800 36596 20806
rect 36544 20742 36596 20748
rect 36648 18766 36676 21508
rect 36728 21490 36780 21496
rect 36912 21412 36964 21418
rect 36912 21354 36964 21360
rect 36728 20460 36780 20466
rect 36728 20402 36780 20408
rect 36740 19514 36768 20402
rect 36820 20324 36872 20330
rect 36820 20266 36872 20272
rect 36832 19854 36860 20266
rect 36820 19848 36872 19854
rect 36820 19790 36872 19796
rect 36728 19508 36780 19514
rect 36728 19450 36780 19456
rect 36924 18970 36952 21354
rect 37004 20936 37056 20942
rect 37004 20878 37056 20884
rect 37016 19854 37044 20878
rect 37108 20398 37136 21966
rect 37476 21894 37504 22714
rect 37844 22658 37872 23530
rect 38212 23322 38240 25162
rect 38292 24744 38344 24750
rect 38292 24686 38344 24692
rect 38304 24274 38332 24686
rect 38292 24268 38344 24274
rect 38292 24210 38344 24216
rect 38304 23730 38332 24210
rect 38396 23866 38424 25230
rect 38660 25152 38712 25158
rect 38660 25094 38712 25100
rect 38672 24818 38700 25094
rect 38660 24812 38712 24818
rect 38660 24754 38712 24760
rect 39040 24614 39068 25434
rect 38568 24608 38620 24614
rect 38568 24550 38620 24556
rect 39028 24608 39080 24614
rect 39028 24550 39080 24556
rect 38580 24426 38608 24550
rect 38580 24410 38792 24426
rect 38580 24404 38804 24410
rect 38580 24398 38752 24404
rect 38752 24346 38804 24352
rect 38752 24200 38804 24206
rect 38752 24142 38804 24148
rect 38384 23860 38436 23866
rect 38384 23802 38436 23808
rect 38292 23724 38344 23730
rect 38292 23666 38344 23672
rect 38200 23316 38252 23322
rect 38028 23276 38200 23304
rect 38028 23118 38056 23276
rect 38200 23258 38252 23264
rect 38660 23248 38712 23254
rect 38660 23190 38712 23196
rect 38016 23112 38068 23118
rect 38016 23054 38068 23060
rect 38568 23112 38620 23118
rect 38568 23054 38620 23060
rect 37752 22630 37872 22658
rect 38028 22642 38056 23054
rect 38580 22817 38608 23054
rect 38566 22808 38622 22817
rect 38566 22743 38622 22752
rect 38384 22704 38436 22710
rect 38384 22646 38436 22652
rect 38016 22636 38068 22642
rect 37556 22092 37608 22098
rect 37556 22034 37608 22040
rect 37464 21888 37516 21894
rect 37464 21830 37516 21836
rect 37372 21480 37424 21486
rect 37372 21422 37424 21428
rect 37188 20460 37240 20466
rect 37188 20402 37240 20408
rect 37096 20392 37148 20398
rect 37096 20334 37148 20340
rect 37004 19848 37056 19854
rect 37004 19790 37056 19796
rect 37108 19360 37136 20334
rect 37200 19553 37228 20402
rect 37186 19544 37242 19553
rect 37186 19479 37242 19488
rect 37280 19440 37332 19446
rect 37280 19382 37332 19388
rect 37016 19332 37136 19360
rect 36912 18964 36964 18970
rect 36912 18906 36964 18912
rect 36924 18834 36952 18906
rect 36912 18828 36964 18834
rect 36912 18770 36964 18776
rect 36636 18760 36688 18766
rect 36636 18702 36688 18708
rect 36544 18216 36596 18222
rect 36544 18158 36596 18164
rect 36084 17206 36136 17212
rect 35992 17196 36044 17202
rect 35992 17138 36044 17144
rect 36188 17190 36492 17218
rect 35900 16992 35952 16998
rect 35900 16934 35952 16940
rect 35912 16658 35940 16934
rect 35900 16652 35952 16658
rect 35900 16594 35952 16600
rect 36004 15910 36032 17138
rect 35992 15904 36044 15910
rect 35992 15846 36044 15852
rect 35716 15496 35768 15502
rect 35716 15438 35768 15444
rect 35728 12918 35756 15438
rect 35900 14340 35952 14346
rect 35900 14282 35952 14288
rect 35808 14068 35860 14074
rect 35808 14010 35860 14016
rect 35716 12912 35768 12918
rect 35716 12854 35768 12860
rect 35636 12406 35756 12434
rect 35624 11008 35676 11014
rect 35624 10950 35676 10956
rect 35532 10804 35584 10810
rect 35532 10746 35584 10752
rect 35348 10600 35400 10606
rect 35348 10542 35400 10548
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35256 10192 35308 10198
rect 35256 10134 35308 10140
rect 34980 10056 35032 10062
rect 34978 10024 34980 10033
rect 35032 10024 35034 10033
rect 34978 9959 35034 9968
rect 35268 9330 35296 10134
rect 35360 9654 35388 10542
rect 35636 10062 35664 10950
rect 35624 10056 35676 10062
rect 35624 9998 35676 10004
rect 35532 9988 35584 9994
rect 35532 9930 35584 9936
rect 35440 9920 35492 9926
rect 35440 9862 35492 9868
rect 35348 9648 35400 9654
rect 35348 9590 35400 9596
rect 35268 9302 35388 9330
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34808 8894 35020 8922
rect 34704 8628 34756 8634
rect 34704 8570 34756 8576
rect 34808 8362 34836 8894
rect 34992 8838 35020 8894
rect 34980 8832 35032 8838
rect 34980 8774 35032 8780
rect 34796 8356 34848 8362
rect 34796 8298 34848 8304
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34612 5568 34664 5574
rect 34612 5510 34664 5516
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34518 4040 34574 4049
rect 34518 3975 34574 3984
rect 34152 3936 34204 3942
rect 34152 3878 34204 3884
rect 34532 3738 34560 3975
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34520 3732 34572 3738
rect 34520 3674 34572 3680
rect 34060 3528 34112 3534
rect 34060 3470 34112 3476
rect 34428 3120 34480 3126
rect 34428 3062 34480 3068
rect 33784 2440 33836 2446
rect 34152 2440 34204 2446
rect 33784 2382 33836 2388
rect 34072 2400 34152 2428
rect 34072 800 34100 2400
rect 34152 2382 34204 2388
rect 34440 800 34468 3062
rect 34532 2378 34560 3674
rect 35360 3670 35388 9302
rect 35452 8498 35480 9862
rect 35544 9722 35572 9930
rect 35532 9716 35584 9722
rect 35532 9658 35584 9664
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 35544 8090 35572 9658
rect 35624 9104 35676 9110
rect 35624 9046 35676 9052
rect 35636 8294 35664 9046
rect 35624 8288 35676 8294
rect 35624 8230 35676 8236
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35728 4282 35756 12406
rect 35820 11150 35848 14010
rect 35912 11898 35940 14282
rect 35992 13728 36044 13734
rect 35992 13670 36044 13676
rect 36004 13258 36032 13670
rect 35992 13252 36044 13258
rect 35992 13194 36044 13200
rect 35900 11892 35952 11898
rect 35900 11834 35952 11840
rect 35992 11756 36044 11762
rect 35992 11698 36044 11704
rect 36004 11354 36032 11698
rect 35992 11348 36044 11354
rect 35992 11290 36044 11296
rect 36084 11280 36136 11286
rect 36084 11222 36136 11228
rect 35808 11144 35860 11150
rect 36096 11121 36124 11222
rect 35808 11086 35860 11092
rect 36082 11112 36138 11121
rect 36082 11047 36138 11056
rect 35808 10668 35860 10674
rect 35808 10610 35860 10616
rect 35820 9178 35848 10610
rect 35992 9376 36044 9382
rect 35992 9318 36044 9324
rect 35808 9172 35860 9178
rect 35808 9114 35860 9120
rect 35900 9104 35952 9110
rect 35900 9046 35952 9052
rect 35912 8673 35940 9046
rect 35898 8664 35954 8673
rect 35898 8599 35954 8608
rect 36004 8566 36032 9318
rect 35992 8560 36044 8566
rect 35992 8502 36044 8508
rect 35900 8288 35952 8294
rect 35900 8230 35952 8236
rect 35912 8090 35940 8230
rect 35900 8084 35952 8090
rect 35900 8026 35952 8032
rect 35912 7546 35940 8026
rect 35900 7540 35952 7546
rect 35900 7482 35952 7488
rect 35716 4276 35768 4282
rect 35716 4218 35768 4224
rect 36188 4214 36216 17190
rect 36452 16788 36504 16794
rect 36556 16776 36584 18158
rect 36820 18148 36872 18154
rect 36820 18090 36872 18096
rect 36636 17536 36688 17542
rect 36636 17478 36688 17484
rect 36504 16748 36584 16776
rect 36452 16730 36504 16736
rect 36648 16658 36676 17478
rect 36832 17134 36860 18090
rect 37016 17898 37044 19332
rect 37096 19236 37148 19242
rect 37096 19178 37148 19184
rect 37108 18970 37136 19178
rect 37096 18964 37148 18970
rect 37096 18906 37148 18912
rect 36924 17870 37044 17898
rect 36924 17338 36952 17870
rect 37004 17808 37056 17814
rect 37292 17796 37320 19382
rect 37384 19310 37412 21422
rect 37476 21350 37504 21830
rect 37464 21344 37516 21350
rect 37464 21286 37516 21292
rect 37476 20602 37504 21286
rect 37568 21146 37596 22034
rect 37646 21448 37702 21457
rect 37646 21383 37702 21392
rect 37660 21350 37688 21383
rect 37648 21344 37700 21350
rect 37648 21286 37700 21292
rect 37556 21140 37608 21146
rect 37556 21082 37608 21088
rect 37464 20596 37516 20602
rect 37464 20538 37516 20544
rect 37462 20088 37518 20097
rect 37462 20023 37518 20032
rect 37476 19990 37504 20023
rect 37464 19984 37516 19990
rect 37464 19926 37516 19932
rect 37372 19304 37424 19310
rect 37568 19281 37596 21082
rect 37372 19246 37424 19252
rect 37554 19272 37610 19281
rect 37554 19207 37610 19216
rect 37056 17768 37320 17796
rect 37004 17750 37056 17756
rect 37464 17672 37516 17678
rect 37568 17660 37596 19207
rect 37648 18284 37700 18290
rect 37648 18226 37700 18232
rect 37516 17632 37596 17660
rect 37464 17614 37516 17620
rect 36912 17332 36964 17338
rect 36912 17274 36964 17280
rect 37556 17332 37608 17338
rect 37556 17274 37608 17280
rect 36820 17128 36872 17134
rect 36820 17070 36872 17076
rect 36924 16998 36952 17274
rect 37280 17128 37332 17134
rect 37280 17070 37332 17076
rect 36912 16992 36964 16998
rect 36964 16940 37044 16946
rect 36912 16934 37044 16940
rect 36924 16918 37044 16934
rect 36636 16652 36688 16658
rect 36636 16594 36688 16600
rect 36360 16584 36412 16590
rect 36360 16526 36412 16532
rect 36372 16250 36400 16526
rect 36544 16516 36596 16522
rect 36544 16458 36596 16464
rect 36360 16244 36412 16250
rect 36360 16186 36412 16192
rect 36452 16176 36504 16182
rect 36452 16118 36504 16124
rect 36464 15502 36492 16118
rect 36556 15638 36584 16458
rect 36912 16108 36964 16114
rect 36912 16050 36964 16056
rect 36924 16017 36952 16050
rect 36910 16008 36966 16017
rect 36910 15943 36966 15952
rect 36544 15632 36596 15638
rect 36544 15574 36596 15580
rect 36452 15496 36504 15502
rect 36452 15438 36504 15444
rect 36268 14408 36320 14414
rect 36268 14350 36320 14356
rect 36280 13938 36308 14350
rect 36268 13932 36320 13938
rect 36268 13874 36320 13880
rect 36280 13394 36308 13874
rect 36544 13864 36596 13870
rect 36544 13806 36596 13812
rect 36360 13796 36412 13802
rect 36360 13738 36412 13744
rect 36268 13388 36320 13394
rect 36268 13330 36320 13336
rect 36372 12850 36400 13738
rect 36556 12986 36584 13806
rect 36726 13152 36782 13161
rect 36726 13087 36782 13096
rect 36544 12980 36596 12986
rect 36544 12922 36596 12928
rect 36360 12844 36412 12850
rect 36360 12786 36412 12792
rect 36268 12776 36320 12782
rect 36268 12718 36320 12724
rect 36280 10266 36308 12718
rect 36372 12442 36400 12786
rect 36360 12436 36412 12442
rect 36360 12378 36412 12384
rect 36740 12238 36768 13087
rect 37016 12238 37044 16918
rect 37292 16590 37320 17070
rect 37464 16788 37516 16794
rect 37464 16730 37516 16736
rect 37476 16590 37504 16730
rect 37280 16584 37332 16590
rect 37280 16526 37332 16532
rect 37464 16584 37516 16590
rect 37464 16526 37516 16532
rect 37372 16516 37424 16522
rect 37372 16458 37424 16464
rect 37280 16244 37332 16250
rect 37280 16186 37332 16192
rect 37292 15065 37320 16186
rect 37278 15056 37334 15065
rect 37278 14991 37334 15000
rect 37096 14816 37148 14822
rect 37096 14758 37148 14764
rect 37108 14414 37136 14758
rect 37096 14408 37148 14414
rect 37096 14350 37148 14356
rect 37108 13326 37136 14350
rect 37384 14278 37412 16458
rect 37464 15904 37516 15910
rect 37464 15846 37516 15852
rect 37476 15434 37504 15846
rect 37568 15706 37596 17274
rect 37660 16522 37688 18226
rect 37648 16516 37700 16522
rect 37648 16458 37700 16464
rect 37556 15700 37608 15706
rect 37556 15642 37608 15648
rect 37464 15428 37516 15434
rect 37464 15370 37516 15376
rect 37462 14920 37518 14929
rect 37462 14855 37464 14864
rect 37516 14855 37518 14864
rect 37464 14826 37516 14832
rect 37476 14414 37504 14826
rect 37464 14408 37516 14414
rect 37464 14350 37516 14356
rect 37372 14272 37424 14278
rect 37372 14214 37424 14220
rect 37280 13524 37332 13530
rect 37280 13466 37332 13472
rect 37096 13320 37148 13326
rect 37096 13262 37148 13268
rect 37108 12306 37136 13262
rect 37292 12434 37320 13466
rect 37384 13394 37412 14214
rect 37556 13728 37608 13734
rect 37556 13670 37608 13676
rect 37372 13388 37424 13394
rect 37372 13330 37424 13336
rect 37384 13190 37412 13330
rect 37568 13326 37596 13670
rect 37752 13530 37780 22630
rect 38016 22578 38068 22584
rect 38200 20868 38252 20874
rect 38200 20810 38252 20816
rect 37832 19984 37884 19990
rect 37832 19926 37884 19932
rect 38106 19952 38162 19961
rect 37844 19514 37872 19926
rect 38106 19887 38162 19896
rect 38120 19718 38148 19887
rect 38108 19712 38160 19718
rect 38108 19654 38160 19660
rect 38120 19514 38148 19654
rect 37832 19508 37884 19514
rect 37832 19450 37884 19456
rect 38108 19508 38160 19514
rect 38108 19450 38160 19456
rect 37844 18834 37872 19450
rect 37832 18828 37884 18834
rect 37832 18770 37884 18776
rect 38108 18624 38160 18630
rect 38108 18566 38160 18572
rect 37832 18420 37884 18426
rect 37832 18362 37884 18368
rect 37844 18086 37872 18362
rect 38120 18329 38148 18566
rect 38106 18320 38162 18329
rect 38106 18255 38162 18264
rect 38108 18216 38160 18222
rect 38108 18158 38160 18164
rect 38120 18086 38148 18158
rect 37832 18080 37884 18086
rect 37832 18022 37884 18028
rect 38108 18080 38160 18086
rect 38108 18022 38160 18028
rect 37844 17785 37872 18022
rect 38016 17808 38068 17814
rect 37830 17776 37886 17785
rect 38016 17750 38068 17756
rect 37830 17711 37886 17720
rect 37924 17672 37976 17678
rect 37924 17614 37976 17620
rect 37936 17513 37964 17614
rect 37922 17504 37978 17513
rect 37922 17439 37978 17448
rect 37832 16652 37884 16658
rect 37832 16594 37884 16600
rect 37844 16153 37872 16594
rect 37830 16144 37886 16153
rect 37830 16079 37886 16088
rect 37936 15706 37964 17439
rect 38028 16794 38056 17750
rect 38108 17740 38160 17746
rect 38108 17682 38160 17688
rect 38016 16788 38068 16794
rect 38016 16730 38068 16736
rect 38120 16522 38148 17682
rect 38108 16516 38160 16522
rect 38108 16458 38160 16464
rect 38120 15978 38148 16458
rect 38212 16182 38240 20810
rect 38292 19304 38344 19310
rect 38290 19272 38292 19281
rect 38344 19272 38346 19281
rect 38290 19207 38346 19216
rect 38292 18760 38344 18766
rect 38290 18728 38292 18737
rect 38344 18728 38346 18737
rect 38290 18663 38346 18672
rect 38292 18624 38344 18630
rect 38292 18566 38344 18572
rect 38304 18426 38332 18566
rect 38292 18420 38344 18426
rect 38292 18362 38344 18368
rect 38290 18184 38346 18193
rect 38290 18119 38346 18128
rect 38304 18086 38332 18119
rect 38292 18080 38344 18086
rect 38292 18022 38344 18028
rect 38304 16794 38332 18022
rect 38292 16788 38344 16794
rect 38292 16730 38344 16736
rect 38200 16176 38252 16182
rect 38200 16118 38252 16124
rect 38396 16130 38424 22646
rect 38672 22642 38700 23190
rect 38764 22778 38792 24142
rect 38936 23520 38988 23526
rect 38936 23462 38988 23468
rect 38752 22772 38804 22778
rect 38752 22714 38804 22720
rect 38660 22636 38712 22642
rect 38660 22578 38712 22584
rect 38948 22574 38976 23462
rect 39040 22982 39068 24550
rect 39304 24064 39356 24070
rect 39304 24006 39356 24012
rect 39316 23866 39344 24006
rect 39304 23860 39356 23866
rect 39304 23802 39356 23808
rect 39028 22976 39080 22982
rect 39028 22918 39080 22924
rect 39212 22636 39264 22642
rect 39212 22578 39264 22584
rect 38936 22568 38988 22574
rect 38936 22510 38988 22516
rect 38658 22264 38714 22273
rect 38658 22199 38714 22208
rect 38672 22166 38700 22199
rect 38660 22160 38712 22166
rect 38660 22102 38712 22108
rect 38752 22160 38804 22166
rect 38752 22102 38804 22108
rect 38614 22024 38666 22030
rect 38764 21978 38792 22102
rect 39028 22024 39080 22030
rect 38666 21972 38792 21978
rect 38614 21966 38792 21972
rect 38626 21950 38792 21966
rect 38856 21984 39028 22012
rect 38660 21888 38712 21894
rect 38856 21842 38884 21984
rect 39028 21966 39080 21972
rect 38712 21836 38884 21842
rect 38660 21830 38884 21836
rect 38672 21814 38884 21830
rect 39224 21690 39252 22578
rect 39212 21684 39264 21690
rect 39212 21626 39264 21632
rect 38568 21548 38620 21554
rect 38568 21490 38620 21496
rect 38844 21548 38896 21554
rect 38844 21490 38896 21496
rect 38580 21146 38608 21490
rect 38568 21140 38620 21146
rect 38568 21082 38620 21088
rect 38750 20904 38806 20913
rect 38750 20839 38752 20848
rect 38804 20839 38806 20848
rect 38752 20810 38804 20816
rect 38752 20392 38804 20398
rect 38752 20334 38804 20340
rect 38474 19816 38530 19825
rect 38474 19751 38530 19760
rect 38488 18306 38516 19751
rect 38764 19514 38792 20334
rect 38856 19922 38884 21490
rect 39120 21480 39172 21486
rect 39120 21422 39172 21428
rect 39132 20874 39160 21422
rect 39224 20890 39252 21626
rect 39304 20912 39356 20918
rect 39120 20868 39172 20874
rect 39120 20810 39172 20816
rect 39224 20862 39304 20890
rect 38936 20392 38988 20398
rect 38936 20334 38988 20340
rect 38844 19916 38896 19922
rect 38844 19858 38896 19864
rect 38752 19508 38804 19514
rect 38752 19450 38804 19456
rect 38660 19168 38712 19174
rect 38660 19110 38712 19116
rect 38672 18834 38700 19110
rect 38660 18828 38712 18834
rect 38660 18770 38712 18776
rect 38844 18760 38896 18766
rect 38844 18702 38896 18708
rect 38660 18692 38712 18698
rect 38712 18652 38792 18680
rect 38660 18634 38712 18640
rect 38566 18320 38622 18329
rect 38488 18278 38566 18306
rect 38566 18255 38622 18264
rect 38476 18148 38528 18154
rect 38476 18090 38528 18096
rect 38488 17610 38516 18090
rect 38476 17604 38528 17610
rect 38476 17546 38528 17552
rect 38580 17338 38608 18255
rect 38660 17672 38712 17678
rect 38764 17660 38792 18652
rect 38856 17762 38884 18702
rect 38948 18290 38976 20334
rect 39224 19242 39252 20862
rect 39304 20854 39356 20860
rect 39304 20800 39356 20806
rect 39304 20742 39356 20748
rect 39316 19378 39344 20742
rect 39396 20324 39448 20330
rect 39396 20266 39448 20272
rect 39408 20058 39436 20266
rect 39488 20256 39540 20262
rect 39488 20198 39540 20204
rect 39396 20052 39448 20058
rect 39396 19994 39448 20000
rect 39500 19854 39528 20198
rect 39488 19848 39540 19854
rect 39488 19790 39540 19796
rect 39304 19372 39356 19378
rect 39304 19314 39356 19320
rect 39212 19236 39264 19242
rect 39212 19178 39264 19184
rect 39224 18766 39252 19178
rect 39304 18896 39356 18902
rect 39304 18838 39356 18844
rect 39316 18766 39344 18838
rect 39212 18760 39264 18766
rect 39212 18702 39264 18708
rect 39304 18760 39356 18766
rect 39304 18702 39356 18708
rect 38936 18284 38988 18290
rect 38936 18226 38988 18232
rect 38856 17734 39068 17762
rect 38844 17672 38896 17678
rect 38764 17632 38844 17660
rect 38660 17614 38712 17620
rect 38844 17614 38896 17620
rect 38672 17354 38700 17614
rect 38568 17332 38620 17338
rect 38672 17326 38792 17354
rect 38568 17274 38620 17280
rect 38660 17264 38712 17270
rect 38660 17206 38712 17212
rect 38672 16590 38700 17206
rect 38660 16584 38712 16590
rect 38660 16526 38712 16532
rect 38764 16454 38792 17326
rect 38856 17218 38884 17614
rect 38936 17604 38988 17610
rect 38936 17546 38988 17552
rect 38948 17338 38976 17546
rect 39040 17542 39068 17734
rect 39224 17660 39252 18702
rect 39304 18216 39356 18222
rect 39302 18184 39304 18193
rect 39356 18184 39358 18193
rect 39302 18119 39358 18128
rect 39304 17672 39356 17678
rect 39224 17632 39304 17660
rect 39304 17614 39356 17620
rect 39316 17542 39344 17614
rect 39028 17536 39080 17542
rect 39028 17478 39080 17484
rect 39120 17536 39172 17542
rect 39120 17478 39172 17484
rect 39304 17536 39356 17542
rect 39304 17478 39356 17484
rect 38936 17332 38988 17338
rect 38936 17274 38988 17280
rect 39040 17270 39068 17301
rect 39028 17264 39080 17270
rect 38856 17212 39028 17218
rect 38856 17206 39080 17212
rect 38856 17190 39068 17206
rect 39132 17202 39160 17478
rect 39040 16522 39068 17190
rect 39120 17196 39172 17202
rect 39120 17138 39172 17144
rect 39212 17128 39264 17134
rect 39212 17070 39264 17076
rect 39028 16516 39080 16522
rect 39028 16458 39080 16464
rect 38752 16448 38804 16454
rect 38752 16390 38804 16396
rect 38396 16114 38608 16130
rect 38396 16108 38620 16114
rect 38396 16102 38568 16108
rect 38108 15972 38160 15978
rect 38108 15914 38160 15920
rect 37924 15700 37976 15706
rect 37924 15642 37976 15648
rect 37936 15076 37964 15642
rect 38016 15088 38068 15094
rect 37936 15048 38016 15076
rect 38016 15030 38068 15036
rect 37832 15020 37884 15026
rect 37832 14962 37884 14968
rect 37844 14550 37872 14962
rect 37832 14544 37884 14550
rect 37832 14486 37884 14492
rect 37740 13524 37792 13530
rect 37740 13466 37792 13472
rect 37832 13388 37884 13394
rect 37832 13330 37884 13336
rect 37556 13320 37608 13326
rect 37556 13262 37608 13268
rect 37372 13184 37424 13190
rect 37372 13126 37424 13132
rect 37740 12912 37792 12918
rect 37740 12854 37792 12860
rect 37648 12640 37700 12646
rect 37648 12582 37700 12588
rect 37556 12436 37608 12442
rect 37292 12406 37504 12434
rect 37096 12300 37148 12306
rect 37096 12242 37148 12248
rect 36544 12232 36596 12238
rect 36544 12174 36596 12180
rect 36728 12232 36780 12238
rect 36728 12174 36780 12180
rect 36912 12232 36964 12238
rect 36912 12174 36964 12180
rect 37004 12232 37056 12238
rect 37004 12174 37056 12180
rect 36452 11280 36504 11286
rect 36450 11248 36452 11257
rect 36504 11248 36506 11257
rect 36450 11183 36506 11192
rect 36452 11008 36504 11014
rect 36452 10950 36504 10956
rect 36464 10674 36492 10950
rect 36360 10668 36412 10674
rect 36360 10610 36412 10616
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36372 10470 36400 10610
rect 36360 10464 36412 10470
rect 36360 10406 36412 10412
rect 36268 10260 36320 10266
rect 36268 10202 36320 10208
rect 36556 9654 36584 12174
rect 36636 12096 36688 12102
rect 36636 12038 36688 12044
rect 36924 12050 36952 12174
rect 37188 12164 37240 12170
rect 37188 12106 37240 12112
rect 36648 11150 36676 12038
rect 36924 12022 37044 12050
rect 36820 11756 36872 11762
rect 36820 11698 36872 11704
rect 36636 11144 36688 11150
rect 36636 11086 36688 11092
rect 36832 10033 36860 11698
rect 37016 11082 37044 12022
rect 37200 11150 37228 12106
rect 37372 12096 37424 12102
rect 37292 12056 37372 12084
rect 37292 11354 37320 12056
rect 37372 12038 37424 12044
rect 37280 11348 37332 11354
rect 37280 11290 37332 11296
rect 37372 11348 37424 11354
rect 37372 11290 37424 11296
rect 37384 11218 37412 11290
rect 37372 11212 37424 11218
rect 37372 11154 37424 11160
rect 37188 11144 37240 11150
rect 37188 11086 37240 11092
rect 37004 11076 37056 11082
rect 37004 11018 37056 11024
rect 36912 10464 36964 10470
rect 36912 10406 36964 10412
rect 36818 10024 36874 10033
rect 36924 9994 36952 10406
rect 36818 9959 36874 9968
rect 36912 9988 36964 9994
rect 36544 9648 36596 9654
rect 36544 9590 36596 9596
rect 36728 8968 36780 8974
rect 36726 8936 36728 8945
rect 36780 8936 36782 8945
rect 36726 8871 36782 8880
rect 36740 8838 36768 8871
rect 36636 8832 36688 8838
rect 36636 8774 36688 8780
rect 36728 8832 36780 8838
rect 36728 8774 36780 8780
rect 36648 8566 36676 8774
rect 36832 8634 36860 9959
rect 36912 9930 36964 9936
rect 37016 9382 37044 11018
rect 37200 10713 37228 11086
rect 37372 11076 37424 11082
rect 37372 11018 37424 11024
rect 37186 10704 37242 10713
rect 37186 10639 37242 10648
rect 37384 9450 37412 11018
rect 37372 9444 37424 9450
rect 37372 9386 37424 9392
rect 37004 9376 37056 9382
rect 37004 9318 37056 9324
rect 36820 8628 36872 8634
rect 36820 8570 36872 8576
rect 36636 8560 36688 8566
rect 36636 8502 36688 8508
rect 36648 8090 36676 8502
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 37476 7954 37504 12406
rect 37556 12378 37608 12384
rect 37568 10810 37596 12378
rect 37660 12102 37688 12582
rect 37752 12442 37780 12854
rect 37740 12436 37792 12442
rect 37740 12378 37792 12384
rect 37738 12336 37794 12345
rect 37738 12271 37740 12280
rect 37792 12271 37794 12280
rect 37740 12242 37792 12248
rect 37648 12096 37700 12102
rect 37648 12038 37700 12044
rect 37752 11898 37780 12242
rect 37740 11892 37792 11898
rect 37740 11834 37792 11840
rect 37648 11756 37700 11762
rect 37648 11698 37700 11704
rect 37660 11558 37688 11698
rect 37648 11552 37700 11558
rect 37648 11494 37700 11500
rect 37844 11354 37872 13330
rect 38120 13326 38148 15914
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38292 15904 38344 15910
rect 38292 15846 38344 15852
rect 38212 15026 38240 15846
rect 38304 15337 38332 15846
rect 38396 15638 38424 16102
rect 38568 16050 38620 16056
rect 39040 15638 39068 16458
rect 38384 15632 38436 15638
rect 38384 15574 38436 15580
rect 39028 15632 39080 15638
rect 39028 15574 39080 15580
rect 38290 15328 38346 15337
rect 38290 15263 38346 15272
rect 38200 15020 38252 15026
rect 38200 14962 38252 14968
rect 38212 14396 38240 14962
rect 38292 14408 38344 14414
rect 38212 14368 38292 14396
rect 38292 14350 38344 14356
rect 38200 13932 38252 13938
rect 38200 13874 38252 13880
rect 38212 13705 38240 13874
rect 38198 13696 38254 13705
rect 38198 13631 38254 13640
rect 38108 13320 38160 13326
rect 38108 13262 38160 13268
rect 38200 12776 38252 12782
rect 38200 12718 38252 12724
rect 38212 11762 38240 12718
rect 38304 12306 38332 14350
rect 38396 14278 38424 15574
rect 38844 15360 38896 15366
rect 38844 15302 38896 15308
rect 38476 15088 38528 15094
rect 38528 15048 38608 15076
rect 38476 15030 38528 15036
rect 38384 14272 38436 14278
rect 38384 14214 38436 14220
rect 38580 13920 38608 15048
rect 38750 14376 38806 14385
rect 38750 14311 38752 14320
rect 38804 14311 38806 14320
rect 38752 14282 38804 14288
rect 38750 14104 38806 14113
rect 38750 14039 38806 14048
rect 38764 13954 38792 14039
rect 38672 13926 38792 13954
rect 38672 13920 38700 13926
rect 38580 13892 38700 13920
rect 38476 13524 38528 13530
rect 38476 13466 38528 13472
rect 38488 13326 38516 13466
rect 38476 13320 38528 13326
rect 38476 13262 38528 13268
rect 38856 12986 38884 15302
rect 39120 14816 39172 14822
rect 39120 14758 39172 14764
rect 38936 14544 38988 14550
rect 38936 14486 38988 14492
rect 38948 13938 38976 14486
rect 39028 14476 39080 14482
rect 39028 14418 39080 14424
rect 38936 13932 38988 13938
rect 38936 13874 38988 13880
rect 39040 13433 39068 14418
rect 39132 14278 39160 14758
rect 39224 14550 39252 17070
rect 39316 16590 39344 17478
rect 39394 16824 39450 16833
rect 39394 16759 39396 16768
rect 39448 16759 39450 16768
rect 39396 16730 39448 16736
rect 39304 16584 39356 16590
rect 39304 16526 39356 16532
rect 39316 15502 39344 16526
rect 39304 15496 39356 15502
rect 39304 15438 39356 15444
rect 39394 15464 39450 15473
rect 39394 15399 39450 15408
rect 39408 15366 39436 15399
rect 39396 15360 39448 15366
rect 39396 15302 39448 15308
rect 39488 15020 39540 15026
rect 39488 14962 39540 14968
rect 39304 14816 39356 14822
rect 39304 14758 39356 14764
rect 39396 14816 39448 14822
rect 39396 14758 39448 14764
rect 39316 14550 39344 14758
rect 39212 14544 39264 14550
rect 39212 14486 39264 14492
rect 39304 14544 39356 14550
rect 39304 14486 39356 14492
rect 39224 14396 39252 14486
rect 39408 14396 39436 14758
rect 39224 14368 39436 14396
rect 39120 14272 39172 14278
rect 39120 14214 39172 14220
rect 39118 14104 39174 14113
rect 39118 14039 39174 14048
rect 39132 13870 39160 14039
rect 39120 13864 39172 13870
rect 39120 13806 39172 13812
rect 39026 13424 39082 13433
rect 38948 13382 39026 13410
rect 38844 12980 38896 12986
rect 38844 12922 38896 12928
rect 38384 12844 38436 12850
rect 38384 12786 38436 12792
rect 38396 12442 38424 12786
rect 38384 12436 38436 12442
rect 38384 12378 38436 12384
rect 38856 12374 38884 12922
rect 38844 12368 38896 12374
rect 38844 12310 38896 12316
rect 38292 12300 38344 12306
rect 38292 12242 38344 12248
rect 38476 12232 38528 12238
rect 38476 12174 38528 12180
rect 38200 11756 38252 11762
rect 38200 11698 38252 11704
rect 37832 11348 37884 11354
rect 37832 11290 37884 11296
rect 37844 11150 37872 11290
rect 37832 11144 37884 11150
rect 37832 11086 37884 11092
rect 38108 11076 38160 11082
rect 38108 11018 38160 11024
rect 37556 10804 37608 10810
rect 37556 10746 37608 10752
rect 37740 10804 37792 10810
rect 37740 10746 37792 10752
rect 37752 10674 37780 10746
rect 37740 10668 37792 10674
rect 37740 10610 37792 10616
rect 37924 10600 37976 10606
rect 37924 10542 37976 10548
rect 37936 9926 37964 10542
rect 37924 9920 37976 9926
rect 37924 9862 37976 9868
rect 38016 9920 38068 9926
rect 38016 9862 38068 9868
rect 37556 9580 37608 9586
rect 37556 9522 37608 9528
rect 37568 8362 37596 9522
rect 37648 9376 37700 9382
rect 37648 9318 37700 9324
rect 37660 8430 37688 9318
rect 37936 9042 37964 9862
rect 38028 9722 38056 9862
rect 38016 9716 38068 9722
rect 38016 9658 38068 9664
rect 38120 9586 38148 11018
rect 38212 10606 38240 11698
rect 38384 11620 38436 11626
rect 38384 11562 38436 11568
rect 38396 11354 38424 11562
rect 38384 11348 38436 11354
rect 38384 11290 38436 11296
rect 38384 11144 38436 11150
rect 38488 11132 38516 12174
rect 38436 11104 38516 11132
rect 38568 11144 38620 11150
rect 38384 11086 38436 11092
rect 38568 11086 38620 11092
rect 38660 11144 38712 11150
rect 38660 11086 38712 11092
rect 38200 10600 38252 10606
rect 38200 10542 38252 10548
rect 38212 10062 38240 10542
rect 38396 10470 38424 11086
rect 38580 10849 38608 11086
rect 38566 10840 38622 10849
rect 38566 10775 38622 10784
rect 38476 10668 38528 10674
rect 38476 10610 38528 10616
rect 38384 10464 38436 10470
rect 38384 10406 38436 10412
rect 38396 10062 38424 10406
rect 38488 10266 38516 10610
rect 38476 10260 38528 10266
rect 38476 10202 38528 10208
rect 38200 10056 38252 10062
rect 38200 9998 38252 10004
rect 38384 10056 38436 10062
rect 38384 9998 38436 10004
rect 38212 9674 38240 9998
rect 38292 9716 38344 9722
rect 38212 9664 38292 9674
rect 38212 9658 38344 9664
rect 38212 9646 38332 9658
rect 38108 9580 38160 9586
rect 38108 9522 38160 9528
rect 37924 9036 37976 9042
rect 37924 8978 37976 8984
rect 38304 8634 38332 9646
rect 38672 9178 38700 11086
rect 38948 10810 38976 13382
rect 39026 13359 39082 13368
rect 39028 13184 39080 13190
rect 39028 13126 39080 13132
rect 39040 12306 39068 13126
rect 39028 12300 39080 12306
rect 39028 12242 39080 12248
rect 39132 11830 39160 13806
rect 39316 12238 39344 14368
rect 39500 13734 39528 14962
rect 39488 13728 39540 13734
rect 39488 13670 39540 13676
rect 39500 13394 39528 13670
rect 39488 13388 39540 13394
rect 39488 13330 39540 13336
rect 39396 13320 39448 13326
rect 39396 13262 39448 13268
rect 39408 12714 39436 13262
rect 39396 12708 39448 12714
rect 39396 12650 39448 12656
rect 39592 12434 39620 26794
rect 42616 26580 42668 26586
rect 42616 26522 42668 26528
rect 42432 26376 42484 26382
rect 42432 26318 42484 26324
rect 40132 25424 40184 25430
rect 40132 25366 40184 25372
rect 39764 25288 39816 25294
rect 39764 25230 39816 25236
rect 39776 22710 39804 25230
rect 40040 24268 40092 24274
rect 40040 24210 40092 24216
rect 40052 23730 40080 24210
rect 40144 24206 40172 25366
rect 41420 25288 41472 25294
rect 41420 25230 41472 25236
rect 40408 24812 40460 24818
rect 40408 24754 40460 24760
rect 40316 24404 40368 24410
rect 40316 24346 40368 24352
rect 40132 24200 40184 24206
rect 40132 24142 40184 24148
rect 40132 24064 40184 24070
rect 40132 24006 40184 24012
rect 40144 23798 40172 24006
rect 40328 23866 40356 24346
rect 40316 23860 40368 23866
rect 40316 23802 40368 23808
rect 40132 23792 40184 23798
rect 40132 23734 40184 23740
rect 40040 23724 40092 23730
rect 40040 23666 40092 23672
rect 40144 23186 40172 23734
rect 40316 23520 40368 23526
rect 40316 23462 40368 23468
rect 40132 23180 40184 23186
rect 40132 23122 40184 23128
rect 39948 22976 40000 22982
rect 39948 22918 40000 22924
rect 39764 22704 39816 22710
rect 39764 22646 39816 22652
rect 39960 22642 39988 22918
rect 39948 22636 40000 22642
rect 39948 22578 40000 22584
rect 40144 22574 40172 23122
rect 40224 23112 40276 23118
rect 40224 23054 40276 23060
rect 40236 22778 40264 23054
rect 40224 22772 40276 22778
rect 40224 22714 40276 22720
rect 40328 22642 40356 23462
rect 40420 23322 40448 24754
rect 40592 24608 40644 24614
rect 40592 24550 40644 24556
rect 40604 23798 40632 24550
rect 41432 24410 41460 25230
rect 42064 24812 42116 24818
rect 42064 24754 42116 24760
rect 41420 24404 41472 24410
rect 41420 24346 41472 24352
rect 40592 23792 40644 23798
rect 40592 23734 40644 23740
rect 40684 23724 40736 23730
rect 40684 23666 40736 23672
rect 40408 23316 40460 23322
rect 40408 23258 40460 23264
rect 40696 23186 40724 23666
rect 40684 23180 40736 23186
rect 40684 23122 40736 23128
rect 40408 22772 40460 22778
rect 40408 22714 40460 22720
rect 40316 22636 40368 22642
rect 40316 22578 40368 22584
rect 40132 22568 40184 22574
rect 40132 22510 40184 22516
rect 40040 22500 40092 22506
rect 40040 22442 40092 22448
rect 39764 22432 39816 22438
rect 39764 22374 39816 22380
rect 39776 21622 39804 22374
rect 40052 22030 40080 22442
rect 40420 22234 40448 22714
rect 40696 22642 40724 23122
rect 41432 22982 41460 24346
rect 42076 23594 42104 24754
rect 42064 23588 42116 23594
rect 42064 23530 42116 23536
rect 42340 23248 42392 23254
rect 42340 23190 42392 23196
rect 41512 23112 41564 23118
rect 41512 23054 41564 23060
rect 41420 22976 41472 22982
rect 41420 22918 41472 22924
rect 40684 22636 40736 22642
rect 40684 22578 40736 22584
rect 40592 22568 40644 22574
rect 40592 22510 40644 22516
rect 40408 22228 40460 22234
rect 40408 22170 40460 22176
rect 40604 22030 40632 22510
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 40408 22024 40460 22030
rect 40408 21966 40460 21972
rect 40592 22024 40644 22030
rect 40592 21966 40644 21972
rect 39948 21956 40000 21962
rect 39948 21898 40000 21904
rect 40224 21956 40276 21962
rect 40224 21898 40276 21904
rect 39960 21622 39988 21898
rect 40132 21888 40184 21894
rect 40132 21830 40184 21836
rect 39764 21616 39816 21622
rect 39764 21558 39816 21564
rect 39948 21616 40000 21622
rect 39948 21558 40000 21564
rect 40144 20942 40172 21830
rect 40236 21486 40264 21898
rect 40420 21554 40448 21966
rect 40408 21548 40460 21554
rect 40460 21508 40540 21536
rect 40408 21490 40460 21496
rect 40224 21480 40276 21486
rect 40224 21422 40276 21428
rect 40132 20936 40184 20942
rect 40236 20924 40264 21422
rect 40236 20896 40448 20924
rect 40132 20878 40184 20884
rect 40316 19780 40368 19786
rect 40316 19722 40368 19728
rect 40132 19712 40184 19718
rect 40132 19654 40184 19660
rect 40144 19553 40172 19654
rect 40130 19544 40186 19553
rect 39856 19508 39908 19514
rect 40130 19479 40186 19488
rect 39856 19450 39908 19456
rect 39868 18290 39896 19450
rect 40040 19236 40092 19242
rect 40040 19178 40092 19184
rect 40052 18970 40080 19178
rect 40132 19168 40184 19174
rect 40132 19110 40184 19116
rect 40040 18964 40092 18970
rect 40040 18906 40092 18912
rect 40052 18834 40080 18906
rect 40040 18828 40092 18834
rect 40040 18770 40092 18776
rect 39948 18624 40000 18630
rect 39948 18566 40000 18572
rect 39960 18290 39988 18566
rect 40144 18426 40172 19110
rect 40224 18692 40276 18698
rect 40224 18634 40276 18640
rect 40236 18426 40264 18634
rect 40328 18630 40356 19722
rect 40420 19310 40448 20896
rect 40512 20398 40540 21508
rect 40696 21486 40724 22578
rect 41052 22160 41104 22166
rect 41052 22102 41104 22108
rect 40960 22024 41012 22030
rect 40960 21966 41012 21972
rect 40684 21480 40736 21486
rect 40684 21422 40736 21428
rect 40696 20942 40724 21422
rect 40684 20936 40736 20942
rect 40684 20878 40736 20884
rect 40696 20602 40724 20878
rect 40684 20596 40736 20602
rect 40684 20538 40736 20544
rect 40500 20392 40552 20398
rect 40500 20334 40552 20340
rect 40972 19718 41000 21966
rect 41064 21894 41092 22102
rect 41524 22098 41552 23054
rect 41512 22092 41564 22098
rect 41512 22034 41564 22040
rect 41144 22024 41196 22030
rect 41328 22024 41380 22030
rect 41196 21984 41328 22012
rect 41144 21966 41196 21972
rect 41328 21966 41380 21972
rect 42064 22024 42116 22030
rect 42064 21966 42116 21972
rect 42248 22024 42300 22030
rect 42248 21966 42300 21972
rect 41052 21888 41104 21894
rect 41052 21830 41104 21836
rect 42076 21690 42104 21966
rect 42260 21690 42288 21966
rect 42352 21962 42380 23190
rect 42340 21956 42392 21962
rect 42340 21898 42392 21904
rect 42064 21684 42116 21690
rect 42064 21626 42116 21632
rect 42248 21684 42300 21690
rect 42248 21626 42300 21632
rect 41696 21412 41748 21418
rect 41696 21354 41748 21360
rect 41512 20460 41564 20466
rect 41708 20448 41736 21354
rect 41788 21344 41840 21350
rect 41788 21286 41840 21292
rect 41800 20466 41828 21286
rect 42340 20936 42392 20942
rect 42340 20878 42392 20884
rect 42248 20800 42300 20806
rect 42248 20742 42300 20748
rect 41564 20420 41736 20448
rect 41788 20460 41840 20466
rect 41512 20402 41564 20408
rect 41788 20402 41840 20408
rect 41328 20324 41380 20330
rect 41248 20284 41328 20312
rect 41144 19780 41196 19786
rect 41144 19722 41196 19728
rect 40776 19712 40828 19718
rect 40776 19654 40828 19660
rect 40960 19712 41012 19718
rect 40960 19654 41012 19660
rect 40788 19446 40816 19654
rect 40776 19440 40828 19446
rect 40776 19382 40828 19388
rect 40408 19304 40460 19310
rect 40408 19246 40460 19252
rect 40316 18624 40368 18630
rect 40316 18566 40368 18572
rect 40132 18420 40184 18426
rect 40132 18362 40184 18368
rect 40224 18420 40276 18426
rect 40224 18362 40276 18368
rect 39856 18284 39908 18290
rect 39856 18226 39908 18232
rect 39948 18284 40000 18290
rect 39948 18226 40000 18232
rect 40420 18222 40448 19246
rect 40972 18698 41000 19654
rect 41156 19378 41184 19722
rect 41144 19372 41196 19378
rect 41144 19314 41196 19320
rect 41248 19310 41276 20284
rect 41328 20266 41380 20272
rect 42064 20052 42116 20058
rect 42064 19994 42116 20000
rect 41420 19780 41472 19786
rect 41420 19722 41472 19728
rect 41432 19514 41460 19722
rect 41510 19544 41566 19553
rect 41420 19508 41472 19514
rect 41510 19479 41566 19488
rect 41420 19450 41472 19456
rect 41236 19304 41288 19310
rect 41236 19246 41288 19252
rect 41524 18902 41552 19479
rect 41604 19372 41656 19378
rect 41604 19314 41656 19320
rect 41512 18896 41564 18902
rect 41512 18838 41564 18844
rect 40500 18692 40552 18698
rect 40500 18634 40552 18640
rect 40960 18692 41012 18698
rect 40960 18634 41012 18640
rect 41420 18692 41472 18698
rect 41420 18634 41472 18640
rect 40512 18222 40540 18634
rect 41328 18284 41380 18290
rect 41328 18226 41380 18232
rect 39764 18216 39816 18222
rect 39764 18158 39816 18164
rect 40408 18216 40460 18222
rect 40500 18216 40552 18222
rect 40408 18158 40460 18164
rect 40498 18184 40500 18193
rect 40552 18184 40554 18193
rect 39776 17270 39804 18158
rect 40498 18119 40554 18128
rect 41340 17814 41368 18226
rect 41432 17814 41460 18634
rect 41512 18420 41564 18426
rect 41512 18362 41564 18368
rect 41524 18170 41552 18362
rect 41616 18290 41644 19314
rect 42076 18766 42104 19994
rect 42260 19854 42288 20742
rect 42248 19848 42300 19854
rect 42248 19790 42300 19796
rect 42352 19174 42380 20878
rect 42340 19168 42392 19174
rect 42340 19110 42392 19116
rect 41880 18760 41932 18766
rect 41880 18702 41932 18708
rect 42064 18760 42116 18766
rect 42064 18702 42116 18708
rect 41696 18420 41748 18426
rect 41696 18362 41748 18368
rect 41708 18329 41736 18362
rect 41694 18320 41750 18329
rect 41604 18284 41656 18290
rect 41892 18290 41920 18702
rect 41694 18255 41750 18264
rect 41880 18284 41932 18290
rect 41604 18226 41656 18232
rect 41880 18226 41932 18232
rect 41524 18142 41644 18170
rect 41512 18080 41564 18086
rect 41512 18022 41564 18028
rect 41328 17808 41380 17814
rect 41328 17750 41380 17756
rect 41420 17808 41472 17814
rect 41420 17750 41472 17756
rect 40132 17740 40184 17746
rect 40132 17682 40184 17688
rect 40224 17740 40276 17746
rect 40224 17682 40276 17688
rect 40144 17610 40172 17682
rect 40236 17649 40264 17682
rect 40316 17672 40368 17678
rect 40222 17640 40278 17649
rect 40132 17604 40184 17610
rect 40316 17614 40368 17620
rect 41144 17672 41196 17678
rect 41144 17614 41196 17620
rect 41328 17672 41380 17678
rect 41524 17626 41552 18022
rect 41616 17814 41644 18142
rect 41696 18148 41748 18154
rect 41696 18090 41748 18096
rect 41604 17808 41656 17814
rect 41604 17750 41656 17756
rect 41380 17620 41552 17626
rect 41328 17614 41552 17620
rect 40222 17575 40278 17584
rect 40132 17546 40184 17552
rect 39764 17264 39816 17270
rect 39764 17206 39816 17212
rect 40328 17134 40356 17614
rect 40868 17196 40920 17202
rect 40868 17138 40920 17144
rect 40316 17128 40368 17134
rect 40316 17070 40368 17076
rect 40880 16833 40908 17138
rect 40866 16824 40922 16833
rect 40866 16759 40922 16768
rect 40408 16652 40460 16658
rect 40408 16594 40460 16600
rect 40420 16561 40448 16594
rect 40406 16552 40462 16561
rect 40406 16487 40462 16496
rect 39672 15632 39724 15638
rect 39672 15574 39724 15580
rect 39684 15366 39712 15574
rect 40500 15428 40552 15434
rect 40500 15370 40552 15376
rect 39672 15360 39724 15366
rect 39672 15302 39724 15308
rect 39684 15094 39712 15302
rect 39672 15088 39724 15094
rect 39672 15030 39724 15036
rect 40512 15026 40540 15370
rect 40500 15020 40552 15026
rect 40500 14962 40552 14968
rect 40040 14952 40092 14958
rect 40040 14894 40092 14900
rect 40224 14952 40276 14958
rect 40408 14952 40460 14958
rect 40224 14894 40276 14900
rect 40328 14912 40408 14940
rect 40052 14278 40080 14894
rect 40236 14822 40264 14894
rect 40224 14816 40276 14822
rect 40224 14758 40276 14764
rect 40224 14408 40276 14414
rect 40224 14350 40276 14356
rect 39856 14272 39908 14278
rect 39856 14214 39908 14220
rect 40040 14272 40092 14278
rect 40040 14214 40092 14220
rect 39868 13938 39896 14214
rect 39948 14068 40000 14074
rect 39948 14010 40000 14016
rect 39764 13932 39816 13938
rect 39764 13874 39816 13880
rect 39856 13932 39908 13938
rect 39856 13874 39908 13880
rect 39776 13190 39804 13874
rect 39856 13728 39908 13734
rect 39856 13670 39908 13676
rect 39868 13530 39896 13670
rect 39856 13524 39908 13530
rect 39856 13466 39908 13472
rect 39764 13184 39816 13190
rect 39764 13126 39816 13132
rect 39960 12986 39988 14010
rect 40236 13841 40264 14350
rect 40222 13832 40278 13841
rect 40222 13767 40278 13776
rect 40038 13424 40094 13433
rect 40038 13359 40094 13368
rect 40052 13326 40080 13359
rect 40040 13320 40092 13326
rect 40040 13262 40092 13268
rect 40132 13252 40184 13258
rect 40132 13194 40184 13200
rect 39948 12980 40000 12986
rect 39948 12922 40000 12928
rect 40144 12850 40172 13194
rect 40132 12844 40184 12850
rect 40132 12786 40184 12792
rect 40038 12608 40094 12617
rect 40038 12543 40094 12552
rect 40052 12442 40080 12543
rect 40040 12436 40092 12442
rect 39592 12406 39712 12434
rect 39304 12232 39356 12238
rect 39304 12174 39356 12180
rect 39396 12096 39448 12102
rect 39224 12044 39396 12050
rect 39224 12038 39448 12044
rect 39224 12022 39436 12038
rect 39224 11898 39252 12022
rect 39212 11892 39264 11898
rect 39212 11834 39264 11840
rect 39304 11892 39356 11898
rect 39304 11834 39356 11840
rect 39120 11824 39172 11830
rect 39120 11766 39172 11772
rect 39212 11552 39264 11558
rect 39212 11494 39264 11500
rect 39224 11150 39252 11494
rect 39212 11144 39264 11150
rect 39212 11086 39264 11092
rect 38936 10804 38988 10810
rect 38936 10746 38988 10752
rect 39316 9994 39344 11834
rect 39580 10464 39632 10470
rect 39580 10406 39632 10412
rect 39592 10130 39620 10406
rect 39580 10124 39632 10130
rect 39580 10066 39632 10072
rect 39304 9988 39356 9994
rect 39304 9930 39356 9936
rect 39120 9376 39172 9382
rect 39120 9318 39172 9324
rect 38660 9172 38712 9178
rect 38660 9114 38712 9120
rect 39132 8974 39160 9318
rect 39120 8968 39172 8974
rect 39120 8910 39172 8916
rect 38660 8900 38712 8906
rect 38660 8842 38712 8848
rect 38672 8634 38700 8842
rect 38292 8628 38344 8634
rect 38292 8570 38344 8576
rect 38660 8628 38712 8634
rect 38660 8570 38712 8576
rect 39132 8498 39160 8910
rect 39120 8492 39172 8498
rect 39120 8434 39172 8440
rect 37648 8424 37700 8430
rect 37648 8366 37700 8372
rect 37556 8356 37608 8362
rect 37556 8298 37608 8304
rect 37464 7948 37516 7954
rect 37464 7890 37516 7896
rect 37464 5636 37516 5642
rect 37464 5578 37516 5584
rect 36176 4208 36228 4214
rect 36176 4150 36228 4156
rect 36636 4208 36688 4214
rect 36636 4150 36688 4156
rect 35348 3664 35400 3670
rect 35348 3606 35400 3612
rect 35900 3392 35952 3398
rect 35900 3334 35952 3340
rect 36268 3392 36320 3398
rect 36268 3334 36320 3340
rect 35532 3052 35584 3058
rect 35532 2994 35584 3000
rect 35348 2984 35400 2990
rect 35348 2926 35400 2932
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34520 2372 34572 2378
rect 34520 2314 34572 2320
rect 34796 2372 34848 2378
rect 34796 2314 34848 2320
rect 34808 800 34836 2314
rect 35360 1578 35388 2926
rect 35176 1550 35388 1578
rect 35176 800 35204 1550
rect 35544 800 35572 2994
rect 35912 800 35940 3334
rect 36280 800 36308 3334
rect 36648 800 36676 4150
rect 37476 4010 37504 5578
rect 37568 5302 37596 8298
rect 39684 7750 39712 12406
rect 40040 12378 40092 12384
rect 39764 12164 39816 12170
rect 39764 12106 39816 12112
rect 39776 11150 39804 12106
rect 40040 11756 40092 11762
rect 40040 11698 40092 11704
rect 40224 11756 40276 11762
rect 40224 11698 40276 11704
rect 40052 11354 40080 11698
rect 40040 11348 40092 11354
rect 40040 11290 40092 11296
rect 39764 11144 39816 11150
rect 39764 11086 39816 11092
rect 40236 11014 40264 11698
rect 40328 11218 40356 14912
rect 40408 14894 40460 14900
rect 41052 14816 41104 14822
rect 41052 14758 41104 14764
rect 40684 14340 40736 14346
rect 40684 14282 40736 14288
rect 40776 14340 40828 14346
rect 40776 14282 40828 14288
rect 40500 13932 40552 13938
rect 40500 13874 40552 13880
rect 40512 12850 40540 13874
rect 40696 13326 40724 14282
rect 40788 13530 40816 14282
rect 40866 13968 40922 13977
rect 41064 13938 41092 14758
rect 41156 13938 41184 17614
rect 41340 17598 41552 17614
rect 41420 17128 41472 17134
rect 41420 17070 41472 17076
rect 41234 16824 41290 16833
rect 41234 16759 41236 16768
rect 41288 16759 41290 16768
rect 41236 16730 41288 16736
rect 41432 16658 41460 17070
rect 41510 16824 41566 16833
rect 41510 16759 41512 16768
rect 41564 16759 41566 16768
rect 41512 16730 41564 16736
rect 41420 16652 41472 16658
rect 41420 16594 41472 16600
rect 41328 16108 41380 16114
rect 41328 16050 41380 16056
rect 41340 15994 41368 16050
rect 41432 16046 41460 16594
rect 41616 16250 41644 17750
rect 41708 17678 41736 18090
rect 41696 17672 41748 17678
rect 41696 17614 41748 17620
rect 42064 16992 42116 16998
rect 42064 16934 42116 16940
rect 41880 16720 41932 16726
rect 41880 16662 41932 16668
rect 41892 16590 41920 16662
rect 42076 16590 42104 16934
rect 41880 16584 41932 16590
rect 41880 16526 41932 16532
rect 42064 16584 42116 16590
rect 42064 16526 42116 16532
rect 41512 16244 41564 16250
rect 41512 16186 41564 16192
rect 41604 16244 41656 16250
rect 41604 16186 41656 16192
rect 41248 15966 41368 15994
rect 41420 16040 41472 16046
rect 41420 15982 41472 15988
rect 41248 15910 41276 15966
rect 41236 15904 41288 15910
rect 41236 15846 41288 15852
rect 41328 15904 41380 15910
rect 41328 15846 41380 15852
rect 41340 15366 41368 15846
rect 41432 15609 41460 15982
rect 41524 15638 41552 16186
rect 41602 15872 41658 15881
rect 41602 15807 41658 15816
rect 41512 15632 41564 15638
rect 41418 15600 41474 15609
rect 41512 15574 41564 15580
rect 41418 15535 41420 15544
rect 41472 15535 41474 15544
rect 41420 15506 41472 15512
rect 41512 15496 41564 15502
rect 41512 15438 41564 15444
rect 41328 15360 41380 15366
rect 41328 15302 41380 15308
rect 41328 15156 41380 15162
rect 41328 15098 41380 15104
rect 41340 14414 41368 15098
rect 41524 14618 41552 15438
rect 41616 14770 41644 15807
rect 42064 15496 42116 15502
rect 42064 15438 42116 15444
rect 41696 15360 41748 15366
rect 41696 15302 41748 15308
rect 41708 14890 41736 15302
rect 42076 15094 42104 15438
rect 41880 15088 41932 15094
rect 41880 15030 41932 15036
rect 42064 15088 42116 15094
rect 42064 15030 42116 15036
rect 41892 14890 41920 15030
rect 41696 14884 41748 14890
rect 41696 14826 41748 14832
rect 41880 14884 41932 14890
rect 41880 14826 41932 14832
rect 42064 14884 42116 14890
rect 42064 14826 42116 14832
rect 41972 14816 42024 14822
rect 41616 14742 41736 14770
rect 41972 14758 42024 14764
rect 41512 14612 41564 14618
rect 41512 14554 41564 14560
rect 41328 14408 41380 14414
rect 41328 14350 41380 14356
rect 41420 14408 41472 14414
rect 41420 14350 41472 14356
rect 41432 14113 41460 14350
rect 41512 14340 41564 14346
rect 41512 14282 41564 14288
rect 41418 14104 41474 14113
rect 41418 14039 41474 14048
rect 40866 13903 40922 13912
rect 41052 13932 41104 13938
rect 40880 13734 40908 13903
rect 41052 13874 41104 13880
rect 41144 13932 41196 13938
rect 41144 13874 41196 13880
rect 40868 13728 40920 13734
rect 40868 13670 40920 13676
rect 40776 13524 40828 13530
rect 40776 13466 40828 13472
rect 40684 13320 40736 13326
rect 40684 13262 40736 13268
rect 41156 13190 41184 13874
rect 41432 13870 41460 14039
rect 41420 13864 41472 13870
rect 41420 13806 41472 13812
rect 41144 13184 41196 13190
rect 41144 13126 41196 13132
rect 41432 12986 41460 13806
rect 41524 13734 41552 14282
rect 41512 13728 41564 13734
rect 41510 13696 41512 13705
rect 41564 13696 41566 13705
rect 41510 13631 41566 13640
rect 41524 13530 41552 13631
rect 41512 13524 41564 13530
rect 41512 13466 41564 13472
rect 41420 12980 41472 12986
rect 41420 12922 41472 12928
rect 40500 12844 40552 12850
rect 40500 12786 40552 12792
rect 41236 12096 41288 12102
rect 41236 12038 41288 12044
rect 41248 11898 41276 12038
rect 41144 11892 41196 11898
rect 41144 11834 41196 11840
rect 41236 11892 41288 11898
rect 41236 11834 41288 11840
rect 40960 11824 41012 11830
rect 40960 11766 41012 11772
rect 40500 11552 40552 11558
rect 40500 11494 40552 11500
rect 40512 11218 40540 11494
rect 40972 11354 41000 11766
rect 41156 11694 41184 11834
rect 41144 11688 41196 11694
rect 41144 11630 41196 11636
rect 40960 11348 41012 11354
rect 40960 11290 41012 11296
rect 40316 11212 40368 11218
rect 40316 11154 40368 11160
rect 40500 11212 40552 11218
rect 40500 11154 40552 11160
rect 40224 11008 40276 11014
rect 40224 10950 40276 10956
rect 40236 10062 40264 10950
rect 40328 10674 40356 11154
rect 41420 10804 41472 10810
rect 41420 10746 41472 10752
rect 41432 10674 41460 10746
rect 40316 10668 40368 10674
rect 40316 10610 40368 10616
rect 41420 10668 41472 10674
rect 41420 10610 41472 10616
rect 41328 10464 41380 10470
rect 41328 10406 41380 10412
rect 41340 10266 41368 10406
rect 41328 10260 41380 10266
rect 41328 10202 41380 10208
rect 40224 10056 40276 10062
rect 40224 9998 40276 10004
rect 40236 8906 40264 9998
rect 40224 8900 40276 8906
rect 40224 8842 40276 8848
rect 39672 7744 39724 7750
rect 39672 7686 39724 7692
rect 37556 5296 37608 5302
rect 37556 5238 37608 5244
rect 38384 5296 38436 5302
rect 38384 5238 38436 5244
rect 38396 4826 38424 5238
rect 41708 4826 41736 14742
rect 41984 14385 42012 14758
rect 41970 14376 42026 14385
rect 41970 14311 42026 14320
rect 41788 12844 41840 12850
rect 41788 12786 41840 12792
rect 41800 12646 41828 12786
rect 41788 12640 41840 12646
rect 41788 12582 41840 12588
rect 41800 12102 41828 12582
rect 41788 12096 41840 12102
rect 41788 12038 41840 12044
rect 42076 10810 42104 14826
rect 42064 10804 42116 10810
rect 42064 10746 42116 10752
rect 42444 4826 42472 26318
rect 42628 21026 42656 26522
rect 43352 26512 43404 26518
rect 43352 26454 43404 26460
rect 42892 24744 42944 24750
rect 42892 24686 42944 24692
rect 42800 23724 42852 23730
rect 42800 23666 42852 23672
rect 42708 22636 42760 22642
rect 42708 22578 42760 22584
rect 42720 21690 42748 22578
rect 42812 22098 42840 23666
rect 42800 22092 42852 22098
rect 42800 22034 42852 22040
rect 42708 21684 42760 21690
rect 42708 21626 42760 21632
rect 42708 21548 42760 21554
rect 42708 21490 42760 21496
rect 42536 20998 42656 21026
rect 42536 18902 42564 20998
rect 42720 20806 42748 21490
rect 42708 20800 42760 20806
rect 42708 20742 42760 20748
rect 42800 20596 42852 20602
rect 42800 20538 42852 20544
rect 42616 20256 42668 20262
rect 42616 20198 42668 20204
rect 42628 19718 42656 20198
rect 42708 19780 42760 19786
rect 42708 19722 42760 19728
rect 42616 19712 42668 19718
rect 42616 19654 42668 19660
rect 42628 19174 42656 19654
rect 42616 19168 42668 19174
rect 42616 19110 42668 19116
rect 42524 18896 42576 18902
rect 42524 18838 42576 18844
rect 42628 18426 42656 19110
rect 42720 18834 42748 19722
rect 42708 18828 42760 18834
rect 42708 18770 42760 18776
rect 42720 18630 42748 18770
rect 42708 18624 42760 18630
rect 42708 18566 42760 18572
rect 42616 18420 42668 18426
rect 42616 18362 42668 18368
rect 42708 16992 42760 16998
rect 42708 16934 42760 16940
rect 42524 16584 42576 16590
rect 42522 16552 42524 16561
rect 42576 16552 42578 16561
rect 42522 16487 42578 16496
rect 42524 16040 42576 16046
rect 42524 15982 42576 15988
rect 42536 15502 42564 15982
rect 42616 15904 42668 15910
rect 42614 15872 42616 15881
rect 42668 15872 42670 15881
rect 42614 15807 42670 15816
rect 42524 15496 42576 15502
rect 42524 15438 42576 15444
rect 42616 15360 42668 15366
rect 42616 15302 42668 15308
rect 42524 15088 42576 15094
rect 42524 15030 42576 15036
rect 42536 13530 42564 15030
rect 42628 14958 42656 15302
rect 42616 14952 42668 14958
rect 42616 14894 42668 14900
rect 42616 14816 42668 14822
rect 42616 14758 42668 14764
rect 42628 14346 42656 14758
rect 42720 14414 42748 16934
rect 42812 16182 42840 20538
rect 42904 16726 42932 24686
rect 43260 23316 43312 23322
rect 43260 23258 43312 23264
rect 43272 22710 43300 23258
rect 43260 22704 43312 22710
rect 43260 22646 43312 22652
rect 43272 18426 43300 22646
rect 43364 22273 43392 26454
rect 44088 26444 44140 26450
rect 44088 26386 44140 26392
rect 44100 24750 44128 26386
rect 44088 24744 44140 24750
rect 44088 24686 44140 24692
rect 44088 24132 44140 24138
rect 44088 24074 44140 24080
rect 43996 23792 44048 23798
rect 43996 23734 44048 23740
rect 43350 22264 43406 22273
rect 43350 22199 43352 22208
rect 43404 22199 43406 22208
rect 43352 22170 43404 22176
rect 43364 22139 43392 22170
rect 43720 21888 43772 21894
rect 43720 21830 43772 21836
rect 43444 20936 43496 20942
rect 43444 20878 43496 20884
rect 43456 20058 43484 20878
rect 43732 20466 43760 21830
rect 44008 21146 44036 23734
rect 44100 23730 44128 24074
rect 44088 23724 44140 23730
rect 44088 23666 44140 23672
rect 43996 21140 44048 21146
rect 43996 21082 44048 21088
rect 44008 20913 44036 21082
rect 43994 20904 44050 20913
rect 43994 20839 44050 20848
rect 43720 20460 43772 20466
rect 43640 20420 43720 20448
rect 43444 20052 43496 20058
rect 43444 19994 43496 20000
rect 43260 18420 43312 18426
rect 43260 18362 43312 18368
rect 43272 18086 43300 18362
rect 43260 18080 43312 18086
rect 43260 18022 43312 18028
rect 43260 17536 43312 17542
rect 43260 17478 43312 17484
rect 43272 16998 43300 17478
rect 43260 16992 43312 16998
rect 43260 16934 43312 16940
rect 42892 16720 42944 16726
rect 42892 16662 42944 16668
rect 42904 16250 42932 16662
rect 43640 16658 43668 20420
rect 43720 20402 43772 20408
rect 44732 19848 44784 19854
rect 44732 19790 44784 19796
rect 44744 19446 44772 19790
rect 44732 19440 44784 19446
rect 44732 19382 44784 19388
rect 44088 18624 44140 18630
rect 44088 18566 44140 18572
rect 44100 18034 44128 18566
rect 44100 18006 44220 18034
rect 44192 16998 44220 18006
rect 44180 16992 44232 16998
rect 44180 16934 44232 16940
rect 44456 16992 44508 16998
rect 44456 16934 44508 16940
rect 43628 16652 43680 16658
rect 43628 16594 43680 16600
rect 42892 16244 42944 16250
rect 42892 16186 42944 16192
rect 42800 16176 42852 16182
rect 42800 16118 42852 16124
rect 42812 15706 42840 16118
rect 42800 15700 42852 15706
rect 42800 15642 42852 15648
rect 42904 15502 42932 16186
rect 42984 15904 43036 15910
rect 42984 15846 43036 15852
rect 42892 15496 42944 15502
rect 42996 15473 43024 15846
rect 43168 15700 43220 15706
rect 43168 15642 43220 15648
rect 42892 15438 42944 15444
rect 42982 15464 43038 15473
rect 42982 15399 43038 15408
rect 43180 15162 43208 15642
rect 43352 15496 43404 15502
rect 43352 15438 43404 15444
rect 43168 15156 43220 15162
rect 43168 15098 43220 15104
rect 43364 15026 43392 15438
rect 43444 15428 43496 15434
rect 43444 15370 43496 15376
rect 43456 15094 43484 15370
rect 43444 15088 43496 15094
rect 43444 15030 43496 15036
rect 43352 15020 43404 15026
rect 43352 14962 43404 14968
rect 43260 14816 43312 14822
rect 43260 14758 43312 14764
rect 42708 14408 42760 14414
rect 42708 14350 42760 14356
rect 42616 14340 42668 14346
rect 42616 14282 42668 14288
rect 43272 14074 43300 14758
rect 43456 14618 43484 15030
rect 43444 14612 43496 14618
rect 43444 14554 43496 14560
rect 43260 14068 43312 14074
rect 43260 14010 43312 14016
rect 42524 13524 42576 13530
rect 42524 13466 42576 13472
rect 42536 12102 42564 13466
rect 42524 12096 42576 12102
rect 42524 12038 42576 12044
rect 42536 8974 42564 12038
rect 43640 11694 43668 16594
rect 43812 16040 43864 16046
rect 43718 16008 43774 16017
rect 43812 15982 43864 15988
rect 43718 15943 43720 15952
rect 43772 15943 43774 15952
rect 43720 15914 43772 15920
rect 43628 11688 43680 11694
rect 43628 11630 43680 11636
rect 43640 9382 43668 11630
rect 43628 9376 43680 9382
rect 43628 9318 43680 9324
rect 42984 9104 43036 9110
rect 42984 9046 43036 9052
rect 42524 8968 42576 8974
rect 42524 8910 42576 8916
rect 42996 4826 43024 9046
rect 43732 6866 43760 15914
rect 43824 14074 43852 15982
rect 44468 15609 44496 16934
rect 44454 15600 44510 15609
rect 44454 15535 44510 15544
rect 44468 15366 44496 15535
rect 44456 15360 44508 15366
rect 44456 15302 44508 15308
rect 44272 14816 44324 14822
rect 44272 14758 44324 14764
rect 44284 14414 44312 14758
rect 44272 14408 44324 14414
rect 44272 14350 44324 14356
rect 43904 14272 43956 14278
rect 43904 14214 43956 14220
rect 43916 14074 43944 14214
rect 43812 14068 43864 14074
rect 43812 14010 43864 14016
rect 43904 14068 43956 14074
rect 43904 14010 43956 14016
rect 44468 9654 44496 15302
rect 44456 9648 44508 9654
rect 44456 9590 44508 9596
rect 43720 6860 43772 6866
rect 43720 6802 43772 6808
rect 44836 6186 44864 30534
rect 47584 29708 47636 29714
rect 47584 29650 47636 29656
rect 44916 26308 44968 26314
rect 44916 26250 44968 26256
rect 44928 6798 44956 26250
rect 46938 12336 46994 12345
rect 46938 12271 46994 12280
rect 46952 11762 46980 12271
rect 46940 11756 46992 11762
rect 46940 11698 46992 11704
rect 46204 9104 46256 9110
rect 46204 9046 46256 9052
rect 46216 8430 46244 9046
rect 46204 8424 46256 8430
rect 46204 8366 46256 8372
rect 44916 6792 44968 6798
rect 44916 6734 44968 6740
rect 44824 6180 44876 6186
rect 44824 6122 44876 6128
rect 38384 4820 38436 4826
rect 38384 4762 38436 4768
rect 41696 4820 41748 4826
rect 41696 4762 41748 4768
rect 42432 4820 42484 4826
rect 42432 4762 42484 4768
rect 42984 4820 43036 4826
rect 42984 4762 43036 4768
rect 37464 4004 37516 4010
rect 37464 3946 37516 3952
rect 37476 3534 37504 3946
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 37924 3392 37976 3398
rect 37924 3334 37976 3340
rect 38108 3392 38160 3398
rect 38108 3334 38160 3340
rect 37740 2848 37792 2854
rect 37740 2790 37792 2796
rect 37372 2576 37424 2582
rect 37372 2518 37424 2524
rect 37004 2304 37056 2310
rect 37004 2246 37056 2252
rect 37016 800 37044 2246
rect 37384 800 37412 2518
rect 37752 800 37780 2790
rect 37936 2446 37964 3334
rect 38120 3058 38148 3334
rect 38396 3058 38424 4762
rect 38660 4480 38712 4486
rect 38660 4422 38712 4428
rect 38672 4010 38700 4422
rect 40040 4140 40092 4146
rect 40040 4082 40092 4088
rect 38660 4004 38712 4010
rect 38660 3946 38712 3952
rect 38108 3052 38160 3058
rect 38108 2994 38160 3000
rect 38384 3052 38436 3058
rect 38384 2994 38436 3000
rect 38476 2848 38528 2854
rect 38476 2790 38528 2796
rect 37924 2440 37976 2446
rect 37924 2382 37976 2388
rect 38108 2304 38160 2310
rect 38108 2246 38160 2252
rect 38120 800 38148 2246
rect 38488 800 38516 2790
rect 38672 2774 38700 3946
rect 38936 3936 38988 3942
rect 38936 3878 38988 3884
rect 39304 3936 39356 3942
rect 39304 3878 39356 3884
rect 38948 3534 38976 3878
rect 38936 3528 38988 3534
rect 38936 3470 38988 3476
rect 38948 3194 38976 3470
rect 39316 3466 39344 3878
rect 40052 3534 40080 4082
rect 41708 3738 41736 4762
rect 41788 3936 41840 3942
rect 41788 3878 41840 3884
rect 41696 3732 41748 3738
rect 41696 3674 41748 3680
rect 41512 3664 41564 3670
rect 41512 3606 41564 3612
rect 40040 3528 40092 3534
rect 40092 3488 40172 3516
rect 40040 3470 40092 3476
rect 39304 3460 39356 3466
rect 39304 3402 39356 3408
rect 38936 3188 38988 3194
rect 38936 3130 38988 3136
rect 39316 3058 39344 3402
rect 40040 3392 40092 3398
rect 40040 3334 40092 3340
rect 39304 3052 39356 3058
rect 39304 2994 39356 3000
rect 38844 2848 38896 2854
rect 38844 2790 38896 2796
rect 39580 2848 39632 2854
rect 39580 2790 39632 2796
rect 38672 2746 38792 2774
rect 38764 2446 38792 2746
rect 38752 2440 38804 2446
rect 38752 2382 38804 2388
rect 38856 800 38884 2790
rect 39212 2304 39264 2310
rect 39212 2246 39264 2252
rect 39224 800 39252 2246
rect 39592 800 39620 2790
rect 39948 2576 40000 2582
rect 39948 2518 40000 2524
rect 39960 800 39988 2518
rect 40052 2446 40080 3334
rect 40144 3194 40172 3488
rect 40776 3392 40828 3398
rect 40776 3334 40828 3340
rect 40132 3188 40184 3194
rect 40132 3130 40184 3136
rect 40316 2848 40368 2854
rect 40316 2790 40368 2796
rect 40040 2440 40092 2446
rect 40040 2382 40092 2388
rect 40328 800 40356 2790
rect 40788 2446 40816 3334
rect 41052 2848 41104 2854
rect 41052 2790 41104 2796
rect 40776 2440 40828 2446
rect 40776 2382 40828 2388
rect 40684 2304 40736 2310
rect 40684 2246 40736 2252
rect 40696 800 40724 2246
rect 41064 800 41092 2790
rect 41420 2576 41472 2582
rect 41420 2518 41472 2524
rect 41432 800 41460 2518
rect 41524 2446 41552 3606
rect 41708 3534 41736 3674
rect 41800 3534 41828 3878
rect 41696 3528 41748 3534
rect 41696 3470 41748 3476
rect 41788 3528 41840 3534
rect 41788 3470 41840 3476
rect 41708 3058 41736 3470
rect 42444 3058 42472 4762
rect 42708 4140 42760 4146
rect 42708 4082 42760 4088
rect 42720 3738 42748 4082
rect 42708 3732 42760 3738
rect 42708 3674 42760 3680
rect 42800 3392 42852 3398
rect 42800 3334 42852 3340
rect 41696 3052 41748 3058
rect 41696 2994 41748 3000
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 42524 2916 42576 2922
rect 42524 2858 42576 2864
rect 41788 2848 41840 2854
rect 41788 2790 41840 2796
rect 41512 2440 41564 2446
rect 41512 2382 41564 2388
rect 41800 800 41828 2790
rect 42156 2304 42208 2310
rect 42156 2246 42208 2252
rect 42168 800 42196 2246
rect 42536 800 42564 2858
rect 42812 2514 42840 3334
rect 42892 2576 42944 2582
rect 42892 2518 42944 2524
rect 42800 2508 42852 2514
rect 42800 2450 42852 2456
rect 42904 800 42932 2518
rect 42996 2446 43024 4762
rect 46940 4752 46992 4758
rect 46940 4694 46992 4700
rect 45560 4616 45612 4622
rect 45560 4558 45612 4564
rect 43628 4480 43680 4486
rect 43628 4422 43680 4428
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 43088 3534 43116 3878
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 43640 3398 43668 4422
rect 45572 4146 45600 4558
rect 45928 4480 45980 4486
rect 45928 4422 45980 4428
rect 45560 4140 45612 4146
rect 45560 4082 45612 4088
rect 43904 4004 43956 4010
rect 43904 3946 43956 3952
rect 45744 4004 45796 4010
rect 45744 3946 45796 3952
rect 43628 3392 43680 3398
rect 43628 3334 43680 3340
rect 43640 3058 43668 3334
rect 43628 3052 43680 3058
rect 43628 2994 43680 3000
rect 43260 2916 43312 2922
rect 43260 2858 43312 2864
rect 42984 2440 43036 2446
rect 42984 2382 43036 2388
rect 43272 800 43300 2858
rect 43916 2446 43944 3946
rect 44640 3936 44692 3942
rect 44640 3878 44692 3884
rect 45652 3936 45704 3942
rect 45652 3878 45704 3884
rect 44088 3392 44140 3398
rect 44088 3334 44140 3340
rect 44100 3058 44128 3334
rect 44652 3058 44680 3878
rect 45192 3392 45244 3398
rect 45192 3334 45244 3340
rect 45560 3392 45612 3398
rect 45560 3334 45612 3340
rect 44088 3052 44140 3058
rect 44088 2994 44140 3000
rect 44640 3052 44692 3058
rect 44640 2994 44692 3000
rect 43996 2916 44048 2922
rect 43996 2858 44048 2864
rect 43904 2440 43956 2446
rect 43904 2382 43956 2388
rect 43628 2304 43680 2310
rect 43628 2246 43680 2252
rect 43640 800 43668 2246
rect 44008 800 44036 2858
rect 44732 2848 44784 2854
rect 44732 2790 44784 2796
rect 44364 2576 44416 2582
rect 44364 2518 44416 2524
rect 44376 800 44404 2518
rect 44744 800 44772 2790
rect 45204 2446 45232 3334
rect 45572 3058 45600 3334
rect 45560 3052 45612 3058
rect 45560 2994 45612 3000
rect 45468 2916 45520 2922
rect 45468 2858 45520 2864
rect 45192 2440 45244 2446
rect 45192 2382 45244 2388
rect 45100 2372 45152 2378
rect 45100 2314 45152 2320
rect 45112 800 45140 2314
rect 45480 800 45508 2858
rect 45664 2514 45692 3878
rect 45652 2508 45704 2514
rect 45652 2450 45704 2456
rect 45756 2446 45784 3946
rect 45940 3534 45968 4422
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 45928 3528 45980 3534
rect 45928 3470 45980 3476
rect 45836 3392 45888 3398
rect 45836 3334 45888 3340
rect 45744 2440 45796 2446
rect 45744 2382 45796 2388
rect 45848 800 45876 3334
rect 46308 3058 46336 3878
rect 46952 3534 46980 4694
rect 46940 3528 46992 3534
rect 46940 3470 46992 3476
rect 46572 3392 46624 3398
rect 46572 3334 46624 3340
rect 46296 3052 46348 3058
rect 46296 2994 46348 3000
rect 46204 2576 46256 2582
rect 46204 2518 46256 2524
rect 46216 800 46244 2518
rect 46584 800 46612 3334
rect 46940 3052 46992 3058
rect 46940 2994 46992 3000
rect 46952 800 46980 2994
rect 47596 2650 47624 29650
rect 47768 3936 47820 3942
rect 47768 3878 47820 3884
rect 47676 3392 47728 3398
rect 47676 3334 47728 3340
rect 47688 3126 47716 3334
rect 47676 3120 47728 3126
rect 47676 3062 47728 3068
rect 47584 2644 47636 2650
rect 47584 2586 47636 2592
rect 47308 2372 47360 2378
rect 47308 2314 47360 2320
rect 47320 800 47348 2314
rect 47688 800 47716 3062
rect 47780 2446 47808 3878
rect 47872 3194 47900 32370
rect 49332 31204 49384 31210
rect 49332 31146 49384 31152
rect 48596 28484 48648 28490
rect 48596 28426 48648 28432
rect 48504 26920 48556 26926
rect 48504 26862 48556 26868
rect 48320 10260 48372 10266
rect 48320 10202 48372 10208
rect 48332 8362 48360 10202
rect 48412 9648 48464 9654
rect 48412 9590 48464 9596
rect 48424 8838 48452 9590
rect 48412 8832 48464 8838
rect 48412 8774 48464 8780
rect 48320 8356 48372 8362
rect 48320 8298 48372 8304
rect 47860 3188 47912 3194
rect 47860 3130 47912 3136
rect 48412 3052 48464 3058
rect 48412 2994 48464 3000
rect 47768 2440 47820 2446
rect 47768 2382 47820 2388
rect 48044 2440 48096 2446
rect 48044 2382 48096 2388
rect 48056 800 48084 2382
rect 48424 800 48452 2994
rect 48516 2582 48544 26862
rect 48608 3194 48636 28426
rect 49056 14272 49108 14278
rect 49056 14214 49108 14220
rect 49068 12434 49096 14214
rect 49068 12406 49188 12434
rect 48964 10736 49016 10742
rect 48964 10678 49016 10684
rect 48780 9580 48832 9586
rect 48780 9522 48832 9528
rect 48792 7546 48820 9522
rect 48976 8974 49004 10678
rect 49056 9580 49108 9586
rect 49056 9522 49108 9528
rect 49068 9178 49096 9522
rect 49160 9178 49188 12406
rect 49056 9172 49108 9178
rect 49056 9114 49108 9120
rect 49148 9172 49200 9178
rect 49148 9114 49200 9120
rect 48964 8968 49016 8974
rect 48964 8910 49016 8916
rect 48780 7540 48832 7546
rect 48780 7482 48832 7488
rect 49056 3936 49108 3942
rect 49056 3878 49108 3884
rect 48872 3392 48924 3398
rect 48872 3334 48924 3340
rect 48596 3188 48648 3194
rect 48596 3130 48648 3136
rect 48504 2576 48556 2582
rect 48504 2518 48556 2524
rect 48884 2378 48912 3334
rect 49068 2446 49096 3878
rect 49344 3194 49372 31146
rect 49884 24676 49936 24682
rect 49884 24618 49936 24624
rect 49700 18692 49752 18698
rect 49700 18634 49752 18640
rect 49712 17814 49740 18634
rect 49896 18290 49924 24618
rect 49884 18284 49936 18290
rect 49884 18226 49936 18232
rect 49700 17808 49752 17814
rect 49700 17750 49752 17756
rect 49700 12232 49752 12238
rect 49700 12174 49752 12180
rect 49712 11801 49740 12174
rect 49698 11792 49754 11801
rect 49698 11727 49754 11736
rect 49700 8832 49752 8838
rect 49700 8774 49752 8780
rect 49712 7478 49740 8774
rect 49700 7472 49752 7478
rect 49700 7414 49752 7420
rect 49976 6792 50028 6798
rect 49976 6734 50028 6740
rect 49424 3392 49476 3398
rect 49424 3334 49476 3340
rect 49608 3392 49660 3398
rect 49608 3334 49660 3340
rect 49332 3188 49384 3194
rect 49332 3130 49384 3136
rect 49436 3058 49464 3334
rect 49424 3052 49476 3058
rect 49424 2994 49476 3000
rect 49620 2990 49648 3334
rect 49148 2984 49200 2990
rect 49148 2926 49200 2932
rect 49608 2984 49660 2990
rect 49608 2926 49660 2932
rect 49056 2440 49108 2446
rect 49056 2382 49108 2388
rect 48872 2372 48924 2378
rect 48872 2314 48924 2320
rect 48964 2372 49016 2378
rect 48964 2314 49016 2320
rect 48976 2258 49004 2314
rect 48792 2230 49004 2258
rect 48792 800 48820 2230
rect 49160 800 49188 2926
rect 49884 2916 49936 2922
rect 49884 2858 49936 2864
rect 49700 2440 49752 2446
rect 49620 2400 49700 2428
rect 49620 2360 49648 2400
rect 49700 2382 49752 2388
rect 49528 2332 49648 2360
rect 49528 800 49556 2332
rect 49896 800 49924 2858
rect 49988 2582 50016 6734
rect 50080 3194 50108 32399
rect 51172 32224 51224 32230
rect 51172 32166 51224 32172
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50804 29640 50856 29646
rect 50804 29582 50856 29588
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50436 9376 50488 9382
rect 50436 9318 50488 9324
rect 50448 8906 50476 9318
rect 50436 8900 50488 8906
rect 50436 8842 50488 8848
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50160 3936 50212 3942
rect 50160 3878 50212 3884
rect 50068 3188 50120 3194
rect 50068 3130 50120 3136
rect 49976 2576 50028 2582
rect 49976 2518 50028 2524
rect 50172 2378 50200 3878
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50816 3194 50844 29582
rect 51080 11824 51132 11830
rect 51080 11766 51132 11772
rect 51092 11150 51120 11766
rect 51080 11144 51132 11150
rect 51080 11086 51132 11092
rect 50896 9580 50948 9586
rect 50896 9522 50948 9528
rect 50908 8634 50936 9522
rect 50896 8628 50948 8634
rect 50896 8570 50948 8576
rect 51080 7744 51132 7750
rect 51080 7686 51132 7692
rect 50988 3936 51040 3942
rect 50988 3878 51040 3884
rect 51000 3466 51028 3878
rect 50988 3460 51040 3466
rect 50988 3402 51040 3408
rect 50804 3188 50856 3194
rect 50804 3130 50856 3136
rect 50620 3120 50672 3126
rect 50620 3062 50672 3068
rect 50160 2372 50212 2378
rect 50160 2314 50212 2320
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50252 2100 50304 2106
rect 50252 2042 50304 2048
rect 50264 800 50292 2042
rect 50632 800 50660 3062
rect 51000 800 51028 3402
rect 51092 2582 51120 7686
rect 51184 3738 51212 32166
rect 52840 31142 52868 43590
rect 52932 43353 52960 43658
rect 52918 43344 52974 43353
rect 52918 43279 52974 43288
rect 53012 42016 53064 42022
rect 53012 41958 53064 41964
rect 53024 41614 53052 41958
rect 53012 41608 53064 41614
rect 53012 41550 53064 41556
rect 53024 41177 53052 41550
rect 53010 41168 53066 41177
rect 53116 41138 53144 44338
rect 53010 41103 53066 41112
rect 53104 41132 53156 41138
rect 53104 41074 53156 41080
rect 52920 40928 52972 40934
rect 52920 40870 52972 40876
rect 52932 40526 52960 40870
rect 53208 40730 53236 47942
rect 53288 47592 53340 47598
rect 53288 47534 53340 47540
rect 53564 47592 53616 47598
rect 53564 47534 53616 47540
rect 53300 41750 53328 47534
rect 53576 47462 53604 47534
rect 53564 47456 53616 47462
rect 53564 47398 53616 47404
rect 53472 46504 53524 46510
rect 53472 46446 53524 46452
rect 53380 45960 53432 45966
rect 53380 45902 53432 45908
rect 53392 44441 53420 45902
rect 53484 44985 53512 46446
rect 53576 46073 53604 47398
rect 53656 47184 53708 47190
rect 53656 47126 53708 47132
rect 53668 47054 53696 47126
rect 53852 47122 53880 47942
rect 53840 47116 53892 47122
rect 53840 47058 53892 47064
rect 53656 47048 53708 47054
rect 53656 46990 53708 46996
rect 53562 46064 53618 46073
rect 53562 45999 53618 46008
rect 53668 45665 53696 46990
rect 53654 45656 53710 45665
rect 53654 45591 53710 45600
rect 53746 45520 53802 45529
rect 53746 45455 53748 45464
rect 53800 45455 53802 45464
rect 53748 45426 53800 45432
rect 53564 45416 53616 45422
rect 53564 45358 53616 45364
rect 53470 44976 53526 44985
rect 53470 44911 53526 44920
rect 53472 44532 53524 44538
rect 53472 44474 53524 44480
rect 53378 44432 53434 44441
rect 53378 44367 53434 44376
rect 53484 44334 53512 44474
rect 53472 44328 53524 44334
rect 53472 44270 53524 44276
rect 53380 43104 53432 43110
rect 53484 43081 53512 44270
rect 53576 43897 53604 45358
rect 53656 44872 53708 44878
rect 53656 44814 53708 44820
rect 53748 44872 53800 44878
rect 53748 44814 53800 44820
rect 53562 43888 53618 43897
rect 53562 43823 53618 43832
rect 53564 43784 53616 43790
rect 53564 43726 53616 43732
rect 53576 43314 53604 43726
rect 53668 43625 53696 44814
rect 53760 43926 53788 44814
rect 53748 43920 53800 43926
rect 53748 43862 53800 43868
rect 53748 43648 53800 43654
rect 53654 43616 53710 43625
rect 53748 43590 53800 43596
rect 53654 43551 53710 43560
rect 53564 43308 53616 43314
rect 53564 43250 53616 43256
rect 53656 43240 53708 43246
rect 53656 43182 53708 43188
rect 53380 43046 53432 43052
rect 53470 43072 53526 43081
rect 53392 42106 53420 43046
rect 53470 43007 53526 43016
rect 53472 42696 53524 42702
rect 53472 42638 53524 42644
rect 53484 42265 53512 42638
rect 53668 42537 53696 43182
rect 53760 42945 53788 43590
rect 53746 42936 53802 42945
rect 53746 42871 53802 42880
rect 53746 42800 53802 42809
rect 53746 42735 53748 42744
rect 53800 42735 53802 42744
rect 53748 42706 53800 42712
rect 53654 42528 53710 42537
rect 53654 42463 53710 42472
rect 53470 42256 53526 42265
rect 53470 42191 53526 42200
rect 53472 42152 53524 42158
rect 53392 42100 53472 42106
rect 53392 42094 53524 42100
rect 53392 42078 53512 42094
rect 53484 41993 53512 42078
rect 53470 41984 53526 41993
rect 53470 41919 53526 41928
rect 53288 41744 53340 41750
rect 53288 41686 53340 41692
rect 53656 41472 53708 41478
rect 53656 41414 53708 41420
rect 53472 41064 53524 41070
rect 53472 41006 53524 41012
rect 53196 40724 53248 40730
rect 53196 40666 53248 40672
rect 53484 40633 53512 41006
rect 53668 40905 53696 41414
rect 53654 40896 53710 40905
rect 53654 40831 53710 40840
rect 53470 40624 53526 40633
rect 53470 40559 53526 40568
rect 52920 40520 52972 40526
rect 52920 40462 52972 40468
rect 53656 40520 53708 40526
rect 53656 40462 53708 40468
rect 52932 39817 52960 40462
rect 53564 39976 53616 39982
rect 53564 39918 53616 39924
rect 53380 39840 53432 39846
rect 52918 39808 52974 39817
rect 53380 39782 53432 39788
rect 52918 39743 52974 39752
rect 53012 39432 53064 39438
rect 53012 39374 53064 39380
rect 53024 39001 53052 39374
rect 53010 38992 53066 39001
rect 53010 38927 53066 38936
rect 53392 38894 53420 39782
rect 53472 39432 53524 39438
rect 53472 39374 53524 39380
rect 53380 38888 53432 38894
rect 53380 38830 53432 38836
rect 53012 38752 53064 38758
rect 53010 38720 53012 38729
rect 53064 38720 53066 38729
rect 53010 38655 53066 38664
rect 53012 37664 53064 37670
rect 53010 37632 53012 37641
rect 53064 37632 53066 37641
rect 53010 37567 53066 37576
rect 53392 37369 53420 38830
rect 53484 37913 53512 39374
rect 53576 38457 53604 39918
rect 53668 39914 53696 40462
rect 53656 39908 53708 39914
rect 53656 39850 53708 39856
rect 53668 39545 53696 39850
rect 53748 39568 53800 39574
rect 53654 39536 53710 39545
rect 53748 39510 53800 39516
rect 53654 39471 53710 39480
rect 53656 39432 53708 39438
rect 53656 39374 53708 39380
rect 53562 38448 53618 38457
rect 53562 38383 53618 38392
rect 53668 38026 53696 39374
rect 53760 38418 53788 39510
rect 53748 38412 53800 38418
rect 53748 38354 53800 38360
rect 53748 38276 53800 38282
rect 53748 38218 53800 38224
rect 53576 37998 53696 38026
rect 53470 37904 53526 37913
rect 53470 37839 53526 37848
rect 53576 37466 53604 37998
rect 53656 37936 53708 37942
rect 53656 37878 53708 37884
rect 53668 37806 53696 37878
rect 53656 37800 53708 37806
rect 53656 37742 53708 37748
rect 53564 37460 53616 37466
rect 53564 37402 53616 37408
rect 53378 37360 53434 37369
rect 53378 37295 53434 37304
rect 53472 37324 53524 37330
rect 53472 37266 53524 37272
rect 53012 37256 53064 37262
rect 53012 37198 53064 37204
rect 53024 37097 53052 37198
rect 53010 37088 53066 37097
rect 53010 37023 53066 37032
rect 53024 36922 53052 37023
rect 53012 36916 53064 36922
rect 53012 36858 53064 36864
rect 53484 36281 53512 37266
rect 53564 37256 53616 37262
rect 53564 37198 53616 37204
rect 53576 36786 53604 37198
rect 53564 36780 53616 36786
rect 53564 36722 53616 36728
rect 53564 36644 53616 36650
rect 53564 36586 53616 36592
rect 53470 36272 53526 36281
rect 53470 36207 53526 36216
rect 53472 36168 53524 36174
rect 53472 36110 53524 36116
rect 53484 35737 53512 36110
rect 53576 36009 53604 36586
rect 53668 36553 53696 37742
rect 53760 36825 53788 38218
rect 53746 36816 53802 36825
rect 53746 36751 53802 36760
rect 53748 36712 53800 36718
rect 53748 36654 53800 36660
rect 53654 36544 53710 36553
rect 53654 36479 53710 36488
rect 53760 36378 53788 36654
rect 53748 36372 53800 36378
rect 53748 36314 53800 36320
rect 53562 36000 53618 36009
rect 53562 35935 53618 35944
rect 53470 35728 53526 35737
rect 53470 35663 53526 35672
rect 53472 35624 53524 35630
rect 53472 35566 53524 35572
rect 53484 35465 53512 35566
rect 53564 35488 53616 35494
rect 53470 35456 53526 35465
rect 53564 35430 53616 35436
rect 53470 35391 53526 35400
rect 53576 35086 53604 35430
rect 53288 35080 53340 35086
rect 53288 35022 53340 35028
rect 53564 35080 53616 35086
rect 53564 35022 53616 35028
rect 53012 34536 53064 34542
rect 53012 34478 53064 34484
rect 53024 34377 53052 34478
rect 53010 34368 53066 34377
rect 53010 34303 53066 34312
rect 53300 34105 53328 35022
rect 53470 34912 53526 34921
rect 53470 34847 53526 34856
rect 53484 34610 53512 34847
rect 53576 34649 53604 35022
rect 53562 34640 53618 34649
rect 53472 34604 53524 34610
rect 53562 34575 53618 34584
rect 53472 34546 53524 34552
rect 53656 34468 53708 34474
rect 53656 34410 53708 34416
rect 53380 34128 53432 34134
rect 53286 34096 53342 34105
rect 53380 34070 53432 34076
rect 53286 34031 53342 34040
rect 53104 33992 53156 33998
rect 53104 33934 53156 33940
rect 53116 33658 53144 33934
rect 53104 33652 53156 33658
rect 53104 33594 53156 33600
rect 53392 33386 53420 34070
rect 53668 33998 53696 34410
rect 53944 33998 53972 50662
rect 54036 35834 54064 52430
rect 54312 52426 54340 55200
rect 54300 52420 54352 52426
rect 54300 52362 54352 52368
rect 54312 52154 54340 52362
rect 54300 52148 54352 52154
rect 54300 52090 54352 52096
rect 54392 51332 54444 51338
rect 54392 51274 54444 51280
rect 54300 51264 54352 51270
rect 54300 51206 54352 51212
rect 54312 50318 54340 51206
rect 54404 50930 54432 51274
rect 54392 50924 54444 50930
rect 54392 50866 54444 50872
rect 54300 50312 54352 50318
rect 54300 50254 54352 50260
rect 54312 48249 54340 50254
rect 54404 49337 54432 50866
rect 54484 50244 54536 50250
rect 54484 50186 54536 50192
rect 54496 49842 54524 50186
rect 54484 49836 54536 49842
rect 54484 49778 54536 49784
rect 54390 49328 54446 49337
rect 54390 49263 54446 49272
rect 54298 48240 54354 48249
rect 54298 48175 54354 48184
rect 54496 47433 54524 49778
rect 54482 47424 54538 47433
rect 54482 47359 54538 47368
rect 54116 46980 54168 46986
rect 54116 46922 54168 46928
rect 54128 40730 54156 46922
rect 54300 42084 54352 42090
rect 54300 42026 54352 42032
rect 54312 41614 54340 42026
rect 54300 41608 54352 41614
rect 54300 41550 54352 41556
rect 54312 41414 54340 41550
rect 54312 41386 54432 41414
rect 54300 40996 54352 41002
rect 54300 40938 54352 40944
rect 54116 40724 54168 40730
rect 54116 40666 54168 40672
rect 54312 40526 54340 40938
rect 54300 40520 54352 40526
rect 54300 40462 54352 40468
rect 54312 39273 54340 40462
rect 54404 40089 54432 41386
rect 54390 40080 54446 40089
rect 54390 40015 54446 40024
rect 54298 39264 54354 39273
rect 54298 39199 54354 39208
rect 54024 35828 54076 35834
rect 54024 35770 54076 35776
rect 53656 33992 53708 33998
rect 53656 33934 53708 33940
rect 53932 33992 53984 33998
rect 53932 33934 53984 33940
rect 53380 33380 53432 33386
rect 53380 33322 53432 33328
rect 54300 33312 54352 33318
rect 54298 33280 54300 33289
rect 54352 33280 54354 33289
rect 54298 33215 54354 33224
rect 54300 32904 54352 32910
rect 54300 32846 54352 32852
rect 54312 32473 54340 32846
rect 54298 32464 54354 32473
rect 54298 32399 54354 32408
rect 54300 31816 54352 31822
rect 54300 31758 54352 31764
rect 54312 31657 54340 31758
rect 54298 31648 54354 31657
rect 54298 31583 54354 31592
rect 52828 31136 52880 31142
rect 52828 31078 52880 31084
rect 54300 31136 54352 31142
rect 54300 31078 54352 31084
rect 54312 30841 54340 31078
rect 54298 30832 54354 30841
rect 54298 30767 54354 30776
rect 54208 30048 54260 30054
rect 54206 30016 54208 30025
rect 54260 30016 54262 30025
rect 54206 29951 54262 29960
rect 54206 29744 54262 29753
rect 54206 29679 54262 29688
rect 54220 29646 54248 29679
rect 54208 29640 54260 29646
rect 54208 29582 54260 29588
rect 53564 29504 53616 29510
rect 53564 29446 53616 29452
rect 53576 29306 53604 29446
rect 53564 29300 53616 29306
rect 53564 29242 53616 29248
rect 54208 29300 54260 29306
rect 54208 29242 54260 29248
rect 54220 29209 54248 29242
rect 54206 29200 54262 29209
rect 54206 29135 54262 29144
rect 54220 28966 54248 28997
rect 54208 28960 54260 28966
rect 54206 28928 54208 28937
rect 54260 28928 54262 28937
rect 54206 28863 54262 28872
rect 54220 28558 54248 28863
rect 54208 28552 54260 28558
rect 54208 28494 54260 28500
rect 53472 28484 53524 28490
rect 53472 28426 53524 28432
rect 53196 28416 53248 28422
rect 53196 28358 53248 28364
rect 52828 28008 52880 28014
rect 52828 27950 52880 27956
rect 52840 27334 52868 27950
rect 52828 27328 52880 27334
rect 52828 27270 52880 27276
rect 52552 26852 52604 26858
rect 52552 26794 52604 26800
rect 52368 26784 52420 26790
rect 52368 26726 52420 26732
rect 52380 26586 52408 26726
rect 52368 26580 52420 26586
rect 52368 26522 52420 26528
rect 52564 26518 52592 26794
rect 52552 26512 52604 26518
rect 52552 26454 52604 26460
rect 52840 25770 52868 27270
rect 52920 26308 52972 26314
rect 52920 26250 52972 26256
rect 52828 25764 52880 25770
rect 52828 25706 52880 25712
rect 52932 25702 52960 26250
rect 52920 25696 52972 25702
rect 52920 25638 52972 25644
rect 52932 24138 52960 25638
rect 52920 24132 52972 24138
rect 52920 24074 52972 24080
rect 53208 18358 53236 28358
rect 53484 28121 53512 28426
rect 53564 28416 53616 28422
rect 53564 28358 53616 28364
rect 54206 28384 54262 28393
rect 53576 28218 53604 28358
rect 54206 28319 54262 28328
rect 54220 28218 54248 28319
rect 53564 28212 53616 28218
rect 53564 28154 53616 28160
rect 54208 28212 54260 28218
rect 54208 28154 54260 28160
rect 53470 28112 53526 28121
rect 53470 28047 53526 28056
rect 53472 27872 53524 27878
rect 53472 27814 53524 27820
rect 53484 27577 53512 27814
rect 53470 27568 53526 27577
rect 53470 27503 53526 27512
rect 53472 27464 53524 27470
rect 53472 27406 53524 27412
rect 53656 27464 53708 27470
rect 53656 27406 53708 27412
rect 53484 27033 53512 27406
rect 53470 27024 53526 27033
rect 53470 26959 53526 26968
rect 53564 26988 53616 26994
rect 53564 26930 53616 26936
rect 53576 26489 53604 26930
rect 53562 26480 53618 26489
rect 53562 26415 53618 26424
rect 53564 26376 53616 26382
rect 53564 26318 53616 26324
rect 53576 26217 53604 26318
rect 53562 26208 53618 26217
rect 53562 26143 53618 26152
rect 53472 25832 53524 25838
rect 53472 25774 53524 25780
rect 53484 25401 53512 25774
rect 53562 25664 53618 25673
rect 53562 25599 53618 25608
rect 53470 25392 53526 25401
rect 53470 25327 53526 25336
rect 53472 25152 53524 25158
rect 53470 25120 53472 25129
rect 53524 25120 53526 25129
rect 53470 25055 53526 25064
rect 53576 24818 53604 25599
rect 53564 24812 53616 24818
rect 53564 24754 53616 24760
rect 53472 24608 53524 24614
rect 53472 24550 53524 24556
rect 53484 24313 53512 24550
rect 53576 24410 53604 24754
rect 53564 24404 53616 24410
rect 53564 24346 53616 24352
rect 53470 24304 53526 24313
rect 53470 24239 53526 24248
rect 53564 23724 53616 23730
rect 53564 23666 53616 23672
rect 53288 23588 53340 23594
rect 53288 23530 53340 23536
rect 53472 23588 53524 23594
rect 53472 23530 53524 23536
rect 53300 22778 53328 23530
rect 53484 22778 53512 23530
rect 53576 23254 53604 23666
rect 53564 23248 53616 23254
rect 53562 23216 53564 23225
rect 53616 23216 53618 23225
rect 53562 23151 53618 23160
rect 53288 22772 53340 22778
rect 53288 22714 53340 22720
rect 53472 22772 53524 22778
rect 53472 22714 53524 22720
rect 53564 22024 53616 22030
rect 53564 21966 53616 21972
rect 53288 21956 53340 21962
rect 53288 21898 53340 21904
rect 53472 21956 53524 21962
rect 53472 21898 53524 21904
rect 53300 21593 53328 21898
rect 53484 21593 53512 21898
rect 53576 21690 53604 21966
rect 53564 21684 53616 21690
rect 53564 21626 53616 21632
rect 53286 21584 53342 21593
rect 53286 21519 53342 21528
rect 53470 21584 53526 21593
rect 53470 21519 53526 21528
rect 53564 20800 53616 20806
rect 53562 20768 53564 20777
rect 53616 20768 53618 20777
rect 53562 20703 53618 20712
rect 53286 20496 53342 20505
rect 53286 20431 53288 20440
rect 53340 20431 53342 20440
rect 53564 20460 53616 20466
rect 53288 20402 53340 20408
rect 53564 20402 53616 20408
rect 53576 19990 53604 20402
rect 53564 19984 53616 19990
rect 53562 19952 53564 19961
rect 53616 19952 53618 19961
rect 53562 19887 53618 19896
rect 53472 18692 53524 18698
rect 53472 18634 53524 18640
rect 53196 18352 53248 18358
rect 53484 18329 53512 18634
rect 53196 18294 53248 18300
rect 53470 18320 53526 18329
rect 53470 18255 53526 18264
rect 53472 18080 53524 18086
rect 53472 18022 53524 18028
rect 53288 17060 53340 17066
rect 53288 17002 53340 17008
rect 53300 16697 53328 17002
rect 53484 16794 53512 18022
rect 53564 17196 53616 17202
rect 53564 17138 53616 17144
rect 53472 16788 53524 16794
rect 53472 16730 53524 16736
rect 53576 16726 53604 17138
rect 53564 16720 53616 16726
rect 53286 16688 53342 16697
rect 53286 16623 53342 16632
rect 53562 16688 53564 16697
rect 53616 16688 53618 16697
rect 53562 16623 53618 16632
rect 53288 15972 53340 15978
rect 53288 15914 53340 15920
rect 53300 15638 53328 15914
rect 53668 15910 53696 27406
rect 54206 27296 54262 27305
rect 54206 27231 54262 27240
rect 54220 27062 54248 27231
rect 54208 27056 54260 27062
rect 54208 26998 54260 27004
rect 54206 26752 54262 26761
rect 54206 26687 54262 26696
rect 54220 26586 54248 26687
rect 54208 26580 54260 26586
rect 54208 26522 54260 26528
rect 54206 25936 54262 25945
rect 54206 25871 54262 25880
rect 53748 25832 53800 25838
rect 53748 25774 53800 25780
rect 53656 15904 53708 15910
rect 53656 15846 53708 15852
rect 53288 15632 53340 15638
rect 53288 15574 53340 15580
rect 53564 15496 53616 15502
rect 53564 15438 53616 15444
rect 53472 15428 53524 15434
rect 53472 15370 53524 15376
rect 53484 15065 53512 15370
rect 53576 15162 53604 15438
rect 53564 15156 53616 15162
rect 53564 15098 53616 15104
rect 53470 15056 53526 15065
rect 53470 14991 53526 15000
rect 53760 14822 53788 25774
rect 54220 25498 54248 25871
rect 54208 25492 54260 25498
rect 54208 25434 54260 25440
rect 54206 24848 54262 24857
rect 54206 24783 54262 24792
rect 54220 24206 54248 24783
rect 54208 24200 54260 24206
rect 54208 24142 54260 24148
rect 54116 24064 54168 24070
rect 54116 24006 54168 24012
rect 54206 24032 54262 24041
rect 54024 23860 54076 23866
rect 54024 23802 54076 23808
rect 54036 23662 54064 23802
rect 54128 23798 54156 24006
rect 54206 23967 54262 23976
rect 54220 23798 54248 23967
rect 54116 23792 54168 23798
rect 54116 23734 54168 23740
rect 54208 23792 54260 23798
rect 54208 23734 54260 23740
rect 54024 23656 54076 23662
rect 54024 23598 54076 23604
rect 54206 23488 54262 23497
rect 54206 23423 54262 23432
rect 54220 23322 54248 23423
rect 54208 23316 54260 23322
rect 54208 23258 54260 23264
rect 54208 22772 54260 22778
rect 54208 22714 54260 22720
rect 54220 22681 54248 22714
rect 54206 22672 54262 22681
rect 54206 22607 54262 22616
rect 54206 22400 54262 22409
rect 54206 22335 54262 22344
rect 54220 22030 54248 22335
rect 54208 22024 54260 22030
rect 54022 21992 54078 22001
rect 54208 21966 54260 21972
rect 54022 21927 54024 21936
rect 54076 21927 54078 21936
rect 54024 21898 54076 21904
rect 54206 21856 54262 21865
rect 54206 21791 54262 21800
rect 54220 21690 54248 21791
rect 54208 21684 54260 21690
rect 54208 21626 54260 21632
rect 54208 21072 54260 21078
rect 54206 21040 54208 21049
rect 54260 21040 54262 21049
rect 54206 20975 54262 20984
rect 54206 20768 54262 20777
rect 54206 20703 54262 20712
rect 54220 20534 54248 20703
rect 54208 20528 54260 20534
rect 54208 20470 54260 20476
rect 54206 20224 54262 20233
rect 54206 20159 54262 20168
rect 54220 20058 54248 20159
rect 54208 20052 54260 20058
rect 54208 19994 54260 20000
rect 54208 19508 54260 19514
rect 54208 19450 54260 19456
rect 54220 19417 54248 19450
rect 54206 19408 54262 19417
rect 54206 19343 54262 19352
rect 54220 19174 54248 19205
rect 54208 19168 54260 19174
rect 54206 19136 54208 19145
rect 54260 19136 54262 19145
rect 54206 19071 54262 19080
rect 54220 18766 54248 19071
rect 54208 18760 54260 18766
rect 54208 18702 54260 18708
rect 54206 18592 54262 18601
rect 54206 18527 54262 18536
rect 54220 18426 54248 18527
rect 54208 18420 54260 18426
rect 54208 18362 54260 18368
rect 54116 17876 54168 17882
rect 54116 17818 54168 17824
rect 54128 17338 54156 17818
rect 54208 17808 54260 17814
rect 54206 17776 54208 17785
rect 54260 17776 54262 17785
rect 54206 17711 54262 17720
rect 54220 17542 54248 17573
rect 54208 17536 54260 17542
rect 54206 17504 54208 17513
rect 54260 17504 54262 17513
rect 54206 17439 54262 17448
rect 54116 17332 54168 17338
rect 54116 17274 54168 17280
rect 54220 17270 54248 17439
rect 54208 17264 54260 17270
rect 54208 17206 54260 17212
rect 54206 16960 54262 16969
rect 54206 16895 54262 16904
rect 54220 16794 54248 16895
rect 54208 16788 54260 16794
rect 54208 16730 54260 16736
rect 54208 16244 54260 16250
rect 54208 16186 54260 16192
rect 54220 16153 54248 16186
rect 54206 16144 54262 16153
rect 54024 16108 54076 16114
rect 54206 16079 54262 16088
rect 54024 16050 54076 16056
rect 54036 15706 54064 16050
rect 54206 15872 54262 15881
rect 54206 15807 54262 15816
rect 54024 15700 54076 15706
rect 54024 15642 54076 15648
rect 54220 15502 54248 15807
rect 54208 15496 54260 15502
rect 54208 15438 54260 15444
rect 54206 15328 54262 15337
rect 54206 15263 54262 15272
rect 54220 15162 54248 15263
rect 54208 15156 54260 15162
rect 54208 15098 54260 15104
rect 54024 15020 54076 15026
rect 54024 14962 54076 14968
rect 54036 14929 54064 14962
rect 54022 14920 54078 14929
rect 54022 14855 54078 14864
rect 53748 14816 53800 14822
rect 53748 14758 53800 14764
rect 54208 14544 54260 14550
rect 54206 14512 54208 14521
rect 54260 14512 54262 14521
rect 54206 14447 54262 14456
rect 54024 14408 54076 14414
rect 54024 14350 54076 14356
rect 54036 14074 54064 14350
rect 54220 14278 54248 14309
rect 54208 14272 54260 14278
rect 54206 14240 54208 14249
rect 54260 14240 54262 14249
rect 54206 14175 54262 14184
rect 54024 14068 54076 14074
rect 54024 14010 54076 14016
rect 54220 14006 54248 14175
rect 54208 14000 54260 14006
rect 54208 13942 54260 13948
rect 53564 13932 53616 13938
rect 53564 13874 53616 13880
rect 53288 13796 53340 13802
rect 53288 13738 53340 13744
rect 53300 13530 53328 13738
rect 53288 13524 53340 13530
rect 53288 13466 53340 13472
rect 53576 13462 53604 13874
rect 53840 13864 53892 13870
rect 53840 13806 53892 13812
rect 53564 13456 53616 13462
rect 53562 13424 53564 13433
rect 53616 13424 53618 13433
rect 53562 13359 53618 13368
rect 53852 12986 53880 13806
rect 54024 13728 54076 13734
rect 54024 13670 54076 13676
rect 54206 13696 54262 13705
rect 54036 13326 54064 13670
rect 54206 13631 54262 13640
rect 54220 13530 54248 13631
rect 54208 13524 54260 13530
rect 54208 13466 54260 13472
rect 54024 13320 54076 13326
rect 54024 13262 54076 13268
rect 53840 12980 53892 12986
rect 53840 12922 53892 12928
rect 54208 12980 54260 12986
rect 54208 12922 54260 12928
rect 54220 12889 54248 12922
rect 54206 12880 54262 12889
rect 54206 12815 54262 12824
rect 54206 12608 54262 12617
rect 54206 12543 54262 12552
rect 54220 12238 54248 12543
rect 54208 12232 54260 12238
rect 54208 12174 54260 12180
rect 53196 12164 53248 12170
rect 53196 12106 53248 12112
rect 53472 12164 53524 12170
rect 53472 12106 53524 12112
rect 53564 12164 53616 12170
rect 53564 12106 53616 12112
rect 53208 9674 53236 12106
rect 53484 11801 53512 12106
rect 53576 11898 53604 12106
rect 54206 12064 54262 12073
rect 54206 11999 54262 12008
rect 54220 11898 54248 11999
rect 53564 11892 53616 11898
rect 53564 11834 53616 11840
rect 54208 11892 54260 11898
rect 54208 11834 54260 11840
rect 53470 11792 53526 11801
rect 53470 11727 53526 11736
rect 54208 11280 54260 11286
rect 54206 11248 54208 11257
rect 54260 11248 54262 11257
rect 54206 11183 54262 11192
rect 54220 11014 54248 11045
rect 54208 11008 54260 11014
rect 54206 10976 54208 10985
rect 54260 10976 54262 10985
rect 54206 10911 54262 10920
rect 54220 10742 54248 10911
rect 54208 10736 54260 10742
rect 54208 10678 54260 10684
rect 53472 10668 53524 10674
rect 53472 10610 53524 10616
rect 53288 10532 53340 10538
rect 53288 10474 53340 10480
rect 53116 9646 53236 9674
rect 53300 9674 53328 10474
rect 53380 10464 53432 10470
rect 53380 10406 53432 10412
rect 53392 9994 53420 10406
rect 53484 10198 53512 10610
rect 54206 10432 54262 10441
rect 54206 10367 54262 10376
rect 54220 10266 54248 10367
rect 54208 10260 54260 10266
rect 54208 10202 54260 10208
rect 53472 10192 53524 10198
rect 53470 10160 53472 10169
rect 53524 10160 53526 10169
rect 53470 10095 53526 10104
rect 53564 10124 53616 10130
rect 53564 10066 53616 10072
rect 53380 9988 53432 9994
rect 53380 9930 53432 9936
rect 53300 9654 53420 9674
rect 53300 9648 53432 9654
rect 53300 9646 53380 9648
rect 53116 9382 53144 9646
rect 53380 9590 53432 9596
rect 53576 9586 53604 10066
rect 54206 9616 54262 9625
rect 53564 9580 53616 9586
rect 54206 9551 54262 9560
rect 53564 9522 53616 9528
rect 51632 9376 51684 9382
rect 51632 9318 51684 9324
rect 52276 9376 52328 9382
rect 52276 9318 52328 9324
rect 52460 9376 52512 9382
rect 52460 9318 52512 9324
rect 53104 9376 53156 9382
rect 53576 9353 53604 9522
rect 54220 9450 54248 9551
rect 54208 9444 54260 9450
rect 54208 9386 54260 9392
rect 53104 9318 53156 9324
rect 53562 9344 53618 9353
rect 51644 8974 51672 9318
rect 52288 9042 52316 9318
rect 52472 9110 52500 9318
rect 53562 9279 53618 9288
rect 52736 9172 52788 9178
rect 52736 9114 52788 9120
rect 52460 9104 52512 9110
rect 52460 9046 52512 9052
rect 52276 9036 52328 9042
rect 52276 8978 52328 8984
rect 52748 8974 52776 9114
rect 51632 8968 51684 8974
rect 51632 8910 51684 8916
rect 52460 8968 52512 8974
rect 52460 8910 52512 8916
rect 52736 8968 52788 8974
rect 52736 8910 52788 8916
rect 52184 8492 52236 8498
rect 52184 8434 52236 8440
rect 52196 7993 52224 8434
rect 52472 8090 52500 8910
rect 53196 8900 53248 8906
rect 53196 8842 53248 8848
rect 52736 8832 52788 8838
rect 52736 8774 52788 8780
rect 52460 8084 52512 8090
rect 52460 8026 52512 8032
rect 52182 7984 52238 7993
rect 52182 7919 52238 7928
rect 52276 7880 52328 7886
rect 52276 7822 52328 7828
rect 52288 7449 52316 7822
rect 52748 7818 52776 8774
rect 52920 7880 52972 7886
rect 52920 7822 52972 7828
rect 52736 7812 52788 7818
rect 52736 7754 52788 7760
rect 52932 7546 52960 7822
rect 53208 7546 53236 8842
rect 53564 8832 53616 8838
rect 53564 8774 53616 8780
rect 54206 8800 54262 8809
rect 53470 8528 53526 8537
rect 53470 8463 53472 8472
rect 53524 8463 53526 8472
rect 53472 8434 53524 8440
rect 53576 8362 53604 8774
rect 54206 8735 54262 8744
rect 54220 8634 54248 8735
rect 54208 8628 54260 8634
rect 54208 8570 54260 8576
rect 53564 8356 53616 8362
rect 53564 8298 53616 8304
rect 54300 7744 54352 7750
rect 53378 7712 53434 7721
rect 54300 7686 54352 7692
rect 53378 7647 53434 7656
rect 52920 7540 52972 7546
rect 52920 7482 52972 7488
rect 53196 7540 53248 7546
rect 53196 7482 53248 7488
rect 52274 7440 52330 7449
rect 53392 7410 53420 7647
rect 52274 7375 52330 7384
rect 53380 7404 53432 7410
rect 53380 7346 53432 7352
rect 53392 7002 53420 7346
rect 54114 7168 54170 7177
rect 54114 7103 54170 7112
rect 54128 7002 54156 7103
rect 53380 6996 53432 7002
rect 53380 6938 53432 6944
rect 54116 6996 54168 7002
rect 54116 6938 54168 6944
rect 51264 6860 51316 6866
rect 51264 6802 51316 6808
rect 51276 6633 51304 6802
rect 54312 6798 54340 7686
rect 54392 7404 54444 7410
rect 54392 7346 54444 7352
rect 54404 6905 54432 7346
rect 54390 6896 54446 6905
rect 54390 6831 54446 6840
rect 54300 6792 54352 6798
rect 54300 6734 54352 6740
rect 51262 6624 51318 6633
rect 51262 6559 51318 6568
rect 54404 6458 54432 6831
rect 54392 6452 54444 6458
rect 54392 6394 54444 6400
rect 51540 6180 51592 6186
rect 51540 6122 51592 6128
rect 51172 3732 51224 3738
rect 51172 3674 51224 3680
rect 51552 3194 51580 6122
rect 51816 3392 51868 3398
rect 51816 3334 51868 3340
rect 52000 3392 52052 3398
rect 52000 3334 52052 3340
rect 51540 3188 51592 3194
rect 51540 3130 51592 3136
rect 51828 3126 51856 3334
rect 51816 3120 51868 3126
rect 51816 3062 51868 3068
rect 51080 2576 51132 2582
rect 51080 2518 51132 2524
rect 51814 2408 51870 2417
rect 52012 2378 52040 3334
rect 51814 2343 51816 2352
rect 51868 2343 51870 2352
rect 52000 2372 52052 2378
rect 51816 2314 51868 2320
rect 52000 2314 52052 2320
rect 52012 2106 52040 2314
rect 52000 2100 52052 2106
rect 52000 2042 52052 2048
rect 19812 734 20024 762
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 34058 0 34114 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 37002 0 37058 800
rect 37370 0 37426 800
rect 37738 0 37794 800
rect 38106 0 38162 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42522 0 42578 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43994 0 44050 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46202 0 46258 800
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47306 0 47362 800
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49146 0 49202 800
rect 49514 0 49570 800
rect 49882 0 49938 800
rect 50250 0 50306 800
rect 50618 0 50674 800
rect 50986 0 51042 800
<< via2 >>
rect 1490 52128 1546 52184
rect 1674 51584 1730 51640
rect 1674 51040 1730 51096
rect 1674 49408 1730 49464
rect 2042 41112 2098 41168
rect 1674 37984 1730 38040
rect 1582 37440 1638 37496
rect 2778 52672 2834 52728
rect 2778 50496 2834 50552
rect 2778 49952 2834 50008
rect 2778 48864 2834 48920
rect 2778 48320 2834 48376
rect 2778 47776 2834 47832
rect 2778 47232 2834 47288
rect 2502 44240 2558 44296
rect 2226 36624 2282 36680
rect 2778 46688 2834 46744
rect 2778 46144 2834 46200
rect 2778 45600 2834 45656
rect 2778 45056 2834 45112
rect 2778 44512 2834 44568
rect 2778 43968 2834 44024
rect 2778 43424 2834 43480
rect 2778 42880 2834 42936
rect 2778 42336 2834 42392
rect 2778 41792 2834 41848
rect 2778 41248 2834 41304
rect 2778 40704 2834 40760
rect 2778 40160 2834 40216
rect 2778 39616 2834 39672
rect 2778 39072 2834 39128
rect 2778 38528 2834 38584
rect 2778 36896 2834 36952
rect 2778 36352 2834 36408
rect 2778 35808 2834 35864
rect 2778 35264 2834 35320
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 3238 34992 3294 35048
rect 1582 34720 1638 34776
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 2778 34176 2834 34232
rect 2778 33632 2834 33688
rect 11610 43152 11666 43208
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 2778 33088 2834 33144
rect 1582 32544 1638 32600
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 2778 32000 2834 32056
rect 2778 31456 2834 31512
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 2778 30912 2834 30968
rect 2778 30368 2834 30424
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 2226 29844 2282 29880
rect 2226 29824 2228 29844
rect 2228 29824 2280 29844
rect 2280 29824 2282 29844
rect 1582 29280 1638 29336
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 2778 28736 2834 28792
rect 2778 28192 2834 28248
rect 2226 27668 2282 27704
rect 2226 27648 2228 27668
rect 2228 27648 2280 27668
rect 2280 27648 2282 27668
rect 1582 27104 1638 27160
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 2778 26560 2834 26616
rect 2226 26036 2282 26072
rect 2226 26016 2228 26036
rect 2228 26016 2280 26036
rect 2280 26016 2282 26036
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 1582 25492 1638 25528
rect 1582 25472 1584 25492
rect 1584 25472 1636 25492
rect 1636 25472 1638 25492
rect 1582 24928 1638 24984
rect 1674 24384 1730 24440
rect 1674 23840 1730 23896
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 1674 23296 1730 23352
rect 1674 22752 1730 22808
rect 1674 22208 1730 22264
rect 1674 21664 1730 21720
rect 1674 21120 1730 21176
rect 1674 20576 1730 20632
rect 1674 20032 1730 20088
rect 1674 19488 1730 19544
rect 1674 18944 1730 19000
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 1674 18400 1730 18456
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1582 17856 1638 17912
rect 1674 17312 1730 17368
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 1674 16768 1730 16824
rect 1674 16224 1730 16280
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1674 15680 1730 15736
rect 1674 15136 1730 15192
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1674 14592 1730 14648
rect 1674 14048 1730 14104
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 1674 13504 1730 13560
rect 1674 12960 1730 13016
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 21270 36100 21326 36136
rect 21270 36080 21272 36100
rect 21272 36080 21324 36100
rect 21324 36080 21326 36100
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 1674 12416 1730 12472
rect 1674 11872 1730 11928
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 1674 11328 1730 11384
rect 1674 10784 1730 10840
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1674 10240 1730 10296
rect 1674 9696 1730 9752
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 1674 9152 1730 9208
rect 1674 8608 1730 8664
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 1674 8064 1730 8120
rect 1674 7520 1730 7576
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1674 6976 1730 7032
rect 1674 6432 1730 6488
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 1674 5888 1730 5944
rect 1674 5344 1730 5400
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 1674 4800 1730 4856
rect 1674 4256 1730 4312
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1674 3712 1730 3768
rect 1674 3168 1730 3224
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10046 3884 10048 3904
rect 10048 3884 10100 3904
rect 10100 3884 10102 3904
rect 10046 3848 10102 3884
rect 10138 3596 10194 3632
rect 10138 3576 10140 3596
rect 10140 3576 10192 3596
rect 10192 3576 10194 3596
rect 9954 3340 9956 3360
rect 9956 3340 10008 3360
rect 10008 3340 10010 3360
rect 9954 3304 10010 3340
rect 10690 3848 10746 3904
rect 10874 3304 10930 3360
rect 12438 5108 12440 5128
rect 12440 5108 12492 5128
rect 12492 5108 12494 5128
rect 12438 5072 12494 5108
rect 14738 15428 14794 15464
rect 14738 15408 14740 15428
rect 14740 15408 14792 15428
rect 14792 15408 14794 15428
rect 14738 15020 14794 15056
rect 14738 15000 14740 15020
rect 14740 15000 14792 15020
rect 14792 15000 14794 15020
rect 14646 14320 14702 14376
rect 14462 13948 14464 13968
rect 14464 13948 14516 13968
rect 14516 13948 14518 13968
rect 14462 13912 14518 13948
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 21178 35264 21234 35320
rect 21178 34992 21234 35048
rect 21730 35028 21732 35048
rect 21732 35028 21784 35048
rect 21784 35028 21786 35048
rect 21730 34992 21786 35028
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 22374 37168 22430 37224
rect 22558 36644 22614 36680
rect 22558 36624 22560 36644
rect 22560 36624 22612 36644
rect 22612 36624 22614 36644
rect 23386 40296 23442 40352
rect 23478 38528 23534 38584
rect 22926 35980 22928 36000
rect 22928 35980 22980 36000
rect 22980 35980 22982 36000
rect 22926 35944 22982 35980
rect 23018 35536 23074 35592
rect 24030 38156 24032 38176
rect 24032 38156 24084 38176
rect 24084 38156 24086 38176
rect 24030 38120 24086 38156
rect 24030 37460 24086 37496
rect 24030 37440 24032 37460
rect 24032 37440 24084 37460
rect 24084 37440 24086 37460
rect 24950 41928 25006 41984
rect 24858 38936 24914 38992
rect 23478 35708 23480 35728
rect 23480 35708 23532 35728
rect 23532 35708 23534 35728
rect 23478 35672 23534 35708
rect 23478 35028 23480 35048
rect 23480 35028 23532 35048
rect 23532 35028 23534 35048
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 15106 16124 15108 16144
rect 15108 16124 15160 16144
rect 15160 16124 15162 16144
rect 15106 16088 15162 16124
rect 15106 14476 15162 14512
rect 15106 14456 15108 14476
rect 15108 14456 15160 14476
rect 15160 14456 15162 14476
rect 14922 13524 14978 13560
rect 14922 13504 14924 13524
rect 14924 13504 14976 13524
rect 14976 13504 14978 13524
rect 12530 2760 12586 2816
rect 12898 2760 12954 2816
rect 15566 15952 15622 16008
rect 13818 5108 13820 5128
rect 13820 5108 13872 5128
rect 13872 5108 13874 5128
rect 13818 5072 13874 5108
rect 14646 8336 14702 8392
rect 14462 3596 14518 3632
rect 14462 3576 14464 3596
rect 14464 3576 14516 3596
rect 14516 3576 14518 3596
rect 15750 9152 15806 9208
rect 16762 16652 16818 16688
rect 16762 16632 16764 16652
rect 16764 16632 16816 16652
rect 16816 16632 16818 16652
rect 16210 9596 16212 9616
rect 16212 9596 16264 9616
rect 16264 9596 16266 9616
rect 16210 9560 16266 9596
rect 18234 17740 18290 17776
rect 18234 17720 18236 17740
rect 18236 17720 18288 17740
rect 18288 17720 18290 17740
rect 17406 15952 17462 16008
rect 17314 8900 17370 8936
rect 17314 8880 17316 8900
rect 17316 8880 17368 8900
rect 17368 8880 17370 8900
rect 17590 13504 17646 13560
rect 18142 14320 18198 14376
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19062 17720 19118 17776
rect 17774 8880 17830 8936
rect 18602 9560 18658 9616
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 20258 16632 20314 16688
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19614 13932 19670 13968
rect 19614 13912 19616 13932
rect 19616 13912 19668 13932
rect 19668 13912 19670 13932
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19798 12316 19800 12336
rect 19800 12316 19852 12336
rect 19852 12316 19854 12336
rect 19798 12280 19854 12316
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 18418 9152 18474 9208
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 20074 12144 20130 12200
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 20902 16108 20958 16144
rect 20902 16088 20904 16108
rect 20904 16088 20956 16108
rect 20956 16088 20958 16108
rect 20810 15408 20866 15464
rect 20718 14456 20774 14512
rect 18602 3848 18658 3904
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 23478 34992 23534 35028
rect 23754 35536 23810 35592
rect 24674 38392 24730 38448
rect 25778 40432 25834 40488
rect 24398 35264 24454 35320
rect 24214 34040 24270 34096
rect 21454 15408 21510 15464
rect 21914 15000 21970 15056
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 23110 21800 23166 21856
rect 23110 16788 23166 16824
rect 23110 16768 23112 16788
rect 23112 16768 23164 16788
rect 23164 16768 23166 16788
rect 22190 12280 22246 12336
rect 22190 12008 22246 12064
rect 23018 12860 23020 12880
rect 23020 12860 23072 12880
rect 23072 12860 23074 12880
rect 23018 12824 23074 12860
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 23570 20984 23626 21040
rect 25410 36488 25466 36544
rect 25502 36352 25558 36408
rect 25042 35708 25044 35728
rect 25044 35708 25096 35728
rect 25096 35708 25098 35728
rect 25042 35672 25098 35708
rect 24030 17484 24032 17504
rect 24032 17484 24084 17504
rect 24084 17484 24086 17504
rect 24030 17448 24086 17484
rect 23754 15036 23756 15056
rect 23756 15036 23808 15056
rect 23808 15036 23810 15056
rect 23754 15000 23810 15036
rect 24398 20440 24454 20496
rect 24950 31864 25006 31920
rect 25594 36116 25596 36136
rect 25596 36116 25648 36136
rect 25648 36116 25650 36136
rect 25594 36080 25650 36116
rect 26054 41656 26110 41712
rect 26238 41248 26294 41304
rect 26514 41520 26570 41576
rect 26146 40704 26202 40760
rect 26146 40568 26202 40624
rect 26422 40024 26478 40080
rect 26054 38800 26110 38856
rect 25870 36624 25926 36680
rect 26054 37304 26110 37360
rect 25410 34448 25466 34504
rect 25042 17720 25098 17776
rect 25134 17584 25190 17640
rect 24674 17196 24730 17232
rect 24674 17176 24676 17196
rect 24676 17176 24728 17196
rect 24728 17176 24730 17196
rect 25042 16652 25098 16688
rect 26238 37576 26294 37632
rect 26146 35400 26202 35456
rect 26882 39480 26938 39536
rect 26606 38292 26608 38312
rect 26608 38292 26660 38312
rect 26660 38292 26662 38312
rect 26606 38256 26662 38292
rect 26514 36896 26570 36952
rect 27066 38936 27122 38992
rect 26790 38664 26846 38720
rect 27526 41964 27528 41984
rect 27528 41964 27580 41984
rect 27580 41964 27582 41984
rect 27526 41928 27582 41964
rect 27434 41248 27490 41304
rect 27526 40568 27582 40624
rect 27342 40160 27398 40216
rect 27986 41812 28042 41848
rect 27986 41792 27988 41812
rect 27988 41792 28040 41812
rect 28040 41792 28042 41812
rect 27986 41656 28042 41712
rect 27986 41384 28042 41440
rect 27710 41248 27766 41304
rect 27802 40704 27858 40760
rect 27434 38936 27490 38992
rect 27618 38956 27674 38992
rect 27618 38936 27620 38956
rect 27620 38936 27672 38956
rect 27672 38936 27674 38956
rect 27526 38528 27582 38584
rect 27158 38392 27214 38448
rect 26698 37848 26754 37904
rect 26698 37612 26700 37632
rect 26700 37612 26752 37632
rect 26752 37612 26754 37632
rect 26698 37576 26754 37612
rect 27158 38120 27214 38176
rect 27342 37460 27398 37496
rect 27342 37440 27344 37460
rect 27344 37440 27396 37460
rect 27396 37440 27398 37460
rect 26790 37188 26846 37224
rect 27066 37204 27068 37224
rect 27068 37204 27120 37224
rect 27120 37204 27122 37224
rect 26790 37168 26792 37188
rect 26792 37168 26844 37188
rect 26844 37168 26846 37188
rect 27066 37168 27122 37204
rect 27066 36896 27122 36952
rect 26698 35672 26754 35728
rect 27618 38256 27674 38312
rect 27526 36216 27582 36272
rect 27434 35944 27490 36000
rect 27526 35808 27582 35864
rect 27434 35536 27490 35592
rect 27618 35536 27674 35592
rect 27342 35264 27398 35320
rect 26422 27548 26424 27568
rect 26424 27548 26476 27568
rect 26476 27548 26478 27568
rect 26422 27512 26478 27548
rect 26790 31728 26846 31784
rect 26974 31864 27030 31920
rect 25042 16632 25044 16652
rect 25044 16632 25096 16652
rect 25096 16632 25098 16652
rect 23570 9460 23572 9480
rect 23572 9460 23624 9480
rect 23624 9460 23626 9480
rect 23570 9424 23626 9460
rect 23754 7384 23810 7440
rect 25318 14900 25320 14920
rect 25320 14900 25372 14920
rect 25372 14900 25374 14920
rect 25318 14864 25374 14900
rect 25318 9560 25374 9616
rect 25226 9424 25282 9480
rect 26238 16768 26294 16824
rect 26054 15156 26110 15192
rect 26054 15136 26056 15156
rect 26056 15136 26108 15156
rect 26108 15136 26110 15156
rect 26330 12144 26386 12200
rect 26514 20984 26570 21040
rect 26146 9288 26202 9344
rect 26422 9036 26478 9072
rect 26422 9016 26424 9036
rect 26424 9016 26476 9036
rect 26476 9016 26478 9036
rect 28078 40452 28134 40488
rect 28078 40432 28080 40452
rect 28080 40432 28132 40452
rect 28132 40432 28134 40452
rect 28262 41656 28318 41712
rect 28538 41384 28594 41440
rect 28814 41928 28870 41984
rect 28722 41792 28778 41848
rect 28722 41520 28778 41576
rect 28078 38800 28134 38856
rect 27894 37712 27950 37768
rect 27894 37188 27950 37224
rect 27894 37168 27896 37188
rect 27896 37168 27948 37188
rect 27948 37168 27950 37188
rect 27894 36660 27896 36680
rect 27896 36660 27948 36680
rect 27948 36660 27950 36680
rect 27894 36624 27950 36660
rect 27894 36488 27950 36544
rect 28538 40160 28594 40216
rect 28262 39480 28318 39536
rect 28446 38392 28502 38448
rect 28262 37984 28318 38040
rect 28262 37612 28264 37632
rect 28264 37612 28316 37632
rect 28316 37612 28318 37632
rect 28262 37576 28318 37612
rect 28170 37032 28226 37088
rect 28262 36896 28318 36952
rect 28078 34448 28134 34504
rect 27986 34040 28042 34096
rect 28722 40588 28778 40624
rect 28722 40568 28724 40588
rect 28724 40568 28776 40588
rect 28776 40568 28778 40588
rect 28814 40296 28870 40352
rect 29366 43152 29422 43208
rect 29642 43188 29644 43208
rect 29644 43188 29696 43208
rect 29696 43188 29698 43208
rect 29642 43152 29698 43188
rect 29090 40840 29146 40896
rect 28998 38528 29054 38584
rect 28998 38428 29006 38448
rect 29006 38428 29054 38448
rect 28998 38392 29054 38428
rect 28814 37848 28870 37904
rect 29458 40876 29460 40896
rect 29460 40876 29512 40896
rect 29512 40876 29514 40896
rect 29458 40840 29514 40876
rect 28722 36660 28724 36680
rect 28724 36660 28776 36680
rect 28776 36660 28778 36680
rect 28722 36624 28778 36660
rect 28722 36352 28778 36408
rect 28998 36488 29054 36544
rect 28814 36236 28870 36272
rect 28814 36216 28816 36236
rect 28816 36216 28868 36236
rect 28868 36216 28870 36236
rect 28630 35808 28686 35864
rect 28538 35692 28594 35728
rect 28538 35672 28540 35692
rect 28540 35672 28592 35692
rect 28592 35672 28594 35692
rect 28814 35536 28870 35592
rect 28722 35264 28778 35320
rect 28998 36100 29054 36136
rect 28998 36080 29000 36100
rect 29000 36080 29052 36100
rect 29052 36080 29054 36100
rect 29090 35436 29092 35456
rect 29092 35436 29144 35456
rect 29144 35436 29146 35456
rect 29090 35400 29146 35436
rect 30286 42744 30342 42800
rect 29826 38700 29828 38720
rect 29828 38700 29880 38720
rect 29880 38700 29882 38720
rect 29274 37712 29330 37768
rect 29274 35944 29330 36000
rect 29458 37984 29514 38040
rect 29826 38664 29882 38700
rect 29734 37984 29790 38040
rect 29458 36352 29514 36408
rect 28998 34992 29054 35048
rect 29366 35400 29422 35456
rect 28262 33088 28318 33144
rect 29090 33360 29146 33416
rect 27434 21528 27490 21584
rect 27526 20340 27528 20360
rect 27528 20340 27580 20360
rect 27580 20340 27582 20360
rect 27526 20304 27582 20340
rect 27710 17740 27766 17776
rect 27710 17720 27712 17740
rect 27712 17720 27764 17740
rect 27764 17720 27766 17740
rect 27434 17176 27490 17232
rect 28630 21428 28632 21448
rect 28632 21428 28684 21448
rect 28684 21428 28686 21448
rect 28630 21392 28686 21428
rect 28354 19488 28410 19544
rect 28814 20304 28870 20360
rect 28630 19292 28686 19348
rect 27986 17484 27988 17504
rect 27988 17484 28040 17504
rect 28040 17484 28042 17504
rect 27986 17448 28042 17484
rect 27710 15272 27766 15328
rect 27618 14900 27620 14920
rect 27620 14900 27672 14920
rect 27672 14900 27674 14920
rect 27618 14864 27674 14900
rect 27710 12824 27766 12880
rect 27434 9424 27490 9480
rect 26790 3732 26846 3768
rect 26790 3712 26792 3732
rect 26792 3712 26844 3732
rect 26844 3712 26846 3732
rect 28354 18300 28356 18320
rect 28356 18300 28408 18320
rect 28408 18300 28410 18320
rect 28354 18264 28410 18300
rect 28722 18808 28778 18864
rect 28630 17312 28686 17368
rect 28078 15544 28134 15600
rect 27894 12416 27950 12472
rect 27986 12008 28042 12064
rect 28262 15136 28318 15192
rect 29642 37868 29698 37904
rect 29642 37848 29644 37868
rect 29644 37848 29696 37868
rect 29696 37848 29698 37868
rect 29642 34604 29698 34640
rect 29642 34584 29644 34604
rect 29644 34584 29696 34604
rect 29696 34584 29698 34604
rect 29090 18264 29146 18320
rect 28906 17584 28962 17640
rect 28814 17312 28870 17368
rect 28998 16224 29054 16280
rect 29458 19896 29514 19952
rect 30102 41676 30158 41712
rect 30102 41656 30104 41676
rect 30104 41656 30156 41676
rect 30156 41656 30158 41676
rect 30378 42236 30380 42256
rect 30380 42236 30432 42256
rect 30432 42236 30434 42256
rect 30378 42200 30434 42236
rect 30286 37168 30342 37224
rect 30378 34720 30434 34776
rect 31022 42744 31078 42800
rect 31482 41656 31538 41712
rect 31482 40044 31538 40080
rect 31482 40024 31484 40044
rect 31484 40024 31536 40044
rect 31536 40024 31538 40044
rect 30562 34892 30564 34912
rect 30564 34892 30616 34912
rect 30616 34892 30618 34912
rect 30562 34856 30618 34892
rect 28446 9560 28502 9616
rect 28630 8780 28632 8800
rect 28632 8780 28684 8800
rect 28684 8780 28686 8800
rect 28630 8744 28686 8780
rect 28630 3732 28686 3768
rect 28630 3712 28632 3732
rect 28632 3712 28684 3732
rect 28684 3712 28686 3732
rect 29090 11636 29092 11656
rect 29092 11636 29144 11656
rect 29144 11636 29146 11656
rect 29090 11600 29146 11636
rect 29090 11328 29146 11384
rect 28906 9288 28962 9344
rect 29826 20576 29882 20632
rect 30470 21392 30526 21448
rect 29550 13504 29606 13560
rect 29458 11328 29514 11384
rect 29366 8336 29422 8392
rect 30286 19760 30342 19816
rect 30286 19660 30288 19680
rect 30288 19660 30340 19680
rect 30340 19660 30342 19680
rect 30286 19624 30342 19660
rect 30010 18264 30066 18320
rect 29826 14476 29882 14512
rect 29826 14456 29828 14476
rect 29828 14456 29880 14476
rect 29880 14456 29882 14476
rect 30010 13776 30066 13832
rect 29918 11772 29920 11792
rect 29920 11772 29972 11792
rect 29972 11772 29974 11792
rect 29918 11736 29974 11772
rect 29826 11600 29882 11656
rect 29918 10784 29974 10840
rect 29918 9696 29974 9752
rect 29734 9424 29790 9480
rect 29642 6976 29698 7032
rect 30194 13776 30250 13832
rect 30470 15272 30526 15328
rect 30838 37884 30840 37904
rect 30840 37884 30892 37904
rect 30892 37884 30894 37904
rect 30838 37848 30894 37884
rect 31482 38276 31538 38312
rect 31482 38256 31484 38276
rect 31484 38256 31536 38276
rect 31536 38256 31538 38276
rect 31022 37984 31078 38040
rect 31206 37984 31262 38040
rect 31206 37032 31262 37088
rect 31206 36352 31262 36408
rect 30930 34720 30986 34776
rect 31114 34468 31170 34504
rect 31114 34448 31116 34468
rect 31116 34448 31168 34468
rect 31168 34448 31170 34468
rect 31298 34584 31354 34640
rect 31482 34992 31538 35048
rect 30930 27648 30986 27704
rect 30838 18572 30840 18592
rect 30840 18572 30892 18592
rect 30892 18572 30894 18592
rect 30838 18536 30894 18572
rect 31390 21836 31392 21856
rect 31392 21836 31444 21856
rect 31444 21836 31446 21856
rect 31390 21800 31446 21836
rect 31022 19760 31078 19816
rect 30746 18300 30748 18320
rect 30748 18300 30800 18320
rect 30800 18300 30802 18320
rect 30746 18264 30802 18300
rect 31114 17720 31170 17776
rect 31390 18420 31446 18456
rect 31390 18400 31392 18420
rect 31392 18400 31444 18420
rect 31444 18400 31446 18420
rect 31390 17720 31446 17776
rect 31298 16088 31354 16144
rect 30562 15136 30618 15192
rect 30286 11328 30342 11384
rect 30654 12416 30710 12472
rect 31574 31728 31630 31784
rect 31758 37848 31814 37904
rect 32310 44260 32366 44296
rect 32310 44240 32312 44260
rect 32312 44240 32364 44260
rect 32364 44240 32366 44260
rect 33322 46996 33324 47016
rect 33324 46996 33376 47016
rect 33376 46996 33378 47016
rect 32586 41556 32588 41576
rect 32588 41556 32640 41576
rect 32640 41556 32642 41576
rect 32586 41520 32642 41556
rect 32770 41148 32772 41168
rect 32772 41148 32824 41168
rect 32824 41148 32826 41168
rect 32770 41112 32826 41148
rect 32678 40840 32734 40896
rect 32586 40468 32588 40488
rect 32588 40468 32640 40488
rect 32640 40468 32642 40488
rect 32586 40432 32642 40468
rect 31942 36216 31998 36272
rect 31758 23860 31814 23896
rect 31758 23840 31760 23860
rect 31760 23840 31812 23860
rect 31812 23840 31814 23860
rect 31758 18284 31814 18320
rect 31758 18264 31760 18284
rect 31760 18264 31812 18284
rect 31812 18264 31814 18284
rect 31022 12844 31078 12880
rect 31022 12824 31024 12844
rect 31024 12824 31076 12844
rect 31076 12824 31078 12844
rect 31022 11328 31078 11384
rect 30746 10668 30802 10704
rect 30746 10648 30748 10668
rect 30748 10648 30800 10668
rect 30800 10648 30802 10668
rect 30378 9868 30380 9888
rect 30380 9868 30432 9888
rect 30432 9868 30434 9888
rect 30378 9832 30434 9868
rect 30746 7420 30748 7440
rect 30748 7420 30800 7440
rect 30800 7420 30802 7440
rect 30746 7384 30802 7420
rect 31390 10784 31446 10840
rect 31850 10684 31852 10704
rect 31852 10684 31904 10704
rect 31904 10684 31906 10704
rect 31850 10648 31906 10684
rect 31850 9036 31906 9072
rect 31850 9016 31852 9036
rect 31852 9016 31904 9036
rect 31904 9016 31906 9036
rect 31850 8608 31906 8664
rect 33322 46960 33378 46996
rect 33322 41792 33378 41848
rect 33598 40840 33654 40896
rect 34334 41792 34390 41848
rect 33966 40060 33968 40080
rect 33968 40060 34020 40080
rect 34020 40060 34022 40080
rect 33966 40024 34022 40060
rect 32218 26016 32274 26072
rect 33230 37868 33286 37904
rect 33230 37848 33232 37868
rect 33232 37848 33284 37868
rect 33284 37848 33286 37868
rect 33230 36524 33232 36544
rect 33232 36524 33284 36544
rect 33284 36524 33286 36544
rect 33230 36488 33286 36524
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 35622 46960 35678 47016
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34702 42200 34758 42256
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 35530 41656 35586 41712
rect 35254 41132 35310 41168
rect 35254 41112 35256 41132
rect 35256 41112 35308 41132
rect 35308 41112 35310 41132
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34426 40432 34482 40488
rect 34610 40432 34666 40488
rect 34334 37712 34390 37768
rect 33782 37168 33838 37224
rect 33506 34892 33508 34912
rect 33508 34892 33560 34912
rect 33560 34892 33562 34912
rect 33506 34856 33562 34892
rect 33230 22072 33286 22128
rect 33598 26036 33654 26072
rect 33598 26016 33600 26036
rect 33600 26016 33652 26036
rect 33652 26016 33654 26036
rect 33598 25236 33600 25256
rect 33600 25236 33652 25256
rect 33652 25236 33654 25256
rect 33598 25200 33654 25236
rect 33506 23976 33562 24032
rect 33506 23840 33562 23896
rect 32126 19624 32182 19680
rect 32034 18672 32090 18728
rect 32402 17584 32458 17640
rect 32310 15952 32366 16008
rect 32494 16108 32550 16144
rect 33506 17040 33562 17096
rect 32494 16088 32496 16108
rect 32496 16088 32548 16108
rect 32548 16088 32550 16108
rect 32402 13640 32458 13696
rect 32402 12724 32404 12744
rect 32404 12724 32456 12744
rect 32456 12724 32458 12744
rect 32402 12688 32458 12724
rect 32034 11228 32036 11248
rect 32036 11228 32088 11248
rect 32088 11228 32090 11248
rect 32034 11192 32090 11228
rect 32310 9036 32366 9072
rect 32310 9016 32312 9036
rect 32312 9016 32364 9036
rect 32364 9016 32366 9036
rect 32586 12844 32642 12880
rect 32586 12824 32588 12844
rect 32588 12824 32640 12844
rect 32640 12824 32642 12844
rect 32586 11076 32642 11112
rect 32586 11056 32588 11076
rect 32588 11056 32640 11076
rect 32640 11056 32642 11076
rect 32770 10668 32826 10704
rect 32770 10648 32772 10668
rect 32772 10648 32824 10668
rect 32824 10648 32826 10668
rect 33414 13504 33470 13560
rect 33690 14456 33746 14512
rect 33046 9968 33102 10024
rect 33598 9036 33654 9072
rect 33598 9016 33600 9036
rect 33600 9016 33652 9036
rect 33652 9016 33654 9036
rect 33874 8780 33876 8800
rect 33876 8780 33928 8800
rect 33928 8780 33930 8800
rect 33874 8744 33930 8780
rect 33322 3732 33378 3768
rect 34334 23432 34390 23488
rect 35622 41520 35678 41576
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35438 23976 35494 24032
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 33322 3712 33324 3732
rect 33324 3712 33376 3732
rect 33376 3712 33378 3732
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35530 22772 35586 22808
rect 35530 22752 35532 22772
rect 35532 22752 35584 22772
rect 35584 22752 35586 22772
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34426 17040 34482 17096
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34978 18400 35034 18456
rect 34702 18264 34758 18320
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35162 16224 35218 16280
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34334 12144 34390 12200
rect 35530 20052 35586 20088
rect 35530 20032 35532 20052
rect 35532 20032 35584 20052
rect 35584 20032 35586 20052
rect 35530 17040 35586 17096
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35530 13132 35532 13152
rect 35532 13132 35584 13152
rect 35584 13132 35586 13152
rect 35530 13096 35586 13132
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35346 12164 35402 12200
rect 35346 12144 35348 12164
rect 35348 12144 35400 12164
rect 35400 12144 35402 12164
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 51998 52556 52054 52592
rect 51998 52536 52000 52556
rect 52000 52536 52052 52556
rect 52052 52536 52054 52556
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50894 46996 50896 47016
rect 50896 46996 50948 47016
rect 50948 46996 50950 47016
rect 50894 46960 50950 46996
rect 51446 47096 51502 47152
rect 51630 46960 51686 47016
rect 51814 46980 51870 47016
rect 51814 46960 51816 46980
rect 51816 46960 51868 46980
rect 51868 46960 51870 46980
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 52366 47912 52422 47968
rect 52182 46824 52238 46880
rect 52642 46552 52698 46608
rect 52182 45736 52238 45792
rect 52458 44940 52514 44976
rect 52458 44920 52460 44940
rect 52460 44920 52512 44940
rect 52512 44920 52514 44940
rect 52182 44648 52238 44704
rect 53470 49000 53526 49056
rect 53562 48728 53618 48784
rect 53654 48456 53710 48512
rect 53102 47640 53158 47696
rect 53010 46316 53012 46336
rect 53012 46316 53064 46336
rect 53064 46316 53066 46336
rect 53010 46280 53066 46316
rect 53010 45228 53012 45248
rect 53012 45228 53064 45248
rect 53064 45228 53066 45248
rect 53010 45192 53066 45228
rect 53010 44140 53012 44160
rect 53012 44140 53064 44160
rect 53064 44140 53066 44160
rect 53010 44104 53066 44140
rect 52366 41656 52422 41712
rect 52366 41384 52422 41440
rect 52366 40296 52422 40352
rect 52090 38956 52146 38992
rect 52090 38936 52092 38956
rect 52092 38936 52144 38956
rect 52144 38936 52146 38956
rect 52182 38120 52238 38176
rect 52366 35128 52422 35184
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50066 32408 50122 32464
rect 36266 23840 36322 23896
rect 36266 19796 36268 19816
rect 36268 19796 36320 19816
rect 36320 19796 36322 19816
rect 36266 19760 36322 19796
rect 36082 17484 36084 17504
rect 36084 17484 36136 17504
rect 36136 17484 36138 17504
rect 36082 17448 36138 17484
rect 36910 22072 36966 22128
rect 38566 22752 38622 22808
rect 37186 19488 37242 19544
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34978 10004 34980 10024
rect 34980 10004 35032 10024
rect 35032 10004 35034 10024
rect 34978 9968 35034 10004
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34518 3984 34574 4040
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 36082 11056 36138 11112
rect 35898 8608 35954 8664
rect 37646 21392 37702 21448
rect 37462 20032 37518 20088
rect 37554 19216 37610 19272
rect 36910 15952 36966 16008
rect 36726 13096 36782 13152
rect 37278 15000 37334 15056
rect 37462 14884 37518 14920
rect 37462 14864 37464 14884
rect 37464 14864 37516 14884
rect 37516 14864 37518 14884
rect 38106 19896 38162 19952
rect 38106 18264 38162 18320
rect 37830 17720 37886 17776
rect 37922 17448 37978 17504
rect 37830 16088 37886 16144
rect 38290 19252 38292 19272
rect 38292 19252 38344 19272
rect 38344 19252 38346 19272
rect 38290 19216 38346 19252
rect 38290 18708 38292 18728
rect 38292 18708 38344 18728
rect 38344 18708 38346 18728
rect 38290 18672 38346 18708
rect 38290 18128 38346 18184
rect 38658 22208 38714 22264
rect 38750 20868 38806 20904
rect 38750 20848 38752 20868
rect 38752 20848 38804 20868
rect 38804 20848 38806 20868
rect 38474 19760 38530 19816
rect 38566 18264 38622 18320
rect 39302 18164 39304 18184
rect 39304 18164 39356 18184
rect 39356 18164 39358 18184
rect 39302 18128 39358 18164
rect 36450 11228 36452 11248
rect 36452 11228 36504 11248
rect 36504 11228 36506 11248
rect 36450 11192 36506 11228
rect 36818 9968 36874 10024
rect 36726 8916 36728 8936
rect 36728 8916 36780 8936
rect 36780 8916 36782 8936
rect 36726 8880 36782 8916
rect 37186 10648 37242 10704
rect 37738 12300 37794 12336
rect 37738 12280 37740 12300
rect 37740 12280 37792 12300
rect 37792 12280 37794 12300
rect 38290 15272 38346 15328
rect 38198 13640 38254 13696
rect 38750 14340 38806 14376
rect 38750 14320 38752 14340
rect 38752 14320 38804 14340
rect 38804 14320 38806 14340
rect 38750 14048 38806 14104
rect 39394 16788 39450 16824
rect 39394 16768 39396 16788
rect 39396 16768 39448 16788
rect 39448 16768 39450 16788
rect 39394 15408 39450 15464
rect 39118 14048 39174 14104
rect 38566 10784 38622 10840
rect 39026 13368 39082 13424
rect 40130 19488 40186 19544
rect 41510 19488 41566 19544
rect 40498 18164 40500 18184
rect 40500 18164 40552 18184
rect 40552 18164 40554 18184
rect 40498 18128 40554 18164
rect 41694 18264 41750 18320
rect 40222 17584 40278 17640
rect 40866 16768 40922 16824
rect 40406 16496 40462 16552
rect 40222 13776 40278 13832
rect 40038 13368 40094 13424
rect 40038 12552 40094 12608
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 40866 13912 40922 13968
rect 41234 16788 41290 16824
rect 41234 16768 41236 16788
rect 41236 16768 41288 16788
rect 41288 16768 41290 16788
rect 41510 16788 41566 16824
rect 41510 16768 41512 16788
rect 41512 16768 41564 16788
rect 41564 16768 41566 16788
rect 41602 15816 41658 15872
rect 41418 15564 41474 15600
rect 41418 15544 41420 15564
rect 41420 15544 41472 15564
rect 41472 15544 41474 15564
rect 41418 14048 41474 14104
rect 41510 13676 41512 13696
rect 41512 13676 41564 13696
rect 41564 13676 41566 13696
rect 41510 13640 41566 13676
rect 41970 14320 42026 14376
rect 42522 16532 42524 16552
rect 42524 16532 42576 16552
rect 42576 16532 42578 16552
rect 42522 16496 42578 16532
rect 42614 15852 42616 15872
rect 42616 15852 42668 15872
rect 42668 15852 42670 15872
rect 42614 15816 42670 15852
rect 43350 22228 43406 22264
rect 43350 22208 43352 22228
rect 43352 22208 43404 22228
rect 43404 22208 43406 22228
rect 43994 20848 44050 20904
rect 42982 15408 43038 15464
rect 43718 15972 43774 16008
rect 43718 15952 43720 15972
rect 43720 15952 43772 15972
rect 43772 15952 43774 15972
rect 44454 15544 44510 15600
rect 46938 12280 46994 12336
rect 49698 11736 49754 11792
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 52918 43288 52974 43344
rect 53010 41112 53066 41168
rect 53562 46008 53618 46064
rect 53654 45600 53710 45656
rect 53746 45484 53802 45520
rect 53746 45464 53748 45484
rect 53748 45464 53800 45484
rect 53800 45464 53802 45484
rect 53470 44920 53526 44976
rect 53378 44376 53434 44432
rect 53562 43832 53618 43888
rect 53654 43560 53710 43616
rect 53470 43016 53526 43072
rect 53746 42880 53802 42936
rect 53746 42764 53802 42800
rect 53746 42744 53748 42764
rect 53748 42744 53800 42764
rect 53800 42744 53802 42764
rect 53654 42472 53710 42528
rect 53470 42200 53526 42256
rect 53470 41928 53526 41984
rect 53654 40840 53710 40896
rect 53470 40568 53526 40624
rect 52918 39752 52974 39808
rect 53010 38936 53066 38992
rect 53010 38700 53012 38720
rect 53012 38700 53064 38720
rect 53064 38700 53066 38720
rect 53010 38664 53066 38700
rect 53010 37612 53012 37632
rect 53012 37612 53064 37632
rect 53064 37612 53066 37632
rect 53010 37576 53066 37612
rect 53654 39480 53710 39536
rect 53562 38392 53618 38448
rect 53470 37848 53526 37904
rect 53378 37304 53434 37360
rect 53010 37032 53066 37088
rect 53470 36216 53526 36272
rect 53746 36760 53802 36816
rect 53654 36488 53710 36544
rect 53562 35944 53618 36000
rect 53470 35672 53526 35728
rect 53470 35400 53526 35456
rect 53010 34312 53066 34368
rect 53470 34856 53526 34912
rect 53562 34584 53618 34640
rect 53286 34040 53342 34096
rect 54390 49272 54446 49328
rect 54298 48184 54354 48240
rect 54482 47368 54538 47424
rect 54390 40024 54446 40080
rect 54298 39208 54354 39264
rect 54298 33260 54300 33280
rect 54300 33260 54352 33280
rect 54352 33260 54354 33280
rect 54298 33224 54354 33260
rect 54298 32408 54354 32464
rect 54298 31592 54354 31648
rect 54298 30776 54354 30832
rect 54206 29996 54208 30016
rect 54208 29996 54260 30016
rect 54260 29996 54262 30016
rect 54206 29960 54262 29996
rect 54206 29688 54262 29744
rect 54206 29144 54262 29200
rect 54206 28908 54208 28928
rect 54208 28908 54260 28928
rect 54260 28908 54262 28928
rect 54206 28872 54262 28908
rect 54206 28328 54262 28384
rect 53470 28056 53526 28112
rect 53470 27512 53526 27568
rect 53470 26968 53526 27024
rect 53562 26424 53618 26480
rect 53562 26152 53618 26208
rect 53562 25608 53618 25664
rect 53470 25336 53526 25392
rect 53470 25100 53472 25120
rect 53472 25100 53524 25120
rect 53524 25100 53526 25120
rect 53470 25064 53526 25100
rect 53470 24248 53526 24304
rect 53562 23196 53564 23216
rect 53564 23196 53616 23216
rect 53616 23196 53618 23216
rect 53562 23160 53618 23196
rect 53286 21528 53342 21584
rect 53470 21528 53526 21584
rect 53562 20748 53564 20768
rect 53564 20748 53616 20768
rect 53616 20748 53618 20768
rect 53562 20712 53618 20748
rect 53286 20460 53342 20496
rect 53286 20440 53288 20460
rect 53288 20440 53340 20460
rect 53340 20440 53342 20460
rect 53562 19932 53564 19952
rect 53564 19932 53616 19952
rect 53616 19932 53618 19952
rect 53562 19896 53618 19932
rect 53470 18264 53526 18320
rect 53286 16632 53342 16688
rect 53562 16668 53564 16688
rect 53564 16668 53616 16688
rect 53616 16668 53618 16688
rect 53562 16632 53618 16668
rect 54206 27240 54262 27296
rect 54206 26696 54262 26752
rect 54206 25880 54262 25936
rect 53470 15000 53526 15056
rect 54206 24792 54262 24848
rect 54206 23976 54262 24032
rect 54206 23432 54262 23488
rect 54206 22616 54262 22672
rect 54206 22344 54262 22400
rect 54022 21956 54078 21992
rect 54022 21936 54024 21956
rect 54024 21936 54076 21956
rect 54076 21936 54078 21956
rect 54206 21800 54262 21856
rect 54206 21020 54208 21040
rect 54208 21020 54260 21040
rect 54260 21020 54262 21040
rect 54206 20984 54262 21020
rect 54206 20712 54262 20768
rect 54206 20168 54262 20224
rect 54206 19352 54262 19408
rect 54206 19116 54208 19136
rect 54208 19116 54260 19136
rect 54260 19116 54262 19136
rect 54206 19080 54262 19116
rect 54206 18536 54262 18592
rect 54206 17756 54208 17776
rect 54208 17756 54260 17776
rect 54260 17756 54262 17776
rect 54206 17720 54262 17756
rect 54206 17484 54208 17504
rect 54208 17484 54260 17504
rect 54260 17484 54262 17504
rect 54206 17448 54262 17484
rect 54206 16904 54262 16960
rect 54206 16088 54262 16144
rect 54206 15816 54262 15872
rect 54206 15272 54262 15328
rect 54022 14864 54078 14920
rect 54206 14492 54208 14512
rect 54208 14492 54260 14512
rect 54260 14492 54262 14512
rect 54206 14456 54262 14492
rect 54206 14220 54208 14240
rect 54208 14220 54260 14240
rect 54260 14220 54262 14240
rect 54206 14184 54262 14220
rect 53562 13404 53564 13424
rect 53564 13404 53616 13424
rect 53616 13404 53618 13424
rect 53562 13368 53618 13404
rect 54206 13640 54262 13696
rect 54206 12824 54262 12880
rect 54206 12552 54262 12608
rect 54206 12008 54262 12064
rect 53470 11736 53526 11792
rect 54206 11228 54208 11248
rect 54208 11228 54260 11248
rect 54260 11228 54262 11248
rect 54206 11192 54262 11228
rect 54206 10956 54208 10976
rect 54208 10956 54260 10976
rect 54260 10956 54262 10976
rect 54206 10920 54262 10956
rect 54206 10376 54262 10432
rect 53470 10140 53472 10160
rect 53472 10140 53524 10160
rect 53524 10140 53526 10160
rect 53470 10104 53526 10140
rect 54206 9560 54262 9616
rect 53562 9288 53618 9344
rect 52182 7928 52238 7984
rect 53470 8492 53526 8528
rect 53470 8472 53472 8492
rect 53472 8472 53524 8492
rect 53524 8472 53526 8492
rect 54206 8744 54262 8800
rect 53378 7656 53434 7712
rect 52274 7384 52330 7440
rect 54114 7112 54170 7168
rect 54390 6840 54446 6896
rect 51262 6568 51318 6624
rect 51814 2372 51870 2408
rect 51814 2352 51816 2372
rect 51816 2352 51868 2372
rect 51868 2352 51870 2372
<< metal3 >>
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 0 52730 800 52760
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 2773 52730 2839 52733
rect 0 52728 2839 52730
rect 0 52672 2778 52728
rect 2834 52672 2839 52728
rect 0 52670 2839 52672
rect 0 52640 800 52670
rect 2773 52667 2839 52670
rect 27838 52532 27844 52596
rect 27908 52594 27914 52596
rect 51993 52594 52059 52597
rect 27908 52592 52059 52594
rect 27908 52536 51998 52592
rect 52054 52536 52059 52592
rect 27908 52534 52059 52536
rect 27908 52532 27914 52534
rect 51993 52531 52059 52534
rect 19570 52256 19886 52257
rect 0 52186 800 52216
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 1485 52186 1551 52189
rect 0 52184 1551 52186
rect 0 52128 1490 52184
rect 1546 52128 1551 52184
rect 0 52126 1551 52128
rect 0 52096 800 52126
rect 1485 52123 1551 52126
rect 4210 51712 4526 51713
rect 0 51642 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 1669 51642 1735 51645
rect 0 51640 1735 51642
rect 0 51584 1674 51640
rect 1730 51584 1735 51640
rect 0 51582 1735 51584
rect 0 51552 800 51582
rect 1669 51579 1735 51582
rect 19570 51168 19886 51169
rect 0 51098 800 51128
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 1669 51098 1735 51101
rect 0 51096 1735 51098
rect 0 51040 1674 51096
rect 1730 51040 1735 51096
rect 0 51038 1735 51040
rect 0 51008 800 51038
rect 1669 51035 1735 51038
rect 4210 50624 4526 50625
rect 0 50554 800 50584
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 2773 50554 2839 50557
rect 0 50552 2839 50554
rect 0 50496 2778 50552
rect 2834 50496 2839 50552
rect 0 50494 2839 50496
rect 0 50464 800 50494
rect 2773 50491 2839 50494
rect 19570 50080 19886 50081
rect 0 50010 800 50040
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 2773 50010 2839 50013
rect 0 50008 2839 50010
rect 0 49952 2778 50008
rect 2834 49952 2839 50008
rect 0 49950 2839 49952
rect 0 49920 800 49950
rect 2773 49947 2839 49950
rect 4210 49536 4526 49537
rect 0 49466 800 49496
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 1669 49466 1735 49469
rect 0 49464 1735 49466
rect 0 49408 1674 49464
rect 1730 49408 1735 49464
rect 0 49406 1735 49408
rect 0 49376 800 49406
rect 1669 49403 1735 49406
rect 54385 49330 54451 49333
rect 55200 49330 56000 49360
rect 54385 49328 56000 49330
rect 54385 49272 54390 49328
rect 54446 49272 56000 49328
rect 54385 49270 56000 49272
rect 54385 49267 54451 49270
rect 55200 49240 56000 49270
rect 53465 49058 53531 49061
rect 55200 49058 56000 49088
rect 53465 49056 56000 49058
rect 53465 49000 53470 49056
rect 53526 49000 56000 49056
rect 53465 48998 56000 49000
rect 53465 48995 53531 48998
rect 19570 48992 19886 48993
rect 0 48922 800 48952
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 55200 48968 56000 48998
rect 50290 48927 50606 48928
rect 2773 48922 2839 48925
rect 0 48920 2839 48922
rect 0 48864 2778 48920
rect 2834 48864 2839 48920
rect 0 48862 2839 48864
rect 0 48832 800 48862
rect 2773 48859 2839 48862
rect 53557 48786 53623 48789
rect 55200 48786 56000 48816
rect 53557 48784 56000 48786
rect 53557 48728 53562 48784
rect 53618 48728 56000 48784
rect 53557 48726 56000 48728
rect 53557 48723 53623 48726
rect 55200 48696 56000 48726
rect 53649 48514 53715 48517
rect 55200 48514 56000 48544
rect 53649 48512 56000 48514
rect 53649 48456 53654 48512
rect 53710 48456 56000 48512
rect 53649 48454 56000 48456
rect 53649 48451 53715 48454
rect 4210 48448 4526 48449
rect 0 48378 800 48408
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 55200 48424 56000 48454
rect 34930 48383 35246 48384
rect 2773 48378 2839 48381
rect 0 48376 2839 48378
rect 0 48320 2778 48376
rect 2834 48320 2839 48376
rect 0 48318 2839 48320
rect 0 48288 800 48318
rect 2773 48315 2839 48318
rect 54293 48242 54359 48245
rect 55200 48242 56000 48272
rect 54293 48240 56000 48242
rect 54293 48184 54298 48240
rect 54354 48184 56000 48240
rect 54293 48182 56000 48184
rect 54293 48179 54359 48182
rect 55200 48152 56000 48182
rect 52361 47970 52427 47973
rect 55200 47970 56000 48000
rect 52361 47968 56000 47970
rect 52361 47912 52366 47968
rect 52422 47912 56000 47968
rect 52361 47910 56000 47912
rect 52361 47907 52427 47910
rect 19570 47904 19886 47905
rect 0 47834 800 47864
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 55200 47880 56000 47910
rect 50290 47839 50606 47840
rect 2773 47834 2839 47837
rect 0 47832 2839 47834
rect 0 47776 2778 47832
rect 2834 47776 2839 47832
rect 0 47774 2839 47776
rect 0 47744 800 47774
rect 2773 47771 2839 47774
rect 53097 47698 53163 47701
rect 55200 47698 56000 47728
rect 53097 47696 56000 47698
rect 53097 47640 53102 47696
rect 53158 47640 56000 47696
rect 53097 47638 56000 47640
rect 53097 47635 53163 47638
rect 55200 47608 56000 47638
rect 54477 47426 54543 47429
rect 55200 47426 56000 47456
rect 54477 47424 56000 47426
rect 54477 47368 54482 47424
rect 54538 47368 56000 47424
rect 54477 47366 56000 47368
rect 54477 47363 54543 47366
rect 4210 47360 4526 47361
rect 0 47290 800 47320
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 55200 47336 56000 47366
rect 34930 47295 35246 47296
rect 2773 47290 2839 47293
rect 0 47288 2839 47290
rect 0 47232 2778 47288
rect 2834 47232 2839 47288
rect 0 47230 2839 47232
rect 0 47200 800 47230
rect 2773 47227 2839 47230
rect 51441 47154 51507 47157
rect 55200 47154 56000 47184
rect 51441 47152 56000 47154
rect 51441 47096 51446 47152
rect 51502 47096 56000 47152
rect 51441 47094 56000 47096
rect 51441 47091 51507 47094
rect 55200 47064 56000 47094
rect 33317 47018 33383 47021
rect 35617 47018 35683 47021
rect 33317 47016 35683 47018
rect 33317 46960 33322 47016
rect 33378 46960 35622 47016
rect 35678 46960 35683 47016
rect 33317 46958 35683 46960
rect 33317 46955 33383 46958
rect 35617 46955 35683 46958
rect 50889 47018 50955 47021
rect 51625 47018 51691 47021
rect 51809 47018 51875 47021
rect 50889 47016 51875 47018
rect 50889 46960 50894 47016
rect 50950 46960 51630 47016
rect 51686 46960 51814 47016
rect 51870 46960 51875 47016
rect 50889 46958 51875 46960
rect 50889 46955 50955 46958
rect 51625 46955 51691 46958
rect 51809 46955 51875 46958
rect 52177 46882 52243 46885
rect 55200 46882 56000 46912
rect 52177 46880 56000 46882
rect 52177 46824 52182 46880
rect 52238 46824 56000 46880
rect 52177 46822 56000 46824
rect 52177 46819 52243 46822
rect 19570 46816 19886 46817
rect 0 46746 800 46776
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 55200 46792 56000 46822
rect 50290 46751 50606 46752
rect 2773 46746 2839 46749
rect 0 46744 2839 46746
rect 0 46688 2778 46744
rect 2834 46688 2839 46744
rect 0 46686 2839 46688
rect 0 46656 800 46686
rect 2773 46683 2839 46686
rect 52637 46610 52703 46613
rect 55200 46610 56000 46640
rect 52637 46608 56000 46610
rect 52637 46552 52642 46608
rect 52698 46552 56000 46608
rect 52637 46550 56000 46552
rect 52637 46547 52703 46550
rect 55200 46520 56000 46550
rect 53005 46338 53071 46341
rect 55200 46338 56000 46368
rect 53005 46336 56000 46338
rect 53005 46280 53010 46336
rect 53066 46280 56000 46336
rect 53005 46278 56000 46280
rect 53005 46275 53071 46278
rect 4210 46272 4526 46273
rect 0 46202 800 46232
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 55200 46248 56000 46278
rect 34930 46207 35246 46208
rect 2773 46202 2839 46205
rect 0 46200 2839 46202
rect 0 46144 2778 46200
rect 2834 46144 2839 46200
rect 0 46142 2839 46144
rect 0 46112 800 46142
rect 2773 46139 2839 46142
rect 53557 46066 53623 46069
rect 55200 46066 56000 46096
rect 53557 46064 56000 46066
rect 53557 46008 53562 46064
rect 53618 46008 56000 46064
rect 53557 46006 56000 46008
rect 53557 46003 53623 46006
rect 55200 45976 56000 46006
rect 52177 45794 52243 45797
rect 55200 45794 56000 45824
rect 52177 45792 56000 45794
rect 52177 45736 52182 45792
rect 52238 45736 56000 45792
rect 52177 45734 56000 45736
rect 52177 45731 52243 45734
rect 19570 45728 19886 45729
rect 0 45658 800 45688
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 55200 45704 56000 45734
rect 50290 45663 50606 45664
rect 2773 45658 2839 45661
rect 0 45656 2839 45658
rect 0 45600 2778 45656
rect 2834 45600 2839 45656
rect 0 45598 2839 45600
rect 0 45568 800 45598
rect 2773 45595 2839 45598
rect 53649 45658 53715 45661
rect 53649 45656 54034 45658
rect 53649 45600 53654 45656
rect 53710 45600 54034 45656
rect 53649 45598 54034 45600
rect 53649 45595 53715 45598
rect 27102 45460 27108 45524
rect 27172 45522 27178 45524
rect 53741 45522 53807 45525
rect 27172 45520 53807 45522
rect 27172 45464 53746 45520
rect 53802 45464 53807 45520
rect 27172 45462 53807 45464
rect 53974 45522 54034 45598
rect 55200 45522 56000 45552
rect 53974 45462 56000 45522
rect 27172 45460 27178 45462
rect 53741 45459 53807 45462
rect 55200 45432 56000 45462
rect 53005 45250 53071 45253
rect 55200 45250 56000 45280
rect 53005 45248 56000 45250
rect 53005 45192 53010 45248
rect 53066 45192 56000 45248
rect 53005 45190 56000 45192
rect 53005 45187 53071 45190
rect 4210 45184 4526 45185
rect 0 45114 800 45144
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 55200 45160 56000 45190
rect 34930 45119 35246 45120
rect 2773 45114 2839 45117
rect 0 45112 2839 45114
rect 0 45056 2778 45112
rect 2834 45056 2839 45112
rect 0 45054 2839 45056
rect 0 45024 800 45054
rect 2773 45051 2839 45054
rect 31334 44916 31340 44980
rect 31404 44978 31410 44980
rect 52453 44978 52519 44981
rect 31404 44976 52519 44978
rect 31404 44920 52458 44976
rect 52514 44920 52519 44976
rect 31404 44918 52519 44920
rect 31404 44916 31410 44918
rect 52453 44915 52519 44918
rect 53465 44978 53531 44981
rect 55200 44978 56000 45008
rect 53465 44976 56000 44978
rect 53465 44920 53470 44976
rect 53526 44920 56000 44976
rect 53465 44918 56000 44920
rect 53465 44915 53531 44918
rect 55200 44888 56000 44918
rect 52177 44706 52243 44709
rect 55200 44706 56000 44736
rect 52177 44704 56000 44706
rect 52177 44648 52182 44704
rect 52238 44648 56000 44704
rect 52177 44646 56000 44648
rect 52177 44643 52243 44646
rect 19570 44640 19886 44641
rect 0 44570 800 44600
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 55200 44616 56000 44646
rect 50290 44575 50606 44576
rect 2773 44570 2839 44573
rect 0 44568 2839 44570
rect 0 44512 2778 44568
rect 2834 44512 2839 44568
rect 0 44510 2839 44512
rect 0 44480 800 44510
rect 2773 44507 2839 44510
rect 53373 44434 53439 44437
rect 55200 44434 56000 44464
rect 53373 44432 56000 44434
rect 53373 44376 53378 44432
rect 53434 44376 56000 44432
rect 53373 44374 56000 44376
rect 53373 44371 53439 44374
rect 55200 44344 56000 44374
rect 2497 44298 2563 44301
rect 32305 44298 32371 44301
rect 2497 44296 32371 44298
rect 2497 44240 2502 44296
rect 2558 44240 32310 44296
rect 32366 44240 32371 44296
rect 2497 44238 32371 44240
rect 2497 44235 2563 44238
rect 32305 44235 32371 44238
rect 53005 44162 53071 44165
rect 55200 44162 56000 44192
rect 53005 44160 56000 44162
rect 53005 44104 53010 44160
rect 53066 44104 56000 44160
rect 53005 44102 56000 44104
rect 53005 44099 53071 44102
rect 4210 44096 4526 44097
rect 0 44026 800 44056
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 55200 44072 56000 44102
rect 34930 44031 35246 44032
rect 2773 44026 2839 44029
rect 0 44024 2839 44026
rect 0 43968 2778 44024
rect 2834 43968 2839 44024
rect 0 43966 2839 43968
rect 0 43936 800 43966
rect 2773 43963 2839 43966
rect 53557 43890 53623 43893
rect 55200 43890 56000 43920
rect 53557 43888 56000 43890
rect 53557 43832 53562 43888
rect 53618 43832 56000 43888
rect 53557 43830 56000 43832
rect 53557 43827 53623 43830
rect 55200 43800 56000 43830
rect 53649 43618 53715 43621
rect 55200 43618 56000 43648
rect 53649 43616 56000 43618
rect 53649 43560 53654 43616
rect 53710 43560 56000 43616
rect 53649 43558 56000 43560
rect 53649 43555 53715 43558
rect 19570 43552 19886 43553
rect 0 43482 800 43512
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 55200 43528 56000 43558
rect 50290 43487 50606 43488
rect 2773 43482 2839 43485
rect 0 43480 2839 43482
rect 0 43424 2778 43480
rect 2834 43424 2839 43480
rect 0 43422 2839 43424
rect 0 43392 800 43422
rect 2773 43419 2839 43422
rect 52913 43346 52979 43349
rect 55200 43346 56000 43376
rect 52913 43344 56000 43346
rect 52913 43288 52918 43344
rect 52974 43288 56000 43344
rect 52913 43286 56000 43288
rect 52913 43283 52979 43286
rect 55200 43256 56000 43286
rect 11605 43210 11671 43213
rect 29361 43210 29427 43213
rect 29637 43210 29703 43213
rect 11605 43208 29703 43210
rect 11605 43152 11610 43208
rect 11666 43152 29366 43208
rect 29422 43152 29642 43208
rect 29698 43152 29703 43208
rect 11605 43150 29703 43152
rect 11605 43147 11671 43150
rect 29361 43147 29427 43150
rect 29637 43147 29703 43150
rect 53465 43074 53531 43077
rect 55200 43074 56000 43104
rect 53465 43072 56000 43074
rect 53465 43016 53470 43072
rect 53526 43016 56000 43072
rect 53465 43014 56000 43016
rect 53465 43011 53531 43014
rect 4210 43008 4526 43009
rect 0 42938 800 42968
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 55200 42984 56000 43014
rect 34930 42943 35246 42944
rect 2773 42938 2839 42941
rect 0 42936 2839 42938
rect 0 42880 2778 42936
rect 2834 42880 2839 42936
rect 0 42878 2839 42880
rect 0 42848 800 42878
rect 2773 42875 2839 42878
rect 53741 42938 53807 42941
rect 53741 42936 54034 42938
rect 53741 42880 53746 42936
rect 53802 42880 54034 42936
rect 53741 42878 54034 42880
rect 53741 42875 53807 42878
rect 30281 42802 30347 42805
rect 31017 42802 31083 42805
rect 53741 42802 53807 42805
rect 30281 42800 53807 42802
rect 30281 42744 30286 42800
rect 30342 42744 31022 42800
rect 31078 42744 53746 42800
rect 53802 42744 53807 42800
rect 30281 42742 53807 42744
rect 53974 42802 54034 42878
rect 55200 42802 56000 42832
rect 53974 42742 56000 42802
rect 30281 42739 30347 42742
rect 31017 42739 31083 42742
rect 53741 42739 53807 42742
rect 55200 42712 56000 42742
rect 53649 42530 53715 42533
rect 55200 42530 56000 42560
rect 53649 42528 56000 42530
rect 53649 42472 53654 42528
rect 53710 42472 56000 42528
rect 53649 42470 56000 42472
rect 53649 42467 53715 42470
rect 19570 42464 19886 42465
rect 0 42394 800 42424
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 55200 42440 56000 42470
rect 50290 42399 50606 42400
rect 2773 42394 2839 42397
rect 0 42392 2839 42394
rect 0 42336 2778 42392
rect 2834 42336 2839 42392
rect 0 42334 2839 42336
rect 0 42304 800 42334
rect 2773 42331 2839 42334
rect 30373 42258 30439 42261
rect 34697 42258 34763 42261
rect 30373 42256 34763 42258
rect 30373 42200 30378 42256
rect 30434 42200 34702 42256
rect 34758 42200 34763 42256
rect 30373 42198 34763 42200
rect 30373 42195 30439 42198
rect 34697 42195 34763 42198
rect 53465 42258 53531 42261
rect 55200 42258 56000 42288
rect 53465 42256 56000 42258
rect 53465 42200 53470 42256
rect 53526 42200 56000 42256
rect 53465 42198 56000 42200
rect 53465 42195 53531 42198
rect 55200 42168 56000 42198
rect 24945 41986 25011 41989
rect 27521 41986 27587 41989
rect 28809 41986 28875 41989
rect 24945 41984 27587 41986
rect 24945 41928 24950 41984
rect 25006 41928 27526 41984
rect 27582 41928 27587 41984
rect 24945 41926 27587 41928
rect 24945 41923 25011 41926
rect 27521 41923 27587 41926
rect 27984 41984 28875 41986
rect 27984 41928 28814 41984
rect 28870 41928 28875 41984
rect 27984 41926 28875 41928
rect 4210 41920 4526 41921
rect 0 41850 800 41880
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 27984 41853 28044 41926
rect 28809 41923 28875 41926
rect 53465 41986 53531 41989
rect 55200 41986 56000 42016
rect 53465 41984 56000 41986
rect 53465 41928 53470 41984
rect 53526 41928 56000 41984
rect 53465 41926 56000 41928
rect 53465 41923 53531 41926
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 55200 41896 56000 41926
rect 34930 41855 35246 41856
rect 2773 41850 2839 41853
rect 0 41848 2839 41850
rect 0 41792 2778 41848
rect 2834 41792 2839 41848
rect 0 41790 2839 41792
rect 0 41760 800 41790
rect 2773 41787 2839 41790
rect 27981 41848 28047 41853
rect 27981 41792 27986 41848
rect 28042 41792 28047 41848
rect 27981 41787 28047 41792
rect 28717 41850 28783 41853
rect 33317 41850 33383 41853
rect 34329 41850 34395 41853
rect 28717 41848 29010 41850
rect 28717 41792 28722 41848
rect 28778 41792 29010 41848
rect 28717 41790 29010 41792
rect 28717 41787 28783 41790
rect 26049 41714 26115 41717
rect 27981 41714 28047 41717
rect 26049 41712 28047 41714
rect 26049 41656 26054 41712
rect 26110 41656 27986 41712
rect 28042 41656 28047 41712
rect 26049 41654 28047 41656
rect 26049 41651 26115 41654
rect 27981 41651 28047 41654
rect 28257 41714 28323 41717
rect 28758 41714 28764 41716
rect 28257 41712 28764 41714
rect 28257 41656 28262 41712
rect 28318 41656 28764 41712
rect 28257 41654 28764 41656
rect 28257 41651 28323 41654
rect 28758 41652 28764 41654
rect 28828 41652 28834 41716
rect 25814 41516 25820 41580
rect 25884 41578 25890 41580
rect 26509 41578 26575 41581
rect 25884 41576 26575 41578
rect 25884 41520 26514 41576
rect 26570 41520 26575 41576
rect 25884 41518 26575 41520
rect 25884 41516 25890 41518
rect 26509 41515 26575 41518
rect 28717 41578 28783 41581
rect 28950 41578 29010 41790
rect 33317 41848 34395 41850
rect 33317 41792 33322 41848
rect 33378 41792 34334 41848
rect 34390 41792 34395 41848
rect 33317 41790 34395 41792
rect 33317 41787 33383 41790
rect 34329 41787 34395 41790
rect 30097 41714 30163 41717
rect 31477 41714 31543 41717
rect 35525 41714 35591 41717
rect 30097 41712 35591 41714
rect 30097 41656 30102 41712
rect 30158 41656 31482 41712
rect 31538 41656 35530 41712
rect 35586 41656 35591 41712
rect 30097 41654 35591 41656
rect 30097 41651 30163 41654
rect 31477 41651 31543 41654
rect 35525 41651 35591 41654
rect 52361 41714 52427 41717
rect 55200 41714 56000 41744
rect 52361 41712 56000 41714
rect 52361 41656 52366 41712
rect 52422 41656 56000 41712
rect 52361 41654 56000 41656
rect 52361 41651 52427 41654
rect 55200 41624 56000 41654
rect 28717 41576 29010 41578
rect 28717 41520 28722 41576
rect 28778 41520 29010 41576
rect 28717 41518 29010 41520
rect 32581 41578 32647 41581
rect 35617 41578 35683 41581
rect 32581 41576 35683 41578
rect 32581 41520 32586 41576
rect 32642 41520 35622 41576
rect 35678 41520 35683 41576
rect 32581 41518 35683 41520
rect 28717 41515 28783 41518
rect 32581 41515 32647 41518
rect 35617 41515 35683 41518
rect 27981 41442 28047 41445
rect 28533 41442 28599 41445
rect 27981 41440 28599 41442
rect 27981 41384 27986 41440
rect 28042 41384 28538 41440
rect 28594 41384 28599 41440
rect 27981 41382 28599 41384
rect 27981 41379 28047 41382
rect 28533 41379 28599 41382
rect 52361 41442 52427 41445
rect 55200 41442 56000 41472
rect 52361 41440 56000 41442
rect 52361 41384 52366 41440
rect 52422 41384 56000 41440
rect 52361 41382 56000 41384
rect 52361 41379 52427 41382
rect 19570 41376 19886 41377
rect 0 41306 800 41336
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 55200 41352 56000 41382
rect 50290 41311 50606 41312
rect 2773 41306 2839 41309
rect 0 41304 2839 41306
rect 0 41248 2778 41304
rect 2834 41248 2839 41304
rect 0 41246 2839 41248
rect 0 41216 800 41246
rect 2773 41243 2839 41246
rect 26233 41306 26299 41309
rect 27429 41306 27495 41309
rect 26233 41304 27495 41306
rect 26233 41248 26238 41304
rect 26294 41248 27434 41304
rect 27490 41248 27495 41304
rect 26233 41246 27495 41248
rect 26233 41243 26299 41246
rect 27429 41243 27495 41246
rect 27705 41306 27771 41309
rect 27838 41306 27844 41308
rect 27705 41304 27844 41306
rect 27705 41248 27710 41304
rect 27766 41248 27844 41304
rect 27705 41246 27844 41248
rect 27705 41243 27771 41246
rect 27838 41244 27844 41246
rect 27908 41244 27914 41308
rect 2037 41170 2103 41173
rect 32765 41170 32831 41173
rect 35249 41170 35315 41173
rect 2037 41168 35315 41170
rect 2037 41112 2042 41168
rect 2098 41112 32770 41168
rect 32826 41112 35254 41168
rect 35310 41112 35315 41168
rect 2037 41110 35315 41112
rect 2037 41107 2103 41110
rect 32765 41107 32831 41110
rect 35249 41107 35315 41110
rect 53005 41170 53071 41173
rect 55200 41170 56000 41200
rect 53005 41168 56000 41170
rect 53005 41112 53010 41168
rect 53066 41112 56000 41168
rect 53005 41110 56000 41112
rect 53005 41107 53071 41110
rect 55200 41080 56000 41110
rect 29085 40898 29151 40901
rect 29310 40898 29316 40900
rect 29085 40896 29316 40898
rect 29085 40840 29090 40896
rect 29146 40840 29316 40896
rect 29085 40838 29316 40840
rect 29085 40835 29151 40838
rect 29310 40836 29316 40838
rect 29380 40836 29386 40900
rect 29453 40898 29519 40901
rect 32673 40898 32739 40901
rect 33593 40898 33659 40901
rect 29453 40896 33659 40898
rect 29453 40840 29458 40896
rect 29514 40840 32678 40896
rect 32734 40840 33598 40896
rect 33654 40840 33659 40896
rect 29453 40838 33659 40840
rect 29453 40835 29519 40838
rect 32673 40835 32739 40838
rect 33593 40835 33659 40838
rect 53649 40898 53715 40901
rect 55200 40898 56000 40928
rect 53649 40896 56000 40898
rect 53649 40840 53654 40896
rect 53710 40840 56000 40896
rect 53649 40838 56000 40840
rect 53649 40835 53715 40838
rect 4210 40832 4526 40833
rect 0 40762 800 40792
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 55200 40808 56000 40838
rect 34930 40767 35246 40768
rect 2773 40762 2839 40765
rect 0 40760 2839 40762
rect 0 40704 2778 40760
rect 2834 40704 2839 40760
rect 0 40702 2839 40704
rect 0 40672 800 40702
rect 2773 40699 2839 40702
rect 26141 40762 26207 40765
rect 27797 40762 27863 40765
rect 26141 40760 27863 40762
rect 26141 40704 26146 40760
rect 26202 40704 27802 40760
rect 27858 40704 27863 40760
rect 26141 40702 27863 40704
rect 26141 40699 26207 40702
rect 27797 40699 27863 40702
rect 26141 40626 26207 40629
rect 27521 40626 27587 40629
rect 28717 40626 28783 40629
rect 26141 40624 28783 40626
rect 26141 40568 26146 40624
rect 26202 40568 27526 40624
rect 27582 40568 28722 40624
rect 28778 40568 28783 40624
rect 26141 40566 28783 40568
rect 26141 40563 26207 40566
rect 27521 40563 27587 40566
rect 28717 40563 28783 40566
rect 53465 40626 53531 40629
rect 55200 40626 56000 40656
rect 53465 40624 56000 40626
rect 53465 40568 53470 40624
rect 53526 40568 56000 40624
rect 53465 40566 56000 40568
rect 53465 40563 53531 40566
rect 55200 40536 56000 40566
rect 25773 40490 25839 40493
rect 28073 40490 28139 40493
rect 25773 40488 28139 40490
rect 25773 40432 25778 40488
rect 25834 40432 28078 40488
rect 28134 40432 28139 40488
rect 25773 40430 28139 40432
rect 25773 40427 25839 40430
rect 28073 40427 28139 40430
rect 32581 40490 32647 40493
rect 34421 40490 34487 40493
rect 34605 40490 34671 40493
rect 32581 40488 34671 40490
rect 32581 40432 32586 40488
rect 32642 40432 34426 40488
rect 34482 40432 34610 40488
rect 34666 40432 34671 40488
rect 32581 40430 34671 40432
rect 32581 40427 32647 40430
rect 34421 40427 34487 40430
rect 34605 40427 34671 40430
rect 23381 40354 23447 40357
rect 28809 40354 28875 40357
rect 23381 40352 28875 40354
rect 23381 40296 23386 40352
rect 23442 40296 28814 40352
rect 28870 40296 28875 40352
rect 23381 40294 28875 40296
rect 23381 40291 23447 40294
rect 28809 40291 28875 40294
rect 52361 40354 52427 40357
rect 55200 40354 56000 40384
rect 52361 40352 56000 40354
rect 52361 40296 52366 40352
rect 52422 40296 56000 40352
rect 52361 40294 56000 40296
rect 52361 40291 52427 40294
rect 19570 40288 19886 40289
rect 0 40218 800 40248
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 55200 40264 56000 40294
rect 50290 40223 50606 40224
rect 2773 40218 2839 40221
rect 0 40216 2839 40218
rect 0 40160 2778 40216
rect 2834 40160 2839 40216
rect 0 40158 2839 40160
rect 0 40128 800 40158
rect 2773 40155 2839 40158
rect 27337 40218 27403 40221
rect 28533 40218 28599 40221
rect 27337 40216 28599 40218
rect 27337 40160 27342 40216
rect 27398 40160 28538 40216
rect 28594 40160 28599 40216
rect 27337 40158 28599 40160
rect 27337 40155 27403 40158
rect 28533 40155 28599 40158
rect 26417 40082 26483 40085
rect 26550 40082 26556 40084
rect 26417 40080 26556 40082
rect 26417 40024 26422 40080
rect 26478 40024 26556 40080
rect 26417 40022 26556 40024
rect 26417 40019 26483 40022
rect 26550 40020 26556 40022
rect 26620 40020 26626 40084
rect 31477 40082 31543 40085
rect 33961 40082 34027 40085
rect 31477 40080 34027 40082
rect 31477 40024 31482 40080
rect 31538 40024 33966 40080
rect 34022 40024 34027 40080
rect 31477 40022 34027 40024
rect 31477 40019 31543 40022
rect 33961 40019 34027 40022
rect 54385 40082 54451 40085
rect 55200 40082 56000 40112
rect 54385 40080 56000 40082
rect 54385 40024 54390 40080
rect 54446 40024 56000 40080
rect 54385 40022 56000 40024
rect 54385 40019 54451 40022
rect 55200 39992 56000 40022
rect 52913 39810 52979 39813
rect 55200 39810 56000 39840
rect 52913 39808 56000 39810
rect 52913 39752 52918 39808
rect 52974 39752 56000 39808
rect 52913 39750 56000 39752
rect 52913 39747 52979 39750
rect 4210 39744 4526 39745
rect 0 39674 800 39704
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 55200 39720 56000 39750
rect 34930 39679 35246 39680
rect 2773 39674 2839 39677
rect 0 39672 2839 39674
rect 0 39616 2778 39672
rect 2834 39616 2839 39672
rect 0 39614 2839 39616
rect 0 39584 800 39614
rect 2773 39611 2839 39614
rect 26877 39538 26943 39541
rect 28257 39538 28323 39541
rect 26877 39536 28323 39538
rect 26877 39480 26882 39536
rect 26938 39480 28262 39536
rect 28318 39480 28323 39536
rect 26877 39478 28323 39480
rect 26877 39475 26943 39478
rect 28257 39475 28323 39478
rect 53649 39538 53715 39541
rect 55200 39538 56000 39568
rect 53649 39536 56000 39538
rect 53649 39480 53654 39536
rect 53710 39480 56000 39536
rect 53649 39478 56000 39480
rect 53649 39475 53715 39478
rect 55200 39448 56000 39478
rect 54293 39266 54359 39269
rect 55200 39266 56000 39296
rect 54293 39264 56000 39266
rect 54293 39208 54298 39264
rect 54354 39208 56000 39264
rect 54293 39206 56000 39208
rect 54293 39203 54359 39206
rect 19570 39200 19886 39201
rect 0 39130 800 39160
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 55200 39176 56000 39206
rect 50290 39135 50606 39136
rect 2773 39130 2839 39133
rect 0 39128 2839 39130
rect 0 39072 2778 39128
rect 2834 39072 2839 39128
rect 0 39070 2839 39072
rect 0 39040 800 39070
rect 2773 39067 2839 39070
rect 24853 38994 24919 38997
rect 27061 38994 27127 38997
rect 27429 38994 27495 38997
rect 27613 38994 27679 38997
rect 24853 38992 27679 38994
rect 24853 38936 24858 38992
rect 24914 38936 27066 38992
rect 27122 38936 27434 38992
rect 27490 38936 27618 38992
rect 27674 38936 27679 38992
rect 24853 38934 27679 38936
rect 24853 38931 24919 38934
rect 27061 38931 27127 38934
rect 27429 38931 27495 38934
rect 27613 38931 27679 38934
rect 29310 38932 29316 38996
rect 29380 38994 29386 38996
rect 52085 38994 52151 38997
rect 29380 38992 52151 38994
rect 29380 38936 52090 38992
rect 52146 38936 52151 38992
rect 29380 38934 52151 38936
rect 29380 38932 29386 38934
rect 52085 38931 52151 38934
rect 53005 38994 53071 38997
rect 55200 38994 56000 39024
rect 53005 38992 56000 38994
rect 53005 38936 53010 38992
rect 53066 38936 56000 38992
rect 53005 38934 56000 38936
rect 53005 38931 53071 38934
rect 55200 38904 56000 38934
rect 26049 38858 26115 38861
rect 28073 38858 28139 38861
rect 26049 38856 28139 38858
rect 26049 38800 26054 38856
rect 26110 38800 28078 38856
rect 28134 38800 28139 38856
rect 26049 38798 28139 38800
rect 26049 38795 26115 38798
rect 28073 38795 28139 38798
rect 26785 38722 26851 38725
rect 26918 38722 26924 38724
rect 26785 38720 26924 38722
rect 26785 38664 26790 38720
rect 26846 38664 26924 38720
rect 26785 38662 26924 38664
rect 26785 38659 26851 38662
rect 26918 38660 26924 38662
rect 26988 38660 26994 38724
rect 29678 38660 29684 38724
rect 29748 38722 29754 38724
rect 29821 38722 29887 38725
rect 29748 38720 29887 38722
rect 29748 38664 29826 38720
rect 29882 38664 29887 38720
rect 29748 38662 29887 38664
rect 29748 38660 29754 38662
rect 29821 38659 29887 38662
rect 53005 38722 53071 38725
rect 55200 38722 56000 38752
rect 53005 38720 56000 38722
rect 53005 38664 53010 38720
rect 53066 38664 56000 38720
rect 53005 38662 56000 38664
rect 53005 38659 53071 38662
rect 4210 38656 4526 38657
rect 0 38586 800 38616
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 55200 38632 56000 38662
rect 34930 38591 35246 38592
rect 2773 38586 2839 38589
rect 0 38584 2839 38586
rect 0 38528 2778 38584
rect 2834 38528 2839 38584
rect 0 38526 2839 38528
rect 0 38496 800 38526
rect 2773 38523 2839 38526
rect 23473 38586 23539 38589
rect 27521 38586 27587 38589
rect 28993 38588 29059 38589
rect 23473 38584 27587 38586
rect 23473 38528 23478 38584
rect 23534 38528 27526 38584
rect 27582 38528 27587 38584
rect 23473 38526 27587 38528
rect 23473 38523 23539 38526
rect 27521 38523 27587 38526
rect 28942 38524 28948 38588
rect 29012 38586 29059 38588
rect 29012 38584 29104 38586
rect 29054 38528 29104 38584
rect 29012 38526 29104 38528
rect 29012 38524 29059 38526
rect 28993 38523 29059 38524
rect 24669 38450 24735 38453
rect 27153 38450 27219 38453
rect 28441 38450 28507 38453
rect 28993 38450 29059 38453
rect 24669 38448 28507 38450
rect 24669 38392 24674 38448
rect 24730 38392 27158 38448
rect 27214 38392 28446 38448
rect 28502 38392 28507 38448
rect 24669 38390 28507 38392
rect 24669 38387 24735 38390
rect 27153 38387 27219 38390
rect 28441 38387 28507 38390
rect 28950 38448 29059 38450
rect 28950 38392 28998 38448
rect 29054 38392 29059 38448
rect 28950 38387 29059 38392
rect 53557 38450 53623 38453
rect 55200 38450 56000 38480
rect 53557 38448 56000 38450
rect 53557 38392 53562 38448
rect 53618 38392 56000 38448
rect 53557 38390 56000 38392
rect 53557 38387 53623 38390
rect 26601 38314 26667 38317
rect 27613 38314 27679 38317
rect 26601 38312 27679 38314
rect 26601 38256 26606 38312
rect 26662 38256 27618 38312
rect 27674 38256 27679 38312
rect 26601 38254 27679 38256
rect 28950 38314 29010 38387
rect 55200 38360 56000 38390
rect 31477 38314 31543 38317
rect 28950 38312 31543 38314
rect 28950 38256 31482 38312
rect 31538 38256 31543 38312
rect 28950 38254 31543 38256
rect 26601 38251 26667 38254
rect 27613 38251 27679 38254
rect 31477 38251 31543 38254
rect 24025 38178 24091 38181
rect 27153 38178 27219 38181
rect 24025 38176 27219 38178
rect 24025 38120 24030 38176
rect 24086 38120 27158 38176
rect 27214 38120 27219 38176
rect 24025 38118 27219 38120
rect 24025 38115 24091 38118
rect 27153 38115 27219 38118
rect 52177 38178 52243 38181
rect 55200 38178 56000 38208
rect 52177 38176 56000 38178
rect 52177 38120 52182 38176
rect 52238 38120 56000 38176
rect 52177 38118 56000 38120
rect 52177 38115 52243 38118
rect 19570 38112 19886 38113
rect 0 38042 800 38072
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 55200 38088 56000 38118
rect 50290 38047 50606 38048
rect 1669 38042 1735 38045
rect 0 38040 1735 38042
rect 0 37984 1674 38040
rect 1730 37984 1735 38040
rect 0 37982 1735 37984
rect 0 37952 800 37982
rect 1669 37979 1735 37982
rect 28257 38042 28323 38045
rect 29453 38042 29519 38045
rect 28257 38040 29519 38042
rect 28257 37984 28262 38040
rect 28318 37984 29458 38040
rect 29514 37984 29519 38040
rect 28257 37982 29519 37984
rect 28257 37979 28323 37982
rect 29453 37979 29519 37982
rect 29729 38042 29795 38045
rect 31017 38042 31083 38045
rect 29729 38040 31083 38042
rect 29729 37984 29734 38040
rect 29790 37984 31022 38040
rect 31078 37984 31083 38040
rect 29729 37982 31083 37984
rect 29729 37979 29795 37982
rect 31017 37979 31083 37982
rect 31201 38042 31267 38045
rect 31334 38042 31340 38044
rect 31201 38040 31340 38042
rect 31201 37984 31206 38040
rect 31262 37984 31340 38040
rect 31201 37982 31340 37984
rect 31201 37979 31267 37982
rect 31334 37980 31340 37982
rect 31404 37980 31410 38044
rect 26366 37844 26372 37908
rect 26436 37906 26442 37908
rect 26693 37906 26759 37909
rect 26436 37904 26759 37906
rect 26436 37848 26698 37904
rect 26754 37848 26759 37904
rect 26436 37846 26759 37848
rect 26436 37844 26442 37846
rect 26693 37843 26759 37846
rect 28809 37906 28875 37909
rect 29637 37906 29703 37909
rect 28809 37904 29703 37906
rect 28809 37848 28814 37904
rect 28870 37848 29642 37904
rect 29698 37848 29703 37904
rect 28809 37846 29703 37848
rect 28809 37843 28875 37846
rect 29637 37843 29703 37846
rect 30833 37906 30899 37909
rect 31753 37906 31819 37909
rect 33225 37906 33291 37909
rect 30833 37904 33291 37906
rect 30833 37848 30838 37904
rect 30894 37848 31758 37904
rect 31814 37848 33230 37904
rect 33286 37848 33291 37904
rect 30833 37846 33291 37848
rect 30833 37843 30899 37846
rect 31753 37843 31819 37846
rect 33225 37843 33291 37846
rect 53465 37906 53531 37909
rect 55200 37906 56000 37936
rect 53465 37904 56000 37906
rect 53465 37848 53470 37904
rect 53526 37848 56000 37904
rect 53465 37846 56000 37848
rect 53465 37843 53531 37846
rect 55200 37816 56000 37846
rect 27889 37770 27955 37773
rect 28206 37770 28212 37772
rect 27889 37768 28212 37770
rect 27889 37712 27894 37768
rect 27950 37712 28212 37768
rect 27889 37710 28212 37712
rect 27889 37707 27955 37710
rect 28206 37708 28212 37710
rect 28276 37708 28282 37772
rect 29269 37770 29335 37773
rect 34329 37770 34395 37773
rect 29269 37768 34395 37770
rect 29269 37712 29274 37768
rect 29330 37712 34334 37768
rect 34390 37712 34395 37768
rect 29269 37710 34395 37712
rect 29269 37707 29335 37710
rect 34329 37707 34395 37710
rect 26233 37634 26299 37637
rect 26693 37634 26759 37637
rect 26233 37632 26759 37634
rect 26233 37576 26238 37632
rect 26294 37576 26698 37632
rect 26754 37576 26759 37632
rect 26233 37574 26759 37576
rect 26233 37571 26299 37574
rect 26693 37571 26759 37574
rect 27654 37572 27660 37636
rect 27724 37634 27730 37636
rect 28257 37634 28323 37637
rect 27724 37632 28323 37634
rect 27724 37576 28262 37632
rect 28318 37576 28323 37632
rect 27724 37574 28323 37576
rect 27724 37572 27730 37574
rect 28257 37571 28323 37574
rect 53005 37634 53071 37637
rect 55200 37634 56000 37664
rect 53005 37632 56000 37634
rect 53005 37576 53010 37632
rect 53066 37576 56000 37632
rect 53005 37574 56000 37576
rect 53005 37571 53071 37574
rect 4210 37568 4526 37569
rect 0 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 55200 37544 56000 37574
rect 34930 37503 35246 37504
rect 1577 37498 1643 37501
rect 0 37496 1643 37498
rect 0 37440 1582 37496
rect 1638 37440 1643 37496
rect 0 37438 1643 37440
rect 0 37408 800 37438
rect 1577 37435 1643 37438
rect 24025 37498 24091 37501
rect 27102 37498 27108 37500
rect 24025 37496 27108 37498
rect 24025 37440 24030 37496
rect 24086 37440 27108 37496
rect 24025 37438 27108 37440
rect 24025 37435 24091 37438
rect 27102 37436 27108 37438
rect 27172 37436 27178 37500
rect 27337 37498 27403 37501
rect 28942 37498 28948 37500
rect 27337 37496 28948 37498
rect 27337 37440 27342 37496
rect 27398 37440 28948 37496
rect 27337 37438 28948 37440
rect 27337 37435 27403 37438
rect 28942 37436 28948 37438
rect 29012 37436 29018 37500
rect 26049 37364 26115 37365
rect 25998 37362 26004 37364
rect 25958 37302 26004 37362
rect 26068 37360 26115 37364
rect 26110 37304 26115 37360
rect 25998 37300 26004 37302
rect 26068 37300 26115 37304
rect 26049 37299 26115 37300
rect 53373 37362 53439 37365
rect 55200 37362 56000 37392
rect 53373 37360 56000 37362
rect 53373 37304 53378 37360
rect 53434 37304 56000 37360
rect 53373 37302 56000 37304
rect 53373 37299 53439 37302
rect 55200 37272 56000 37302
rect 22369 37226 22435 37229
rect 26785 37226 26851 37229
rect 27061 37228 27127 37229
rect 27061 37226 27108 37228
rect 22369 37224 26851 37226
rect 22369 37168 22374 37224
rect 22430 37168 26790 37224
rect 26846 37168 26851 37224
rect 22369 37166 26851 37168
rect 27016 37224 27108 37226
rect 27016 37168 27066 37224
rect 27016 37166 27108 37168
rect 22369 37163 22435 37166
rect 26785 37163 26851 37166
rect 27061 37164 27108 37166
rect 27172 37164 27178 37228
rect 27889 37226 27955 37229
rect 29678 37226 29684 37228
rect 27889 37224 29684 37226
rect 27889 37168 27894 37224
rect 27950 37168 29684 37224
rect 27889 37166 29684 37168
rect 27061 37163 27127 37164
rect 27889 37163 27955 37166
rect 29678 37164 29684 37166
rect 29748 37164 29754 37228
rect 30281 37226 30347 37229
rect 33777 37226 33843 37229
rect 30281 37224 33843 37226
rect 30281 37168 30286 37224
rect 30342 37168 33782 37224
rect 33838 37168 33843 37224
rect 30281 37166 33843 37168
rect 30281 37163 30347 37166
rect 33777 37163 33843 37166
rect 28165 37090 28231 37093
rect 31201 37090 31267 37093
rect 28165 37088 31267 37090
rect 28165 37032 28170 37088
rect 28226 37032 31206 37088
rect 31262 37032 31267 37088
rect 28165 37030 31267 37032
rect 28165 37027 28231 37030
rect 31201 37027 31267 37030
rect 53005 37090 53071 37093
rect 55200 37090 56000 37120
rect 53005 37088 56000 37090
rect 53005 37032 53010 37088
rect 53066 37032 56000 37088
rect 53005 37030 56000 37032
rect 53005 37027 53071 37030
rect 19570 37024 19886 37025
rect 0 36954 800 36984
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 55200 37000 56000 37030
rect 50290 36959 50606 36960
rect 2773 36954 2839 36957
rect 0 36952 2839 36954
rect 0 36896 2778 36952
rect 2834 36896 2839 36952
rect 0 36894 2839 36896
rect 0 36864 800 36894
rect 2773 36891 2839 36894
rect 26509 36954 26575 36957
rect 27061 36954 27127 36957
rect 28257 36954 28323 36957
rect 26509 36952 28323 36954
rect 26509 36896 26514 36952
rect 26570 36896 27066 36952
rect 27122 36896 28262 36952
rect 28318 36896 28323 36952
rect 26509 36894 28323 36896
rect 26509 36891 26575 36894
rect 27061 36891 27127 36894
rect 28257 36891 28323 36894
rect 53741 36818 53807 36821
rect 55200 36818 56000 36848
rect 53741 36816 56000 36818
rect 53741 36760 53746 36816
rect 53802 36760 56000 36816
rect 53741 36758 56000 36760
rect 53741 36755 53807 36758
rect 55200 36728 56000 36758
rect 2221 36682 2287 36685
rect 22553 36682 22619 36685
rect 25865 36682 25931 36685
rect 2221 36680 25931 36682
rect 2221 36624 2226 36680
rect 2282 36624 22558 36680
rect 22614 36624 25870 36680
rect 25926 36624 25931 36680
rect 2221 36622 25931 36624
rect 2221 36619 2287 36622
rect 22553 36619 22619 36622
rect 25865 36619 25931 36622
rect 27889 36682 27955 36685
rect 28717 36682 28783 36685
rect 27889 36680 28783 36682
rect 27889 36624 27894 36680
rect 27950 36624 28722 36680
rect 28778 36624 28783 36680
rect 27889 36622 28783 36624
rect 27889 36619 27955 36622
rect 28717 36619 28783 36622
rect 25405 36546 25471 36549
rect 27889 36546 27955 36549
rect 25405 36544 27955 36546
rect 25405 36488 25410 36544
rect 25466 36488 27894 36544
rect 27950 36488 27955 36544
rect 25405 36486 27955 36488
rect 25405 36483 25471 36486
rect 27889 36483 27955 36486
rect 28993 36546 29059 36549
rect 33225 36546 33291 36549
rect 28993 36544 33291 36546
rect 28993 36488 28998 36544
rect 29054 36488 33230 36544
rect 33286 36488 33291 36544
rect 28993 36486 33291 36488
rect 28993 36483 29059 36486
rect 33225 36483 33291 36486
rect 53649 36546 53715 36549
rect 55200 36546 56000 36576
rect 53649 36544 56000 36546
rect 53649 36488 53654 36544
rect 53710 36488 56000 36544
rect 53649 36486 56000 36488
rect 53649 36483 53715 36486
rect 4210 36480 4526 36481
rect 0 36410 800 36440
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 55200 36456 56000 36486
rect 34930 36415 35246 36416
rect 2773 36410 2839 36413
rect 0 36408 2839 36410
rect 0 36352 2778 36408
rect 2834 36352 2839 36408
rect 0 36350 2839 36352
rect 0 36320 800 36350
rect 2773 36347 2839 36350
rect 25497 36410 25563 36413
rect 28717 36410 28783 36413
rect 25497 36408 28783 36410
rect 25497 36352 25502 36408
rect 25558 36352 28722 36408
rect 28778 36352 28783 36408
rect 25497 36350 28783 36352
rect 25497 36347 25563 36350
rect 28717 36347 28783 36350
rect 29453 36410 29519 36413
rect 31201 36410 31267 36413
rect 29453 36408 31267 36410
rect 29453 36352 29458 36408
rect 29514 36352 31206 36408
rect 31262 36352 31267 36408
rect 29453 36350 31267 36352
rect 29453 36347 29519 36350
rect 31201 36347 31267 36350
rect 27521 36274 27587 36277
rect 28809 36274 28875 36277
rect 31937 36274 32003 36277
rect 27521 36272 28875 36274
rect 27521 36216 27526 36272
rect 27582 36216 28814 36272
rect 28870 36216 28875 36272
rect 27521 36214 28875 36216
rect 27521 36211 27587 36214
rect 28809 36211 28875 36214
rect 29134 36272 32003 36274
rect 29134 36216 31942 36272
rect 31998 36216 32003 36272
rect 29134 36214 32003 36216
rect 21265 36138 21331 36141
rect 25589 36138 25655 36141
rect 21265 36136 25655 36138
rect 21265 36080 21270 36136
rect 21326 36080 25594 36136
rect 25650 36080 25655 36136
rect 21265 36078 25655 36080
rect 21265 36075 21331 36078
rect 25589 36075 25655 36078
rect 28993 36138 29059 36141
rect 29134 36138 29194 36214
rect 31937 36211 32003 36214
rect 53465 36274 53531 36277
rect 55200 36274 56000 36304
rect 53465 36272 56000 36274
rect 53465 36216 53470 36272
rect 53526 36216 56000 36272
rect 53465 36214 56000 36216
rect 53465 36211 53531 36214
rect 55200 36184 56000 36214
rect 28993 36136 29194 36138
rect 28993 36080 28998 36136
rect 29054 36080 29194 36136
rect 28993 36078 29194 36080
rect 28993 36075 29059 36078
rect 22921 36002 22987 36005
rect 27429 36002 27495 36005
rect 22921 36000 27495 36002
rect 22921 35944 22926 36000
rect 22982 35944 27434 36000
rect 27490 35944 27495 36000
rect 22921 35942 27495 35944
rect 22921 35939 22987 35942
rect 27429 35939 27495 35942
rect 29269 36004 29335 36005
rect 29269 36000 29316 36004
rect 29380 36002 29386 36004
rect 53557 36002 53623 36005
rect 55200 36002 56000 36032
rect 29269 35944 29274 36000
rect 29269 35940 29316 35944
rect 29380 35942 29426 36002
rect 53557 36000 56000 36002
rect 53557 35944 53562 36000
rect 53618 35944 56000 36000
rect 53557 35942 56000 35944
rect 29380 35940 29386 35942
rect 29269 35939 29335 35940
rect 53557 35939 53623 35942
rect 19570 35936 19886 35937
rect 0 35866 800 35896
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 55200 35912 56000 35942
rect 50290 35871 50606 35872
rect 2773 35866 2839 35869
rect 0 35864 2839 35866
rect 0 35808 2778 35864
rect 2834 35808 2839 35864
rect 0 35806 2839 35808
rect 0 35776 800 35806
rect 2773 35803 2839 35806
rect 27521 35866 27587 35869
rect 28625 35866 28691 35869
rect 27521 35864 28691 35866
rect 27521 35808 27526 35864
rect 27582 35808 28630 35864
rect 28686 35808 28691 35864
rect 27521 35806 28691 35808
rect 27521 35803 27587 35806
rect 28625 35803 28691 35806
rect 23473 35730 23539 35733
rect 25037 35730 25103 35733
rect 23473 35728 25103 35730
rect 23473 35672 23478 35728
rect 23534 35672 25042 35728
rect 25098 35672 25103 35728
rect 23473 35670 25103 35672
rect 23473 35667 23539 35670
rect 25037 35667 25103 35670
rect 26693 35730 26759 35733
rect 28533 35730 28599 35733
rect 26693 35728 28599 35730
rect 26693 35672 26698 35728
rect 26754 35672 28538 35728
rect 28594 35672 28599 35728
rect 26693 35670 28599 35672
rect 26693 35667 26759 35670
rect 28533 35667 28599 35670
rect 53465 35730 53531 35733
rect 55200 35730 56000 35760
rect 53465 35728 56000 35730
rect 53465 35672 53470 35728
rect 53526 35672 56000 35728
rect 53465 35670 56000 35672
rect 53465 35667 53531 35670
rect 55200 35640 56000 35670
rect 23013 35594 23079 35597
rect 23749 35594 23815 35597
rect 27429 35596 27495 35597
rect 27429 35594 27476 35596
rect 23013 35592 23815 35594
rect 23013 35536 23018 35592
rect 23074 35536 23754 35592
rect 23810 35536 23815 35592
rect 23013 35534 23815 35536
rect 27384 35592 27476 35594
rect 27384 35536 27434 35592
rect 27384 35534 27476 35536
rect 23013 35531 23079 35534
rect 23749 35531 23815 35534
rect 27429 35532 27476 35534
rect 27540 35532 27546 35596
rect 27613 35594 27679 35597
rect 28809 35594 28875 35597
rect 27613 35592 28875 35594
rect 27613 35536 27618 35592
rect 27674 35536 28814 35592
rect 28870 35536 28875 35592
rect 27613 35534 28875 35536
rect 27429 35531 27495 35532
rect 27613 35531 27679 35534
rect 28809 35531 28875 35534
rect 26141 35458 26207 35461
rect 26366 35458 26372 35460
rect 26141 35456 26372 35458
rect 26141 35400 26146 35456
rect 26202 35400 26372 35456
rect 26141 35398 26372 35400
rect 26141 35395 26207 35398
rect 26366 35396 26372 35398
rect 26436 35396 26442 35460
rect 29085 35458 29151 35461
rect 29361 35458 29427 35461
rect 29085 35456 29427 35458
rect 29085 35400 29090 35456
rect 29146 35400 29366 35456
rect 29422 35400 29427 35456
rect 29085 35398 29427 35400
rect 29085 35395 29151 35398
rect 29361 35395 29427 35398
rect 53465 35458 53531 35461
rect 55200 35458 56000 35488
rect 53465 35456 56000 35458
rect 53465 35400 53470 35456
rect 53526 35400 56000 35456
rect 53465 35398 56000 35400
rect 53465 35395 53531 35398
rect 4210 35392 4526 35393
rect 0 35322 800 35352
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 55200 35368 56000 35398
rect 34930 35327 35246 35328
rect 2773 35322 2839 35325
rect 0 35320 2839 35322
rect 0 35264 2778 35320
rect 2834 35264 2839 35320
rect 0 35262 2839 35264
rect 0 35232 800 35262
rect 2773 35259 2839 35262
rect 21173 35322 21239 35325
rect 24393 35322 24459 35325
rect 21173 35320 24459 35322
rect 21173 35264 21178 35320
rect 21234 35264 24398 35320
rect 24454 35264 24459 35320
rect 21173 35262 24459 35264
rect 21173 35259 21239 35262
rect 24393 35259 24459 35262
rect 27337 35322 27403 35325
rect 28717 35322 28783 35325
rect 27337 35320 28783 35322
rect 27337 35264 27342 35320
rect 27398 35264 28722 35320
rect 28778 35264 28783 35320
rect 27337 35262 28783 35264
rect 27337 35259 27403 35262
rect 28717 35259 28783 35262
rect 52361 35186 52427 35189
rect 55200 35186 56000 35216
rect 52361 35184 56000 35186
rect 52361 35128 52366 35184
rect 52422 35128 56000 35184
rect 52361 35126 56000 35128
rect 52361 35123 52427 35126
rect 55200 35096 56000 35126
rect 3233 35050 3299 35053
rect 21173 35050 21239 35053
rect 3233 35048 21239 35050
rect 3233 34992 3238 35048
rect 3294 34992 21178 35048
rect 21234 34992 21239 35048
rect 3233 34990 21239 34992
rect 3233 34987 3299 34990
rect 21173 34987 21239 34990
rect 21725 35050 21791 35053
rect 23473 35050 23539 35053
rect 21725 35048 23539 35050
rect 21725 34992 21730 35048
rect 21786 34992 23478 35048
rect 23534 34992 23539 35048
rect 21725 34990 23539 34992
rect 21725 34987 21791 34990
rect 23473 34987 23539 34990
rect 28993 35050 29059 35053
rect 31477 35050 31543 35053
rect 28993 35048 31543 35050
rect 28993 34992 28998 35048
rect 29054 34992 31482 35048
rect 31538 34992 31543 35048
rect 28993 34990 31543 34992
rect 28993 34987 29059 34990
rect 31477 34987 31543 34990
rect 26366 34852 26372 34916
rect 26436 34914 26442 34916
rect 30557 34914 30623 34917
rect 33501 34914 33567 34917
rect 26436 34854 27630 34914
rect 26436 34852 26442 34854
rect 19570 34848 19886 34849
rect 0 34778 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 1577 34778 1643 34781
rect 0 34776 1643 34778
rect 0 34720 1582 34776
rect 1638 34720 1643 34776
rect 0 34718 1643 34720
rect 0 34688 800 34718
rect 1577 34715 1643 34718
rect 27570 34642 27630 34854
rect 30557 34912 33567 34914
rect 30557 34856 30562 34912
rect 30618 34856 33506 34912
rect 33562 34856 33567 34912
rect 30557 34854 33567 34856
rect 30557 34851 30623 34854
rect 33501 34851 33567 34854
rect 53465 34914 53531 34917
rect 55200 34914 56000 34944
rect 53465 34912 56000 34914
rect 53465 34856 53470 34912
rect 53526 34856 56000 34912
rect 53465 34854 56000 34856
rect 53465 34851 53531 34854
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 55200 34824 56000 34854
rect 50290 34783 50606 34784
rect 30373 34778 30439 34781
rect 30925 34778 30991 34781
rect 30373 34776 30991 34778
rect 30373 34720 30378 34776
rect 30434 34720 30930 34776
rect 30986 34720 30991 34776
rect 30373 34718 30991 34720
rect 30373 34715 30439 34718
rect 30925 34715 30991 34718
rect 29637 34642 29703 34645
rect 31293 34642 31359 34645
rect 27570 34582 29562 34642
rect 25405 34506 25471 34509
rect 28073 34506 28139 34509
rect 25405 34504 28139 34506
rect 25405 34448 25410 34504
rect 25466 34448 28078 34504
rect 28134 34448 28139 34504
rect 25405 34446 28139 34448
rect 29502 34506 29562 34582
rect 29637 34640 31359 34642
rect 29637 34584 29642 34640
rect 29698 34584 31298 34640
rect 31354 34584 31359 34640
rect 29637 34582 31359 34584
rect 29637 34579 29703 34582
rect 31293 34579 31359 34582
rect 53557 34642 53623 34645
rect 55200 34642 56000 34672
rect 53557 34640 56000 34642
rect 53557 34584 53562 34640
rect 53618 34584 56000 34640
rect 53557 34582 56000 34584
rect 53557 34579 53623 34582
rect 55200 34552 56000 34582
rect 31109 34506 31175 34509
rect 29502 34504 31175 34506
rect 29502 34448 31114 34504
rect 31170 34448 31175 34504
rect 29502 34446 31175 34448
rect 25405 34443 25471 34446
rect 28073 34443 28139 34446
rect 31109 34443 31175 34446
rect 53005 34370 53071 34373
rect 55200 34370 56000 34400
rect 53005 34368 56000 34370
rect 53005 34312 53010 34368
rect 53066 34312 56000 34368
rect 53005 34310 56000 34312
rect 53005 34307 53071 34310
rect 4210 34304 4526 34305
rect 0 34234 800 34264
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 55200 34280 56000 34310
rect 34930 34239 35246 34240
rect 2773 34234 2839 34237
rect 0 34232 2839 34234
rect 0 34176 2778 34232
rect 2834 34176 2839 34232
rect 0 34174 2839 34176
rect 0 34144 800 34174
rect 2773 34171 2839 34174
rect 24209 34098 24275 34101
rect 27981 34098 28047 34101
rect 24209 34096 28047 34098
rect 24209 34040 24214 34096
rect 24270 34040 27986 34096
rect 28042 34040 28047 34096
rect 24209 34038 28047 34040
rect 24209 34035 24275 34038
rect 27981 34035 28047 34038
rect 53281 34098 53347 34101
rect 55200 34098 56000 34128
rect 53281 34096 56000 34098
rect 53281 34040 53286 34096
rect 53342 34040 56000 34096
rect 53281 34038 56000 34040
rect 53281 34035 53347 34038
rect 55200 34008 56000 34038
rect 19570 33760 19886 33761
rect 0 33690 800 33720
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 55200 33736 56000 33856
rect 50290 33695 50606 33696
rect 2773 33690 2839 33693
rect 0 33688 2839 33690
rect 0 33632 2778 33688
rect 2834 33632 2839 33688
rect 0 33630 2839 33632
rect 0 33600 800 33630
rect 2773 33627 2839 33630
rect 55200 33464 56000 33584
rect 29085 33420 29151 33421
rect 29085 33416 29132 33420
rect 29196 33418 29202 33420
rect 29085 33360 29090 33416
rect 29085 33356 29132 33360
rect 29196 33358 29242 33418
rect 29196 33356 29202 33358
rect 29085 33355 29151 33356
rect 54293 33282 54359 33285
rect 55200 33282 56000 33312
rect 54293 33280 56000 33282
rect 54293 33224 54298 33280
rect 54354 33224 56000 33280
rect 54293 33222 56000 33224
rect 54293 33219 54359 33222
rect 4210 33216 4526 33217
rect 0 33146 800 33176
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 55200 33192 56000 33222
rect 34930 33151 35246 33152
rect 2773 33146 2839 33149
rect 28257 33148 28323 33149
rect 0 33144 2839 33146
rect 0 33088 2778 33144
rect 2834 33088 2839 33144
rect 0 33086 2839 33088
rect 0 33056 800 33086
rect 2773 33083 2839 33086
rect 28206 33084 28212 33148
rect 28276 33146 28323 33148
rect 28276 33144 28368 33146
rect 28318 33088 28368 33144
rect 28276 33086 28368 33088
rect 28276 33084 28323 33086
rect 28257 33083 28323 33084
rect 55200 32920 56000 33040
rect 19570 32672 19886 32673
rect 0 32602 800 32632
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 55200 32648 56000 32768
rect 50290 32607 50606 32608
rect 1577 32602 1643 32605
rect 0 32600 1643 32602
rect 0 32544 1582 32600
rect 1638 32544 1643 32600
rect 0 32542 1643 32544
rect 0 32512 800 32542
rect 1577 32539 1643 32542
rect 28942 32404 28948 32468
rect 29012 32466 29018 32468
rect 50061 32466 50127 32469
rect 29012 32464 50127 32466
rect 29012 32408 50066 32464
rect 50122 32408 50127 32464
rect 29012 32406 50127 32408
rect 29012 32404 29018 32406
rect 50061 32403 50127 32406
rect 54293 32466 54359 32469
rect 55200 32466 56000 32496
rect 54293 32464 56000 32466
rect 54293 32408 54298 32464
rect 54354 32408 56000 32464
rect 54293 32406 56000 32408
rect 54293 32403 54359 32406
rect 55200 32376 56000 32406
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 55200 32104 56000 32224
rect 34930 32063 35246 32064
rect 2773 32058 2839 32061
rect 0 32056 2839 32058
rect 0 32000 2778 32056
rect 2834 32000 2839 32056
rect 0 31998 2839 32000
rect 0 31968 800 31998
rect 2773 31995 2839 31998
rect 24945 31922 25011 31925
rect 26969 31922 27035 31925
rect 24945 31920 27035 31922
rect 24945 31864 24950 31920
rect 25006 31864 26974 31920
rect 27030 31864 27035 31920
rect 24945 31862 27035 31864
rect 24945 31859 25011 31862
rect 26969 31859 27035 31862
rect 55200 31832 56000 31952
rect 26366 31724 26372 31788
rect 26436 31786 26442 31788
rect 26785 31786 26851 31789
rect 26436 31784 26851 31786
rect 26436 31728 26790 31784
rect 26846 31728 26851 31784
rect 26436 31726 26851 31728
rect 26436 31724 26442 31726
rect 26785 31723 26851 31726
rect 31569 31786 31635 31789
rect 32622 31786 32628 31788
rect 31569 31784 32628 31786
rect 31569 31728 31574 31784
rect 31630 31728 32628 31784
rect 31569 31726 32628 31728
rect 31569 31723 31635 31726
rect 32622 31724 32628 31726
rect 32692 31724 32698 31788
rect 54293 31650 54359 31653
rect 55200 31650 56000 31680
rect 54293 31648 56000 31650
rect 54293 31592 54298 31648
rect 54354 31592 56000 31648
rect 54293 31590 56000 31592
rect 54293 31587 54359 31590
rect 19570 31584 19886 31585
rect 0 31514 800 31544
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 55200 31560 56000 31590
rect 50290 31519 50606 31520
rect 2773 31514 2839 31517
rect 0 31512 2839 31514
rect 0 31456 2778 31512
rect 2834 31456 2839 31512
rect 0 31454 2839 31456
rect 0 31424 800 31454
rect 2773 31451 2839 31454
rect 55200 31288 56000 31408
rect 4210 31040 4526 31041
rect 0 30970 800 31000
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 55200 31016 56000 31136
rect 34930 30975 35246 30976
rect 2773 30970 2839 30973
rect 0 30968 2839 30970
rect 0 30912 2778 30968
rect 2834 30912 2839 30968
rect 0 30910 2839 30912
rect 0 30880 800 30910
rect 2773 30907 2839 30910
rect 54293 30834 54359 30837
rect 55200 30834 56000 30864
rect 54293 30832 56000 30834
rect 54293 30776 54298 30832
rect 54354 30776 56000 30832
rect 54293 30774 56000 30776
rect 54293 30771 54359 30774
rect 55200 30744 56000 30774
rect 19570 30496 19886 30497
rect 0 30426 800 30456
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 55200 30472 56000 30592
rect 50290 30431 50606 30432
rect 2773 30426 2839 30429
rect 0 30424 2839 30426
rect 0 30368 2778 30424
rect 2834 30368 2839 30424
rect 0 30366 2839 30368
rect 0 30336 800 30366
rect 2773 30363 2839 30366
rect 55200 30200 56000 30320
rect 54201 30018 54267 30021
rect 55200 30018 56000 30048
rect 54201 30016 56000 30018
rect 54201 29960 54206 30016
rect 54262 29960 56000 30016
rect 54201 29958 56000 29960
rect 54201 29955 54267 29958
rect 4210 29952 4526 29953
rect 0 29882 800 29912
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 55200 29928 56000 29958
rect 34930 29887 35246 29888
rect 2221 29882 2287 29885
rect 0 29880 2287 29882
rect 0 29824 2226 29880
rect 2282 29824 2287 29880
rect 0 29822 2287 29824
rect 0 29792 800 29822
rect 2221 29819 2287 29822
rect 54201 29746 54267 29749
rect 55200 29746 56000 29776
rect 54201 29744 56000 29746
rect 54201 29688 54206 29744
rect 54262 29688 56000 29744
rect 54201 29686 56000 29688
rect 54201 29683 54267 29686
rect 55200 29656 56000 29686
rect 19570 29408 19886 29409
rect 0 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 55200 29384 56000 29504
rect 50290 29343 50606 29344
rect 1577 29338 1643 29341
rect 0 29336 1643 29338
rect 0 29280 1582 29336
rect 1638 29280 1643 29336
rect 0 29278 1643 29280
rect 0 29248 800 29278
rect 1577 29275 1643 29278
rect 54201 29202 54267 29205
rect 55200 29202 56000 29232
rect 54201 29200 56000 29202
rect 54201 29144 54206 29200
rect 54262 29144 56000 29200
rect 54201 29142 56000 29144
rect 54201 29139 54267 29142
rect 55200 29112 56000 29142
rect 54201 28930 54267 28933
rect 55200 28930 56000 28960
rect 54201 28928 56000 28930
rect 54201 28872 54206 28928
rect 54262 28872 56000 28928
rect 54201 28870 56000 28872
rect 54201 28867 54267 28870
rect 4210 28864 4526 28865
rect 0 28794 800 28824
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 55200 28840 56000 28870
rect 34930 28799 35246 28800
rect 2773 28794 2839 28797
rect 0 28792 2839 28794
rect 0 28736 2778 28792
rect 2834 28736 2839 28792
rect 0 28734 2839 28736
rect 0 28704 800 28734
rect 2773 28731 2839 28734
rect 55200 28568 56000 28688
rect 54201 28386 54267 28389
rect 55200 28386 56000 28416
rect 54201 28384 56000 28386
rect 54201 28328 54206 28384
rect 54262 28328 56000 28384
rect 54201 28326 56000 28328
rect 54201 28323 54267 28326
rect 19570 28320 19886 28321
rect 0 28250 800 28280
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 55200 28296 56000 28326
rect 50290 28255 50606 28256
rect 2773 28250 2839 28253
rect 0 28248 2839 28250
rect 0 28192 2778 28248
rect 2834 28192 2839 28248
rect 0 28190 2839 28192
rect 0 28160 800 28190
rect 2773 28187 2839 28190
rect 53465 28114 53531 28117
rect 55200 28114 56000 28144
rect 53465 28112 56000 28114
rect 53465 28056 53470 28112
rect 53526 28056 56000 28112
rect 53465 28054 56000 28056
rect 53465 28051 53531 28054
rect 55200 28024 56000 28054
rect 4210 27776 4526 27777
rect 0 27706 800 27736
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 55200 27752 56000 27872
rect 34930 27711 35246 27712
rect 2221 27706 2287 27709
rect 0 27704 2287 27706
rect 0 27648 2226 27704
rect 2282 27648 2287 27704
rect 0 27646 2287 27648
rect 0 27616 800 27646
rect 2221 27643 2287 27646
rect 30046 27644 30052 27708
rect 30116 27706 30122 27708
rect 30925 27706 30991 27709
rect 30116 27704 30991 27706
rect 30116 27648 30930 27704
rect 30986 27648 30991 27704
rect 30116 27646 30991 27648
rect 30116 27644 30122 27646
rect 30925 27643 30991 27646
rect 26417 27570 26483 27573
rect 26550 27570 26556 27572
rect 26417 27568 26556 27570
rect 26417 27512 26422 27568
rect 26478 27512 26556 27568
rect 26417 27510 26556 27512
rect 26417 27507 26483 27510
rect 26550 27508 26556 27510
rect 26620 27508 26626 27572
rect 53465 27570 53531 27573
rect 55200 27570 56000 27600
rect 53465 27568 56000 27570
rect 53465 27512 53470 27568
rect 53526 27512 56000 27568
rect 53465 27510 56000 27512
rect 53465 27507 53531 27510
rect 55200 27480 56000 27510
rect 54201 27298 54267 27301
rect 55200 27298 56000 27328
rect 54201 27296 56000 27298
rect 54201 27240 54206 27296
rect 54262 27240 56000 27296
rect 54201 27238 56000 27240
rect 54201 27235 54267 27238
rect 19570 27232 19886 27233
rect 0 27162 800 27192
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 55200 27208 56000 27238
rect 50290 27167 50606 27168
rect 1577 27162 1643 27165
rect 0 27160 1643 27162
rect 0 27104 1582 27160
rect 1638 27104 1643 27160
rect 0 27102 1643 27104
rect 0 27072 800 27102
rect 1577 27099 1643 27102
rect 53465 27026 53531 27029
rect 55200 27026 56000 27056
rect 53465 27024 56000 27026
rect 53465 26968 53470 27024
rect 53526 26968 56000 27024
rect 53465 26966 56000 26968
rect 53465 26963 53531 26966
rect 55200 26936 56000 26966
rect 54201 26754 54267 26757
rect 55200 26754 56000 26784
rect 54201 26752 56000 26754
rect 54201 26696 54206 26752
rect 54262 26696 56000 26752
rect 54201 26694 56000 26696
rect 54201 26691 54267 26694
rect 4210 26688 4526 26689
rect 0 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 55200 26664 56000 26694
rect 34930 26623 35246 26624
rect 2773 26618 2839 26621
rect 0 26616 2839 26618
rect 0 26560 2778 26616
rect 2834 26560 2839 26616
rect 0 26558 2839 26560
rect 0 26528 800 26558
rect 2773 26555 2839 26558
rect 53557 26482 53623 26485
rect 55200 26482 56000 26512
rect 53557 26480 56000 26482
rect 53557 26424 53562 26480
rect 53618 26424 56000 26480
rect 53557 26422 56000 26424
rect 53557 26419 53623 26422
rect 55200 26392 56000 26422
rect 53557 26210 53623 26213
rect 55200 26210 56000 26240
rect 53557 26208 56000 26210
rect 53557 26152 53562 26208
rect 53618 26152 56000 26208
rect 53557 26150 56000 26152
rect 53557 26147 53623 26150
rect 19570 26144 19886 26145
rect 0 26074 800 26104
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 55200 26120 56000 26150
rect 50290 26079 50606 26080
rect 2221 26074 2287 26077
rect 0 26072 2287 26074
rect 0 26016 2226 26072
rect 2282 26016 2287 26072
rect 0 26014 2287 26016
rect 0 25984 800 26014
rect 2221 26011 2287 26014
rect 32213 26074 32279 26077
rect 33593 26074 33659 26077
rect 32213 26072 33659 26074
rect 32213 26016 32218 26072
rect 32274 26016 33598 26072
rect 33654 26016 33659 26072
rect 32213 26014 33659 26016
rect 32213 26011 32279 26014
rect 33593 26011 33659 26014
rect 54201 25938 54267 25941
rect 55200 25938 56000 25968
rect 54201 25936 56000 25938
rect 54201 25880 54206 25936
rect 54262 25880 56000 25936
rect 54201 25878 56000 25880
rect 54201 25875 54267 25878
rect 55200 25848 56000 25878
rect 53557 25666 53623 25669
rect 55200 25666 56000 25696
rect 53557 25664 56000 25666
rect 53557 25608 53562 25664
rect 53618 25608 56000 25664
rect 53557 25606 56000 25608
rect 53557 25603 53623 25606
rect 4210 25600 4526 25601
rect 0 25530 800 25560
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 55200 25576 56000 25606
rect 34930 25535 35246 25536
rect 1577 25530 1643 25533
rect 0 25528 1643 25530
rect 0 25472 1582 25528
rect 1638 25472 1643 25528
rect 0 25470 1643 25472
rect 0 25440 800 25470
rect 1577 25467 1643 25470
rect 53465 25394 53531 25397
rect 55200 25394 56000 25424
rect 53465 25392 56000 25394
rect 53465 25336 53470 25392
rect 53526 25336 56000 25392
rect 53465 25334 56000 25336
rect 53465 25331 53531 25334
rect 55200 25304 56000 25334
rect 33358 25196 33364 25260
rect 33428 25258 33434 25260
rect 33593 25258 33659 25261
rect 33428 25256 33659 25258
rect 33428 25200 33598 25256
rect 33654 25200 33659 25256
rect 33428 25198 33659 25200
rect 33428 25196 33434 25198
rect 33593 25195 33659 25198
rect 53465 25122 53531 25125
rect 55200 25122 56000 25152
rect 53465 25120 56000 25122
rect 53465 25064 53470 25120
rect 53526 25064 56000 25120
rect 53465 25062 56000 25064
rect 53465 25059 53531 25062
rect 19570 25056 19886 25057
rect 0 24986 800 25016
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 55200 25032 56000 25062
rect 50290 24991 50606 24992
rect 1577 24986 1643 24989
rect 0 24984 1643 24986
rect 0 24928 1582 24984
rect 1638 24928 1643 24984
rect 0 24926 1643 24928
rect 0 24896 800 24926
rect 1577 24923 1643 24926
rect 54201 24850 54267 24853
rect 55200 24850 56000 24880
rect 54201 24848 56000 24850
rect 54201 24792 54206 24848
rect 54262 24792 56000 24848
rect 54201 24790 56000 24792
rect 54201 24787 54267 24790
rect 55200 24760 56000 24790
rect 4210 24512 4526 24513
rect 0 24442 800 24472
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 55200 24488 56000 24608
rect 34930 24447 35246 24448
rect 1669 24442 1735 24445
rect 0 24440 1735 24442
rect 0 24384 1674 24440
rect 1730 24384 1735 24440
rect 0 24382 1735 24384
rect 0 24352 800 24382
rect 1669 24379 1735 24382
rect 53465 24306 53531 24309
rect 55200 24306 56000 24336
rect 53465 24304 56000 24306
rect 53465 24248 53470 24304
rect 53526 24248 56000 24304
rect 53465 24246 56000 24248
rect 53465 24243 53531 24246
rect 55200 24216 56000 24246
rect 33501 24034 33567 24037
rect 35433 24034 35499 24037
rect 33501 24032 35499 24034
rect 33501 23976 33506 24032
rect 33562 23976 35438 24032
rect 35494 23976 35499 24032
rect 33501 23974 35499 23976
rect 33501 23971 33567 23974
rect 35433 23971 35499 23974
rect 54201 24034 54267 24037
rect 55200 24034 56000 24064
rect 54201 24032 56000 24034
rect 54201 23976 54206 24032
rect 54262 23976 56000 24032
rect 54201 23974 56000 23976
rect 54201 23971 54267 23974
rect 19570 23968 19886 23969
rect 0 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 55200 23944 56000 23974
rect 50290 23903 50606 23904
rect 1669 23898 1735 23901
rect 0 23896 1735 23898
rect 0 23840 1674 23896
rect 1730 23840 1735 23896
rect 0 23838 1735 23840
rect 0 23808 800 23838
rect 1669 23835 1735 23838
rect 31753 23898 31819 23901
rect 33501 23898 33567 23901
rect 36261 23898 36327 23901
rect 31753 23896 36327 23898
rect 31753 23840 31758 23896
rect 31814 23840 33506 23896
rect 33562 23840 36266 23896
rect 36322 23840 36327 23896
rect 31753 23838 36327 23840
rect 31753 23835 31819 23838
rect 33501 23835 33567 23838
rect 36261 23835 36327 23838
rect 55200 23672 56000 23792
rect 34094 23428 34100 23492
rect 34164 23490 34170 23492
rect 34329 23490 34395 23493
rect 34164 23488 34395 23490
rect 34164 23432 34334 23488
rect 34390 23432 34395 23488
rect 34164 23430 34395 23432
rect 34164 23428 34170 23430
rect 34329 23427 34395 23430
rect 54201 23490 54267 23493
rect 55200 23490 56000 23520
rect 54201 23488 56000 23490
rect 54201 23432 54206 23488
rect 54262 23432 56000 23488
rect 54201 23430 56000 23432
rect 54201 23427 54267 23430
rect 4210 23424 4526 23425
rect 0 23354 800 23384
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 55200 23400 56000 23430
rect 34930 23359 35246 23360
rect 1669 23354 1735 23357
rect 0 23352 1735 23354
rect 0 23296 1674 23352
rect 1730 23296 1735 23352
rect 0 23294 1735 23296
rect 0 23264 800 23294
rect 1669 23291 1735 23294
rect 53557 23218 53623 23221
rect 55200 23218 56000 23248
rect 53557 23216 56000 23218
rect 53557 23160 53562 23216
rect 53618 23160 56000 23216
rect 53557 23158 56000 23160
rect 53557 23155 53623 23158
rect 55200 23128 56000 23158
rect 19570 22880 19886 22881
rect 0 22810 800 22840
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 55200 22856 56000 22976
rect 50290 22815 50606 22816
rect 1669 22810 1735 22813
rect 0 22808 1735 22810
rect 0 22752 1674 22808
rect 1730 22752 1735 22808
rect 0 22750 1735 22752
rect 0 22720 800 22750
rect 1669 22747 1735 22750
rect 35525 22810 35591 22813
rect 38561 22810 38627 22813
rect 35525 22808 38627 22810
rect 35525 22752 35530 22808
rect 35586 22752 38566 22808
rect 38622 22752 38627 22808
rect 35525 22750 38627 22752
rect 35525 22747 35591 22750
rect 38561 22747 38627 22750
rect 54201 22674 54267 22677
rect 55200 22674 56000 22704
rect 54201 22672 56000 22674
rect 54201 22616 54206 22672
rect 54262 22616 56000 22672
rect 54201 22614 56000 22616
rect 54201 22611 54267 22614
rect 55200 22584 56000 22614
rect 54201 22402 54267 22405
rect 55200 22402 56000 22432
rect 54201 22400 56000 22402
rect 54201 22344 54206 22400
rect 54262 22344 56000 22400
rect 54201 22342 56000 22344
rect 54201 22339 54267 22342
rect 4210 22336 4526 22337
rect 0 22266 800 22296
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 55200 22312 56000 22342
rect 34930 22271 35246 22272
rect 1669 22266 1735 22269
rect 0 22264 1735 22266
rect 0 22208 1674 22264
rect 1730 22208 1735 22264
rect 0 22206 1735 22208
rect 0 22176 800 22206
rect 1669 22203 1735 22206
rect 38653 22266 38719 22269
rect 43345 22266 43411 22269
rect 38653 22264 43411 22266
rect 38653 22208 38658 22264
rect 38714 22208 43350 22264
rect 43406 22208 43411 22264
rect 38653 22206 43411 22208
rect 38653 22203 38719 22206
rect 43345 22203 43411 22206
rect 33225 22130 33291 22133
rect 36905 22130 36971 22133
rect 33225 22128 36971 22130
rect 33225 22072 33230 22128
rect 33286 22072 36910 22128
rect 36966 22072 36971 22128
rect 33225 22070 36971 22072
rect 33225 22067 33291 22070
rect 36905 22067 36971 22070
rect 55200 22040 56000 22160
rect 54017 21994 54083 21997
rect 31710 21992 54083 21994
rect 31710 21936 54022 21992
rect 54078 21936 54083 21992
rect 31710 21934 54083 21936
rect 23105 21858 23171 21861
rect 31385 21858 31451 21861
rect 31710 21858 31770 21934
rect 54017 21931 54083 21934
rect 23105 21856 31770 21858
rect 23105 21800 23110 21856
rect 23166 21800 31390 21856
rect 31446 21800 31770 21856
rect 23105 21798 31770 21800
rect 54201 21858 54267 21861
rect 55200 21858 56000 21888
rect 54201 21856 56000 21858
rect 54201 21800 54206 21856
rect 54262 21800 56000 21856
rect 54201 21798 56000 21800
rect 23105 21795 23171 21798
rect 31385 21795 31451 21798
rect 54201 21795 54267 21798
rect 19570 21792 19886 21793
rect 0 21722 800 21752
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 55200 21768 56000 21798
rect 50290 21727 50606 21728
rect 1669 21722 1735 21725
rect 0 21720 1735 21722
rect 0 21664 1674 21720
rect 1730 21664 1735 21720
rect 0 21662 1735 21664
rect 0 21632 800 21662
rect 1669 21659 1735 21662
rect 27429 21586 27495 21589
rect 53281 21586 53347 21589
rect 27429 21584 53347 21586
rect 27429 21528 27434 21584
rect 27490 21528 53286 21584
rect 53342 21528 53347 21584
rect 27429 21526 53347 21528
rect 27429 21523 27495 21526
rect 53281 21523 53347 21526
rect 53465 21586 53531 21589
rect 55200 21586 56000 21616
rect 53465 21584 56000 21586
rect 53465 21528 53470 21584
rect 53526 21528 56000 21584
rect 53465 21526 56000 21528
rect 53465 21523 53531 21526
rect 55200 21496 56000 21526
rect 28625 21450 28691 21453
rect 28758 21450 28764 21452
rect 28625 21448 28764 21450
rect 28625 21392 28630 21448
rect 28686 21392 28764 21448
rect 28625 21390 28764 21392
rect 28625 21387 28691 21390
rect 28758 21388 28764 21390
rect 28828 21388 28834 21452
rect 30465 21450 30531 21453
rect 37641 21450 37707 21453
rect 30465 21448 37707 21450
rect 30465 21392 30470 21448
rect 30526 21392 37646 21448
rect 37702 21392 37707 21448
rect 30465 21390 37707 21392
rect 30465 21387 30531 21390
rect 37641 21387 37707 21390
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 55200 21224 56000 21344
rect 34930 21183 35246 21184
rect 1669 21178 1735 21181
rect 0 21176 1735 21178
rect 0 21120 1674 21176
rect 1730 21120 1735 21176
rect 0 21118 1735 21120
rect 0 21088 800 21118
rect 1669 21115 1735 21118
rect 23565 21042 23631 21045
rect 26509 21042 26575 21045
rect 23565 21040 26575 21042
rect 23565 20984 23570 21040
rect 23626 20984 26514 21040
rect 26570 20984 26575 21040
rect 23565 20982 26575 20984
rect 23565 20979 23631 20982
rect 26509 20979 26575 20982
rect 54201 21042 54267 21045
rect 55200 21042 56000 21072
rect 54201 21040 56000 21042
rect 54201 20984 54206 21040
rect 54262 20984 56000 21040
rect 54201 20982 56000 20984
rect 54201 20979 54267 20982
rect 55200 20952 56000 20982
rect 38745 20906 38811 20909
rect 43989 20906 44055 20909
rect 38745 20904 44055 20906
rect 38745 20848 38750 20904
rect 38806 20848 43994 20904
rect 44050 20848 44055 20904
rect 38745 20846 44055 20848
rect 38745 20843 38811 20846
rect 43989 20843 44055 20846
rect 53557 20770 53623 20773
rect 54201 20770 54267 20773
rect 55200 20770 56000 20800
rect 53557 20768 56000 20770
rect 53557 20712 53562 20768
rect 53618 20712 54206 20768
rect 54262 20712 56000 20768
rect 53557 20710 56000 20712
rect 53557 20707 53623 20710
rect 54201 20707 54267 20710
rect 19570 20704 19886 20705
rect 0 20634 800 20664
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 55200 20680 56000 20710
rect 50290 20639 50606 20640
rect 1669 20634 1735 20637
rect 0 20632 1735 20634
rect 0 20576 1674 20632
rect 1730 20576 1735 20632
rect 0 20574 1735 20576
rect 0 20544 800 20574
rect 1669 20571 1735 20574
rect 29494 20572 29500 20636
rect 29564 20634 29570 20636
rect 29821 20634 29887 20637
rect 29564 20632 29887 20634
rect 29564 20576 29826 20632
rect 29882 20576 29887 20632
rect 29564 20574 29887 20576
rect 29564 20572 29570 20574
rect 29821 20571 29887 20574
rect 24393 20498 24459 20501
rect 53281 20498 53347 20501
rect 24393 20496 53347 20498
rect 24393 20440 24398 20496
rect 24454 20440 53286 20496
rect 53342 20440 53347 20496
rect 24393 20438 53347 20440
rect 24393 20435 24459 20438
rect 53281 20435 53347 20438
rect 55200 20408 56000 20528
rect 27521 20362 27587 20365
rect 28809 20362 28875 20365
rect 27521 20360 28875 20362
rect 27521 20304 27526 20360
rect 27582 20304 28814 20360
rect 28870 20304 28875 20360
rect 27521 20302 28875 20304
rect 27521 20299 27587 20302
rect 28809 20299 28875 20302
rect 54201 20226 54267 20229
rect 55200 20226 56000 20256
rect 54201 20224 56000 20226
rect 54201 20168 54206 20224
rect 54262 20168 56000 20224
rect 54201 20166 56000 20168
rect 54201 20163 54267 20166
rect 4210 20160 4526 20161
rect 0 20090 800 20120
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 55200 20136 56000 20166
rect 34930 20095 35246 20096
rect 1669 20090 1735 20093
rect 0 20088 1735 20090
rect 0 20032 1674 20088
rect 1730 20032 1735 20088
rect 0 20030 1735 20032
rect 0 20000 800 20030
rect 1669 20027 1735 20030
rect 35525 20090 35591 20093
rect 37457 20090 37523 20093
rect 35525 20088 37523 20090
rect 35525 20032 35530 20088
rect 35586 20032 37462 20088
rect 37518 20032 37523 20088
rect 35525 20030 37523 20032
rect 35525 20027 35591 20030
rect 37457 20027 37523 20030
rect 29453 19954 29519 19957
rect 38101 19954 38167 19957
rect 29453 19952 38167 19954
rect 29453 19896 29458 19952
rect 29514 19896 38106 19952
rect 38162 19896 38167 19952
rect 29453 19894 38167 19896
rect 29453 19891 29519 19894
rect 38101 19891 38167 19894
rect 53557 19954 53623 19957
rect 55200 19954 56000 19984
rect 53557 19952 56000 19954
rect 53557 19896 53562 19952
rect 53618 19896 56000 19952
rect 53557 19894 56000 19896
rect 53557 19891 53623 19894
rect 55200 19864 56000 19894
rect 30281 19818 30347 19821
rect 31017 19818 31083 19821
rect 30281 19816 31083 19818
rect 30281 19760 30286 19816
rect 30342 19760 31022 19816
rect 31078 19760 31083 19816
rect 30281 19758 31083 19760
rect 30281 19755 30347 19758
rect 31017 19755 31083 19758
rect 36261 19818 36327 19821
rect 38469 19818 38535 19821
rect 36261 19816 38535 19818
rect 36261 19760 36266 19816
rect 36322 19760 38474 19816
rect 38530 19760 38535 19816
rect 36261 19758 38535 19760
rect 36261 19755 36327 19758
rect 38469 19755 38535 19758
rect 30281 19682 30347 19685
rect 32121 19682 32187 19685
rect 30281 19680 32187 19682
rect 30281 19624 30286 19680
rect 30342 19624 32126 19680
rect 32182 19624 32187 19680
rect 30281 19622 32187 19624
rect 30281 19619 30347 19622
rect 32121 19619 32187 19622
rect 19570 19616 19886 19617
rect 0 19546 800 19576
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 55200 19592 56000 19712
rect 50290 19551 50606 19552
rect 1669 19546 1735 19549
rect 0 19544 1735 19546
rect 0 19488 1674 19544
rect 1730 19488 1735 19544
rect 0 19486 1735 19488
rect 0 19456 800 19486
rect 1669 19483 1735 19486
rect 28349 19546 28415 19549
rect 37181 19546 37247 19549
rect 28349 19544 37247 19546
rect 28349 19488 28354 19544
rect 28410 19488 37186 19544
rect 37242 19488 37247 19544
rect 28349 19486 37247 19488
rect 28349 19483 28415 19486
rect 37181 19483 37247 19486
rect 40125 19546 40191 19549
rect 41505 19546 41571 19549
rect 40125 19544 41571 19546
rect 40125 19488 40130 19544
rect 40186 19488 41510 19544
rect 41566 19488 41571 19544
rect 40125 19486 41571 19488
rect 40125 19483 40191 19486
rect 41505 19483 41571 19486
rect 54201 19410 54267 19413
rect 55200 19410 56000 19440
rect 54201 19408 56000 19410
rect 28625 19350 28691 19353
rect 28582 19348 28691 19350
rect 28582 19292 28630 19348
rect 28686 19292 28691 19348
rect 54201 19352 54206 19408
rect 54262 19352 56000 19408
rect 54201 19350 56000 19352
rect 54201 19347 54267 19350
rect 55200 19320 56000 19350
rect 28582 19287 28691 19292
rect 4210 19072 4526 19073
rect 0 19002 800 19032
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 1669 19002 1735 19005
rect 0 19000 1735 19002
rect 0 18944 1674 19000
rect 1730 18944 1735 19000
rect 0 18942 1735 18944
rect 0 18912 800 18942
rect 1669 18939 1735 18942
rect 28582 18866 28642 19287
rect 37549 19274 37615 19277
rect 38285 19276 38351 19277
rect 38285 19274 38332 19276
rect 37549 19272 38332 19274
rect 37549 19216 37554 19272
rect 37610 19216 38290 19272
rect 37549 19214 38332 19216
rect 37549 19211 37615 19214
rect 38285 19212 38332 19214
rect 38396 19212 38402 19276
rect 38285 19211 38351 19212
rect 54201 19138 54267 19141
rect 55200 19138 56000 19168
rect 54201 19136 56000 19138
rect 54201 19080 54206 19136
rect 54262 19080 56000 19136
rect 54201 19078 56000 19080
rect 54201 19075 54267 19078
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 55200 19048 56000 19078
rect 34930 19007 35246 19008
rect 28717 18866 28783 18869
rect 28582 18864 28783 18866
rect 28582 18808 28722 18864
rect 28778 18808 28783 18864
rect 28582 18806 28783 18808
rect 28717 18803 28783 18806
rect 55200 18776 56000 18896
rect 32029 18730 32095 18733
rect 38285 18730 38351 18733
rect 32029 18728 38351 18730
rect 32029 18672 32034 18728
rect 32090 18672 38290 18728
rect 38346 18672 38351 18728
rect 32029 18670 38351 18672
rect 32029 18667 32095 18670
rect 38285 18667 38351 18670
rect 30833 18594 30899 18597
rect 30966 18594 30972 18596
rect 30833 18592 30972 18594
rect 30833 18536 30838 18592
rect 30894 18536 30972 18592
rect 30833 18534 30972 18536
rect 30833 18531 30899 18534
rect 30966 18532 30972 18534
rect 31036 18532 31042 18596
rect 54201 18594 54267 18597
rect 55200 18594 56000 18624
rect 54201 18592 56000 18594
rect 54201 18536 54206 18592
rect 54262 18536 56000 18592
rect 54201 18534 56000 18536
rect 54201 18531 54267 18534
rect 19570 18528 19886 18529
rect 0 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 55200 18504 56000 18534
rect 50290 18463 50606 18464
rect 1669 18458 1735 18461
rect 0 18456 1735 18458
rect 0 18400 1674 18456
rect 1730 18400 1735 18456
rect 0 18398 1735 18400
rect 0 18368 800 18398
rect 1669 18395 1735 18398
rect 31385 18458 31451 18461
rect 34973 18458 35039 18461
rect 31385 18456 35039 18458
rect 31385 18400 31390 18456
rect 31446 18400 34978 18456
rect 35034 18400 35039 18456
rect 31385 18398 35039 18400
rect 31385 18395 31451 18398
rect 34973 18395 35039 18398
rect 28349 18322 28415 18325
rect 29085 18322 29151 18325
rect 30005 18322 30071 18325
rect 28349 18320 30071 18322
rect 28349 18264 28354 18320
rect 28410 18264 29090 18320
rect 29146 18264 30010 18320
rect 30066 18264 30071 18320
rect 28349 18262 30071 18264
rect 28349 18259 28415 18262
rect 29085 18259 29151 18262
rect 30005 18259 30071 18262
rect 30741 18322 30807 18325
rect 31753 18322 31819 18325
rect 30741 18320 31819 18322
rect 30741 18264 30746 18320
rect 30802 18264 31758 18320
rect 31814 18264 31819 18320
rect 30741 18262 31819 18264
rect 30741 18259 30807 18262
rect 31753 18259 31819 18262
rect 34697 18322 34763 18325
rect 38101 18322 38167 18325
rect 34697 18320 38167 18322
rect 34697 18264 34702 18320
rect 34758 18264 38106 18320
rect 38162 18264 38167 18320
rect 34697 18262 38167 18264
rect 34697 18259 34763 18262
rect 38101 18259 38167 18262
rect 38561 18322 38627 18325
rect 41689 18322 41755 18325
rect 38561 18320 41755 18322
rect 38561 18264 38566 18320
rect 38622 18264 41694 18320
rect 41750 18264 41755 18320
rect 38561 18262 41755 18264
rect 38561 18259 38627 18262
rect 41689 18259 41755 18262
rect 53465 18322 53531 18325
rect 55200 18322 56000 18352
rect 53465 18320 56000 18322
rect 53465 18264 53470 18320
rect 53526 18264 56000 18320
rect 53465 18262 56000 18264
rect 53465 18259 53531 18262
rect 55200 18232 56000 18262
rect 38285 18186 38351 18189
rect 39297 18186 39363 18189
rect 40493 18186 40559 18189
rect 38285 18184 40559 18186
rect 38285 18128 38290 18184
rect 38346 18128 39302 18184
rect 39358 18128 40498 18184
rect 40554 18128 40559 18184
rect 38285 18126 40559 18128
rect 38285 18123 38351 18126
rect 39297 18123 39363 18126
rect 40493 18123 40559 18126
rect 4210 17984 4526 17985
rect 0 17914 800 17944
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 55200 17960 56000 18080
rect 34930 17919 35246 17920
rect 1577 17914 1643 17917
rect 0 17912 1643 17914
rect 0 17856 1582 17912
rect 1638 17856 1643 17912
rect 0 17854 1643 17856
rect 0 17824 800 17854
rect 1577 17851 1643 17854
rect 18229 17778 18295 17781
rect 19057 17778 19123 17781
rect 25037 17778 25103 17781
rect 18229 17776 25103 17778
rect 18229 17720 18234 17776
rect 18290 17720 19062 17776
rect 19118 17720 25042 17776
rect 25098 17720 25103 17776
rect 18229 17718 25103 17720
rect 18229 17715 18295 17718
rect 19057 17715 19123 17718
rect 25037 17715 25103 17718
rect 27705 17778 27771 17781
rect 27838 17778 27844 17780
rect 27705 17776 27844 17778
rect 27705 17720 27710 17776
rect 27766 17720 27844 17776
rect 27705 17718 27844 17720
rect 27705 17715 27771 17718
rect 27838 17716 27844 17718
rect 27908 17778 27914 17780
rect 29310 17778 29316 17780
rect 27908 17718 29316 17778
rect 27908 17716 27914 17718
rect 29310 17716 29316 17718
rect 29380 17716 29386 17780
rect 31109 17778 31175 17781
rect 31385 17778 31451 17781
rect 37825 17778 37891 17781
rect 31109 17776 37891 17778
rect 31109 17720 31114 17776
rect 31170 17720 31390 17776
rect 31446 17720 37830 17776
rect 37886 17720 37891 17776
rect 31109 17718 37891 17720
rect 31109 17715 31175 17718
rect 31385 17715 31451 17718
rect 37825 17715 37891 17718
rect 54201 17778 54267 17781
rect 55200 17778 56000 17808
rect 54201 17776 56000 17778
rect 54201 17720 54206 17776
rect 54262 17720 56000 17776
rect 54201 17718 56000 17720
rect 54201 17715 54267 17718
rect 55200 17688 56000 17718
rect 25129 17642 25195 17645
rect 28901 17642 28967 17645
rect 25129 17640 28967 17642
rect 25129 17584 25134 17640
rect 25190 17584 28906 17640
rect 28962 17584 28967 17640
rect 25129 17582 28967 17584
rect 25129 17579 25195 17582
rect 28901 17579 28967 17582
rect 32397 17642 32463 17645
rect 40217 17642 40283 17645
rect 32397 17640 40283 17642
rect 32397 17584 32402 17640
rect 32458 17584 40222 17640
rect 40278 17584 40283 17640
rect 32397 17582 40283 17584
rect 32397 17579 32463 17582
rect 40217 17579 40283 17582
rect 24025 17506 24091 17509
rect 27981 17506 28047 17509
rect 24025 17504 28047 17506
rect 24025 17448 24030 17504
rect 24086 17448 27986 17504
rect 28042 17448 28047 17504
rect 24025 17446 28047 17448
rect 24025 17443 24091 17446
rect 27981 17443 28047 17446
rect 36077 17506 36143 17509
rect 37917 17506 37983 17509
rect 36077 17504 37983 17506
rect 36077 17448 36082 17504
rect 36138 17448 37922 17504
rect 37978 17448 37983 17504
rect 36077 17446 37983 17448
rect 36077 17443 36143 17446
rect 37917 17443 37983 17446
rect 54201 17506 54267 17509
rect 55200 17506 56000 17536
rect 54201 17504 56000 17506
rect 54201 17448 54206 17504
rect 54262 17448 56000 17504
rect 54201 17446 56000 17448
rect 54201 17443 54267 17446
rect 19570 17440 19886 17441
rect 0 17370 800 17400
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 55200 17416 56000 17446
rect 50290 17375 50606 17376
rect 1669 17370 1735 17373
rect 0 17368 1735 17370
rect 0 17312 1674 17368
rect 1730 17312 1735 17368
rect 0 17310 1735 17312
rect 0 17280 800 17310
rect 1669 17307 1735 17310
rect 28625 17370 28691 17373
rect 28809 17370 28875 17373
rect 28625 17368 28875 17370
rect 28625 17312 28630 17368
rect 28686 17312 28814 17368
rect 28870 17312 28875 17368
rect 28625 17310 28875 17312
rect 28625 17307 28691 17310
rect 28809 17307 28875 17310
rect 24669 17234 24735 17237
rect 27429 17234 27495 17237
rect 24669 17232 27495 17234
rect 24669 17176 24674 17232
rect 24730 17176 27434 17232
rect 27490 17176 27495 17232
rect 24669 17174 27495 17176
rect 24669 17171 24735 17174
rect 27429 17171 27495 17174
rect 55200 17144 56000 17264
rect 33501 17098 33567 17101
rect 34421 17098 34487 17101
rect 35525 17098 35591 17101
rect 33501 17096 35591 17098
rect 33501 17040 33506 17096
rect 33562 17040 34426 17096
rect 34482 17040 35530 17096
rect 35586 17040 35591 17096
rect 33501 17038 35591 17040
rect 33501 17035 33567 17038
rect 34421 17035 34487 17038
rect 35525 17035 35591 17038
rect 54201 16962 54267 16965
rect 55200 16962 56000 16992
rect 54201 16960 56000 16962
rect 54201 16904 54206 16960
rect 54262 16904 56000 16960
rect 54201 16902 56000 16904
rect 54201 16899 54267 16902
rect 4210 16896 4526 16897
rect 0 16826 800 16856
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 55200 16872 56000 16902
rect 34930 16831 35246 16832
rect 1669 16826 1735 16829
rect 0 16824 1735 16826
rect 0 16768 1674 16824
rect 1730 16768 1735 16824
rect 0 16766 1735 16768
rect 0 16736 800 16766
rect 1669 16763 1735 16766
rect 23105 16826 23171 16829
rect 26233 16826 26299 16829
rect 23105 16824 26299 16826
rect 23105 16768 23110 16824
rect 23166 16768 26238 16824
rect 26294 16768 26299 16824
rect 23105 16766 26299 16768
rect 23105 16763 23171 16766
rect 26233 16763 26299 16766
rect 39389 16826 39455 16829
rect 40861 16826 40927 16829
rect 39389 16824 40927 16826
rect 39389 16768 39394 16824
rect 39450 16768 40866 16824
rect 40922 16768 40927 16824
rect 39389 16766 40927 16768
rect 39389 16763 39455 16766
rect 40861 16763 40927 16766
rect 41229 16826 41295 16829
rect 41505 16826 41571 16829
rect 41229 16824 41571 16826
rect 41229 16768 41234 16824
rect 41290 16768 41510 16824
rect 41566 16768 41571 16824
rect 41229 16766 41571 16768
rect 41229 16763 41295 16766
rect 41505 16763 41571 16766
rect 16757 16690 16823 16693
rect 20253 16690 20319 16693
rect 25037 16690 25103 16693
rect 53281 16690 53347 16693
rect 16757 16688 53347 16690
rect 16757 16632 16762 16688
rect 16818 16632 20258 16688
rect 20314 16632 25042 16688
rect 25098 16632 53286 16688
rect 53342 16632 53347 16688
rect 16757 16630 53347 16632
rect 16757 16627 16823 16630
rect 20253 16627 20319 16630
rect 25037 16627 25103 16630
rect 53281 16627 53347 16630
rect 53557 16690 53623 16693
rect 55200 16690 56000 16720
rect 53557 16688 56000 16690
rect 53557 16632 53562 16688
rect 53618 16632 56000 16688
rect 53557 16630 56000 16632
rect 53557 16627 53623 16630
rect 55200 16600 56000 16630
rect 40401 16554 40467 16557
rect 42517 16554 42583 16557
rect 40401 16552 42583 16554
rect 40401 16496 40406 16552
rect 40462 16496 42522 16552
rect 42578 16496 42583 16552
rect 40401 16494 42583 16496
rect 40401 16491 40467 16494
rect 42517 16491 42583 16494
rect 19570 16352 19886 16353
rect 0 16282 800 16312
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 55200 16328 56000 16448
rect 50290 16287 50606 16288
rect 1669 16282 1735 16285
rect 0 16280 1735 16282
rect 0 16224 1674 16280
rect 1730 16224 1735 16280
rect 0 16222 1735 16224
rect 0 16192 800 16222
rect 1669 16219 1735 16222
rect 28993 16282 29059 16285
rect 35157 16282 35223 16285
rect 28993 16280 35223 16282
rect 28993 16224 28998 16280
rect 29054 16224 35162 16280
rect 35218 16224 35223 16280
rect 28993 16222 35223 16224
rect 28993 16219 29059 16222
rect 35157 16219 35223 16222
rect 15101 16146 15167 16149
rect 20897 16146 20963 16149
rect 15101 16144 20963 16146
rect 15101 16088 15106 16144
rect 15162 16088 20902 16144
rect 20958 16088 20963 16144
rect 15101 16086 20963 16088
rect 15101 16083 15167 16086
rect 20897 16083 20963 16086
rect 31293 16146 31359 16149
rect 32489 16146 32555 16149
rect 37825 16146 37891 16149
rect 31293 16144 37891 16146
rect 31293 16088 31298 16144
rect 31354 16088 32494 16144
rect 32550 16088 37830 16144
rect 37886 16088 37891 16144
rect 31293 16086 37891 16088
rect 31293 16083 31359 16086
rect 32489 16083 32555 16086
rect 37825 16083 37891 16086
rect 54201 16146 54267 16149
rect 55200 16146 56000 16176
rect 54201 16144 56000 16146
rect 54201 16088 54206 16144
rect 54262 16088 56000 16144
rect 54201 16086 56000 16088
rect 54201 16083 54267 16086
rect 55200 16056 56000 16086
rect 15561 16010 15627 16013
rect 17401 16010 17467 16013
rect 15561 16008 17467 16010
rect 15561 15952 15566 16008
rect 15622 15952 17406 16008
rect 17462 15952 17467 16008
rect 15561 15950 17467 15952
rect 15561 15947 15627 15950
rect 17401 15947 17467 15950
rect 32305 16010 32371 16013
rect 36905 16010 36971 16013
rect 43713 16010 43779 16013
rect 32305 16008 35404 16010
rect 32305 15952 32310 16008
rect 32366 15952 35404 16008
rect 32305 15950 35404 15952
rect 32305 15947 32371 15950
rect 35344 15874 35404 15950
rect 36905 16008 43779 16010
rect 36905 15952 36910 16008
rect 36966 15952 43718 16008
rect 43774 15952 43779 16008
rect 36905 15950 43779 15952
rect 36905 15947 36971 15950
rect 43713 15947 43779 15950
rect 41597 15874 41663 15877
rect 42609 15874 42675 15877
rect 35344 15872 42675 15874
rect 35344 15816 41602 15872
rect 41658 15816 42614 15872
rect 42670 15816 42675 15872
rect 35344 15814 42675 15816
rect 41597 15811 41663 15814
rect 42609 15811 42675 15814
rect 54201 15874 54267 15877
rect 55200 15874 56000 15904
rect 54201 15872 56000 15874
rect 54201 15816 54206 15872
rect 54262 15816 56000 15872
rect 54201 15814 56000 15816
rect 54201 15811 54267 15814
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 55200 15784 56000 15814
rect 34930 15743 35246 15744
rect 1669 15738 1735 15741
rect 0 15736 1735 15738
rect 0 15680 1674 15736
rect 1730 15680 1735 15736
rect 0 15678 1735 15680
rect 0 15648 800 15678
rect 1669 15675 1735 15678
rect 26918 15540 26924 15604
rect 26988 15602 26994 15604
rect 28073 15602 28139 15605
rect 26988 15600 28139 15602
rect 26988 15544 28078 15600
rect 28134 15544 28139 15600
rect 26988 15542 28139 15544
rect 26988 15540 26994 15542
rect 28073 15539 28139 15542
rect 41413 15602 41479 15605
rect 44449 15602 44515 15605
rect 41413 15600 44515 15602
rect 41413 15544 41418 15600
rect 41474 15544 44454 15600
rect 44510 15544 44515 15600
rect 41413 15542 44515 15544
rect 41413 15539 41479 15542
rect 44449 15539 44515 15542
rect 55200 15512 56000 15632
rect 14733 15466 14799 15469
rect 20805 15466 20871 15469
rect 21449 15466 21515 15469
rect 14733 15464 21515 15466
rect 14733 15408 14738 15464
rect 14794 15408 20810 15464
rect 20866 15408 21454 15464
rect 21510 15408 21515 15464
rect 14733 15406 21515 15408
rect 14733 15403 14799 15406
rect 20805 15403 20871 15406
rect 21449 15403 21515 15406
rect 39389 15466 39455 15469
rect 42977 15466 43043 15469
rect 39389 15464 43043 15466
rect 39389 15408 39394 15464
rect 39450 15408 42982 15464
rect 43038 15408 43043 15464
rect 39389 15406 43043 15408
rect 39389 15403 39455 15406
rect 42977 15403 43043 15406
rect 25998 15268 26004 15332
rect 26068 15330 26074 15332
rect 27705 15330 27771 15333
rect 26068 15328 27771 15330
rect 26068 15272 27710 15328
rect 27766 15272 27771 15328
rect 26068 15270 27771 15272
rect 26068 15268 26074 15270
rect 27705 15267 27771 15270
rect 30465 15330 30531 15333
rect 38285 15330 38351 15333
rect 30465 15328 38351 15330
rect 30465 15272 30470 15328
rect 30526 15272 38290 15328
rect 38346 15272 38351 15328
rect 30465 15270 38351 15272
rect 30465 15267 30531 15270
rect 38285 15267 38351 15270
rect 54201 15330 54267 15333
rect 55200 15330 56000 15360
rect 54201 15328 56000 15330
rect 54201 15272 54206 15328
rect 54262 15272 56000 15328
rect 54201 15270 56000 15272
rect 54201 15267 54267 15270
rect 19570 15264 19886 15265
rect 0 15194 800 15224
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 55200 15240 56000 15270
rect 50290 15199 50606 15200
rect 1669 15194 1735 15197
rect 0 15192 1735 15194
rect 0 15136 1674 15192
rect 1730 15136 1735 15192
rect 0 15134 1735 15136
rect 0 15104 800 15134
rect 1669 15131 1735 15134
rect 25814 15132 25820 15196
rect 25884 15194 25890 15196
rect 26049 15194 26115 15197
rect 28257 15194 28323 15197
rect 30557 15196 30623 15197
rect 30557 15194 30604 15196
rect 25884 15192 28323 15194
rect 25884 15136 26054 15192
rect 26110 15136 28262 15192
rect 28318 15136 28323 15192
rect 25884 15134 28323 15136
rect 30512 15192 30604 15194
rect 30512 15136 30562 15192
rect 30512 15134 30604 15136
rect 25884 15132 25890 15134
rect 26049 15131 26115 15134
rect 28257 15131 28323 15134
rect 30557 15132 30604 15134
rect 30668 15132 30674 15196
rect 30557 15131 30623 15132
rect 14733 15058 14799 15061
rect 21909 15058 21975 15061
rect 23749 15058 23815 15061
rect 37273 15058 37339 15061
rect 14733 15056 37339 15058
rect 14733 15000 14738 15056
rect 14794 15000 21914 15056
rect 21970 15000 23754 15056
rect 23810 15000 37278 15056
rect 37334 15000 37339 15056
rect 14733 14998 37339 15000
rect 14733 14995 14799 14998
rect 21909 14995 21975 14998
rect 23749 14995 23815 14998
rect 37273 14995 37339 14998
rect 53465 15058 53531 15061
rect 55200 15058 56000 15088
rect 53465 15056 56000 15058
rect 53465 15000 53470 15056
rect 53526 15000 56000 15056
rect 53465 14998 56000 15000
rect 53465 14995 53531 14998
rect 55200 14968 56000 14998
rect 25313 14922 25379 14925
rect 27613 14922 27679 14925
rect 25313 14920 27679 14922
rect 25313 14864 25318 14920
rect 25374 14864 27618 14920
rect 27674 14864 27679 14920
rect 25313 14862 27679 14864
rect 25313 14859 25379 14862
rect 27613 14859 27679 14862
rect 37457 14922 37523 14925
rect 54017 14922 54083 14925
rect 37457 14920 54083 14922
rect 37457 14864 37462 14920
rect 37518 14864 54022 14920
rect 54078 14864 54083 14920
rect 37457 14862 54083 14864
rect 37457 14859 37523 14862
rect 54017 14859 54083 14862
rect 4210 14720 4526 14721
rect 0 14650 800 14680
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 55200 14696 56000 14816
rect 34930 14655 35246 14656
rect 1669 14650 1735 14653
rect 0 14648 1735 14650
rect 0 14592 1674 14648
rect 1730 14592 1735 14648
rect 0 14590 1735 14592
rect 0 14560 800 14590
rect 1669 14587 1735 14590
rect 15101 14514 15167 14517
rect 20713 14514 20779 14517
rect 15101 14512 20779 14514
rect 15101 14456 15106 14512
rect 15162 14456 20718 14512
rect 20774 14456 20779 14512
rect 15101 14454 20779 14456
rect 15101 14451 15167 14454
rect 20713 14451 20779 14454
rect 29821 14514 29887 14517
rect 33685 14514 33751 14517
rect 29821 14512 33751 14514
rect 29821 14456 29826 14512
rect 29882 14456 33690 14512
rect 33746 14456 33751 14512
rect 29821 14454 33751 14456
rect 29821 14451 29887 14454
rect 33685 14451 33751 14454
rect 54201 14514 54267 14517
rect 55200 14514 56000 14544
rect 54201 14512 56000 14514
rect 54201 14456 54206 14512
rect 54262 14456 56000 14512
rect 54201 14454 56000 14456
rect 54201 14451 54267 14454
rect 55200 14424 56000 14454
rect 14641 14378 14707 14381
rect 18137 14378 18203 14381
rect 14641 14376 18203 14378
rect 14641 14320 14646 14376
rect 14702 14320 18142 14376
rect 18198 14320 18203 14376
rect 14641 14318 18203 14320
rect 14641 14315 14707 14318
rect 18137 14315 18203 14318
rect 38745 14378 38811 14381
rect 41965 14378 42031 14381
rect 38745 14376 42031 14378
rect 38745 14320 38750 14376
rect 38806 14320 41970 14376
rect 42026 14320 42031 14376
rect 38745 14318 42031 14320
rect 38745 14315 38811 14318
rect 41965 14315 42031 14318
rect 54201 14242 54267 14245
rect 55200 14242 56000 14272
rect 54201 14240 56000 14242
rect 54201 14184 54206 14240
rect 54262 14184 56000 14240
rect 54201 14182 56000 14184
rect 54201 14179 54267 14182
rect 19570 14176 19886 14177
rect 0 14106 800 14136
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 55200 14152 56000 14182
rect 50290 14111 50606 14112
rect 1669 14106 1735 14109
rect 0 14104 1735 14106
rect 0 14048 1674 14104
rect 1730 14048 1735 14104
rect 0 14046 1735 14048
rect 0 14016 800 14046
rect 1669 14043 1735 14046
rect 38745 14106 38811 14109
rect 39113 14106 39179 14109
rect 41413 14106 41479 14109
rect 38745 14104 41479 14106
rect 38745 14048 38750 14104
rect 38806 14048 39118 14104
rect 39174 14048 41418 14104
rect 41474 14048 41479 14104
rect 38745 14046 41479 14048
rect 38745 14043 38811 14046
rect 39113 14043 39179 14046
rect 41413 14043 41479 14046
rect 14457 13970 14523 13973
rect 19609 13970 19675 13973
rect 14457 13968 19675 13970
rect 14457 13912 14462 13968
rect 14518 13912 19614 13968
rect 19670 13912 19675 13968
rect 14457 13910 19675 13912
rect 14457 13907 14523 13910
rect 19609 13907 19675 13910
rect 38326 13908 38332 13972
rect 38396 13970 38402 13972
rect 40861 13970 40927 13973
rect 38396 13968 40927 13970
rect 38396 13912 40866 13968
rect 40922 13912 40927 13968
rect 38396 13910 40927 13912
rect 38396 13908 38402 13910
rect 40861 13907 40927 13910
rect 55200 13880 56000 14000
rect 30005 13834 30071 13837
rect 30189 13834 30255 13837
rect 40217 13834 40283 13837
rect 30005 13832 40283 13834
rect 30005 13776 30010 13832
rect 30066 13776 30194 13832
rect 30250 13776 40222 13832
rect 40278 13776 40283 13832
rect 30005 13774 40283 13776
rect 30005 13771 30071 13774
rect 30189 13771 30255 13774
rect 40217 13771 40283 13774
rect 32397 13698 32463 13701
rect 32622 13698 32628 13700
rect 32397 13696 32628 13698
rect 32397 13640 32402 13696
rect 32458 13640 32628 13696
rect 32397 13638 32628 13640
rect 32397 13635 32463 13638
rect 32622 13636 32628 13638
rect 32692 13636 32698 13700
rect 38193 13698 38259 13701
rect 41505 13698 41571 13701
rect 38193 13696 41571 13698
rect 38193 13640 38198 13696
rect 38254 13640 41510 13696
rect 41566 13640 41571 13696
rect 38193 13638 41571 13640
rect 38193 13635 38259 13638
rect 41505 13635 41571 13638
rect 54201 13698 54267 13701
rect 55200 13698 56000 13728
rect 54201 13696 56000 13698
rect 54201 13640 54206 13696
rect 54262 13640 56000 13696
rect 54201 13638 56000 13640
rect 54201 13635 54267 13638
rect 4210 13632 4526 13633
rect 0 13562 800 13592
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 55200 13608 56000 13638
rect 34930 13567 35246 13568
rect 1669 13562 1735 13565
rect 0 13560 1735 13562
rect 0 13504 1674 13560
rect 1730 13504 1735 13560
rect 0 13502 1735 13504
rect 0 13472 800 13502
rect 1669 13499 1735 13502
rect 14917 13562 14983 13565
rect 17585 13562 17651 13565
rect 14917 13560 17651 13562
rect 14917 13504 14922 13560
rect 14978 13504 17590 13560
rect 17646 13504 17651 13560
rect 14917 13502 17651 13504
rect 14917 13499 14983 13502
rect 17585 13499 17651 13502
rect 29545 13562 29611 13565
rect 33409 13562 33475 13565
rect 29545 13560 33475 13562
rect 29545 13504 29550 13560
rect 29606 13504 33414 13560
rect 33470 13504 33475 13560
rect 29545 13502 33475 13504
rect 29545 13499 29611 13502
rect 33409 13499 33475 13502
rect 39021 13426 39087 13429
rect 40033 13426 40099 13429
rect 39021 13424 40099 13426
rect 39021 13368 39026 13424
rect 39082 13368 40038 13424
rect 40094 13368 40099 13424
rect 39021 13366 40099 13368
rect 39021 13363 39087 13366
rect 40033 13363 40099 13366
rect 53557 13426 53623 13429
rect 55200 13426 56000 13456
rect 53557 13424 56000 13426
rect 53557 13368 53562 13424
rect 53618 13368 56000 13424
rect 53557 13366 56000 13368
rect 53557 13363 53623 13366
rect 55200 13336 56000 13366
rect 35525 13154 35591 13157
rect 36721 13154 36787 13157
rect 35525 13152 36787 13154
rect 35525 13096 35530 13152
rect 35586 13096 36726 13152
rect 36782 13096 36787 13152
rect 35525 13094 36787 13096
rect 35525 13091 35591 13094
rect 36721 13091 36787 13094
rect 19570 13088 19886 13089
rect 0 13018 800 13048
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 55200 13064 56000 13184
rect 50290 13023 50606 13024
rect 1669 13018 1735 13021
rect 0 13016 1735 13018
rect 0 12960 1674 13016
rect 1730 12960 1735 13016
rect 0 12958 1735 12960
rect 0 12928 800 12958
rect 1669 12955 1735 12958
rect 23013 12882 23079 12885
rect 27705 12882 27771 12885
rect 23013 12880 27771 12882
rect 23013 12824 23018 12880
rect 23074 12824 27710 12880
rect 27766 12824 27771 12880
rect 23013 12822 27771 12824
rect 23013 12819 23079 12822
rect 27705 12819 27771 12822
rect 31017 12882 31083 12885
rect 32581 12882 32647 12885
rect 31017 12880 32647 12882
rect 31017 12824 31022 12880
rect 31078 12824 32586 12880
rect 32642 12824 32647 12880
rect 31017 12822 32647 12824
rect 31017 12819 31083 12822
rect 32581 12819 32647 12822
rect 54201 12882 54267 12885
rect 55200 12882 56000 12912
rect 54201 12880 56000 12882
rect 54201 12824 54206 12880
rect 54262 12824 56000 12880
rect 54201 12822 56000 12824
rect 54201 12819 54267 12822
rect 55200 12792 56000 12822
rect 32397 12746 32463 12749
rect 32397 12744 40050 12746
rect 32397 12688 32402 12744
rect 32458 12688 40050 12744
rect 32397 12686 40050 12688
rect 32397 12683 32463 12686
rect 39990 12613 40050 12686
rect 39990 12608 40099 12613
rect 39990 12552 40038 12608
rect 40094 12552 40099 12608
rect 39990 12550 40099 12552
rect 40033 12547 40099 12550
rect 54201 12610 54267 12613
rect 55200 12610 56000 12640
rect 54201 12608 56000 12610
rect 54201 12552 54206 12608
rect 54262 12552 56000 12608
rect 54201 12550 56000 12552
rect 54201 12547 54267 12550
rect 4210 12544 4526 12545
rect 0 12474 800 12504
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 55200 12520 56000 12550
rect 34930 12479 35246 12480
rect 1669 12474 1735 12477
rect 0 12472 1735 12474
rect 0 12416 1674 12472
rect 1730 12416 1735 12472
rect 0 12414 1735 12416
rect 0 12384 800 12414
rect 1669 12411 1735 12414
rect 27889 12474 27955 12477
rect 30649 12474 30715 12477
rect 27889 12472 30715 12474
rect 27889 12416 27894 12472
rect 27950 12416 30654 12472
rect 30710 12416 30715 12472
rect 27889 12414 30715 12416
rect 27889 12411 27955 12414
rect 30649 12411 30715 12414
rect 19793 12338 19859 12341
rect 22185 12338 22251 12341
rect 19793 12336 22251 12338
rect 19793 12280 19798 12336
rect 19854 12280 22190 12336
rect 22246 12280 22251 12336
rect 19793 12278 22251 12280
rect 19793 12275 19859 12278
rect 22185 12275 22251 12278
rect 37733 12338 37799 12341
rect 46933 12338 46999 12341
rect 37733 12336 46999 12338
rect 37733 12280 37738 12336
rect 37794 12280 46938 12336
rect 46994 12280 46999 12336
rect 37733 12278 46999 12280
rect 37733 12275 37799 12278
rect 46933 12275 46999 12278
rect 55200 12248 56000 12368
rect 20069 12202 20135 12205
rect 26325 12202 26391 12205
rect 20069 12200 26391 12202
rect 20069 12144 20074 12200
rect 20130 12144 26330 12200
rect 26386 12144 26391 12200
rect 20069 12142 26391 12144
rect 20069 12139 20135 12142
rect 26325 12139 26391 12142
rect 34329 12202 34395 12205
rect 35341 12202 35407 12205
rect 34329 12200 35407 12202
rect 34329 12144 34334 12200
rect 34390 12144 35346 12200
rect 35402 12144 35407 12200
rect 34329 12142 35407 12144
rect 34329 12139 34395 12142
rect 35341 12139 35407 12142
rect 22185 12066 22251 12069
rect 27981 12066 28047 12069
rect 22185 12064 28047 12066
rect 22185 12008 22190 12064
rect 22246 12008 27986 12064
rect 28042 12008 28047 12064
rect 22185 12006 28047 12008
rect 22185 12003 22251 12006
rect 27981 12003 28047 12006
rect 54201 12066 54267 12069
rect 55200 12066 56000 12096
rect 54201 12064 56000 12066
rect 54201 12008 54206 12064
rect 54262 12008 56000 12064
rect 54201 12006 56000 12008
rect 54201 12003 54267 12006
rect 19570 12000 19886 12001
rect 0 11930 800 11960
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 55200 11976 56000 12006
rect 50290 11935 50606 11936
rect 1669 11930 1735 11933
rect 0 11928 1735 11930
rect 0 11872 1674 11928
rect 1730 11872 1735 11928
rect 0 11870 1735 11872
rect 0 11840 800 11870
rect 1669 11867 1735 11870
rect 29913 11794 29979 11797
rect 49693 11794 49759 11797
rect 29913 11792 49759 11794
rect 29913 11736 29918 11792
rect 29974 11736 49698 11792
rect 49754 11736 49759 11792
rect 29913 11734 49759 11736
rect 29913 11731 29979 11734
rect 49693 11731 49759 11734
rect 53465 11794 53531 11797
rect 55200 11794 56000 11824
rect 53465 11792 56000 11794
rect 53465 11736 53470 11792
rect 53526 11736 56000 11792
rect 53465 11734 56000 11736
rect 53465 11731 53531 11734
rect 55200 11704 56000 11734
rect 29085 11658 29151 11661
rect 29821 11658 29887 11661
rect 29085 11656 29887 11658
rect 29085 11600 29090 11656
rect 29146 11600 29826 11656
rect 29882 11600 29887 11656
rect 29085 11598 29887 11600
rect 29085 11595 29151 11598
rect 29821 11595 29887 11598
rect 4210 11456 4526 11457
rect 0 11386 800 11416
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 55200 11432 56000 11552
rect 34930 11391 35246 11392
rect 1669 11386 1735 11389
rect 0 11384 1735 11386
rect 0 11328 1674 11384
rect 1730 11328 1735 11384
rect 0 11326 1735 11328
rect 0 11296 800 11326
rect 1669 11323 1735 11326
rect 29085 11386 29151 11389
rect 29453 11386 29519 11389
rect 29085 11384 29519 11386
rect 29085 11328 29090 11384
rect 29146 11328 29458 11384
rect 29514 11328 29519 11384
rect 29085 11326 29519 11328
rect 29085 11323 29151 11326
rect 29453 11323 29519 11326
rect 30281 11386 30347 11389
rect 31017 11386 31083 11389
rect 30281 11384 31083 11386
rect 30281 11328 30286 11384
rect 30342 11328 31022 11384
rect 31078 11328 31083 11384
rect 30281 11326 31083 11328
rect 30281 11323 30347 11326
rect 31017 11323 31083 11326
rect 32029 11250 32095 11253
rect 36445 11250 36511 11253
rect 32029 11248 36511 11250
rect 32029 11192 32034 11248
rect 32090 11192 36450 11248
rect 36506 11192 36511 11248
rect 32029 11190 36511 11192
rect 32029 11187 32095 11190
rect 36445 11187 36511 11190
rect 54201 11250 54267 11253
rect 55200 11250 56000 11280
rect 54201 11248 56000 11250
rect 54201 11192 54206 11248
rect 54262 11192 56000 11248
rect 54201 11190 56000 11192
rect 54201 11187 54267 11190
rect 55200 11160 56000 11190
rect 32581 11114 32647 11117
rect 36077 11114 36143 11117
rect 32581 11112 36143 11114
rect 32581 11056 32586 11112
rect 32642 11056 36082 11112
rect 36138 11056 36143 11112
rect 32581 11054 36143 11056
rect 32581 11051 32647 11054
rect 36077 11051 36143 11054
rect 54201 10978 54267 10981
rect 55200 10978 56000 11008
rect 54201 10976 56000 10978
rect 54201 10920 54206 10976
rect 54262 10920 56000 10976
rect 54201 10918 56000 10920
rect 54201 10915 54267 10918
rect 19570 10912 19886 10913
rect 0 10842 800 10872
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 55200 10888 56000 10918
rect 50290 10847 50606 10848
rect 1669 10842 1735 10845
rect 0 10840 1735 10842
rect 0 10784 1674 10840
rect 1730 10784 1735 10840
rect 0 10782 1735 10784
rect 0 10752 800 10782
rect 1669 10779 1735 10782
rect 29913 10842 29979 10845
rect 30046 10842 30052 10844
rect 29913 10840 30052 10842
rect 29913 10784 29918 10840
rect 29974 10784 30052 10840
rect 29913 10782 30052 10784
rect 29913 10779 29979 10782
rect 30046 10780 30052 10782
rect 30116 10780 30122 10844
rect 31385 10842 31451 10845
rect 38561 10842 38627 10845
rect 31385 10840 38627 10842
rect 31385 10784 31390 10840
rect 31446 10784 38566 10840
rect 38622 10784 38627 10840
rect 31385 10782 38627 10784
rect 31385 10779 31451 10782
rect 38561 10779 38627 10782
rect 30741 10706 30807 10709
rect 31845 10706 31911 10709
rect 30741 10704 31911 10706
rect 30741 10648 30746 10704
rect 30802 10648 31850 10704
rect 31906 10648 31911 10704
rect 30741 10646 31911 10648
rect 30741 10643 30807 10646
rect 31845 10643 31911 10646
rect 32765 10706 32831 10709
rect 37181 10706 37247 10709
rect 32765 10704 37247 10706
rect 32765 10648 32770 10704
rect 32826 10648 37186 10704
rect 37242 10648 37247 10704
rect 32765 10646 37247 10648
rect 32765 10643 32831 10646
rect 37181 10643 37247 10646
rect 55200 10616 56000 10736
rect 54201 10434 54267 10437
rect 55200 10434 56000 10464
rect 54201 10432 56000 10434
rect 54201 10376 54206 10432
rect 54262 10376 56000 10432
rect 54201 10374 56000 10376
rect 54201 10371 54267 10374
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 55200 10344 56000 10374
rect 34930 10303 35246 10304
rect 1669 10298 1735 10301
rect 0 10296 1735 10298
rect 0 10240 1674 10296
rect 1730 10240 1735 10296
rect 0 10238 1735 10240
rect 0 10208 800 10238
rect 1669 10235 1735 10238
rect 53465 10162 53531 10165
rect 55200 10162 56000 10192
rect 53465 10160 56000 10162
rect 53465 10104 53470 10160
rect 53526 10104 56000 10160
rect 53465 10102 56000 10104
rect 53465 10099 53531 10102
rect 55200 10072 56000 10102
rect 33041 10026 33107 10029
rect 34973 10026 35039 10029
rect 36813 10026 36879 10029
rect 33041 10024 36879 10026
rect 33041 9968 33046 10024
rect 33102 9968 34978 10024
rect 35034 9968 36818 10024
rect 36874 9968 36879 10024
rect 33041 9966 36879 9968
rect 33041 9963 33107 9966
rect 34973 9963 35039 9966
rect 36813 9963 36879 9966
rect 30373 9892 30439 9893
rect 30373 9890 30420 9892
rect 30328 9888 30420 9890
rect 30328 9832 30378 9888
rect 30328 9830 30420 9832
rect 30373 9828 30420 9830
rect 30484 9828 30490 9892
rect 30373 9827 30439 9828
rect 19570 9824 19886 9825
rect 0 9754 800 9784
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 55200 9800 56000 9920
rect 50290 9759 50606 9760
rect 1669 9754 1735 9757
rect 0 9752 1735 9754
rect 0 9696 1674 9752
rect 1730 9696 1735 9752
rect 0 9694 1735 9696
rect 0 9664 800 9694
rect 1669 9691 1735 9694
rect 29494 9692 29500 9756
rect 29564 9754 29570 9756
rect 29913 9754 29979 9757
rect 29564 9752 29979 9754
rect 29564 9696 29918 9752
rect 29974 9696 29979 9752
rect 29564 9694 29979 9696
rect 29564 9692 29570 9694
rect 29913 9691 29979 9694
rect 16205 9618 16271 9621
rect 18597 9618 18663 9621
rect 16205 9616 18663 9618
rect 16205 9560 16210 9616
rect 16266 9560 18602 9616
rect 18658 9560 18663 9616
rect 16205 9558 18663 9560
rect 16205 9555 16271 9558
rect 18597 9555 18663 9558
rect 25313 9618 25379 9621
rect 28441 9618 28507 9621
rect 25313 9616 28507 9618
rect 25313 9560 25318 9616
rect 25374 9560 28446 9616
rect 28502 9560 28507 9616
rect 25313 9558 28507 9560
rect 25313 9555 25379 9558
rect 28441 9555 28507 9558
rect 54201 9618 54267 9621
rect 55200 9618 56000 9648
rect 54201 9616 56000 9618
rect 54201 9560 54206 9616
rect 54262 9560 56000 9616
rect 54201 9558 56000 9560
rect 54201 9555 54267 9558
rect 55200 9528 56000 9558
rect 23565 9482 23631 9485
rect 25221 9482 25287 9485
rect 23565 9480 25287 9482
rect 23565 9424 23570 9480
rect 23626 9424 25226 9480
rect 25282 9424 25287 9480
rect 23565 9422 25287 9424
rect 23565 9419 23631 9422
rect 25221 9419 25287 9422
rect 27429 9482 27495 9485
rect 29729 9482 29795 9485
rect 27429 9480 29795 9482
rect 27429 9424 27434 9480
rect 27490 9424 29734 9480
rect 29790 9424 29795 9480
rect 27429 9422 29795 9424
rect 27429 9419 27495 9422
rect 29729 9419 29795 9422
rect 26141 9346 26207 9349
rect 28901 9346 28967 9349
rect 26141 9344 28967 9346
rect 26141 9288 26146 9344
rect 26202 9288 28906 9344
rect 28962 9288 28967 9344
rect 26141 9286 28967 9288
rect 26141 9283 26207 9286
rect 28901 9283 28967 9286
rect 53557 9346 53623 9349
rect 55200 9346 56000 9376
rect 53557 9344 56000 9346
rect 53557 9288 53562 9344
rect 53618 9288 56000 9344
rect 53557 9286 56000 9288
rect 53557 9283 53623 9286
rect 4210 9280 4526 9281
rect 0 9210 800 9240
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 55200 9256 56000 9286
rect 34930 9215 35246 9216
rect 1669 9210 1735 9213
rect 0 9208 1735 9210
rect 0 9152 1674 9208
rect 1730 9152 1735 9208
rect 0 9150 1735 9152
rect 0 9120 800 9150
rect 1669 9147 1735 9150
rect 15745 9210 15811 9213
rect 18413 9210 18479 9213
rect 15745 9208 18479 9210
rect 15745 9152 15750 9208
rect 15806 9152 18418 9208
rect 18474 9152 18479 9208
rect 15745 9150 18479 9152
rect 15745 9147 15811 9150
rect 18413 9147 18479 9150
rect 26417 9074 26483 9077
rect 31845 9074 31911 9077
rect 32305 9074 32371 9077
rect 33593 9074 33659 9077
rect 26417 9072 32138 9074
rect 26417 9016 26422 9072
rect 26478 9016 31850 9072
rect 31906 9016 32138 9072
rect 26417 9014 32138 9016
rect 26417 9011 26483 9014
rect 31845 9011 31911 9014
rect 17309 8938 17375 8941
rect 17769 8938 17835 8941
rect 17309 8936 17835 8938
rect 17309 8880 17314 8936
rect 17370 8880 17774 8936
rect 17830 8880 17835 8936
rect 17309 8878 17835 8880
rect 32078 8938 32138 9014
rect 32305 9072 33659 9074
rect 32305 9016 32310 9072
rect 32366 9016 33598 9072
rect 33654 9016 33659 9072
rect 32305 9014 33659 9016
rect 32305 9011 32371 9014
rect 33593 9011 33659 9014
rect 55200 8984 56000 9104
rect 36721 8938 36787 8941
rect 32078 8936 36787 8938
rect 32078 8880 36726 8936
rect 36782 8880 36787 8936
rect 32078 8878 36787 8880
rect 17309 8875 17375 8878
rect 17769 8875 17835 8878
rect 36721 8875 36787 8878
rect 28625 8802 28691 8805
rect 33869 8802 33935 8805
rect 28625 8800 33935 8802
rect 28625 8744 28630 8800
rect 28686 8744 33874 8800
rect 33930 8744 33935 8800
rect 28625 8742 33935 8744
rect 28625 8739 28691 8742
rect 33869 8739 33935 8742
rect 54201 8802 54267 8805
rect 55200 8802 56000 8832
rect 54201 8800 56000 8802
rect 54201 8744 54206 8800
rect 54262 8744 56000 8800
rect 54201 8742 56000 8744
rect 54201 8739 54267 8742
rect 19570 8736 19886 8737
rect 0 8666 800 8696
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 55200 8712 56000 8742
rect 50290 8671 50606 8672
rect 1669 8666 1735 8669
rect 0 8664 1735 8666
rect 0 8608 1674 8664
rect 1730 8608 1735 8664
rect 0 8606 1735 8608
rect 0 8576 800 8606
rect 1669 8603 1735 8606
rect 31845 8666 31911 8669
rect 35893 8666 35959 8669
rect 31845 8664 35959 8666
rect 31845 8608 31850 8664
rect 31906 8608 35898 8664
rect 35954 8608 35959 8664
rect 31845 8606 35959 8608
rect 31845 8603 31911 8606
rect 35893 8603 35959 8606
rect 53465 8530 53531 8533
rect 55200 8530 56000 8560
rect 53465 8528 56000 8530
rect 53465 8472 53470 8528
rect 53526 8472 56000 8528
rect 53465 8470 56000 8472
rect 53465 8467 53531 8470
rect 55200 8440 56000 8470
rect 14641 8394 14707 8397
rect 29361 8394 29427 8397
rect 14641 8392 29427 8394
rect 14641 8336 14646 8392
rect 14702 8336 29366 8392
rect 29422 8336 29427 8392
rect 14641 8334 29427 8336
rect 14641 8331 14707 8334
rect 29361 8331 29427 8334
rect 4210 8192 4526 8193
rect 0 8122 800 8152
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 55200 8168 56000 8288
rect 34930 8127 35246 8128
rect 1669 8122 1735 8125
rect 0 8120 1735 8122
rect 0 8064 1674 8120
rect 1730 8064 1735 8120
rect 0 8062 1735 8064
rect 0 8032 800 8062
rect 1669 8059 1735 8062
rect 52177 7986 52243 7989
rect 55200 7986 56000 8016
rect 52177 7984 56000 7986
rect 52177 7928 52182 7984
rect 52238 7928 56000 7984
rect 52177 7926 56000 7928
rect 52177 7923 52243 7926
rect 55200 7896 56000 7926
rect 53373 7714 53439 7717
rect 55200 7714 56000 7744
rect 53373 7712 56000 7714
rect 53373 7656 53378 7712
rect 53434 7656 56000 7712
rect 53373 7654 56000 7656
rect 53373 7651 53439 7654
rect 19570 7648 19886 7649
rect 0 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 55200 7624 56000 7654
rect 50290 7583 50606 7584
rect 1669 7578 1735 7581
rect 0 7576 1735 7578
rect 0 7520 1674 7576
rect 1730 7520 1735 7576
rect 0 7518 1735 7520
rect 0 7488 800 7518
rect 1669 7515 1735 7518
rect 23749 7442 23815 7445
rect 30414 7442 30420 7444
rect 23749 7440 30420 7442
rect 23749 7384 23754 7440
rect 23810 7384 30420 7440
rect 23749 7382 30420 7384
rect 23749 7379 23815 7382
rect 30414 7380 30420 7382
rect 30484 7442 30490 7444
rect 30741 7442 30807 7445
rect 30484 7440 30807 7442
rect 30484 7384 30746 7440
rect 30802 7384 30807 7440
rect 30484 7382 30807 7384
rect 30484 7380 30490 7382
rect 30741 7379 30807 7382
rect 52269 7442 52335 7445
rect 55200 7442 56000 7472
rect 52269 7440 56000 7442
rect 52269 7384 52274 7440
rect 52330 7384 56000 7440
rect 52269 7382 56000 7384
rect 52269 7379 52335 7382
rect 55200 7352 56000 7382
rect 54109 7170 54175 7173
rect 55200 7170 56000 7200
rect 54109 7168 56000 7170
rect 54109 7112 54114 7168
rect 54170 7112 56000 7168
rect 54109 7110 56000 7112
rect 54109 7107 54175 7110
rect 4210 7104 4526 7105
rect 0 7034 800 7064
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 55200 7080 56000 7110
rect 34930 7039 35246 7040
rect 1669 7034 1735 7037
rect 0 7032 1735 7034
rect 0 6976 1674 7032
rect 1730 6976 1735 7032
rect 0 6974 1735 6976
rect 0 6944 800 6974
rect 1669 6971 1735 6974
rect 29637 7034 29703 7037
rect 30966 7034 30972 7036
rect 29637 7032 30972 7034
rect 29637 6976 29642 7032
rect 29698 6976 30972 7032
rect 29637 6974 30972 6976
rect 29637 6971 29703 6974
rect 30966 6972 30972 6974
rect 31036 6972 31042 7036
rect 54385 6898 54451 6901
rect 55200 6898 56000 6928
rect 54385 6896 56000 6898
rect 54385 6840 54390 6896
rect 54446 6840 56000 6896
rect 54385 6838 56000 6840
rect 54385 6835 54451 6838
rect 55200 6808 56000 6838
rect 51257 6626 51323 6629
rect 55200 6626 56000 6656
rect 51257 6624 56000 6626
rect 51257 6568 51262 6624
rect 51318 6568 56000 6624
rect 51257 6566 56000 6568
rect 51257 6563 51323 6566
rect 19570 6560 19886 6561
rect 0 6490 800 6520
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 55200 6536 56000 6566
rect 50290 6495 50606 6496
rect 1669 6490 1735 6493
rect 0 6488 1735 6490
rect 0 6432 1674 6488
rect 1730 6432 1735 6488
rect 0 6430 1735 6432
rect 0 6400 800 6430
rect 1669 6427 1735 6430
rect 4210 6016 4526 6017
rect 0 5946 800 5976
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 1669 5946 1735 5949
rect 0 5944 1735 5946
rect 0 5888 1674 5944
rect 1730 5888 1735 5944
rect 0 5886 1735 5888
rect 0 5856 800 5886
rect 1669 5883 1735 5886
rect 19570 5472 19886 5473
rect 0 5402 800 5432
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 1669 5402 1735 5405
rect 0 5400 1735 5402
rect 0 5344 1674 5400
rect 1730 5344 1735 5400
rect 0 5342 1735 5344
rect 0 5312 800 5342
rect 1669 5339 1735 5342
rect 12433 5130 12499 5133
rect 13813 5130 13879 5133
rect 12433 5128 13879 5130
rect 12433 5072 12438 5128
rect 12494 5072 13818 5128
rect 13874 5072 13879 5128
rect 12433 5070 13879 5072
rect 12433 5067 12499 5070
rect 13813 5067 13879 5070
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1669 4858 1735 4861
rect 0 4856 1735 4858
rect 0 4800 1674 4856
rect 1730 4800 1735 4856
rect 0 4798 1735 4800
rect 0 4768 800 4798
rect 1669 4795 1735 4798
rect 19570 4384 19886 4385
rect 0 4314 800 4344
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 1669 4314 1735 4317
rect 0 4312 1735 4314
rect 0 4256 1674 4312
rect 1730 4256 1735 4312
rect 0 4254 1735 4256
rect 0 4224 800 4254
rect 1669 4251 1735 4254
rect 34094 3980 34100 4044
rect 34164 4042 34170 4044
rect 34513 4042 34579 4045
rect 34164 4040 34579 4042
rect 34164 3984 34518 4040
rect 34574 3984 34579 4040
rect 34164 3982 34579 3984
rect 34164 3980 34170 3982
rect 34513 3979 34579 3982
rect 10041 3906 10107 3909
rect 10685 3906 10751 3909
rect 18597 3906 18663 3909
rect 10041 3904 18663 3906
rect 10041 3848 10046 3904
rect 10102 3848 10690 3904
rect 10746 3848 18602 3904
rect 18658 3848 18663 3904
rect 10041 3846 18663 3848
rect 10041 3843 10107 3846
rect 10685 3843 10751 3846
rect 18597 3843 18663 3846
rect 4210 3840 4526 3841
rect 0 3770 800 3800
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 1669 3770 1735 3773
rect 0 3768 1735 3770
rect 0 3712 1674 3768
rect 1730 3712 1735 3768
rect 0 3710 1735 3712
rect 0 3680 800 3710
rect 1669 3707 1735 3710
rect 26785 3770 26851 3773
rect 27838 3770 27844 3772
rect 26785 3768 27844 3770
rect 26785 3712 26790 3768
rect 26846 3712 27844 3768
rect 26785 3710 27844 3712
rect 26785 3707 26851 3710
rect 27838 3708 27844 3710
rect 27908 3708 27914 3772
rect 28625 3770 28691 3773
rect 33317 3772 33383 3773
rect 28758 3770 28764 3772
rect 28625 3768 28764 3770
rect 28625 3712 28630 3768
rect 28686 3712 28764 3768
rect 28625 3710 28764 3712
rect 28625 3707 28691 3710
rect 28758 3708 28764 3710
rect 28828 3708 28834 3772
rect 33317 3770 33364 3772
rect 33272 3768 33364 3770
rect 33272 3712 33322 3768
rect 33272 3710 33364 3712
rect 33317 3708 33364 3710
rect 33428 3708 33434 3772
rect 33317 3707 33383 3708
rect 10133 3634 10199 3637
rect 14457 3634 14523 3637
rect 10133 3632 14523 3634
rect 10133 3576 10138 3632
rect 10194 3576 14462 3632
rect 14518 3576 14523 3632
rect 10133 3574 14523 3576
rect 10133 3571 10199 3574
rect 14457 3571 14523 3574
rect 9949 3362 10015 3365
rect 10869 3362 10935 3365
rect 9949 3360 10935 3362
rect 9949 3304 9954 3360
rect 10010 3304 10874 3360
rect 10930 3304 10935 3360
rect 9949 3302 10935 3304
rect 9949 3299 10015 3302
rect 10869 3299 10935 3302
rect 19570 3296 19886 3297
rect 0 3226 800 3256
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 1669 3226 1735 3229
rect 0 3224 1735 3226
rect 0 3168 1674 3224
rect 1730 3168 1735 3224
rect 0 3166 1735 3168
rect 0 3136 800 3166
rect 1669 3163 1735 3166
rect 12525 2818 12591 2821
rect 12893 2818 12959 2821
rect 12525 2816 12959 2818
rect 12525 2760 12530 2816
rect 12586 2760 12898 2816
rect 12954 2760 12959 2816
rect 12525 2758 12959 2760
rect 12525 2755 12591 2758
rect 12893 2755 12959 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 27470 2348 27476 2412
rect 27540 2410 27546 2412
rect 51809 2410 51875 2413
rect 27540 2408 51875 2410
rect 27540 2352 51814 2408
rect 51870 2352 51875 2408
rect 27540 2350 51875 2352
rect 27540 2348 27546 2350
rect 51809 2347 51875 2350
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
<< via3 >>
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 27844 52532 27908 52596
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 27108 45460 27172 45524
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 31340 44916 31404 44980
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 28764 41652 28828 41716
rect 25820 41516 25884 41580
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 27844 41244 27908 41308
rect 29316 40836 29380 40900
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 26556 40020 26620 40084
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 29316 38932 29380 38996
rect 26924 38660 26988 38724
rect 29684 38660 29748 38724
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 28948 38584 29012 38588
rect 28948 38528 28998 38584
rect 28998 38528 29012 38584
rect 28948 38524 29012 38528
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 31340 37980 31404 38044
rect 26372 37844 26436 37908
rect 28212 37708 28276 37772
rect 27660 37572 27724 37636
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 27108 37436 27172 37500
rect 28948 37436 29012 37500
rect 26004 37360 26068 37364
rect 26004 37304 26054 37360
rect 26054 37304 26068 37360
rect 26004 37300 26068 37304
rect 27108 37224 27172 37228
rect 27108 37168 27122 37224
rect 27122 37168 27172 37224
rect 27108 37164 27172 37168
rect 29684 37164 29748 37228
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 29316 36000 29380 36004
rect 29316 35944 29330 36000
rect 29330 35944 29380 36000
rect 29316 35940 29380 35944
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 27476 35592 27540 35596
rect 27476 35536 27490 35592
rect 27490 35536 27540 35592
rect 27476 35532 27540 35536
rect 26372 35396 26436 35460
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 26372 34852 26436 34916
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 29132 33416 29196 33420
rect 29132 33360 29146 33416
rect 29146 33360 29196 33416
rect 29132 33356 29196 33360
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 28212 33144 28276 33148
rect 28212 33088 28262 33144
rect 28262 33088 28276 33144
rect 28212 33084 28276 33088
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 28948 32404 29012 32468
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 26372 31724 26436 31788
rect 32628 31724 32692 31788
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 30052 27644 30116 27708
rect 26556 27508 26620 27572
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 33364 25196 33428 25260
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 34100 23428 34164 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 28764 21388 28828 21452
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 29500 20572 29564 20636
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 38332 19272 38396 19276
rect 38332 19216 38346 19272
rect 38346 19216 38396 19272
rect 38332 19212 38396 19216
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 30972 18532 31036 18596
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 27844 17716 27908 17780
rect 29316 17716 29380 17780
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 26924 15540 26988 15604
rect 26004 15268 26068 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 25820 15132 25884 15196
rect 30604 15192 30668 15196
rect 30604 15136 30618 15192
rect 30618 15136 30668 15192
rect 30604 15132 30668 15136
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 38332 13908 38396 13972
rect 32628 13636 32692 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 30052 10780 30116 10844
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 30420 9888 30484 9892
rect 30420 9832 30434 9888
rect 30434 9832 30484 9888
rect 30420 9828 30484 9832
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 29500 9692 29564 9756
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 30420 7380 30484 7444
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 30972 6972 31036 7036
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 34100 3980 34164 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 27844 3708 27908 3772
rect 28764 3708 28828 3772
rect 33364 3768 33428 3772
rect 33364 3712 33378 3768
rect 33378 3712 33428 3768
rect 33364 3708 33428 3712
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 27476 2348 27540 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 52800 4528 53360
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 53344 19888 53360
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 34928 52800 35248 53360
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 27843 52596 27909 52597
rect 27843 52532 27844 52596
rect 27908 52532 27909 52596
rect 27843 52531 27909 52532
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 27107 45524 27173 45525
rect 27107 45460 27108 45524
rect 27172 45460 27173 45524
rect 27107 45459 27173 45460
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 25819 41580 25885 41581
rect 25819 41516 25820 41580
rect 25884 41516 25885 41580
rect 25819 41515 25885 41516
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 25822 15197 25882 41515
rect 26555 40084 26621 40085
rect 26555 40020 26556 40084
rect 26620 40020 26621 40084
rect 26555 40019 26621 40020
rect 26371 37908 26437 37909
rect 26371 37844 26372 37908
rect 26436 37844 26437 37908
rect 26371 37843 26437 37844
rect 26003 37364 26069 37365
rect 26003 37300 26004 37364
rect 26068 37300 26069 37364
rect 26003 37299 26069 37300
rect 26006 15333 26066 37299
rect 26374 35461 26434 37843
rect 26371 35460 26437 35461
rect 26371 35396 26372 35460
rect 26436 35396 26437 35460
rect 26371 35395 26437 35396
rect 26374 34917 26434 35395
rect 26371 34916 26437 34917
rect 26371 34852 26372 34916
rect 26436 34852 26437 34916
rect 26371 34851 26437 34852
rect 26374 31789 26434 34851
rect 26371 31788 26437 31789
rect 26371 31724 26372 31788
rect 26436 31724 26437 31788
rect 26371 31723 26437 31724
rect 26558 27573 26618 40019
rect 26923 38724 26989 38725
rect 26923 38660 26924 38724
rect 26988 38660 26989 38724
rect 26923 38659 26989 38660
rect 26555 27572 26621 27573
rect 26555 27508 26556 27572
rect 26620 27508 26621 27572
rect 26555 27507 26621 27508
rect 26926 15605 26986 38659
rect 27110 37501 27170 45459
rect 27846 41309 27906 52531
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 31339 44980 31405 44981
rect 31339 44916 31340 44980
rect 31404 44916 31405 44980
rect 31339 44915 31405 44916
rect 28763 41716 28829 41717
rect 28763 41652 28764 41716
rect 28828 41652 28829 41716
rect 28763 41651 28829 41652
rect 27843 41308 27909 41309
rect 27843 41244 27844 41308
rect 27908 41244 27909 41308
rect 27843 41243 27909 41244
rect 28211 37772 28277 37773
rect 28211 37708 28212 37772
rect 28276 37708 28277 37772
rect 28211 37707 28277 37708
rect 27659 37636 27725 37637
rect 27659 37572 27660 37636
rect 27724 37572 27725 37636
rect 27659 37571 27725 37572
rect 27107 37500 27173 37501
rect 27107 37436 27108 37500
rect 27172 37436 27173 37500
rect 27107 37435 27173 37436
rect 27110 37229 27170 37435
rect 27107 37228 27173 37229
rect 27107 37164 27108 37228
rect 27172 37164 27173 37228
rect 27107 37163 27173 37164
rect 27662 35730 27722 37571
rect 27478 35670 27722 35730
rect 27478 35597 27538 35670
rect 27475 35596 27541 35597
rect 27475 35532 27476 35596
rect 27540 35532 27541 35596
rect 27475 35531 27541 35532
rect 26923 15604 26989 15605
rect 26923 15540 26924 15604
rect 26988 15540 26989 15604
rect 26923 15539 26989 15540
rect 26003 15332 26069 15333
rect 26003 15268 26004 15332
rect 26068 15268 26069 15332
rect 26003 15267 26069 15268
rect 25819 15196 25885 15197
rect 25819 15132 25820 15196
rect 25884 15132 25885 15196
rect 25819 15131 25885 15132
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 27478 2413 27538 35531
rect 28214 33149 28274 37707
rect 28211 33148 28277 33149
rect 28211 33084 28212 33148
rect 28276 33084 28277 33148
rect 28211 33083 28277 33084
rect 28766 21453 28826 41651
rect 29315 40900 29381 40901
rect 29315 40836 29316 40900
rect 29380 40836 29381 40900
rect 29315 40835 29381 40836
rect 29318 38997 29378 40835
rect 29315 38996 29381 38997
rect 29315 38932 29316 38996
rect 29380 38932 29381 38996
rect 29315 38931 29381 38932
rect 29683 38724 29749 38725
rect 29683 38660 29684 38724
rect 29748 38660 29749 38724
rect 29683 38659 29749 38660
rect 28947 38588 29013 38589
rect 28947 38524 28948 38588
rect 29012 38524 29013 38588
rect 28947 38523 29013 38524
rect 28950 38450 29010 38523
rect 28950 38390 29194 38450
rect 28947 37500 29013 37501
rect 28947 37436 28948 37500
rect 29012 37436 29013 37500
rect 28947 37435 29013 37436
rect 28950 32469 29010 37435
rect 29134 33421 29194 38390
rect 29686 37229 29746 38659
rect 31342 38045 31402 44915
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 31339 38044 31405 38045
rect 31339 37980 31340 38044
rect 31404 37980 31405 38044
rect 31339 37979 31405 37980
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 29683 37228 29749 37229
rect 29683 37164 29684 37228
rect 29748 37164 29749 37228
rect 29683 37163 29749 37164
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 29315 36004 29381 36005
rect 29315 35940 29316 36004
rect 29380 35940 29381 36004
rect 29315 35939 29381 35940
rect 29131 33420 29197 33421
rect 29131 33356 29132 33420
rect 29196 33356 29197 33420
rect 29131 33355 29197 33356
rect 28947 32468 29013 32469
rect 28947 32404 28948 32468
rect 29012 32404 29013 32468
rect 28947 32403 29013 32404
rect 28763 21452 28829 21453
rect 28763 21388 28764 21452
rect 28828 21388 28829 21452
rect 28763 21387 28829 21388
rect 27843 17780 27909 17781
rect 27843 17716 27844 17780
rect 27908 17716 27909 17780
rect 27843 17715 27909 17716
rect 27846 3773 27906 17715
rect 28766 3773 28826 21387
rect 29318 17781 29378 35939
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 32627 31788 32693 31789
rect 32627 31724 32628 31788
rect 32692 31724 32693 31788
rect 32627 31723 32693 31724
rect 30051 27708 30117 27709
rect 30051 27644 30052 27708
rect 30116 27644 30117 27708
rect 30051 27643 30117 27644
rect 29499 20636 29565 20637
rect 29499 20572 29500 20636
rect 29564 20572 29565 20636
rect 29499 20571 29565 20572
rect 29315 17780 29381 17781
rect 29315 17716 29316 17780
rect 29380 17716 29381 17780
rect 29315 17715 29381 17716
rect 29502 9757 29562 20571
rect 30054 10845 30114 27643
rect 30971 18596 31037 18597
rect 30971 18532 30972 18596
rect 31036 18532 31037 18596
rect 30971 18531 31037 18532
rect 30603 15196 30669 15197
rect 30603 15132 30604 15196
rect 30668 15132 30669 15196
rect 30603 15131 30669 15132
rect 30606 12450 30666 15131
rect 30422 12390 30666 12450
rect 30051 10844 30117 10845
rect 30051 10780 30052 10844
rect 30116 10780 30117 10844
rect 30051 10779 30117 10780
rect 30422 9893 30482 12390
rect 30419 9892 30485 9893
rect 30419 9828 30420 9892
rect 30484 9828 30485 9892
rect 30419 9827 30485 9828
rect 29499 9756 29565 9757
rect 29499 9692 29500 9756
rect 29564 9692 29565 9756
rect 29499 9691 29565 9692
rect 30422 7445 30482 9827
rect 30419 7444 30485 7445
rect 30419 7380 30420 7444
rect 30484 7380 30485 7444
rect 30419 7379 30485 7380
rect 30974 7037 31034 18531
rect 32630 13701 32690 31723
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 33363 25260 33429 25261
rect 33363 25196 33364 25260
rect 33428 25196 33429 25260
rect 33363 25195 33429 25196
rect 32627 13700 32693 13701
rect 32627 13636 32628 13700
rect 32692 13636 32693 13700
rect 32627 13635 32693 13636
rect 30971 7036 31037 7037
rect 30971 6972 30972 7036
rect 31036 6972 31037 7036
rect 30971 6971 31037 6972
rect 33366 3773 33426 25195
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34099 23492 34165 23493
rect 34099 23428 34100 23492
rect 34164 23428 34165 23492
rect 34099 23427 34165 23428
rect 34102 4045 34162 23427
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 50288 53344 50608 53360
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 38331 19276 38397 19277
rect 38331 19212 38332 19276
rect 38396 19212 38397 19276
rect 38331 19211 38397 19212
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 38334 13973 38394 19211
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 38331 13972 38397 13973
rect 38331 13908 38332 13972
rect 38396 13908 38397 13972
rect 38331 13907 38397 13908
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34099 4044 34165 4045
rect 34099 3980 34100 4044
rect 34164 3980 34165 4044
rect 34099 3979 34165 3980
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 27843 3772 27909 3773
rect 27843 3708 27844 3772
rect 27908 3708 27909 3772
rect 27843 3707 27909 3708
rect 28763 3772 28829 3773
rect 28763 3708 28764 3772
rect 28828 3708 28829 3772
rect 28763 3707 28829 3708
rect 33363 3772 33429 3773
rect 33363 3708 33364 3772
rect 33428 3708 33429 3772
rect 33363 3707 33429 3708
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 27475 2412 27541 2413
rect 27475 2348 27476 2412
rect 27540 2348 27541 2412
rect 27475 2347 27541 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__A0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23920 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__A
timestamp 1666464484
transform 1 0 33396 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__A
timestamp 1666464484
transform 1 0 34868 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__A
timestamp 1666464484
transform 1 0 14536 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__B_N
timestamp 1666464484
transform -1 0 14904 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__A
timestamp 1666464484
transform 1 0 20700 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__B_N
timestamp 1666464484
transform -1 0 20884 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__A
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__B_N
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__C
timestamp 1666464484
transform 1 0 23000 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__A
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__B_N
timestamp 1666464484
transform -1 0 21068 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__A
timestamp 1666464484
transform 1 0 15456 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__B_N
timestamp 1666464484
transform 1 0 15824 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__A
timestamp 1666464484
transform 1 0 31648 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__A
timestamp 1666464484
transform 1 0 23368 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A
timestamp 1666464484
transform 1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__B_N
timestamp 1666464484
transform -1 0 21988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__B
timestamp 1666464484
transform 1 0 22908 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__B
timestamp 1666464484
transform 1 0 22448 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A
timestamp 1666464484
transform 1 0 21988 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__A2
timestamp 1666464484
transform 1 0 53084 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__B1
timestamp 1666464484
transform 1 0 52716 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__A1
timestamp 1666464484
transform -1 0 28520 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__A2
timestamp 1666464484
transform 1 0 29716 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__B1
timestamp 1666464484
transform -1 0 31648 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A1
timestamp 1666464484
transform 1 0 27324 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__B1
timestamp 1666464484
transform 1 0 28888 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__A1
timestamp 1666464484
transform 1 0 30544 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__B1
timestamp 1666464484
transform -1 0 29072 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__A
timestamp 1666464484
transform -1 0 30728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__A
timestamp 1666464484
transform 1 0 21528 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__B
timestamp 1666464484
transform 1 0 22540 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__A
timestamp 1666464484
transform -1 0 11960 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__B
timestamp 1666464484
transform -1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A1
timestamp 1666464484
transform -1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A2
timestamp 1666464484
transform -1 0 12696 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__B1
timestamp 1666464484
transform -1 0 12696 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A
timestamp 1666464484
transform -1 0 31004 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__A
timestamp 1666464484
transform 1 0 34040 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__A
timestamp 1666464484
transform -1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__A
timestamp 1666464484
transform 1 0 28796 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__B
timestamp 1666464484
transform 1 0 27784 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__A
timestamp 1666464484
transform -1 0 42688 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__B
timestamp 1666464484
transform -1 0 42780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__A
timestamp 1666464484
transform 1 0 25024 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 1666464484
transform 1 0 24380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A
timestamp 1666464484
transform 1 0 14444 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__B
timestamp 1666464484
transform -1 0 12328 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A
timestamp 1666464484
transform -1 0 15180 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__B
timestamp 1666464484
transform -1 0 15732 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A
timestamp 1666464484
transform -1 0 23828 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__A1
timestamp 1666464484
transform 1 0 32476 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__A2
timestamp 1666464484
transform -1 0 32476 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__B1
timestamp 1666464484
transform 1 0 33212 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__B2
timestamp 1666464484
transform -1 0 29900 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__A
timestamp 1666464484
transform 1 0 26496 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A1
timestamp 1666464484
transform -1 0 31740 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A2
timestamp 1666464484
transform -1 0 30452 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__B2
timestamp 1666464484
transform -1 0 31188 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A1
timestamp 1666464484
transform -1 0 29808 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A2
timestamp 1666464484
transform 1 0 30728 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B1
timestamp 1666464484
transform 1 0 29072 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B2
timestamp 1666464484
transform -1 0 30912 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__A1
timestamp 1666464484
transform 1 0 29716 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__A2
timestamp 1666464484
transform -1 0 30544 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__B1
timestamp 1666464484
transform 1 0 31832 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__B2
timestamp 1666464484
transform -1 0 31096 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__A
timestamp 1666464484
transform 1 0 32844 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__A1
timestamp 1666464484
transform 1 0 29716 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__A2
timestamp 1666464484
transform 1 0 30268 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__B1
timestamp 1666464484
transform 1 0 25116 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__B2
timestamp 1666464484
transform -1 0 24748 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A1
timestamp 1666464484
transform -1 0 31556 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A2
timestamp 1666464484
transform 1 0 29716 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__B2
timestamp 1666464484
transform -1 0 32476 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A1
timestamp 1666464484
transform 1 0 31096 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A2
timestamp 1666464484
transform 1 0 30820 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A1
timestamp 1666464484
transform -1 0 24932 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A1
timestamp 1666464484
transform -1 0 34316 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A2
timestamp 1666464484
transform 1 0 30912 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__B1
timestamp 1666464484
transform 1 0 30360 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__B2
timestamp 1666464484
transform -1 0 31004 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A2
timestamp 1666464484
transform 1 0 14628 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__B1
timestamp 1666464484
transform 1 0 14996 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__B2
timestamp 1666464484
transform 1 0 13432 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A1
timestamp 1666464484
transform -1 0 33488 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A2
timestamp 1666464484
transform 1 0 31372 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__B1
timestamp 1666464484
transform -1 0 32384 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__B2
timestamp 1666464484
transform 1 0 32752 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A1
timestamp 1666464484
transform -1 0 32108 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A1
timestamp 1666464484
transform -1 0 34776 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A2
timestamp 1666464484
transform -1 0 30452 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__B1
timestamp 1666464484
transform 1 0 31280 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__B2
timestamp 1666464484
transform 1 0 32292 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A1
timestamp 1666464484
transform -1 0 22356 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A2
timestamp 1666464484
transform 1 0 21620 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__B1
timestamp 1666464484
transform -1 0 22540 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__B2
timestamp 1666464484
transform -1 0 22448 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A1
timestamp 1666464484
transform -1 0 16100 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A2
timestamp 1666464484
transform 1 0 15548 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B1
timestamp 1666464484
transform 1 0 16468 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B2
timestamp 1666464484
transform -1 0 14444 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A1
timestamp 1666464484
transform -1 0 33028 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A1
timestamp 1666464484
transform 1 0 25300 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A2
timestamp 1666464484
transform 1 0 31924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__B2
timestamp 1666464484
transform -1 0 31280 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A1
timestamp 1666464484
transform -1 0 25760 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A2
timestamp 1666464484
transform 1 0 25208 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__B1
timestamp 1666464484
transform -1 0 29256 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__B2
timestamp 1666464484
transform -1 0 24840 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A1
timestamp 1666464484
transform 1 0 31464 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A2
timestamp 1666464484
transform 1 0 27692 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__B1
timestamp 1666464484
transform 1 0 29256 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__B2
timestamp 1666464484
transform -1 0 27324 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A1
timestamp 1666464484
transform -1 0 33948 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A2
timestamp 1666464484
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__B1
timestamp 1666464484
transform 1 0 31556 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__B2
timestamp 1666464484
transform -1 0 33028 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A1
timestamp 1666464484
transform 1 0 22816 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A2
timestamp 1666464484
transform -1 0 23552 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__B2
timestamp 1666464484
transform -1 0 24840 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A1
timestamp 1666464484
transform -1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A2
timestamp 1666464484
transform 1 0 25484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__B1
timestamp 1666464484
transform 1 0 24932 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__B2
timestamp 1666464484
transform 1 0 28060 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A1
timestamp 1666464484
transform -1 0 26128 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A2
timestamp 1666464484
transform 1 0 26496 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B1
timestamp 1666464484
transform 1 0 26772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B2
timestamp 1666464484
transform -1 0 28336 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A1
timestamp 1666464484
transform -1 0 25024 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A2
timestamp 1666464484
transform 1 0 25852 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B1
timestamp 1666464484
transform 1 0 28152 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B2
timestamp 1666464484
transform 1 0 24472 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A2
timestamp 1666464484
transform 1 0 14444 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B1
timestamp 1666464484
transform 1 0 14812 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A1
timestamp 1666464484
transform -1 0 34500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A2
timestamp 1666464484
transform 1 0 30452 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__B1
timestamp 1666464484
transform -1 0 32476 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__B2
timestamp 1666464484
transform -1 0 33948 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__C1
timestamp 1666464484
transform -1 0 26036 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A1
timestamp 1666464484
transform 1 0 23920 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A2
timestamp 1666464484
transform 1 0 25668 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__B1
timestamp 1666464484
transform 1 0 24104 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__B2
timestamp 1666464484
transform -1 0 24840 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A1
timestamp 1666464484
transform 1 0 23092 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A2
timestamp 1666464484
transform 1 0 25300 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__B2
timestamp 1666464484
transform -1 0 24380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A1
timestamp 1666464484
transform 1 0 25208 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A2
timestamp 1666464484
transform 1 0 29072 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A1
timestamp 1666464484
transform 1 0 22448 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A2
timestamp 1666464484
transform 1 0 23000 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__B1
timestamp 1666464484
transform 1 0 23920 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__B2
timestamp 1666464484
transform -1 0 24932 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A1
timestamp 1666464484
transform -1 0 22448 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A2
timestamp 1666464484
transform -1 0 23000 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__B1
timestamp 1666464484
transform 1 0 24748 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__B2
timestamp 1666464484
transform -1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A1
timestamp 1666464484
transform -1 0 25668 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__B2
timestamp 1666464484
transform 1 0 28796 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A1
timestamp 1666464484
transform -1 0 24104 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A2
timestamp 1666464484
transform 1 0 26036 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__B2
timestamp 1666464484
transform -1 0 25208 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A1
timestamp 1666464484
transform 1 0 23368 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A2
timestamp 1666464484
transform 1 0 26588 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A1
timestamp 1666464484
transform -1 0 23644 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B1
timestamp 1666464484
transform 1 0 23920 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B2
timestamp 1666464484
transform -1 0 23552 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__A1
timestamp 1666464484
transform 1 0 21344 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__A2
timestamp 1666464484
transform 1 0 21344 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B1
timestamp 1666464484
transform -1 0 23000 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B2
timestamp 1666464484
transform -1 0 20424 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__A1
timestamp 1666464484
transform 1 0 32844 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__A2
timestamp 1666464484
transform -1 0 31004 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__B2
timestamp 1666464484
transform -1 0 32108 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A2
timestamp 1666464484
transform 1 0 23736 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A1
timestamp 1666464484
transform -1 0 24472 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A2
timestamp 1666464484
transform -1 0 25116 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B1
timestamp 1666464484
transform 1 0 25944 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B2
timestamp 1666464484
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A2
timestamp 1666464484
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B1
timestamp 1666464484
transform 1 0 27324 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B2
timestamp 1666464484
transform 1 0 26772 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A1
timestamp 1666464484
transform 1 0 20792 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A2
timestamp 1666464484
transform 1 0 22908 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B1
timestamp 1666464484
transform 1 0 22724 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B2
timestamp 1666464484
transform -1 0 21252 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A1
timestamp 1666464484
transform -1 0 21344 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A2
timestamp 1666464484
transform 1 0 22264 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__B1
timestamp 1666464484
transform 1 0 23368 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__B2
timestamp 1666464484
transform 1 0 21712 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A1
timestamp 1666464484
transform -1 0 28520 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__B2
timestamp 1666464484
transform -1 0 32476 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A1
timestamp 1666464484
transform -1 0 26496 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A2
timestamp 1666464484
transform 1 0 26128 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__B2
timestamp 1666464484
transform -1 0 27876 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A
timestamp 1666464484
transform 1 0 24932 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A2
timestamp 1666464484
transform -1 0 25944 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B1
timestamp 1666464484
transform 1 0 25944 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B2
timestamp 1666464484
transform -1 0 24748 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A1
timestamp 1666464484
transform 1 0 21988 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B2
timestamp 1666464484
transform -1 0 22724 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A1
timestamp 1666464484
transform 1 0 29900 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B1
timestamp 1666464484
transform -1 0 24840 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B2
timestamp 1666464484
transform 1 0 31188 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A1
timestamp 1666464484
transform -1 0 23736 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A2
timestamp 1666464484
transform -1 0 22632 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B1
timestamp 1666464484
transform 1 0 23000 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B2
timestamp 1666464484
transform 1 0 22816 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A1
timestamp 1666464484
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A2
timestamp 1666464484
transform 1 0 25484 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B1
timestamp 1666464484
transform 1 0 26036 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B2
timestamp 1666464484
transform -1 0 27968 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A1
timestamp 1666464484
transform -1 0 22908 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A2
timestamp 1666464484
transform -1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__B1
timestamp 1666464484
transform -1 0 23000 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__B2
timestamp 1666464484
transform -1 0 23092 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A2
timestamp 1666464484
transform -1 0 25760 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B1
timestamp 1666464484
transform 1 0 24380 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B2
timestamp 1666464484
transform 1 0 28244 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A1
timestamp 1666464484
transform 1 0 23092 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__B1
timestamp 1666464484
transform 1 0 24564 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__B2
timestamp 1666464484
transform -1 0 23460 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A1
timestamp 1666464484
transform -1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A2
timestamp 1666464484
transform 1 0 23460 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__B2
timestamp 1666464484
transform -1 0 23552 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A1
timestamp 1666464484
transform 1 0 28796 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A2
timestamp 1666464484
transform 1 0 24012 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A2
timestamp 1666464484
transform 1 0 23828 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__B1
timestamp 1666464484
transform 1 0 23276 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__B2
timestamp 1666464484
transform 1 0 22264 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A2
timestamp 1666464484
transform 1 0 17480 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__B1
timestamp 1666464484
transform 1 0 17848 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__B2
timestamp 1666464484
transform -1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A2
timestamp 1666464484
transform -1 0 23552 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__B2
timestamp 1666464484
transform -1 0 25576 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A1
timestamp 1666464484
transform 1 0 25944 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A2
timestamp 1666464484
transform 1 0 26496 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__B1
timestamp 1666464484
transform 1 0 27968 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__B2
timestamp 1666464484
transform 1 0 28520 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A2
timestamp 1666464484
transform 1 0 27324 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B1
timestamp 1666464484
transform -1 0 27324 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B2
timestamp 1666464484
transform -1 0 26680 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A1
timestamp 1666464484
transform -1 0 31464 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B1
timestamp 1666464484
transform -1 0 30360 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B2
timestamp 1666464484
transform 1 0 31372 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A1
timestamp 1666464484
transform 1 0 26404 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A2
timestamp 1666464484
transform 1 0 27600 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A2
timestamp 1666464484
transform 1 0 31188 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B2
timestamp 1666464484
transform -1 0 29256 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A1
timestamp 1666464484
transform 1 0 28428 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A2
timestamp 1666464484
transform -1 0 27692 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B1
timestamp 1666464484
transform 1 0 25484 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B2
timestamp 1666464484
transform 1 0 27140 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A1
timestamp 1666464484
transform -1 0 29164 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A2
timestamp 1666464484
transform -1 0 28152 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A2
timestamp 1666464484
transform 1 0 29624 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__B1
timestamp 1666464484
transform 1 0 29440 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__B2
timestamp 1666464484
transform 1 0 29072 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A1
timestamp 1666464484
transform 1 0 35788 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__B1
timestamp 1666464484
transform 1 0 34684 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__B2
timestamp 1666464484
transform -1 0 35788 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A2
timestamp 1666464484
transform 1 0 50968 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B1
timestamp 1666464484
transform 1 0 52900 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A2
timestamp 1666464484
transform 1 0 31556 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B1
timestamp 1666464484
transform 1 0 30636 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B2
timestamp 1666464484
transform -1 0 30636 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__C1
timestamp 1666464484
transform -1 0 31924 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A1
timestamp 1666464484
transform -1 0 31832 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A2
timestamp 1666464484
transform 1 0 32844 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__B1
timestamp 1666464484
transform 1 0 31096 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__B2
timestamp 1666464484
transform -1 0 33580 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A2
timestamp 1666464484
transform -1 0 35788 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__B2
timestamp 1666464484
transform -1 0 36340 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A2
timestamp 1666464484
transform 1 0 50876 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B1
timestamp 1666464484
transform -1 0 53084 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A2
timestamp 1666464484
transform 1 0 34224 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B1
timestamp 1666464484
transform -1 0 32476 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B2
timestamp 1666464484
transform -1 0 32476 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__C1
timestamp 1666464484
transform 1 0 34868 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A2
timestamp 1666464484
transform -1 0 34960 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B1
timestamp 1666464484
transform 1 0 33948 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B2
timestamp 1666464484
transform -1 0 35512 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A1
timestamp 1666464484
transform -1 0 35420 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A2
timestamp 1666464484
transform -1 0 35972 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B2
timestamp 1666464484
transform -1 0 35328 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A2
timestamp 1666464484
transform 1 0 50324 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__B1
timestamp 1666464484
transform 1 0 50876 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A2
timestamp 1666464484
transform -1 0 33948 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B1
timestamp 1666464484
transform 1 0 33212 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B2
timestamp 1666464484
transform 1 0 32660 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__C1
timestamp 1666464484
transform 1 0 35696 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A1
timestamp 1666464484
transform 1 0 31832 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A2
timestamp 1666464484
transform 1 0 32292 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__B1
timestamp 1666464484
transform 1 0 31280 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__B2
timestamp 1666464484
transform -1 0 33580 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A2
timestamp 1666464484
transform 1 0 35144 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B1
timestamp 1666464484
transform -1 0 35604 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B2
timestamp 1666464484
transform -1 0 35052 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A2
timestamp 1666464484
transform -1 0 51796 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__B1
timestamp 1666464484
transform 1 0 51428 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A2
timestamp 1666464484
transform 1 0 33212 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__B1
timestamp 1666464484
transform -1 0 32844 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__B2
timestamp 1666464484
transform -1 0 34316 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__C1
timestamp 1666464484
transform -1 0 35604 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A2
timestamp 1666464484
transform 1 0 34868 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B1
timestamp 1666464484
transform -1 0 34500 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B2
timestamp 1666464484
transform -1 0 36432 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A1
timestamp 1666464484
transform 1 0 32476 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A2
timestamp 1666464484
transform -1 0 35880 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__B2
timestamp 1666464484
transform -1 0 34132 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A1
timestamp 1666464484
transform -1 0 35236 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B1
timestamp 1666464484
transform 1 0 33580 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B2
timestamp 1666464484
transform -1 0 36432 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A1
timestamp 1666464484
transform 1 0 34500 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A2
timestamp 1666464484
transform -1 0 35880 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__B1
timestamp 1666464484
transform 1 0 33028 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__B2
timestamp 1666464484
transform -1 0 33580 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A1
timestamp 1666464484
transform 1 0 36248 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B1
timestamp 1666464484
transform 1 0 34868 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B2
timestamp 1666464484
transform 1 0 36800 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A1
timestamp 1666464484
transform 1 0 34132 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A2
timestamp 1666464484
transform 1 0 35420 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B1
timestamp 1666464484
transform -1 0 33028 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B2
timestamp 1666464484
transform 1 0 32292 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A0
timestamp 1666464484
transform 1 0 22080 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__S
timestamp 1666464484
transform -1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A
timestamp 1666464484
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A3
timestamp 1666464484
transform -1 0 15272 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A
timestamp 1666464484
transform 1 0 15088 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A2
timestamp 1666464484
transform -1 0 8648 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A3
timestamp 1666464484
transform -1 0 9200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A3
timestamp 1666464484
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A3
timestamp 1666464484
transform 1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A3
timestamp 1666464484
transform 1 0 14352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A3
timestamp 1666464484
transform 1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A3
timestamp 1666464484
transform 1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A3
timestamp 1666464484
transform 1 0 13984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A3
timestamp 1666464484
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A3
timestamp 1666464484
transform 1 0 13616 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A3
timestamp 1666464484
transform 1 0 14536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A3
timestamp 1666464484
transform -1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A3
timestamp 1666464484
transform 1 0 15640 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A3
timestamp 1666464484
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A3
timestamp 1666464484
transform 1 0 13432 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A3
timestamp 1666464484
transform -1 0 13248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A3
timestamp 1666464484
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A3
timestamp 1666464484
transform 1 0 13064 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A3
timestamp 1666464484
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A3
timestamp 1666464484
transform -1 0 12696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A3
timestamp 1666464484
transform 1 0 13064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A_N
timestamp 1666464484
transform -1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A3
timestamp 1666464484
transform 1 0 13064 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A_N
timestamp 1666464484
transform 1 0 16192 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A3
timestamp 1666464484
transform -1 0 12696 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__A_N
timestamp 1666464484
transform 1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A3
timestamp 1666464484
transform 1 0 12696 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A_N
timestamp 1666464484
transform -1 0 17388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A3
timestamp 1666464484
transform 1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A_N
timestamp 1666464484
transform 1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A_N
timestamp 1666464484
transform -1 0 17940 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B_N
timestamp 1666464484
transform -1 0 42044 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A
timestamp 1666464484
transform 1 0 44804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__B
timestamp 1666464484
transform -1 0 43884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 1666464484
transform 1 0 43148 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A
timestamp 1666464484
transform 1 0 44252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A
timestamp 1666464484
transform 1 0 43056 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1666464484
transform -1 0 29900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A1
timestamp 1666464484
transform 1 0 40572 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A2
timestamp 1666464484
transform -1 0 40940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A3
timestamp 1666464484
transform -1 0 40204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A1
timestamp 1666464484
transform -1 0 32108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A
timestamp 1666464484
transform 1 0 42504 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1666464484
transform 1 0 32476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__C
timestamp 1666464484
transform 1 0 30728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__D
timestamp 1666464484
transform -1 0 32476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A1
timestamp 1666464484
transform -1 0 37996 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A1
timestamp 1666464484
transform -1 0 31096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A2
timestamp 1666464484
transform 1 0 29808 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A3
timestamp 1666464484
transform -1 0 33028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A1
timestamp 1666464484
transform 1 0 31556 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A2
timestamp 1666464484
transform 1 0 30820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A3
timestamp 1666464484
transform -1 0 32292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__B
timestamp 1666464484
transform 1 0 37444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__B
timestamp 1666464484
transform -1 0 43884 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__B1
timestamp 1666464484
transform -1 0 34316 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__B1
timestamp 1666464484
transform 1 0 41124 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__B
timestamp 1666464484
transform 1 0 28520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__B1
timestamp 1666464484
transform -1 0 30452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__B
timestamp 1666464484
transform 1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A1_N
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__B2
timestamp 1666464484
transform 1 0 26312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A
timestamp 1666464484
transform 1 0 41676 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B1
timestamp 1666464484
transform -1 0 22172 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__B
timestamp 1666464484
transform 1 0 25484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__B1
timestamp 1666464484
transform -1 0 17756 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A
timestamp 1666464484
transform -1 0 45356 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1666464484
transform 1 0 43148 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__B1
timestamp 1666464484
transform -1 0 20332 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1666464484
transform 1 0 30452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A3
timestamp 1666464484
transform -1 0 23092 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A1
timestamp 1666464484
transform -1 0 22172 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A3
timestamp 1666464484
transform -1 0 23092 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A2
timestamp 1666464484
transform -1 0 32476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__B
timestamp 1666464484
transform -1 0 43332 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__B2
timestamp 1666464484
transform 1 0 44160 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A1
timestamp 1666464484
transform -1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__S
timestamp 1666464484
transform 1 0 27508 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A
timestamp 1666464484
transform 1 0 31648 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1666464484
transform -1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A1
timestamp 1666464484
transform -1 0 27968 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A1
timestamp 1666464484
transform -1 0 33672 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A1
timestamp 1666464484
transform 1 0 30820 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A1
timestamp 1666464484
transform 1 0 32476 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A1
timestamp 1666464484
transform 1 0 32384 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A1
timestamp 1666464484
transform -1 0 36156 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A2
timestamp 1666464484
transform 1 0 40020 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A1
timestamp 1666464484
transform -1 0 36708 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A1
timestamp 1666464484
transform -1 0 38916 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A2
timestamp 1666464484
transform 1 0 38180 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A1
timestamp 1666464484
transform -1 0 42780 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A1
timestamp 1666464484
transform -1 0 42872 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A2
timestamp 1666464484
transform 1 0 43240 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A1
timestamp 1666464484
transform 1 0 35788 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A1
timestamp 1666464484
transform 1 0 37076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A2
timestamp 1666464484
transform 1 0 37444 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A
timestamp 1666464484
transform -1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A
timestamp 1666464484
transform 1 0 41124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A1
timestamp 1666464484
transform 1 0 36340 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A2
timestamp 1666464484
transform 1 0 34224 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B2
timestamp 1666464484
transform -1 0 34684 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A
timestamp 1666464484
transform 1 0 33028 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1666464484
transform 1 0 35420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A2
timestamp 1666464484
transform 1 0 35788 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B2
timestamp 1666464484
transform 1 0 33580 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1666464484
transform 1 0 36984 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A1
timestamp 1666464484
transform 1 0 37536 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A2
timestamp 1666464484
transform -1 0 35236 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__B2
timestamp 1666464484
transform -1 0 40296 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1666464484
transform -1 0 35052 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__B
timestamp 1666464484
transform 1 0 42964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__B
timestamp 1666464484
transform 1 0 39284 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A_N
timestamp 1666464484
transform 1 0 41308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A_N
timestamp 1666464484
transform -1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__B
timestamp 1666464484
transform 1 0 29072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A
timestamp 1666464484
transform -1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A2
timestamp 1666464484
transform -1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1666464484
transform -1 0 17756 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A2
timestamp 1666464484
transform 1 0 15272 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__B
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B
timestamp 1666464484
transform -1 0 30544 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A0
timestamp 1666464484
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A
timestamp 1666464484
transform 1 0 28612 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A
timestamp 1666464484
transform -1 0 28612 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A1
timestamp 1666464484
transform -1 0 23552 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A0
timestamp 1666464484
transform -1 0 27876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1666464484
transform -1 0 27324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A0
timestamp 1666464484
transform 1 0 31464 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A
timestamp 1666464484
transform 1 0 34868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A0
timestamp 1666464484
transform -1 0 30176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A
timestamp 1666464484
transform -1 0 29440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A0
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A
timestamp 1666464484
transform 1 0 27508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__B1
timestamp 1666464484
transform 1 0 33396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A1
timestamp 1666464484
transform 1 0 28980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A1
timestamp 1666464484
transform -1 0 26404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A
timestamp 1666464484
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1666464484
transform 1 0 44804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__C
timestamp 1666464484
transform 1 0 44068 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A1
timestamp 1666464484
transform 1 0 36524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__S
timestamp 1666464484
transform -1 0 36156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A
timestamp 1666464484
transform 1 0 33764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A1
timestamp 1666464484
transform 1 0 37260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__S
timestamp 1666464484
transform 1 0 35052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1666464484
transform 1 0 36432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A1
timestamp 1666464484
transform 1 0 35420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__S
timestamp 1666464484
transform 1 0 34500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A
timestamp 1666464484
transform 1 0 33028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A1
timestamp 1666464484
transform 1 0 36708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__S
timestamp 1666464484
transform 1 0 35880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A
timestamp 1666464484
transform 1 0 32292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A1
timestamp 1666464484
transform 1 0 37444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__S
timestamp 1666464484
transform 1 0 33948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__A
timestamp 1666464484
transform -1 0 41860 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A1
timestamp 1666464484
transform 1 0 31372 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__S
timestamp 1666464484
transform 1 0 32660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A
timestamp 1666464484
transform 1 0 29256 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A1
timestamp 1666464484
transform -1 0 19596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__S
timestamp 1666464484
transform -1 0 26588 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A
timestamp 1666464484
transform -1 0 24748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1666464484
transform 1 0 25760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__S
timestamp 1666464484
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__A1
timestamp 1666464484
transform -1 0 14536 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__S
timestamp 1666464484
transform -1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A
timestamp 1666464484
transform -1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A1
timestamp 1666464484
transform -1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__S
timestamp 1666464484
transform 1 0 14996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A
timestamp 1666464484
transform 1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A1
timestamp 1666464484
transform 1 0 16652 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1666464484
transform -1 0 18400 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A1
timestamp 1666464484
transform -1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A
timestamp 1666464484
transform -1 0 20424 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A1
timestamp 1666464484
transform 1 0 42688 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A
timestamp 1666464484
transform -1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A1
timestamp 1666464484
transform 1 0 31556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A
timestamp 1666464484
transform -1 0 42320 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A1
timestamp 1666464484
transform -1 0 21620 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A
timestamp 1666464484
transform 1 0 20792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A1
timestamp 1666464484
transform 1 0 20792 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A
timestamp 1666464484
transform 1 0 22356 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A1
timestamp 1666464484
transform -1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A
timestamp 1666464484
transform 1 0 27784 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A1
timestamp 1666464484
transform -1 0 30176 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1666464484
transform 1 0 28980 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A1
timestamp 1666464484
transform 1 0 29440 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A
timestamp 1666464484
transform 1 0 31372 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A1
timestamp 1666464484
transform -1 0 31464 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A
timestamp 1666464484
transform 1 0 31832 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A1
timestamp 1666464484
transform 1 0 43884 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1666464484
transform -1 0 33488 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A1
timestamp 1666464484
transform 1 0 42596 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A
timestamp 1666464484
transform 1 0 43608 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A1
timestamp 1666464484
transform -1 0 42688 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A
timestamp 1666464484
transform 1 0 43700 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A1
timestamp 1666464484
transform 1 0 43240 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1666464484
transform 1 0 43792 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A
timestamp 1666464484
transform -1 0 50600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__C
timestamp 1666464484
transform 1 0 31004 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__D_N
timestamp 1666464484
transform 1 0 31556 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A0
timestamp 1666464484
transform 1 0 22816 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A0
timestamp 1666464484
transform -1 0 26312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A1
timestamp 1666464484
transform 1 0 24932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A0
timestamp 1666464484
transform 1 0 21344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A0
timestamp 1666464484
transform 1 0 22356 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__A0
timestamp 1666464484
transform -1 0 26220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__A0
timestamp 1666464484
transform -1 0 18308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A0
timestamp 1666464484
transform -1 0 24564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A0
timestamp 1666464484
transform -1 0 25208 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__A0
timestamp 1666464484
transform -1 0 20240 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A0
timestamp 1666464484
transform -1 0 20792 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A0
timestamp 1666464484
transform -1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A0
timestamp 1666464484
transform -1 0 14628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A0
timestamp 1666464484
transform -1 0 16192 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A0
timestamp 1666464484
transform -1 0 14352 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A0
timestamp 1666464484
transform -1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A0
timestamp 1666464484
transform -1 0 13432 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A0
timestamp 1666464484
transform -1 0 14628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A0
timestamp 1666464484
transform -1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A0
timestamp 1666464484
transform -1 0 13800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A0
timestamp 1666464484
transform -1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__A0
timestamp 1666464484
transform -1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A0
timestamp 1666464484
transform -1 0 17204 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A0
timestamp 1666464484
transform -1 0 18308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A0
timestamp 1666464484
transform -1 0 19964 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A0
timestamp 1666464484
transform -1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A0
timestamp 1666464484
transform -1 0 17848 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A0
timestamp 1666464484
transform -1 0 15180 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A0
timestamp 1666464484
transform 1 0 25484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__S
timestamp 1666464484
transform -1 0 24012 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A0
timestamp 1666464484
transform 1 0 25576 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__S
timestamp 1666464484
transform 1 0 24748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A0
timestamp 1666464484
transform 1 0 25668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__S
timestamp 1666464484
transform 1 0 28336 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__A0
timestamp 1666464484
transform 1 0 26956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__S
timestamp 1666464484
transform 1 0 28336 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__CLK
timestamp 1666464484
transform 1 0 39836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__CLK
timestamp 1666464484
transform -1 0 38732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__CLK
timestamp 1666464484
transform -1 0 38180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__CLK
timestamp 1666464484
transform 1 0 40940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__CLK
timestamp 1666464484
transform 1 0 41860 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__CLK
timestamp 1666464484
transform 1 0 42596 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__CLK
timestamp 1666464484
transform 1 0 43516 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__CLK
timestamp 1666464484
transform -1 0 44436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__CLK
timestamp 1666464484
transform 1 0 44344 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__CLK
timestamp 1666464484
transform 1 0 44252 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__CLK
timestamp 1666464484
transform 1 0 43700 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__CLK
timestamp 1666464484
transform 1 0 43240 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__CLK
timestamp 1666464484
transform 1 0 43056 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__CLK
timestamp 1666464484
transform -1 0 43608 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__CLK
timestamp 1666464484
transform 1 0 41400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__CLK
timestamp 1666464484
transform 1 0 41952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__CLK
timestamp 1666464484
transform 1 0 42412 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__CLK
timestamp 1666464484
transform -1 0 42780 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__CLK
timestamp 1666464484
transform 1 0 41492 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__CLK
timestamp 1666464484
transform 1 0 41860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__CLK
timestamp 1666464484
transform -1 0 27140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__CLK
timestamp 1666464484
transform 1 0 24564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__CLK
timestamp 1666464484
transform -1 0 15180 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__CLK
timestamp 1666464484
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__CLK
timestamp 1666464484
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__CLK
timestamp 1666464484
transform 1 0 18768 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__CLK
timestamp 1666464484
transform 1 0 35880 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__CLK
timestamp 1666464484
transform -1 0 29072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__CLK
timestamp 1666464484
transform 1 0 21344 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__CLK
timestamp 1666464484
transform 1 0 22632 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__CLK
timestamp 1666464484
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__CLK
timestamp 1666464484
transform 1 0 34224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__CLK
timestamp 1666464484
transform 1 0 37444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__CLK
timestamp 1666464484
transform 1 0 23368 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__CLK
timestamp 1666464484
transform 1 0 42596 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__CLK
timestamp 1666464484
transform 1 0 41952 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__CLK
timestamp 1666464484
transform -1 0 43056 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__CLK
timestamp 1666464484
transform 1 0 42596 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__CLK
timestamp 1666464484
transform 1 0 48208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__CLK
timestamp 1666464484
transform 1 0 42596 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__CLK
timestamp 1666464484
transform 1 0 36064 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__CLK
timestamp 1666464484
transform 1 0 43148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__CLK
timestamp 1666464484
transform -1 0 52440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__A
timestamp 1666464484
transform 1 0 37444 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__A
timestamp 1666464484
transform 1 0 37996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__A
timestamp 1666464484
transform 1 0 38732 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__A
timestamp 1666464484
transform 1 0 39836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__A
timestamp 1666464484
transform 1 0 41308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__A
timestamp 1666464484
transform 1 0 41676 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1666464484
transform 1 0 43700 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_wb_clk_i_A
timestamp 1666464484
transform -1 0 25300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_wb_clk_i_A
timestamp 1666464484
transform -1 0 28060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_wb_clk_i_A
timestamp 1666464484
transform -1 0 14536 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_wb_clk_i_A
timestamp 1666464484
transform 1 0 16100 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_wb_clk_i_A
timestamp 1666464484
transform 1 0 43148 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_wb_clk_i_A
timestamp 1666464484
transform 1 0 43792 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_wb_clk_i_A
timestamp 1666464484
transform 1 0 43148 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_wb_clk_i_A
timestamp 1666464484
transform -1 0 44436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout355_A
timestamp 1666464484
transform -1 0 43516 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout356_A
timestamp 1666464484
transform -1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 53084 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 53084 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform 1 0 52900 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 51888 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 51796 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 51888 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform 1 0 52900 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 52440 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 52440 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 52440 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 53084 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1666464484
transform -1 0 51796 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1666464484
transform -1 0 51888 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1666464484
transform -1 0 51796 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1666464484
transform -1 0 51888 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1666464484
transform -1 0 52440 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1666464484
transform -1 0 53084 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1666464484
transform -1 0 51796 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1666464484
transform -1 0 52440 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1666464484
transform -1 0 52440 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1666464484
transform -1 0 52440 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1666464484
transform -1 0 51888 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1666464484
transform -1 0 52440 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1666464484
transform -1 0 51796 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1666464484
transform -1 0 51152 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1666464484
transform -1 0 51244 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1666464484
transform -1 0 53084 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1666464484
transform -1 0 2484 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1666464484
transform -1 0 2484 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1666464484
transform -1 0 2944 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1666464484
transform -1 0 2392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1666464484
transform -1 0 2392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1666464484
transform -1 0 3036 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1666464484
transform -1 0 2944 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1666464484
transform -1 0 2392 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1666464484
transform -1 0 53084 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1666464484
transform -1 0 51796 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1666464484
transform -1 0 50600 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1666464484
transform 1 0 52900 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1666464484
transform -1 0 49864 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1666464484
transform -1 0 51796 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1666464484
transform -1 0 50232 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1666464484
transform 1 0 52900 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1666464484
transform -1 0 52440 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1666464484
transform -1 0 53084 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1666464484
transform -1 0 50784 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1666464484
transform -1 0 51888 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1666464484
transform -1 0 52716 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1666464484
transform -1 0 53268 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1666464484
transform -1 0 51888 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1666464484
transform -1 0 54372 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1666464484
transform -1 0 52440 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1666464484
transform -1 0 53728 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1666464484
transform -1 0 51244 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1666464484
transform -1 0 52440 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1666464484
transform -1 0 51796 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1666464484
transform -1 0 51152 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1666464484
transform -1 0 52348 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1666464484
transform -1 0 51244 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1666464484
transform -1 0 51152 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1666464484
transform 1 0 52900 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1666464484
transform -1 0 51244 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1666464484
transform -1 0 3036 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1666464484
transform -1 0 3036 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1666464484
transform -1 0 3036 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1666464484
transform -1 0 3036 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1666464484
transform -1 0 3036 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1666464484
transform -1 0 3036 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1666464484
transform -1 0 3036 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1666464484
transform -1 0 3036 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1666464484
transform -1 0 3036 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1666464484
transform -1 0 3036 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1666464484
transform -1 0 3036 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1666464484
transform -1 0 3036 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1666464484
transform -1 0 2484 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1666464484
transform -1 0 3036 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1666464484
transform -1 0 3036 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1666464484
transform -1 0 2484 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1666464484
transform -1 0 3036 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1666464484
transform -1 0 3036 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1666464484
transform -1 0 2484 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1666464484
transform -1 0 3036 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1666464484
transform -1 0 3036 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1666464484
transform -1 0 3036 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1666464484
transform -1 0 3036 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1666464484
transform -1 0 3036 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1666464484
transform -1 0 3036 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1666464484
transform -1 0 3036 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1666464484
transform -1 0 3036 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1666464484
transform -1 0 10948 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1666464484
transform -1 0 22908 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1666464484
transform -1 0 24104 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1666464484
transform -1 0 26496 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1666464484
transform -1 0 26680 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1666464484
transform -1 0 28060 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1666464484
transform -1 0 29256 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1666464484
transform -1 0 31280 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1666464484
transform -1 0 31832 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1666464484
transform -1 0 32936 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1666464484
transform -1 0 34040 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1666464484
transform -1 0 12144 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1666464484
transform -1 0 36064 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1666464484
transform -1 0 36432 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1666464484
transform -1 0 38456 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1666464484
transform -1 0 38824 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1666464484
transform -1 0 40848 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1666464484
transform -1 0 42044 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1666464484
transform -1 0 42596 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1666464484
transform 1 0 13616 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1666464484
transform -1 0 15272 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1666464484
transform -1 0 17020 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1666464484
transform -1 0 16928 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1666464484
transform -1 0 18952 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1666464484
transform -1 0 19688 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1666464484
transform -1 0 20516 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1666464484
transform -1 0 22080 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1666464484
transform 1 0 47104 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1666464484
transform -1 0 51980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1666464484
transform -1 0 51060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1666464484
transform -1 0 49036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input121_A
timestamp 1666464484
transform -1 0 48484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input122_A
timestamp 1666464484
transform -1 0 49220 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input123_A
timestamp 1666464484
transform -1 0 49588 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input124_A
timestamp 1666464484
transform -1 0 50324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input125_A
timestamp 1666464484
transform -1 0 50508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input126_A
timestamp 1666464484
transform -1 0 53084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input127_A
timestamp 1666464484
transform -1 0 52348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input128_A
timestamp 1666464484
transform -1 0 52532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input129_A
timestamp 1666464484
transform -1 0 45356 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input130_A
timestamp 1666464484
transform -1 0 46000 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input131_A
timestamp 1666464484
transform -1 0 47288 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_A
timestamp 1666464484
transform -1 0 48024 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_A
timestamp 1666464484
transform -1 0 49864 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_A
timestamp 1666464484
transform -1 0 51612 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_A
timestamp 1666464484
transform -1 0 51612 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input136_A
timestamp 1666464484
transform -1 0 53176 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input137_A
timestamp 1666464484
transform -1 0 3036 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input138_A
timestamp 1666464484
transform -1 0 3036 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input139_A
timestamp 1666464484
transform -1 0 2944 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input140_A
timestamp 1666464484
transform -1 0 2392 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input141_A
timestamp 1666464484
transform -1 0 3036 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input142_A
timestamp 1666464484
transform -1 0 3036 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input143_A
timestamp 1666464484
transform -1 0 3036 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input144_A
timestamp 1666464484
transform -1 0 2392 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input145_A
timestamp 1666464484
transform -1 0 2944 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input146_A
timestamp 1666464484
transform -1 0 3588 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input147_A
timestamp 1666464484
transform -1 0 3220 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input148_A
timestamp 1666464484
transform -1 0 4140 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input149_A
timestamp 1666464484
transform -1 0 4968 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input150_A
timestamp 1666464484
transform -1 0 6532 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input151_A
timestamp 1666464484
transform -1 0 7728 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input152_A
timestamp 1666464484
transform -1 0 8648 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input153_A
timestamp 1666464484
transform -1 0 10120 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input154_A
timestamp 1666464484
transform -1 0 3036 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input155_A
timestamp 1666464484
transform -1 0 2392 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input156_A
timestamp 1666464484
transform -1 0 2944 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input157_A
timestamp 1666464484
transform -1 0 3036 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input158_A
timestamp 1666464484
transform -1 0 3036 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input159_A
timestamp 1666464484
transform -1 0 3036 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input160_A
timestamp 1666464484
transform -1 0 2392 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input161_A
timestamp 1666464484
transform -1 0 2944 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input162_A
timestamp 1666464484
transform -1 0 54372 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input163_A
timestamp 1666464484
transform -1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input164_A
timestamp 1666464484
transform -1 0 8096 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input165_A
timestamp 1666464484
transform -1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input166_A
timestamp 1666464484
transform -1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input167_A
timestamp 1666464484
transform -1 0 10028 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input168_A
timestamp 1666464484
transform -1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input169_A
timestamp 1666464484
transform -1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input170_A
timestamp 1666464484
transform -1 0 10764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input171_A
timestamp 1666464484
transform -1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input172_A
timestamp 1666464484
transform -1 0 10672 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input173_A
timestamp 1666464484
transform -1 0 11684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input174_A
timestamp 1666464484
transform -1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input175_A
timestamp 1666464484
transform -1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input176_A
timestamp 1666464484
transform -1 0 13524 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input177_A
timestamp 1666464484
transform -1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input178_A
timestamp 1666464484
transform -1 0 15088 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input179_A
timestamp 1666464484
transform -1 0 14168 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input180_A
timestamp 1666464484
transform -1 0 15456 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input181_A
timestamp 1666464484
transform -1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input182_A
timestamp 1666464484
transform -1 0 14720 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input183_A
timestamp 1666464484
transform -1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input184_A
timestamp 1666464484
transform -1 0 16560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input185_A
timestamp 1666464484
transform -1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input186_A
timestamp 1666464484
transform -1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input187_A
timestamp 1666464484
transform -1 0 17572 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input188_A
timestamp 1666464484
transform -1 0 17848 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input189_A
timestamp 1666464484
transform -1 0 18308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input190_A
timestamp 1666464484
transform -1 0 19596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input191_A
timestamp 1666464484
transform -1 0 6900 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input192_A
timestamp 1666464484
transform -1 0 6532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input193_A
timestamp 1666464484
transform -1 0 4968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input194_A
timestamp 1666464484
transform -1 0 8188 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input195_A
timestamp 1666464484
transform -1 0 7544 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input196_A
timestamp 1666464484
transform 1 0 52900 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input197_A
timestamp 1666464484
transform -1 0 53820 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input198_A
timestamp 1666464484
transform -1 0 2484 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input199_A
timestamp 1666464484
transform -1 0 43608 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input200_A
timestamp 1666464484
transform -1 0 3036 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input201_A
timestamp 1666464484
transform -1 0 54372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input202_A
timestamp 1666464484
transform -1 0 52440 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input203_A
timestamp 1666464484
transform -1 0 52900 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input204_A
timestamp 1666464484
transform -1 0 52532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input205_A
timestamp 1666464484
transform -1 0 51888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input206_A
timestamp 1666464484
transform -1 0 51244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input207_A
timestamp 1666464484
transform -1 0 53636 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input208_A
timestamp 1666464484
transform -1 0 53636 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input209_A
timestamp 1666464484
transform -1 0 52900 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input210_A
timestamp 1666464484
transform -1 0 53636 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input211_A
timestamp 1666464484
transform -1 0 53636 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input212_A
timestamp 1666464484
transform -1 0 53636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input213_A
timestamp 1666464484
transform -1 0 52900 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input214_A
timestamp 1666464484
transform -1 0 53636 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input215_A
timestamp 1666464484
transform -1 0 53636 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input216_A
timestamp 1666464484
transform -1 0 53636 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input217_A
timestamp 1666464484
transform -1 0 53084 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input218_A
timestamp 1666464484
transform -1 0 53084 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input219_A
timestamp 1666464484
transform -1 0 53636 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input220_A
timestamp 1666464484
transform -1 0 52440 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input221_A
timestamp 1666464484
transform -1 0 51888 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input222_A
timestamp 1666464484
transform -1 0 52900 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input223_A
timestamp 1666464484
transform -1 0 53084 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input224_A
timestamp 1666464484
transform -1 0 53636 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input225_A
timestamp 1666464484
transform -1 0 53636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input226_A
timestamp 1666464484
transform -1 0 53636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input227_A
timestamp 1666464484
transform -1 0 52900 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input228_A
timestamp 1666464484
transform -1 0 53636 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input229_A
timestamp 1666464484
transform -1 0 53636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input230_A
timestamp 1666464484
transform -1 0 53636 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input231_A
timestamp 1666464484
transform -1 0 52900 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input232_A
timestamp 1666464484
transform -1 0 53636 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input233_A
timestamp 1666464484
transform -1 0 53636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input234_A
timestamp 1666464484
transform -1 0 51796 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output235_A
timestamp 1666464484
transform 1 0 2208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output263_A
timestamp 1666464484
transform 1 0 36800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output266_A
timestamp 1666464484
transform -1 0 39100 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output267_A
timestamp 1666464484
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output268_A
timestamp 1666464484
transform -1 0 39468 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output270_A
timestamp 1666464484
transform -1 0 40572 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output272_A
timestamp 1666464484
transform -1 0 41124 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output274_A
timestamp 1666464484
transform 1 0 41308 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output275_A
timestamp 1666464484
transform -1 0 43148 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output276_A
timestamp 1666464484
transform 1 0 42412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output278_A
timestamp 1666464484
transform -1 0 43700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output289_A
timestamp 1666464484
transform -1 0 47564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output290_A
timestamp 1666464484
transform 1 0 22632 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output291_A
timestamp 1666464484
transform 1 0 23736 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output292_A
timestamp 1666464484
transform 1 0 23184 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output293_A
timestamp 1666464484
transform -1 0 23828 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output294_A
timestamp 1666464484
transform -1 0 23276 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output295_A
timestamp 1666464484
transform 1 0 25300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output296_A
timestamp 1666464484
transform -1 0 24932 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output297_A
timestamp 1666464484
transform 1 0 24196 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output298_A
timestamp 1666464484
transform 1 0 25944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output299_A
timestamp 1666464484
transform 1 0 26496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output300_A
timestamp 1666464484
transform 1 0 26680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output301_A
timestamp 1666464484
transform 1 0 26128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output302_A
timestamp 1666464484
transform 1 0 27324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output303_A
timestamp 1666464484
transform 1 0 27876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output304_A
timestamp 1666464484
transform -1 0 29164 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output305_A
timestamp 1666464484
transform 1 0 28520 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output306_A
timestamp 1666464484
transform 1 0 31556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output307_A
timestamp 1666464484
transform 1 0 29532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output308_A
timestamp 1666464484
transform 1 0 30820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output309_A
timestamp 1666464484
transform 1 0 30452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output310_A
timestamp 1666464484
transform 1 0 31740 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output311_A
timestamp 1666464484
transform 1 0 31188 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output312_A
timestamp 1666464484
transform 1 0 32660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output313_A
timestamp 1666464484
transform 1 0 32660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output314_A
timestamp 1666464484
transform 1 0 33764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output315_A
timestamp 1666464484
transform 1 0 33212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output316_A
timestamp 1666464484
transform 1 0 34868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output317_A
timestamp 1666464484
transform 1 0 2300 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output319_A
timestamp 1666464484
transform 1 0 2300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output320_A
timestamp 1666464484
transform -1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output322_A
timestamp 1666464484
transform 1 0 2300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output323_A
timestamp 1666464484
transform -1 0 2484 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output324_A
timestamp 1666464484
transform -1 0 2484 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output326_A
timestamp 1666464484
transform -1 0 2484 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output331_A
timestamp 1666464484
transform 1 0 53452 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output339_A
timestamp 1666464484
transform 1 0 52256 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output341_A
timestamp 1666464484
transform 1 0 52716 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output342_A
timestamp 1666464484
transform 1 0 52900 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output343_A
timestamp 1666464484
transform 1 0 52256 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output344_A
timestamp 1666464484
transform 1 0 52900 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output345_A
timestamp 1666464484
transform 1 0 53452 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output346_A
timestamp 1666464484
transform 1 0 53452 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48
timestamp 1666464484
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1666464484
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1666464484
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1666464484
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1666464484
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1666464484
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1666464484
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1666464484
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1666464484
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1666464484
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1666464484
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145
timestamp 1666464484
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 1666464484
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp 1666464484
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666464484
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1666464484
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 1666464484
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1666464484
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666464484
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1666464484
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_208
timestamp 1666464484
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1666464484
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666464484
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_229
timestamp 1666464484
transform 1 0 22172 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_234
timestamp 1666464484
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_242
timestamp 1666464484
transform 1 0 23368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1666464484
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_257
timestamp 1666464484
transform 1 0 24748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1666464484
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_270
timestamp 1666464484
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1666464484
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_285
timestamp 1666464484
transform 1 0 27324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1666464484
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_298
timestamp 1666464484
transform 1 0 28520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1666464484
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1666464484
transform 1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_323
timestamp 1666464484
transform 1 0 30820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_331
timestamp 1666464484
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1666464484
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_343
timestamp 1666464484
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_351
timestamp 1666464484
transform 1 0 33396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1666464484
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1666464484
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1666464484
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_370
timestamp 1666464484
transform 1 0 35144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1666464484
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_384
timestamp 1666464484
transform 1 0 36432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1666464484
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1666464484
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_399
timestamp 1666464484
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_407
timestamp 1666464484
transform 1 0 38548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415
timestamp 1666464484
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1666464484
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666464484
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_427
timestamp 1666464484
transform 1 0 40388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_435
timestamp 1666464484
transform 1 0 41124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_443
timestamp 1666464484
transform 1 0 41860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1666464484
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666464484
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_455
timestamp 1666464484
transform 1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_463
timestamp 1666464484
transform 1 0 43700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1666464484
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1666464484
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1666464484
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_483
timestamp 1666464484
transform 1 0 45540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_491
timestamp 1666464484
transform 1 0 46276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_499
timestamp 1666464484
transform 1 0 47012 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1666464484
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1666464484
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_511
timestamp 1666464484
transform 1 0 48116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_519
timestamp 1666464484
transform 1 0 48852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_527
timestamp 1666464484
transform 1 0 49588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1666464484
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1666464484
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_539
timestamp 1666464484
transform 1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_547
timestamp 1666464484
transform 1 0 51428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_555
timestamp 1666464484
transform 1 0 52164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1666464484
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_561
timestamp 1666464484
transform 1 0 52716 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_565
timestamp 1666464484
transform 1 0 53084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_577
timestamp 1666464484
transform 1 0 54188 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1666464484
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_63
timestamp 1666464484
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_67
timestamp 1666464484
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1666464484
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_88
timestamp 1666464484
transform 1 0 9200 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_95
timestamp 1666464484
transform 1 0 9844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1666464484
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_126
timestamp 1666464484
transform 1 0 12696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1666464484
transform 1 0 13340 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1666464484
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_150
timestamp 1666464484
transform 1 0 14904 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_154
timestamp 1666464484
transform 1 0 15272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1666464484
transform 1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_162
timestamp 1666464484
transform 1 0 16008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1666464484
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_175
timestamp 1666464484
transform 1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_182
timestamp 1666464484
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_186
timestamp 1666464484
transform 1 0 18216 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_190
timestamp 1666464484
transform 1 0 18584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_194
timestamp 1666464484
transform 1 0 18952 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_198
timestamp 1666464484
transform 1 0 19320 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1666464484
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_214
timestamp 1666464484
transform 1 0 20792 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_218
timestamp 1666464484
transform 1 0 21160 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1666464484
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1666464484
transform 1 0 22356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_238
timestamp 1666464484
transform 1 0 23000 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_246
timestamp 1666464484
transform 1 0 23736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_254
timestamp 1666464484
transform 1 0 24472 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1666464484
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_270
timestamp 1666464484
transform 1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1666464484
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_291
timestamp 1666464484
transform 1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_299
timestamp 1666464484
transform 1 0 28612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_305
timestamp 1666464484
transform 1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_311
timestamp 1666464484
transform 1 0 29716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_319
timestamp 1666464484
transform 1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_327
timestamp 1666464484
transform 1 0 31188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1666464484
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_343
timestamp 1666464484
transform 1 0 32660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_351
timestamp 1666464484
transform 1 0 33396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_358
timestamp 1666464484
transform 1 0 34040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_365
timestamp 1666464484
transform 1 0 34684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_372
timestamp 1666464484
transform 1 0 35328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_379
timestamp 1666464484
transform 1 0 35972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp 1666464484
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1666464484
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1666464484
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_411
timestamp 1666464484
transform 1 0 38916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1666464484
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_427
timestamp 1666464484
transform 1 0 40388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_435
timestamp 1666464484
transform 1 0 41124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_443
timestamp 1666464484
transform 1 0 41860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1666464484
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1666464484
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_455
timestamp 1666464484
transform 1 0 42964 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_463
timestamp 1666464484
transform 1 0 43700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_471
timestamp 1666464484
transform 1 0 44436 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_479
timestamp 1666464484
transform 1 0 45172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1666464484
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_495
timestamp 1666464484
transform 1 0 46644 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_499
timestamp 1666464484
transform 1 0 47012 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1666464484
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1666464484
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_511
timestamp 1666464484
transform 1 0 48116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_519
timestamp 1666464484
transform 1 0 48852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_527
timestamp 1666464484
transform 1 0 49588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_535
timestamp 1666464484
transform 1 0 50324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1666464484
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_551
timestamp 1666464484
transform 1 0 51796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_557
timestamp 1666464484
transform 1 0 52348 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1666464484
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_573
timestamp 1666464484
transform 1 0 53820 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_9
timestamp 1666464484
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1666464484
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_59
timestamp 1666464484
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_66
timestamp 1666464484
transform 1 0 7176 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1666464484
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1666464484
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1666464484
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_115
timestamp 1666464484
transform 1 0 11684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_126
timestamp 1666464484
transform 1 0 12696 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_134
timestamp 1666464484
transform 1 0 13432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1666464484
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_152
timestamp 1666464484
transform 1 0 15088 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_162
timestamp 1666464484
transform 1 0 16008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_168
timestamp 1666464484
transform 1 0 16560 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_176
timestamp 1666464484
transform 1 0 17296 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_179
timestamp 1666464484
transform 1 0 17572 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1666464484
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_206
timestamp 1666464484
transform 1 0 20056 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_218
timestamp 1666464484
transform 1 0 21160 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_224
timestamp 1666464484
transform 1 0 21712 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_233
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1666464484
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1666464484
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_263
timestamp 1666464484
transform 1 0 25300 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_271
timestamp 1666464484
transform 1 0 26036 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_274
timestamp 1666464484
transform 1 0 26312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_280
timestamp 1666464484
transform 1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_284
timestamp 1666464484
transform 1 0 27232 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_287
timestamp 1666464484
transform 1 0 27508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_293
timestamp 1666464484
transform 1 0 28060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_297
timestamp 1666464484
transform 1 0 28428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1666464484
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_317
timestamp 1666464484
transform 1 0 30268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_321
timestamp 1666464484
transform 1 0 30636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_329
timestamp 1666464484
transform 1 0 31372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_335
timestamp 1666464484
transform 1 0 31924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_345
timestamp 1666464484
transform 1 0 32844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_351
timestamp 1666464484
transform 1 0 33396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1666464484
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1666464484
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1666464484
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_369
timestamp 1666464484
transform 1 0 35052 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_377
timestamp 1666464484
transform 1 0 35788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_382
timestamp 1666464484
transform 1 0 36248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_389
timestamp 1666464484
transform 1 0 36892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_396
timestamp 1666464484
transform 1 0 37536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_403
timestamp 1666464484
transform 1 0 38180 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_414
timestamp 1666464484
transform 1 0 39192 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1666464484
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_426
timestamp 1666464484
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 1666464484
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_439
timestamp 1666464484
transform 1 0 41492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_446
timestamp 1666464484
transform 1 0 42136 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_458
timestamp 1666464484
transform 1 0 43240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_465
timestamp 1666464484
transform 1 0 43884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1666464484
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1666464484
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_482
timestamp 1666464484
transform 1 0 45448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_486
timestamp 1666464484
transform 1 0 45816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_491
timestamp 1666464484
transform 1 0 46276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_499
timestamp 1666464484
transform 1 0 47012 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_505
timestamp 1666464484
transform 1 0 47564 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_515
timestamp 1666464484
transform 1 0 48484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_521
timestamp 1666464484
transform 1 0 49036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_527
timestamp 1666464484
transform 1 0 49588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1666464484
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1666464484
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_537
timestamp 1666464484
transform 1 0 50508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_547
timestamp 1666464484
transform 1 0 51428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_553
timestamp 1666464484
transform 1 0 51980 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_559
timestamp 1666464484
transform 1 0 52532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_571
timestamp 1666464484
transform 1 0 53636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_579
timestamp 1666464484
transform 1 0 54372 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_9
timestamp 1666464484
transform 1 0 1932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_21
timestamp 1666464484
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_33
timestamp 1666464484
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_45
timestamp 1666464484
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1666464484
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_63
timestamp 1666464484
transform 1 0 6900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_67
timestamp 1666464484
transform 1 0 7268 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_70
timestamp 1666464484
transform 1 0 7544 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_76
timestamp 1666464484
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_82
timestamp 1666464484
transform 1 0 8648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_88
timestamp 1666464484
transform 1 0 9200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1666464484
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1666464484
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_117
timestamp 1666464484
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_124
timestamp 1666464484
transform 1 0 12512 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_132
timestamp 1666464484
transform 1 0 13248 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1666464484
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_139
timestamp 1666464484
transform 1 0 13892 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_142
timestamp 1666464484
transform 1 0 14168 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_148
timestamp 1666464484
transform 1 0 14720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_154
timestamp 1666464484
transform 1 0 15272 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1666464484
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_177
timestamp 1666464484
transform 1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_182
timestamp 1666464484
transform 1 0 17848 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_194
timestamp 1666464484
transform 1 0 18952 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_206
timestamp 1666464484
transform 1 0 20056 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1666464484
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1666464484
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_241
timestamp 1666464484
transform 1 0 23276 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_247
timestamp 1666464484
transform 1 0 23828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_253
timestamp 1666464484
transform 1 0 24380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_259
timestamp 1666464484
transform 1 0 24932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_265
timestamp 1666464484
transform 1 0 25484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_269
timestamp 1666464484
transform 1 0 25852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_272
timestamp 1666464484
transform 1 0 26128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1666464484
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1666464484
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1666464484
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_317
timestamp 1666464484
transform 1 0 30268 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_325
timestamp 1666464484
transform 1 0 31004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_333
timestamp 1666464484
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_345
timestamp 1666464484
transform 1 0 32844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_357
timestamp 1666464484
transform 1 0 33948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_369
timestamp 1666464484
transform 1 0 35052 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_381
timestamp 1666464484
transform 1 0 36156 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_390
timestamp 1666464484
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1666464484
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_397
timestamp 1666464484
transform 1 0 37628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_403
timestamp 1666464484
transform 1 0 38180 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_411
timestamp 1666464484
transform 1 0 38916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_417
timestamp 1666464484
transform 1 0 39468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_423
timestamp 1666464484
transform 1 0 40020 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_429
timestamp 1666464484
transform 1 0 40572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_435
timestamp 1666464484
transform 1 0 41124 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_443
timestamp 1666464484
transform 1 0 41860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1666464484
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_449
timestamp 1666464484
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_455
timestamp 1666464484
transform 1 0 42964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_461
timestamp 1666464484
transform 1 0 43516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_468
timestamp 1666464484
transform 1 0 44160 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_475
timestamp 1666464484
transform 1 0 44804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_482
timestamp 1666464484
transform 1 0 45448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_489
timestamp 1666464484
transform 1 0 46092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_496
timestamp 1666464484
transform 1 0 46736 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1666464484
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_517
timestamp 1666464484
transform 1 0 48668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_523
timestamp 1666464484
transform 1 0 49220 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_531
timestamp 1666464484
transform 1 0 49956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_535
timestamp 1666464484
transform 1 0 50324 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_543
timestamp 1666464484
transform 1 0 51060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_555
timestamp 1666464484
transform 1 0 52164 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1666464484
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1666464484
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_573
timestamp 1666464484
transform 1 0 53820 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_9
timestamp 1666464484
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1666464484
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_69
timestamp 1666464484
transform 1 0 7452 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp 1666464484
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_92
timestamp 1666464484
transform 1 0 9568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_98
timestamp 1666464484
transform 1 0 10120 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_115
timestamp 1666464484
transform 1 0 11684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_125
timestamp 1666464484
transform 1 0 12604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1666464484
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1666464484
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_150
timestamp 1666464484
transform 1 0 14904 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_156
timestamp 1666464484
transform 1 0 15456 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_168
timestamp 1666464484
transform 1 0 16560 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_180
timestamp 1666464484
transform 1 0 17664 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1666464484
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_233
timestamp 1666464484
transform 1 0 22540 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_236
timestamp 1666464484
transform 1 0 22816 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_242
timestamp 1666464484
transform 1 0 23368 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1666464484
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_259
timestamp 1666464484
transform 1 0 24932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_262
timestamp 1666464484
transform 1 0 25208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_268
timestamp 1666464484
transform 1 0 25760 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_274
timestamp 1666464484
transform 1 0 26312 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_286
timestamp 1666464484
transform 1 0 27416 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_298
timestamp 1666464484
transform 1 0 28520 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1666464484
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1666464484
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1666464484
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1666464484
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1666464484
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1666464484
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1666464484
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1666464484
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1666464484
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_401
timestamp 1666464484
transform 1 0 37996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_407
timestamp 1666464484
transform 1 0 38548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1666464484
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1666464484
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1666464484
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_433
timestamp 1666464484
transform 1 0 40940 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_439
timestamp 1666464484
transform 1 0 41492 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_447
timestamp 1666464484
transform 1 0 42228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_451
timestamp 1666464484
transform 1 0 42596 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_457
timestamp 1666464484
transform 1 0 43148 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_463
timestamp 1666464484
transform 1 0 43700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1666464484
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_477
timestamp 1666464484
transform 1 0 44988 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_486
timestamp 1666464484
transform 1 0 45816 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_498
timestamp 1666464484
transform 1 0 46920 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_510
timestamp 1666464484
transform 1 0 48024 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_522
timestamp 1666464484
transform 1 0 49128 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_530
timestamp 1666464484
transform 1 0 49864 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1666464484
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1666464484
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1666464484
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1666464484
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1666464484
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1666464484
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1666464484
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1666464484
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1666464484
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 1666464484
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_90
timestamp 1666464484
transform 1 0 9384 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_94
timestamp 1666464484
transform 1 0 9752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_97
timestamp 1666464484
transform 1 0 10028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_101
timestamp 1666464484
transform 1 0 10396 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_104
timestamp 1666464484
transform 1 0 10672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1666464484
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_117
timestamp 1666464484
transform 1 0 11868 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_130
timestamp 1666464484
transform 1 0 13064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_140
timestamp 1666464484
transform 1 0 13984 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_146
timestamp 1666464484
transform 1 0 14536 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_152
timestamp 1666464484
transform 1 0 15088 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1666464484
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_255
timestamp 1666464484
transform 1 0 24564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_267
timestamp 1666464484
transform 1 0 25668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1666464484
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_285
timestamp 1666464484
transform 1 0 27324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_291
timestamp 1666464484
transform 1 0 27876 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_299
timestamp 1666464484
transform 1 0 28612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_305
timestamp 1666464484
transform 1 0 29164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_308
timestamp 1666464484
transform 1 0 29440 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_316
timestamp 1666464484
transform 1 0 30176 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_322
timestamp 1666464484
transform 1 0 30728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1666464484
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666464484
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1666464484
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1666464484
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1666464484
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1666464484
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1666464484
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1666464484
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1666464484
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1666464484
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1666464484
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1666464484
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1666464484
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1666464484
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1666464484
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1666464484
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1666464484
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1666464484
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1666464484
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1666464484
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1666464484
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1666464484
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1666464484
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1666464484
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1666464484
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_573
timestamp 1666464484
transform 1 0 53820 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_9
timestamp 1666464484
transform 1 0 1932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1666464484
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_105
timestamp 1666464484
transform 1 0 10764 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_116
timestamp 1666464484
transform 1 0 11776 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_126
timestamp 1666464484
transform 1 0 12696 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 1666464484
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_145
timestamp 1666464484
transform 1 0 14444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_157
timestamp 1666464484
transform 1 0 15548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_169
timestamp 1666464484
transform 1 0 16652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_181
timestamp 1666464484
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1666464484
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_238
timestamp 1666464484
transform 1 0 23000 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_244
timestamp 1666464484
transform 1 0 23552 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1666464484
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_257
timestamp 1666464484
transform 1 0 24748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_263
timestamp 1666464484
transform 1 0 25300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_269
timestamp 1666464484
transform 1 0 25852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_275
timestamp 1666464484
transform 1 0 26404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_283
timestamp 1666464484
transform 1 0 27140 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_293
timestamp 1666464484
transform 1 0 28060 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_299
timestamp 1666464484
transform 1 0 28612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_305
timestamp 1666464484
transform 1 0 29164 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_313
timestamp 1666464484
transform 1 0 29900 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_318
timestamp 1666464484
transform 1 0 30360 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_324
timestamp 1666464484
transform 1 0 30912 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_336
timestamp 1666464484
transform 1 0 32016 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_348
timestamp 1666464484
transform 1 0 33120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1666464484
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1666464484
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1666464484
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1666464484
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1666464484
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1666464484
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1666464484
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1666464484
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1666464484
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1666464484
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1666464484
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1666464484
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1666464484
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1666464484
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1666464484
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1666464484
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1666464484
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1666464484
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1666464484
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1666464484
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1666464484
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1666464484
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_9
timestamp 1666464484
transform 1 0 1932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_21
timestamp 1666464484
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_33
timestamp 1666464484
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_45
timestamp 1666464484
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1666464484
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1666464484
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1666464484
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_148
timestamp 1666464484
transform 1 0 14720 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1666464484
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_177
timestamp 1666464484
transform 1 0 17388 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_183
timestamp 1666464484
transform 1 0 17940 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_194
timestamp 1666464484
transform 1 0 18952 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1666464484
transform 1 0 19596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 1666464484
transform 1 0 20240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_214
timestamp 1666464484
transform 1 0 20792 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1666464484
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_233
timestamp 1666464484
transform 1 0 22540 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_239
timestamp 1666464484
transform 1 0 23092 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_246
timestamp 1666464484
transform 1 0 23736 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_254
timestamp 1666464484
transform 1 0 24472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_264
timestamp 1666464484
transform 1 0 25392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_270
timestamp 1666464484
transform 1 0 25944 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1666464484
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_289
timestamp 1666464484
transform 1 0 27692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_295
timestamp 1666464484
transform 1 0 28244 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_301
timestamp 1666464484
transform 1 0 28796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_305
timestamp 1666464484
transform 1 0 29164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_308
timestamp 1666464484
transform 1 0 29440 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_314
timestamp 1666464484
transform 1 0 29992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_320
timestamp 1666464484
transform 1 0 30544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_326
timestamp 1666464484
transform 1 0 31096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1666464484
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_341
timestamp 1666464484
transform 1 0 32476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_353
timestamp 1666464484
transform 1 0 33580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_365
timestamp 1666464484
transform 1 0 34684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_377
timestamp 1666464484
transform 1 0 35788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_389
timestamp 1666464484
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1666464484
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1666464484
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1666464484
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1666464484
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1666464484
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1666464484
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1666464484
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1666464484
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1666464484
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1666464484
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1666464484
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666464484
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1666464484
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1666464484
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1666464484
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1666464484
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1666464484
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1666464484
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1666464484
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_573
timestamp 1666464484
transform 1 0 53820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_579
timestamp 1666464484
transform 1 0 54372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_9
timestamp 1666464484
transform 1 0 1932 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1666464484
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_129
timestamp 1666464484
transform 1 0 12972 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1666464484
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1666464484
transform 1 0 14720 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_154
timestamp 1666464484
transform 1 0 15272 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_166
timestamp 1666464484
transform 1 0 16376 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_172
timestamp 1666464484
transform 1 0 16928 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_179
timestamp 1666464484
transform 1 0 17572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_187
timestamp 1666464484
transform 1 0 18308 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1666464484
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_215
timestamp 1666464484
transform 1 0 20884 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_224
timestamp 1666464484
transform 1 0 21712 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1666464484
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1666464484
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_264
timestamp 1666464484
transform 1 0 25392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_271
timestamp 1666464484
transform 1 0 26036 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_283
timestamp 1666464484
transform 1 0 27140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_291
timestamp 1666464484
transform 1 0 27876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_297
timestamp 1666464484
transform 1 0 28428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_300
timestamp 1666464484
transform 1 0 28704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1666464484
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_313
timestamp 1666464484
transform 1 0 29900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_319
timestamp 1666464484
transform 1 0 30452 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_325
timestamp 1666464484
transform 1 0 31004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_331
timestamp 1666464484
transform 1 0 31556 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_337
timestamp 1666464484
transform 1 0 32108 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_343
timestamp 1666464484
transform 1 0 32660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_349
timestamp 1666464484
transform 1 0 33212 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1666464484
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666464484
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1666464484
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1666464484
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1666464484
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1666464484
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1666464484
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1666464484
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1666464484
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1666464484
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1666464484
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1666464484
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1666464484
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1666464484
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1666464484
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1666464484
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1666464484
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1666464484
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1666464484
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1666464484
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1666464484
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1666464484
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1666464484
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_571
timestamp 1666464484
transform 1 0 53636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_579
timestamp 1666464484
transform 1 0 54372 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1666464484
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1666464484
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1666464484
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1666464484
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1666464484
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1666464484
transform 1 0 13248 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_138
timestamp 1666464484
transform 1 0 13800 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_150
timestamp 1666464484
transform 1 0 14904 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_160
timestamp 1666464484
transform 1 0 15824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1666464484
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1666464484
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_202
timestamp 1666464484
transform 1 0 19688 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1666464484
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_236
timestamp 1666464484
transform 1 0 22816 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_244
timestamp 1666464484
transform 1 0 23552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_261
timestamp 1666464484
transform 1 0 25116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_267
timestamp 1666464484
transform 1 0 25668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1666464484
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1666464484
transform 1 0 27416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_290
timestamp 1666464484
transform 1 0 27784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_294
timestamp 1666464484
transform 1 0 28152 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_301
timestamp 1666464484
transform 1 0 28796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_314
timestamp 1666464484
transform 1 0 29992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_321
timestamp 1666464484
transform 1 0 30636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_327
timestamp 1666464484
transform 1 0 31188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1666464484
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_341
timestamp 1666464484
transform 1 0 32476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_347
timestamp 1666464484
transform 1 0 33028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_353
timestamp 1666464484
transform 1 0 33580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_359
timestamp 1666464484
transform 1 0 34132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_365
timestamp 1666464484
transform 1 0 34684 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_371
timestamp 1666464484
transform 1 0 35236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_383
timestamp 1666464484
transform 1 0 36340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1666464484
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1666464484
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1666464484
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1666464484
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1666464484
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1666464484
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1666464484
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1666464484
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1666464484
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1666464484
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1666464484
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1666464484
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1666464484
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1666464484
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1666464484
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1666464484
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1666464484
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_553
timestamp 1666464484
transform 1 0 51980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_558
timestamp 1666464484
transform 1 0 52440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_561
timestamp 1666464484
transform 1 0 52716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_565
timestamp 1666464484
transform 1 0 53084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_569
timestamp 1666464484
transform 1 0 53452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_579
timestamp 1666464484
transform 1 0 54372 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_9
timestamp 1666464484
transform 1 0 1932 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1666464484
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_130
timestamp 1666464484
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1666464484
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1666464484
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1666464484
transform 1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1666464484
transform 1 0 15272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_160
timestamp 1666464484
transform 1 0 15824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_168
timestamp 1666464484
transform 1 0 16560 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_171
timestamp 1666464484
transform 1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1666464484
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1666464484
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_203
timestamp 1666464484
transform 1 0 19780 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_220
timestamp 1666464484
transform 1 0 21344 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_226
timestamp 1666464484
transform 1 0 21896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1666464484
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1666464484
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_257
timestamp 1666464484
transform 1 0 24748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_270
timestamp 1666464484
transform 1 0 25944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_276
timestamp 1666464484
transform 1 0 26496 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_289
timestamp 1666464484
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_293
timestamp 1666464484
transform 1 0 28060 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_297
timestamp 1666464484
transform 1 0 28428 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1666464484
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_327
timestamp 1666464484
transform 1 0 31188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_333
timestamp 1666464484
transform 1 0 31740 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_339
timestamp 1666464484
transform 1 0 32292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_345
timestamp 1666464484
transform 1 0 32844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_349
timestamp 1666464484
transform 1 0 33212 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_355
timestamp 1666464484
transform 1 0 33764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp 1666464484
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1666464484
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_369
timestamp 1666464484
transform 1 0 35052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_375
timestamp 1666464484
transform 1 0 35604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_381
timestamp 1666464484
transform 1 0 36156 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_387
timestamp 1666464484
transform 1 0 36708 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_399
timestamp 1666464484
transform 1 0 37812 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_411
timestamp 1666464484
transform 1 0 38916 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1666464484
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1666464484
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1666464484
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1666464484
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1666464484
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1666464484
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1666464484
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1666464484
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1666464484
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1666464484
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1666464484
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1666464484
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1666464484
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1666464484
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_545
timestamp 1666464484
transform 1 0 51244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_549
timestamp 1666464484
transform 1 0 51612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_552
timestamp 1666464484
transform 1 0 51888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_559
timestamp 1666464484
transform 1 0 52532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_579
timestamp 1666464484
transform 1 0 54372 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_9
timestamp 1666464484
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_21
timestamp 1666464484
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_33
timestamp 1666464484
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_45
timestamp 1666464484
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1666464484
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_140
timestamp 1666464484
transform 1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_150
timestamp 1666464484
transform 1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_160
timestamp 1666464484
transform 1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1666464484
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_177
timestamp 1666464484
transform 1 0 17388 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_185
timestamp 1666464484
transform 1 0 18124 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 1666464484
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1666464484
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_236
timestamp 1666464484
transform 1 0 22816 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_240
timestamp 1666464484
transform 1 0 23184 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_257
timestamp 1666464484
transform 1 0 24748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_264
timestamp 1666464484
transform 1 0 25392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1666464484
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_299
timestamp 1666464484
transform 1 0 28612 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_323
timestamp 1666464484
transform 1 0 30820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1666464484
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_342
timestamp 1666464484
transform 1 0 32568 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_350
timestamp 1666464484
transform 1 0 33304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_367
timestamp 1666464484
transform 1 0 34868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_374
timestamp 1666464484
transform 1 0 35512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_380
timestamp 1666464484
transform 1 0 36064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_386
timestamp 1666464484
transform 1 0 36616 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1666464484
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_397
timestamp 1666464484
transform 1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1666464484
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_409
timestamp 1666464484
transform 1 0 38732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_421
timestamp 1666464484
transform 1 0 39836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_433
timestamp 1666464484
transform 1 0 40940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_445
timestamp 1666464484
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1666464484
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1666464484
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1666464484
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1666464484
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1666464484
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1666464484
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1666464484
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1666464484
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1666464484
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_541
timestamp 1666464484
transform 1 0 50876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_545
timestamp 1666464484
transform 1 0 51244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_551
timestamp 1666464484
transform 1 0 51796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_558
timestamp 1666464484
transform 1 0 52440 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_561
timestamp 1666464484
transform 1 0 52716 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_571
timestamp 1666464484
transform 1 0 53636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_579
timestamp 1666464484
transform 1 0 54372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_9
timestamp 1666464484
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1666464484
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_129
timestamp 1666464484
transform 1 0 12972 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1666464484
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_150
timestamp 1666464484
transform 1 0 14904 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 1666464484
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1666464484
transform 1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_175
timestamp 1666464484
transform 1 0 17204 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_183
timestamp 1666464484
transform 1 0 17940 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_187
timestamp 1666464484
transform 1 0 18308 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1666464484
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_208
timestamp 1666464484
transform 1 0 20240 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_225
timestamp 1666464484
transform 1 0 21804 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_234
timestamp 1666464484
transform 1 0 22632 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_241
timestamp 1666464484
transform 1 0 23276 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1666464484
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_264
timestamp 1666464484
transform 1 0 25392 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_270
timestamp 1666464484
transform 1 0 25944 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_288
timestamp 1666464484
transform 1 0 27600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1666464484
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1666464484
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_327
timestamp 1666464484
transform 1 0 31188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_331
timestamp 1666464484
transform 1 0 31556 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_341
timestamp 1666464484
transform 1 0 32476 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_348
timestamp 1666464484
transform 1 0 33120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_352
timestamp 1666464484
transform 1 0 33488 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1666464484
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1666464484
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_376
timestamp 1666464484
transform 1 0 35696 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_383
timestamp 1666464484
transform 1 0 36340 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_389
timestamp 1666464484
transform 1 0 36892 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_395
timestamp 1666464484
transform 1 0 37444 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_401
timestamp 1666464484
transform 1 0 37996 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_414
timestamp 1666464484
transform 1 0 39192 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1666464484
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1666464484
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1666464484
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1666464484
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1666464484
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1666464484
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1666464484
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1666464484
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1666464484
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_513
timestamp 1666464484
transform 1 0 48300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_517
timestamp 1666464484
transform 1 0 48668 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_521
timestamp 1666464484
transform 1 0 49036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_527
timestamp 1666464484
transform 1 0 49588 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1666464484
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_533
timestamp 1666464484
transform 1 0 50140 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_538
timestamp 1666464484
transform 1 0 50600 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_546
timestamp 1666464484
transform 1 0 51336 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_552
timestamp 1666464484
transform 1 0 51888 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_560
timestamp 1666464484
transform 1 0 52624 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_564
timestamp 1666464484
transform 1 0 52992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_574
timestamp 1666464484
transform 1 0 53912 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_580
timestamp 1666464484
transform 1 0 54464 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_9
timestamp 1666464484
transform 1 0 1932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_21
timestamp 1666464484
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_33
timestamp 1666464484
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1666464484
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1666464484
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1666464484
transform 1 0 12972 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_136
timestamp 1666464484
transform 1 0 13616 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_147
timestamp 1666464484
transform 1 0 14628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_158
timestamp 1666464484
transform 1 0 15640 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1666464484
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_177
timestamp 1666464484
transform 1 0 17388 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_185
timestamp 1666464484
transform 1 0 18124 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1666464484
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_206
timestamp 1666464484
transform 1 0 20056 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1666464484
transform 1 0 20884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1666464484
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_232
timestamp 1666464484
transform 1 0 22448 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_245
timestamp 1666464484
transform 1 0 23644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_262
timestamp 1666464484
transform 1 0 25208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_266
timestamp 1666464484
transform 1 0 25576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1666464484
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_292
timestamp 1666464484
transform 1 0 27968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_296
timestamp 1666464484
transform 1 0 28336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_303
timestamp 1666464484
transform 1 0 28980 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_316
timestamp 1666464484
transform 1 0 30176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_324
timestamp 1666464484
transform 1 0 30912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_328
timestamp 1666464484
transform 1 0 31280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1666464484
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_355
timestamp 1666464484
transform 1 0 33764 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_363
timestamp 1666464484
transform 1 0 34500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_380
timestamp 1666464484
transform 1 0 36064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_387
timestamp 1666464484
transform 1 0 36708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1666464484
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1666464484
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_397
timestamp 1666464484
transform 1 0 37628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_417
timestamp 1666464484
transform 1 0 39468 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_423
timestamp 1666464484
transform 1 0 40020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_435
timestamp 1666464484
transform 1 0 41124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1666464484
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1666464484
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1666464484
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1666464484
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1666464484
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1666464484
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1666464484
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_505
timestamp 1666464484
transform 1 0 47564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_511
timestamp 1666464484
transform 1 0 48116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_514
timestamp 1666464484
transform 1 0 48392 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_534
timestamp 1666464484
transform 1 0 50232 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_543
timestamp 1666464484
transform 1 0 51060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_555
timestamp 1666464484
transform 1 0 52164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_558
timestamp 1666464484
transform 1 0 52440 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_561
timestamp 1666464484
transform 1 0 52716 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_571
timestamp 1666464484
transform 1 0 53636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_579
timestamp 1666464484
transform 1 0 54372 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_9
timestamp 1666464484
transform 1 0 1932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1666464484
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_129
timestamp 1666464484
transform 1 0 12972 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1666464484
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_147
timestamp 1666464484
transform 1 0 14628 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_158
timestamp 1666464484
transform 1 0 15640 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_164
timestamp 1666464484
transform 1 0 16192 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_174
timestamp 1666464484
transform 1 0 17112 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1666464484
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1666464484
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_208
timestamp 1666464484
transform 1 0 20240 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1666464484
transform 1 0 20884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_225
timestamp 1666464484
transform 1 0 21804 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666464484
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666464484
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_264
timestamp 1666464484
transform 1 0 25392 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_270
timestamp 1666464484
transform 1 0 25944 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_291
timestamp 1666464484
transform 1 0 27876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_298
timestamp 1666464484
transform 1 0 28520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_302
timestamp 1666464484
transform 1 0 28888 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1666464484
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_315
timestamp 1666464484
transform 1 0 30084 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_323
timestamp 1666464484
transform 1 0 30820 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_330
timestamp 1666464484
transform 1 0 31464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_339
timestamp 1666464484
transform 1 0 32292 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_349
timestamp 1666464484
transform 1 0 33212 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1666464484
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1666464484
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_372
timestamp 1666464484
transform 1 0 35328 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_379
timestamp 1666464484
transform 1 0 35972 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_401
timestamp 1666464484
transform 1 0 37996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_411
timestamp 1666464484
transform 1 0 38916 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_417
timestamp 1666464484
transform 1 0 39468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1666464484
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_428
timestamp 1666464484
transform 1 0 40480 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_440
timestamp 1666464484
transform 1 0 41584 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_452
timestamp 1666464484
transform 1 0 42688 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_464
timestamp 1666464484
transform 1 0 43792 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1666464484
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1666464484
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1666464484
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1666464484
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1666464484
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1666464484
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1666464484
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1666464484
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_557
timestamp 1666464484
transform 1 0 52348 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_565
timestamp 1666464484
transform 1 0 53084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_571
timestamp 1666464484
transform 1 0 53636 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_579
timestamp 1666464484
transform 1 0 54372 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_9
timestamp 1666464484
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1666464484
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1666464484
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1666464484
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1666464484
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_133
timestamp 1666464484
transform 1 0 13340 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_136
timestamp 1666464484
transform 1 0 13616 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_146
timestamp 1666464484
transform 1 0 14536 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_157
timestamp 1666464484
transform 1 0 15548 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1666464484
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_177
timestamp 1666464484
transform 1 0 17388 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_201
timestamp 1666464484
transform 1 0 19596 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_208
timestamp 1666464484
transform 1 0 20240 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1666464484
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_229
timestamp 1666464484
transform 1 0 22172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_238
timestamp 1666464484
transform 1 0 23000 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_262
timestamp 1666464484
transform 1 0 25208 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_268
timestamp 1666464484
transform 1 0 25760 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1666464484
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_288
timestamp 1666464484
transform 1 0 27600 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_297
timestamp 1666464484
transform 1 0 28428 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_306
timestamp 1666464484
transform 1 0 29256 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_317
timestamp 1666464484
transform 1 0 30268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1666464484
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666464484
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_341
timestamp 1666464484
transform 1 0 32476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_348
timestamp 1666464484
transform 1 0 33120 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_356
timestamp 1666464484
transform 1 0 33856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_373
timestamp 1666464484
transform 1 0 35420 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1666464484
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1666464484
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_399
timestamp 1666464484
transform 1 0 37812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_419
timestamp 1666464484
transform 1 0 39652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_429
timestamp 1666464484
transform 1 0 40572 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_439
timestamp 1666464484
transform 1 0 41492 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_445
timestamp 1666464484
transform 1 0 42044 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1666464484
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1666464484
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1666464484
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1666464484
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1666464484
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666464484
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1666464484
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1666464484
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1666464484
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1666464484
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1666464484
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1666464484
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_561
timestamp 1666464484
transform 1 0 52716 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_571
timestamp 1666464484
transform 1 0 53636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_579
timestamp 1666464484
transform 1 0 54372 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_9
timestamp 1666464484
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1666464484
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_129
timestamp 1666464484
transform 1 0 12972 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_132
timestamp 1666464484
transform 1 0 13248 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1666464484
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1666464484
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1666464484
transform 1 0 15272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_164
timestamp 1666464484
transform 1 0 16192 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_174
timestamp 1666464484
transform 1 0 17112 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1666464484
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_201
timestamp 1666464484
transform 1 0 19596 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_229
timestamp 1666464484
transform 1 0 22172 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1666464484
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_259
timestamp 1666464484
transform 1 0 24932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_268
timestamp 1666464484
transform 1 0 25760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_277
timestamp 1666464484
transform 1 0 26588 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_283
timestamp 1666464484
transform 1 0 27140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_293
timestamp 1666464484
transform 1 0 28060 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_299
timestamp 1666464484
transform 1 0 28612 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1666464484
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_316
timestamp 1666464484
transform 1 0 30176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_328
timestamp 1666464484
transform 1 0 31280 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_340
timestamp 1666464484
transform 1 0 32384 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_355
timestamp 1666464484
transform 1 0 33764 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1666464484
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1666464484
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_375
timestamp 1666464484
transform 1 0 35604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_387
timestamp 1666464484
transform 1 0 36708 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_399
timestamp 1666464484
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_409
timestamp 1666464484
transform 1 0 38732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_416
timestamp 1666464484
transform 1 0 39376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1666464484
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_429
timestamp 1666464484
transform 1 0 40572 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_435
timestamp 1666464484
transform 1 0 41124 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_447
timestamp 1666464484
transform 1 0 42228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_459
timestamp 1666464484
transform 1 0 43332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_471
timestamp 1666464484
transform 1 0 44436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1666464484
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1666464484
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1666464484
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1666464484
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1666464484
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1666464484
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1666464484
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1666464484
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1666464484
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1666464484
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_571
timestamp 1666464484
transform 1 0 53636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_579
timestamp 1666464484
transform 1 0 54372 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_9
timestamp 1666464484
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_21
timestamp 1666464484
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_33
timestamp 1666464484
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_45
timestamp 1666464484
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1666464484
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_121
timestamp 1666464484
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_126
timestamp 1666464484
transform 1 0 12696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1666464484
transform 1 0 13248 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_138
timestamp 1666464484
transform 1 0 13800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1666464484
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_155
timestamp 1666464484
transform 1 0 15364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1666464484
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_175
timestamp 1666464484
transform 1 0 17204 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_198
timestamp 1666464484
transform 1 0 19320 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1666464484
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_229
timestamp 1666464484
transform 1 0 22172 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_239
timestamp 1666464484
transform 1 0 23092 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_247
timestamp 1666464484
transform 1 0 23828 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_253
timestamp 1666464484
transform 1 0 24380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_299
timestamp 1666464484
transform 1 0 28612 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1666464484
transform 1 0 29256 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_319
timestamp 1666464484
transform 1 0 30452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_331
timestamp 1666464484
transform 1 0 31556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1666464484
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_341
timestamp 1666464484
transform 1 0 32476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_361
timestamp 1666464484
transform 1 0 34316 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_365
timestamp 1666464484
transform 1 0 34684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_369
timestamp 1666464484
transform 1 0 35052 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_389
timestamp 1666464484
transform 1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1666464484
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_400
timestamp 1666464484
transform 1 0 37904 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_422
timestamp 1666464484
transform 1 0 39928 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_431
timestamp 1666464484
transform 1 0 40756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_437
timestamp 1666464484
transform 1 0 41308 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1666464484
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1666464484
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1666464484
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1666464484
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1666464484
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1666464484
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1666464484
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1666464484
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1666464484
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1666464484
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1666464484
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1666464484
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1666464484
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1666464484
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_561
timestamp 1666464484
transform 1 0 52716 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_571
timestamp 1666464484
transform 1 0 53636 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_579
timestamp 1666464484
transform 1 0 54372 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_9
timestamp 1666464484
transform 1 0 1932 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1666464484
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_117
timestamp 1666464484
transform 1 0 11868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_120
timestamp 1666464484
transform 1 0 12144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1666464484
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_132
timestamp 1666464484
transform 1 0 13248 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1666464484
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_147
timestamp 1666464484
transform 1 0 14628 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_156
timestamp 1666464484
transform 1 0 15456 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_167
timestamp 1666464484
transform 1 0 16468 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_177
timestamp 1666464484
transform 1 0 17388 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1666464484
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_203
timestamp 1666464484
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_207
timestamp 1666464484
transform 1 0 20148 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_220
timestamp 1666464484
transform 1 0 21344 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_237
timestamp 1666464484
transform 1 0 22908 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1666464484
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_271
timestamp 1666464484
transform 1 0 26036 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_280
timestamp 1666464484
transform 1 0 26864 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_292
timestamp 1666464484
transform 1 0 27968 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_300
timestamp 1666464484
transform 1 0 28704 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1666464484
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_327
timestamp 1666464484
transform 1 0 31188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_333
timestamp 1666464484
transform 1 0 31740 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_345
timestamp 1666464484
transform 1 0 32844 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_353
timestamp 1666464484
transform 1 0 33580 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1666464484
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1666464484
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_373
timestamp 1666464484
transform 1 0 35420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_389
timestamp 1666464484
transform 1 0 36892 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_399
timestamp 1666464484
transform 1 0 37812 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_403
timestamp 1666464484
transform 1 0 38180 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_410
timestamp 1666464484
transform 1 0 38824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_417
timestamp 1666464484
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1666464484
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_425
timestamp 1666464484
transform 1 0 40204 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_431
timestamp 1666464484
transform 1 0 40756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_437
timestamp 1666464484
transform 1 0 41308 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_443
timestamp 1666464484
transform 1 0 41860 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_455
timestamp 1666464484
transform 1 0 42964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_467
timestamp 1666464484
transform 1 0 44068 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1666464484
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1666464484
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1666464484
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1666464484
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1666464484
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1666464484
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1666464484
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1666464484
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1666464484
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_557
timestamp 1666464484
transform 1 0 52348 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_563
timestamp 1666464484
transform 1 0 52900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_571
timestamp 1666464484
transform 1 0 53636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_579
timestamp 1666464484
transform 1 0 54372 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1666464484
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_21
timestamp 1666464484
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_33
timestamp 1666464484
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1666464484
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1666464484
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1666464484
transform 1 0 11960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_124
timestamp 1666464484
transform 1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1666464484
transform 1 0 13064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1666464484
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1666464484
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_155
timestamp 1666464484
transform 1 0 15364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_174
timestamp 1666464484
transform 1 0 17112 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_182
timestamp 1666464484
transform 1 0 17848 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_202
timestamp 1666464484
transform 1 0 19688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1666464484
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_233
timestamp 1666464484
transform 1 0 22540 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_239
timestamp 1666464484
transform 1 0 23092 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_251
timestamp 1666464484
transform 1 0 24196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_264
timestamp 1666464484
transform 1 0 25392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1666464484
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_293
timestamp 1666464484
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_304
timestamp 1666464484
transform 1 0 29072 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_318
timestamp 1666464484
transform 1 0 30360 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1666464484
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1666464484
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_346
timestamp 1666464484
transform 1 0 32936 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_352
timestamp 1666464484
transform 1 0 33488 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_361
timestamp 1666464484
transform 1 0 34316 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_373
timestamp 1666464484
transform 1 0 35420 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_386
timestamp 1666464484
transform 1 0 36616 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1666464484
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_400
timestamp 1666464484
transform 1 0 37904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_420
timestamp 1666464484
transform 1 0 39744 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_427
timestamp 1666464484
transform 1 0 40388 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_433
timestamp 1666464484
transform 1 0 40940 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_439
timestamp 1666464484
transform 1 0 41492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_445
timestamp 1666464484
transform 1 0 42044 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1666464484
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1666464484
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1666464484
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1666464484
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1666464484
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1666464484
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1666464484
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1666464484
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1666464484
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1666464484
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1666464484
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1666464484
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1666464484
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_573
timestamp 1666464484
transform 1 0 53820 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_579
timestamp 1666464484
transform 1 0 54372 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_9
timestamp 1666464484
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1666464484
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1666464484
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_132
timestamp 1666464484
transform 1 0 13248 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1666464484
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_150
timestamp 1666464484
transform 1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_158
timestamp 1666464484
transform 1 0 15640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_169
timestamp 1666464484
transform 1 0 16652 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_177
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1666464484
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_202
timestamp 1666464484
transform 1 0 19688 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1666464484
transform 1 0 20424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_234
timestamp 1666464484
transform 1 0 22632 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1666464484
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_260
timestamp 1666464484
transform 1 0 25024 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_272
timestamp 1666464484
transform 1 0 26128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_278
timestamp 1666464484
transform 1 0 26680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_287
timestamp 1666464484
transform 1 0 27508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_299
timestamp 1666464484
transform 1 0 28612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1666464484
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_318
timestamp 1666464484
transform 1 0 30360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_328
timestamp 1666464484
transform 1 0 31280 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_340
timestamp 1666464484
transform 1 0 32384 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_354
timestamp 1666464484
transform 1 0 33672 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1666464484
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1666464484
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_383
timestamp 1666464484
transform 1 0 36340 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_399
timestamp 1666464484
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_407
timestamp 1666464484
transform 1 0 38548 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_411
timestamp 1666464484
transform 1 0 38916 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_417
timestamp 1666464484
transform 1 0 39468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1666464484
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_427
timestamp 1666464484
transform 1 0 40388 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_434
timestamp 1666464484
transform 1 0 41032 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_440
timestamp 1666464484
transform 1 0 41584 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_446
timestamp 1666464484
transform 1 0 42136 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_452
timestamp 1666464484
transform 1 0 42688 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_464
timestamp 1666464484
transform 1 0 43792 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1666464484
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1666464484
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1666464484
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1666464484
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1666464484
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1666464484
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1666464484
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1666464484
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1666464484
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_571
timestamp 1666464484
transform 1 0 53636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_579
timestamp 1666464484
transform 1 0 54372 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_9
timestamp 1666464484
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1666464484
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1666464484
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1666464484
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1666464484
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1666464484
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_122
timestamp 1666464484
transform 1 0 12328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_128
timestamp 1666464484
transform 1 0 12880 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1666464484
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1666464484
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_146
timestamp 1666464484
transform 1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_155
timestamp 1666464484
transform 1 0 15364 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1666464484
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_178
timestamp 1666464484
transform 1 0 17480 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_186
timestamp 1666464484
transform 1 0 18216 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1666464484
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_209
timestamp 1666464484
transform 1 0 20332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1666464484
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_231
timestamp 1666464484
transform 1 0 22356 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1666464484
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1666464484
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_258
timestamp 1666464484
transform 1 0 24840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1666464484
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_299
timestamp 1666464484
transform 1 0 28612 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_315
timestamp 1666464484
transform 1 0 30084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_321
timestamp 1666464484
transform 1 0 30636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1666464484
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_347
timestamp 1666464484
transform 1 0 33028 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_355
timestamp 1666464484
transform 1 0 33764 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_375
timestamp 1666464484
transform 1 0 35604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_387
timestamp 1666464484
transform 1 0 36708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1666464484
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1666464484
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_411
timestamp 1666464484
transform 1 0 38916 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_419
timestamp 1666464484
transform 1 0 39652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_427
timestamp 1666464484
transform 1 0 40388 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_435
timestamp 1666464484
transform 1 0 41124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1666464484
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1666464484
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_449
timestamp 1666464484
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_453
timestamp 1666464484
transform 1 0 42780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_459
timestamp 1666464484
transform 1 0 43332 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_465
timestamp 1666464484
transform 1 0 43884 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_477
timestamp 1666464484
transform 1 0 44988 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_489
timestamp 1666464484
transform 1 0 46092 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_501
timestamp 1666464484
transform 1 0 47196 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1666464484
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1666464484
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1666464484
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1666464484
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1666464484
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1666464484
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_561
timestamp 1666464484
transform 1 0 52716 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_571
timestamp 1666464484
transform 1 0 53636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_579
timestamp 1666464484
transform 1 0 54372 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_9
timestamp 1666464484
transform 1 0 1932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1666464484
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_126
timestamp 1666464484
transform 1 0 12696 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_132
timestamp 1666464484
transform 1 0 13248 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1666464484
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_147
timestamp 1666464484
transform 1 0 14628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1666464484
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1666464484
transform 1 0 17204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1666464484
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1666464484
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1666464484
transform 1 0 20884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_228
timestamp 1666464484
transform 1 0 22080 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_232
timestamp 1666464484
transform 1 0 22448 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1666464484
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_258
timestamp 1666464484
transform 1 0 24840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_278
timestamp 1666464484
transform 1 0 26680 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_286
timestamp 1666464484
transform 1 0 27416 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_294
timestamp 1666464484
transform 1 0 28152 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1666464484
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_328
timestamp 1666464484
transform 1 0 31280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_339
timestamp 1666464484
transform 1 0 32292 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_350
timestamp 1666464484
transform 1 0 33304 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1666464484
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1666464484
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_383
timestamp 1666464484
transform 1 0 36340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_397
timestamp 1666464484
transform 1 0 37628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_406
timestamp 1666464484
transform 1 0 38456 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_412
timestamp 1666464484
transform 1 0 39008 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1666464484
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1666464484
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_439
timestamp 1666464484
transform 1 0 41492 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_445
timestamp 1666464484
transform 1 0 42044 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_451
timestamp 1666464484
transform 1 0 42596 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_457
timestamp 1666464484
transform 1 0 43148 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_463
timestamp 1666464484
transform 1 0 43700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1666464484
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1666464484
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1666464484
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1666464484
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1666464484
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1666464484
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1666464484
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1666464484
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1666464484
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1666464484
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1666464484
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_571
timestamp 1666464484
transform 1 0 53636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_579
timestamp 1666464484
transform 1 0 54372 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_9
timestamp 1666464484
transform 1 0 1932 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_21
timestamp 1666464484
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_33
timestamp 1666464484
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1666464484
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1666464484
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_129
timestamp 1666464484
transform 1 0 12972 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1666464484
transform 1 0 13248 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1666464484
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_144
timestamp 1666464484
transform 1 0 14352 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_150
timestamp 1666464484
transform 1 0 14904 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_156
timestamp 1666464484
transform 1 0 15456 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1666464484
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_178
timestamp 1666464484
transform 1 0 17480 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_206
timestamp 1666464484
transform 1 0 20056 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1666464484
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_231
timestamp 1666464484
transform 1 0 22356 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_237
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_250
timestamp 1666464484
transform 1 0 24104 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_264
timestamp 1666464484
transform 1 0 25392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1666464484
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_290
timestamp 1666464484
transform 1 0 27784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_300
timestamp 1666464484
transform 1 0 28704 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_310
timestamp 1666464484
transform 1 0 29624 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_314
timestamp 1666464484
transform 1 0 29992 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_321
timestamp 1666464484
transform 1 0 30636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1666464484
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_355
timestamp 1666464484
transform 1 0 33764 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_367
timestamp 1666464484
transform 1 0 34868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_378
timestamp 1666464484
transform 1 0 35880 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_384
timestamp 1666464484
transform 1 0 36432 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1666464484
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1666464484
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_411
timestamp 1666464484
transform 1 0 38916 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_422
timestamp 1666464484
transform 1 0 39928 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_431
timestamp 1666464484
transform 1 0 40756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_440
timestamp 1666464484
transform 1 0 41584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1666464484
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_449
timestamp 1666464484
transform 1 0 42412 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_453
timestamp 1666464484
transform 1 0 42780 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_459
timestamp 1666464484
transform 1 0 43332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_465
timestamp 1666464484
transform 1 0 43884 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_471
timestamp 1666464484
transform 1 0 44436 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_477
timestamp 1666464484
transform 1 0 44988 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_489
timestamp 1666464484
transform 1 0 46092 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_501
timestamp 1666464484
transform 1 0 47196 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1666464484
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1666464484
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1666464484
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1666464484
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1666464484
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1666464484
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_561
timestamp 1666464484
transform 1 0 52716 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_571
timestamp 1666464484
transform 1 0 53636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_579
timestamp 1666464484
transform 1 0 54372 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_9
timestamp 1666464484
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1666464484
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1666464484
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_147
timestamp 1666464484
transform 1 0 14628 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1666464484
transform 1 0 15732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_166
timestamp 1666464484
transform 1 0 16376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1666464484
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1666464484
transform 1 0 20884 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1666464484
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1666464484
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1666464484
transform 1 0 26036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_283
timestamp 1666464484
transform 1 0 27140 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_289
timestamp 1666464484
transform 1 0 27692 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_299
timestamp 1666464484
transform 1 0 28612 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1666464484
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_316
timestamp 1666464484
transform 1 0 30176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_325
timestamp 1666464484
transform 1 0 31004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_345
timestamp 1666464484
transform 1 0 32844 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1666464484
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666464484
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1666464484
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_374
timestamp 1666464484
transform 1 0 35512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_380
timestamp 1666464484
transform 1 0 36064 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_404
timestamp 1666464484
transform 1 0 38272 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_410
timestamp 1666464484
transform 1 0 38824 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_418
timestamp 1666464484
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1666464484
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_439
timestamp 1666464484
transform 1 0 41492 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_446
timestamp 1666464484
transform 1 0 42136 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_453
timestamp 1666464484
transform 1 0 42780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_460
timestamp 1666464484
transform 1 0 43424 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_466
timestamp 1666464484
transform 1 0 43976 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_472
timestamp 1666464484
transform 1 0 44528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_477
timestamp 1666464484
transform 1 0 44988 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_481
timestamp 1666464484
transform 1 0 45356 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_493
timestamp 1666464484
transform 1 0 46460 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_505
timestamp 1666464484
transform 1 0 47564 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_517
timestamp 1666464484
transform 1 0 48668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_529
timestamp 1666464484
transform 1 0 49772 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1666464484
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1666464484
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_557
timestamp 1666464484
transform 1 0 52348 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_563
timestamp 1666464484
transform 1 0 52900 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_571
timestamp 1666464484
transform 1 0 53636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_579
timestamp 1666464484
transform 1 0 54372 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1666464484
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1666464484
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1666464484
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1666464484
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1666464484
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_147
timestamp 1666464484
transform 1 0 14628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1666464484
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1666464484
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1666464484
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_178
timestamp 1666464484
transform 1 0 17480 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1666464484
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_210
timestamp 1666464484
transform 1 0 20424 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1666464484
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_229
timestamp 1666464484
transform 1 0 22172 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_238
timestamp 1666464484
transform 1 0 23000 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_262
timestamp 1666464484
transform 1 0 25208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1666464484
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_290
timestamp 1666464484
transform 1 0 27784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_300
timestamp 1666464484
transform 1 0 28704 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_307
timestamp 1666464484
transform 1 0 29348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_318
timestamp 1666464484
transform 1 0 30360 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_324
timestamp 1666464484
transform 1 0 30912 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_330
timestamp 1666464484
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_342
timestamp 1666464484
transform 1 0 32568 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_351
timestamp 1666464484
transform 1 0 33396 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_355
timestamp 1666464484
transform 1 0 33764 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_362
timestamp 1666464484
transform 1 0 34408 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1666464484
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1666464484
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_398
timestamp 1666464484
transform 1 0 37720 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_408
timestamp 1666464484
transform 1 0 38640 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_432
timestamp 1666464484
transform 1 0 40848 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_440
timestamp 1666464484
transform 1 0 41584 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_446
timestamp 1666464484
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_449
timestamp 1666464484
transform 1 0 42412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_453
timestamp 1666464484
transform 1 0 42780 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_459
timestamp 1666464484
transform 1 0 43332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_465
timestamp 1666464484
transform 1 0 43884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_471
timestamp 1666464484
transform 1 0 44436 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_477
timestamp 1666464484
transform 1 0 44988 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_489
timestamp 1666464484
transform 1 0 46092 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_501
timestamp 1666464484
transform 1 0 47196 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1666464484
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1666464484
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1666464484
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1666464484
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1666464484
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1666464484
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1666464484
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_573
timestamp 1666464484
transform 1 0 53820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_579
timestamp 1666464484
transform 1 0 54372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_9
timestamp 1666464484
transform 1 0 1932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1666464484
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1666464484
transform 1 0 14812 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_159
timestamp 1666464484
transform 1 0 15732 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_171
timestamp 1666464484
transform 1 0 16836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_178
timestamp 1666464484
transform 1 0 17480 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1666464484
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1666464484
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1666464484
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_220
timestamp 1666464484
transform 1 0 21344 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_228
timestamp 1666464484
transform 1 0 22080 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_232
timestamp 1666464484
transform 1 0 22448 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1666464484
transform 1 0 23276 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1666464484
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_264
timestamp 1666464484
transform 1 0 25392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_276
timestamp 1666464484
transform 1 0 26496 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_287
timestamp 1666464484
transform 1 0 27508 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_293
timestamp 1666464484
transform 1 0 28060 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1666464484
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1666464484
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_314
timestamp 1666464484
transform 1 0 29992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_326
timestamp 1666464484
transform 1 0 31096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_342
timestamp 1666464484
transform 1 0 32568 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_346
timestamp 1666464484
transform 1 0 32936 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_353
timestamp 1666464484
transform 1 0 33580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_361
timestamp 1666464484
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1666464484
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_372
timestamp 1666464484
transform 1 0 35328 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_380
timestamp 1666464484
transform 1 0 36064 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_389
timestamp 1666464484
transform 1 0 36892 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_398
timestamp 1666464484
transform 1 0 37720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_406
timestamp 1666464484
transform 1 0 38456 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_417
timestamp 1666464484
transform 1 0 39468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1666464484
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_439
timestamp 1666464484
transform 1 0 41492 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_446
timestamp 1666464484
transform 1 0 42136 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_452
timestamp 1666464484
transform 1 0 42688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_458
timestamp 1666464484
transform 1 0 43240 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_464
timestamp 1666464484
transform 1 0 43792 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_470
timestamp 1666464484
transform 1 0 44344 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1666464484
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1666464484
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1666464484
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1666464484
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1666464484
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1666464484
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1666464484
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1666464484
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1666464484
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_571
timestamp 1666464484
transform 1 0 53636 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_579
timestamp 1666464484
transform 1 0 54372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_9
timestamp 1666464484
transform 1 0 1932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1666464484
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1666464484
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1666464484
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1666464484
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1666464484
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_177
timestamp 1666464484
transform 1 0 17388 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_183
timestamp 1666464484
transform 1 0 17940 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_207
timestamp 1666464484
transform 1 0 20148 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1666464484
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_231
timestamp 1666464484
transform 1 0 22356 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_251
timestamp 1666464484
transform 1 0 24196 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_258
timestamp 1666464484
transform 1 0 24840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1666464484
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_291
timestamp 1666464484
transform 1 0 27876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_295
timestamp 1666464484
transform 1 0 28244 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_312
timestamp 1666464484
transform 1 0 29808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1666464484
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_355
timestamp 1666464484
transform 1 0 33764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_361
timestamp 1666464484
transform 1 0 34316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_378
timestamp 1666464484
transform 1 0 35880 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_382
timestamp 1666464484
transform 1 0 36248 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1666464484
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1666464484
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_397
timestamp 1666464484
transform 1 0 37628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_406
timestamp 1666464484
transform 1 0 38456 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_426
timestamp 1666464484
transform 1 0 40296 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_435
timestamp 1666464484
transform 1 0 41124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_442
timestamp 1666464484
transform 1 0 41768 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1666464484
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_453
timestamp 1666464484
transform 1 0 42780 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_459
timestamp 1666464484
transform 1 0 43332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_465
timestamp 1666464484
transform 1 0 43884 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_471
timestamp 1666464484
transform 1 0 44436 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_483
timestamp 1666464484
transform 1 0 45540 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_495
timestamp 1666464484
transform 1 0 46644 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1666464484
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1666464484
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1666464484
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1666464484
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1666464484
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1666464484
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1666464484
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_561
timestamp 1666464484
transform 1 0 52716 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_571
timestamp 1666464484
transform 1 0 53636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_579
timestamp 1666464484
transform 1 0 54372 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_9
timestamp 1666464484
transform 1 0 1932 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1666464484
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_175
timestamp 1666464484
transform 1 0 17204 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 1666464484
transform 1 0 17756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_187
timestamp 1666464484
transform 1 0 18308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1666464484
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1666464484
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1666464484
transform 1 0 22080 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_235
timestamp 1666464484
transform 1 0 22724 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_244
timestamp 1666464484
transform 1 0 23552 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1666464484
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1666464484
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_276
timestamp 1666464484
transform 1 0 26496 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_284
timestamp 1666464484
transform 1 0 27232 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_292
timestamp 1666464484
transform 1 0 27968 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_296
timestamp 1666464484
transform 1 0 28336 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1666464484
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_320
timestamp 1666464484
transform 1 0 30544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_329
timestamp 1666464484
transform 1 0 31372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_333
timestamp 1666464484
transform 1 0 31740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_343
timestamp 1666464484
transform 1 0 32660 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1666464484
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1666464484
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_376
timestamp 1666464484
transform 1 0 35696 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_382
timestamp 1666464484
transform 1 0 36248 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_402
timestamp 1666464484
transform 1 0 38088 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_415
timestamp 1666464484
transform 1 0 39284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1666464484
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_421
timestamp 1666464484
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_427
timestamp 1666464484
transform 1 0 40388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_435
timestamp 1666464484
transform 1 0 41124 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_442
timestamp 1666464484
transform 1 0 41768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_448
timestamp 1666464484
transform 1 0 42320 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_454
timestamp 1666464484
transform 1 0 42872 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_460
timestamp 1666464484
transform 1 0 43424 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1666464484
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1666464484
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1666464484
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1666464484
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1666464484
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1666464484
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1666464484
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1666464484
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1666464484
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1666464484
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_571
timestamp 1666464484
transform 1 0 53636 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_579
timestamp 1666464484
transform 1 0 54372 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_8
timestamp 1666464484
transform 1 0 1840 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_14
timestamp 1666464484
transform 1 0 2392 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_26
timestamp 1666464484
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_38
timestamp 1666464484
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1666464484
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_177
timestamp 1666464484
transform 1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_182
timestamp 1666464484
transform 1 0 17848 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_188
timestamp 1666464484
transform 1 0 18400 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_208
timestamp 1666464484
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1666464484
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_231
timestamp 1666464484
transform 1 0 22356 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_235
timestamp 1666464484
transform 1 0 22724 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_255
timestamp 1666464484
transform 1 0 24564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_275
timestamp 1666464484
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1666464484
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_287
timestamp 1666464484
transform 1 0 27508 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_298
timestamp 1666464484
transform 1 0 28520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_318
timestamp 1666464484
transform 1 0 30360 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_327
timestamp 1666464484
transform 1 0 31188 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1666464484
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_346
timestamp 1666464484
transform 1 0 32936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_350
timestamp 1666464484
transform 1 0 33304 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_358
timestamp 1666464484
transform 1 0 34040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_378
timestamp 1666464484
transform 1 0 35880 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1666464484
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1666464484
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_399
timestamp 1666464484
transform 1 0 37812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_408
timestamp 1666464484
transform 1 0 38640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_415
timestamp 1666464484
transform 1 0 39284 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_424
timestamp 1666464484
transform 1 0 40112 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_433
timestamp 1666464484
transform 1 0 40940 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_440
timestamp 1666464484
transform 1 0 41584 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1666464484
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1666464484
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_453
timestamp 1666464484
transform 1 0 42780 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_459
timestamp 1666464484
transform 1 0 43332 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_471
timestamp 1666464484
transform 1 0 44436 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_483
timestamp 1666464484
transform 1 0 45540 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_495
timestamp 1666464484
transform 1 0 46644 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1666464484
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1666464484
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1666464484
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1666464484
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1666464484
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1666464484
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1666464484
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_561
timestamp 1666464484
transform 1 0 52716 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_571
timestamp 1666464484
transform 1 0 53636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_579
timestamp 1666464484
transform 1 0 54372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_9
timestamp 1666464484
transform 1 0 1932 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_185
timestamp 1666464484
transform 1 0 18124 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_188
timestamp 1666464484
transform 1 0 18400 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1666464484
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_202
timestamp 1666464484
transform 1 0 19688 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1666464484
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_233
timestamp 1666464484
transform 1 0 22540 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_239
timestamp 1666464484
transform 1 0 23092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_259
timestamp 1666464484
transform 1 0 24932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1666464484
transform 1 0 26036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_282
timestamp 1666464484
transform 1 0 27048 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_286
timestamp 1666464484
transform 1 0 27416 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_290
timestamp 1666464484
transform 1 0 27784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_302
timestamp 1666464484
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_319
timestamp 1666464484
transform 1 0 30452 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_325
timestamp 1666464484
transform 1 0 31004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_345
timestamp 1666464484
transform 1 0 32844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_356
timestamp 1666464484
transform 1 0 33856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1666464484
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1666464484
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_375
timestamp 1666464484
transform 1 0 35604 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_386
timestamp 1666464484
transform 1 0 36616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_398
timestamp 1666464484
transform 1 0 37720 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_405
timestamp 1666464484
transform 1 0 38364 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_416
timestamp 1666464484
transform 1 0 39376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1666464484
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_439
timestamp 1666464484
transform 1 0 41492 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_446
timestamp 1666464484
transform 1 0 42136 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_452
timestamp 1666464484
transform 1 0 42688 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_458
timestamp 1666464484
transform 1 0 43240 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_470
timestamp 1666464484
transform 1 0 44344 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1666464484
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1666464484
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1666464484
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1666464484
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1666464484
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1666464484
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1666464484
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1666464484
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_557
timestamp 1666464484
transform 1 0 52348 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_563
timestamp 1666464484
transform 1 0 52900 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_571
timestamp 1666464484
transform 1 0 53636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_579
timestamp 1666464484
transform 1 0 54372 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_9
timestamp 1666464484
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_21
timestamp 1666464484
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1666464484
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1666464484
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1666464484
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_187
timestamp 1666464484
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_207
timestamp 1666464484
transform 1 0 20148 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1666464484
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_243
timestamp 1666464484
transform 1 0 23460 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_247
timestamp 1666464484
transform 1 0 23828 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_253
timestamp 1666464484
transform 1 0 24380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_265
timestamp 1666464484
transform 1 0 25484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_269
timestamp 1666464484
transform 1 0 25852 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1666464484
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_292
timestamp 1666464484
transform 1 0 27968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_303
timestamp 1666464484
transform 1 0 28980 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_310
timestamp 1666464484
transform 1 0 29624 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_320
timestamp 1666464484
transform 1 0 30544 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1666464484
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_347
timestamp 1666464484
transform 1 0 33028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_356
timestamp 1666464484
transform 1 0 33856 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_360
timestamp 1666464484
transform 1 0 34224 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_377
timestamp 1666464484
transform 1 0 35788 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1666464484
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_393
timestamp 1666464484
transform 1 0 37260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_406
timestamp 1666464484
transform 1 0 38456 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_416
timestamp 1666464484
transform 1 0 39376 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_423
timestamp 1666464484
transform 1 0 40020 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_427
timestamp 1666464484
transform 1 0 40388 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_435
timestamp 1666464484
transform 1 0 41124 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_442
timestamp 1666464484
transform 1 0 41768 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_449
timestamp 1666464484
transform 1 0 42412 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_453
timestamp 1666464484
transform 1 0 42780 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_465
timestamp 1666464484
transform 1 0 43884 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_477
timestamp 1666464484
transform 1 0 44988 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_489
timestamp 1666464484
transform 1 0 46092 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_501
timestamp 1666464484
transform 1 0 47196 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1666464484
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1666464484
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1666464484
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1666464484
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1666464484
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1666464484
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_561
timestamp 1666464484
transform 1 0 52716 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_571
timestamp 1666464484
transform 1 0 53636 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_579
timestamp 1666464484
transform 1 0 54372 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1666464484
transform 1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_146
timestamp 1666464484
transform 1 0 14536 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_158
timestamp 1666464484
transform 1 0 15640 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_170
timestamp 1666464484
transform 1 0 16744 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_182
timestamp 1666464484
transform 1 0 17848 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_190
timestamp 1666464484
transform 1 0 18584 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1666464484
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_210
timestamp 1666464484
transform 1 0 20424 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_216
timestamp 1666464484
transform 1 0 20976 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_223
timestamp 1666464484
transform 1 0 21620 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_236
timestamp 1666464484
transform 1 0 22816 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_244
timestamp 1666464484
transform 1 0 23552 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1666464484
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_264
timestamp 1666464484
transform 1 0 25392 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_284
timestamp 1666464484
transform 1 0 27232 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_294
timestamp 1666464484
transform 1 0 28152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1666464484
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_319
timestamp 1666464484
transform 1 0 30452 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_339
timestamp 1666464484
transform 1 0 32292 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_359
timestamp 1666464484
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1666464484
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1666464484
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_383
timestamp 1666464484
transform 1 0 36340 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_390
timestamp 1666464484
transform 1 0 36984 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_394
timestamp 1666464484
transform 1 0 37352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_411
timestamp 1666464484
transform 1 0 38916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_418
timestamp 1666464484
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_421
timestamp 1666464484
transform 1 0 39836 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_441
timestamp 1666464484
transform 1 0 41676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_450
timestamp 1666464484
transform 1 0 42504 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_456
timestamp 1666464484
transform 1 0 43056 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_462
timestamp 1666464484
transform 1 0 43608 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_474
timestamp 1666464484
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1666464484
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1666464484
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1666464484
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1666464484
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1666464484
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1666464484
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1666464484
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1666464484
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1666464484
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_571
timestamp 1666464484
transform 1 0 53636 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_579
timestamp 1666464484
transform 1 0 54372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_9
timestamp 1666464484
transform 1 0 1932 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666464484
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_200
timestamp 1666464484
transform 1 0 19504 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_210
timestamp 1666464484
transform 1 0 20424 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_216
timestamp 1666464484
transform 1 0 20976 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1666464484
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_230
timestamp 1666464484
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1666464484
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_245
timestamp 1666464484
transform 1 0 23644 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_258
timestamp 1666464484
transform 1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1666464484
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_286
timestamp 1666464484
transform 1 0 27416 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_306
timestamp 1666464484
transform 1 0 29256 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_310
timestamp 1666464484
transform 1 0 29624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_318
timestamp 1666464484
transform 1 0 30360 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_322
timestamp 1666464484
transform 1 0 30728 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_331
timestamp 1666464484
transform 1 0 31556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1666464484
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_347
timestamp 1666464484
transform 1 0 33028 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_361
timestamp 1666464484
transform 1 0 34316 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_381
timestamp 1666464484
transform 1 0 36156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1666464484
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1666464484
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_403
timestamp 1666464484
transform 1 0 38180 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_411
timestamp 1666464484
transform 1 0 38916 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_432
timestamp 1666464484
transform 1 0 40848 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_443
timestamp 1666464484
transform 1 0 41860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1666464484
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_449
timestamp 1666464484
transform 1 0 42412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_453
timestamp 1666464484
transform 1 0 42780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_459
timestamp 1666464484
transform 1 0 43332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_465
timestamp 1666464484
transform 1 0 43884 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_471
timestamp 1666464484
transform 1 0 44436 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_483
timestamp 1666464484
transform 1 0 45540 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_495
timestamp 1666464484
transform 1 0 46644 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1666464484
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1666464484
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1666464484
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1666464484
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1666464484
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1666464484
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1666464484
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_561
timestamp 1666464484
transform 1 0 52716 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_571
timestamp 1666464484
transform 1 0 53636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_579
timestamp 1666464484
transform 1 0 54372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_9
timestamp 1666464484
transform 1 0 1932 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_205
timestamp 1666464484
transform 1 0 19964 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_211
timestamp 1666464484
transform 1 0 20516 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_217
timestamp 1666464484
transform 1 0 21068 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1666464484
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1666464484
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_240
timestamp 1666464484
transform 1 0 23184 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_246
timestamp 1666464484
transform 1 0 23736 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1666464484
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_271
timestamp 1666464484
transform 1 0 26036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_285
timestamp 1666464484
transform 1 0 27324 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_289
timestamp 1666464484
transform 1 0 27692 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_292
timestamp 1666464484
transform 1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1666464484
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_319
timestamp 1666464484
transform 1 0 30452 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_335
timestamp 1666464484
transform 1 0 31924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_347
timestamp 1666464484
transform 1 0 33028 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_353
timestamp 1666464484
transform 1 0 33580 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1666464484
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1666464484
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_376
timestamp 1666464484
transform 1 0 35696 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_404
timestamp 1666464484
transform 1 0 38272 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_410
timestamp 1666464484
transform 1 0 38824 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_418
timestamp 1666464484
transform 1 0 39560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1666464484
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_426
timestamp 1666464484
transform 1 0 40296 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_430
timestamp 1666464484
transform 1 0 40664 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_447
timestamp 1666464484
transform 1 0 42228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_454
timestamp 1666464484
transform 1 0 42872 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_461
timestamp 1666464484
transform 1 0 43516 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_467
timestamp 1666464484
transform 1 0 44068 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1666464484
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1666464484
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1666464484
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1666464484
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1666464484
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1666464484
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1666464484
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1666464484
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1666464484
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1666464484
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_571
timestamp 1666464484
transform 1 0 53636 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_579
timestamp 1666464484
transform 1 0 54372 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_9
timestamp 1666464484
transform 1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1666464484
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1666464484
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666464484
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_142
timestamp 1666464484
transform 1 0 14168 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_154
timestamp 1666464484
transform 1 0 15272 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1666464484
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_205
timestamp 1666464484
transform 1 0 19964 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_215
timestamp 1666464484
transform 1 0 20884 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1666464484
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_233
timestamp 1666464484
transform 1 0 22540 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_244
timestamp 1666464484
transform 1 0 23552 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_264
timestamp 1666464484
transform 1 0 25392 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1666464484
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1666464484
transform 1 0 27968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1666464484
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_317
timestamp 1666464484
transform 1 0 30268 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_331
timestamp 1666464484
transform 1 0 31556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1666464484
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_348
timestamp 1666464484
transform 1 0 33120 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_354
timestamp 1666464484
transform 1 0 33672 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_366
timestamp 1666464484
transform 1 0 34776 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_379
timestamp 1666464484
transform 1 0 35972 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1666464484
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1666464484
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_411
timestamp 1666464484
transform 1 0 38916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_424
timestamp 1666464484
transform 1 0 40112 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1666464484
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1666464484
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_453
timestamp 1666464484
transform 1 0 42780 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_465
timestamp 1666464484
transform 1 0 43884 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_477
timestamp 1666464484
transform 1 0 44988 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_489
timestamp 1666464484
transform 1 0 46092 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_501
timestamp 1666464484
transform 1 0 47196 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1666464484
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1666464484
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1666464484
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1666464484
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1666464484
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1666464484
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_561
timestamp 1666464484
transform 1 0 52716 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_571
timestamp 1666464484
transform 1 0 53636 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_579
timestamp 1666464484
transform 1 0 54372 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_9
timestamp 1666464484
transform 1 0 1932 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_147
timestamp 1666464484
transform 1 0 14628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_150
timestamp 1666464484
transform 1 0 14904 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_158
timestamp 1666464484
transform 1 0 15640 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_170
timestamp 1666464484
transform 1 0 16744 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_182
timestamp 1666464484
transform 1 0 17848 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1666464484
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_209
timestamp 1666464484
transform 1 0 20332 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_215
timestamp 1666464484
transform 1 0 20884 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_221
timestamp 1666464484
transform 1 0 21436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_227
timestamp 1666464484
transform 1 0 21988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_237
timestamp 1666464484
transform 1 0 22908 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_243
timestamp 1666464484
transform 1 0 23460 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_247
timestamp 1666464484
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666464484
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_260
timestamp 1666464484
transform 1 0 25024 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_271
timestamp 1666464484
transform 1 0 26036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_280
timestamp 1666464484
transform 1 0 26864 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 1666464484
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_320
timestamp 1666464484
transform 1 0 30544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_333
timestamp 1666464484
transform 1 0 31740 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_346
timestamp 1666464484
transform 1 0 32936 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_358
timestamp 1666464484
transform 1 0 34040 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1666464484
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_383
timestamp 1666464484
transform 1 0 36340 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_390
timestamp 1666464484
transform 1 0 36984 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_394
timestamp 1666464484
transform 1 0 37352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_404
timestamp 1666464484
transform 1 0 38272 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1666464484
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1666464484
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1666464484
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_430
timestamp 1666464484
transform 1 0 40664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_439
timestamp 1666464484
transform 1 0 41492 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_448
timestamp 1666464484
transform 1 0 42320 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_454
timestamp 1666464484
transform 1 0 42872 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_460
timestamp 1666464484
transform 1 0 43424 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_466
timestamp 1666464484
transform 1 0 43976 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_474
timestamp 1666464484
transform 1 0 44712 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1666464484
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1666464484
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1666464484
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1666464484
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1666464484
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1666464484
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1666464484
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1666464484
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_557
timestamp 1666464484
transform 1 0 52348 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_563
timestamp 1666464484
transform 1 0 52900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_571
timestamp 1666464484
transform 1 0 53636 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_579
timestamp 1666464484
transform 1 0 54372 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_9
timestamp 1666464484
transform 1 0 1932 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_16
timestamp 1666464484
transform 1 0 2576 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_28
timestamp 1666464484
transform 1 0 3680 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_40
timestamp 1666464484
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1666464484
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_146
timestamp 1666464484
transform 1 0 14536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1666464484
transform 1 0 15456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_162
timestamp 1666464484
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666464484
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666464484
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1666464484
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1666464484
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_233
timestamp 1666464484
transform 1 0 22540 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_239
timestamp 1666464484
transform 1 0 23092 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_253
timestamp 1666464484
transform 1 0 24380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1666464484
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_272
timestamp 1666464484
transform 1 0 26128 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1666464484
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_290
timestamp 1666464484
transform 1 0 27784 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_297
timestamp 1666464484
transform 1 0 28428 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_305
timestamp 1666464484
transform 1 0 29164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_314
timestamp 1666464484
transform 1 0 29992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1666464484
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_348
timestamp 1666464484
transform 1 0 33120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_361
timestamp 1666464484
transform 1 0 34316 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_365
timestamp 1666464484
transform 1 0 34684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_375
timestamp 1666464484
transform 1 0 35604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1666464484
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1666464484
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_402
timestamp 1666464484
transform 1 0 38088 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_408
timestamp 1666464484
transform 1 0 38640 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_416
timestamp 1666464484
transform 1 0 39376 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_425
timestamp 1666464484
transform 1 0 40204 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_429
timestamp 1666464484
transform 1 0 40572 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_446
timestamp 1666464484
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1666464484
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_454
timestamp 1666464484
transform 1 0 42872 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_460
timestamp 1666464484
transform 1 0 43424 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_472
timestamp 1666464484
transform 1 0 44528 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_484
timestamp 1666464484
transform 1 0 45632 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_496
timestamp 1666464484
transform 1 0 46736 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1666464484
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1666464484
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1666464484
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1666464484
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1666464484
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1666464484
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_561
timestamp 1666464484
transform 1 0 52716 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_571
timestamp 1666464484
transform 1 0 53636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_579
timestamp 1666464484
transform 1 0 54372 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_9
timestamp 1666464484
transform 1 0 1932 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1666464484
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_145
timestamp 1666464484
transform 1 0 14444 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_148
timestamp 1666464484
transform 1 0 14720 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_160
timestamp 1666464484
transform 1 0 15824 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_172
timestamp 1666464484
transform 1 0 16928 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_184
timestamp 1666464484
transform 1 0 18032 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666464484
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_221
timestamp 1666464484
transform 1 0 21436 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_229
timestamp 1666464484
transform 1 0 22172 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_234
timestamp 1666464484
transform 1 0 22632 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_241
timestamp 1666464484
transform 1 0 23276 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1666464484
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_260
timestamp 1666464484
transform 1 0 25024 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_268
timestamp 1666464484
transform 1 0 25760 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_278
timestamp 1666464484
transform 1 0 26680 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_285
timestamp 1666464484
transform 1 0 27324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_289
timestamp 1666464484
transform 1 0 27692 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_292
timestamp 1666464484
transform 1 0 27968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_298
timestamp 1666464484
transform 1 0 28520 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1666464484
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_328
timestamp 1666464484
transform 1 0 31280 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_348
timestamp 1666464484
transform 1 0 33120 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_354
timestamp 1666464484
transform 1 0 33672 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1666464484
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1666464484
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_376
timestamp 1666464484
transform 1 0 35696 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_392
timestamp 1666464484
transform 1 0 37168 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1666464484
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_414
timestamp 1666464484
transform 1 0 39192 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1666464484
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_428
timestamp 1666464484
transform 1 0 40480 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_432
timestamp 1666464484
transform 1 0 40848 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_449
timestamp 1666464484
transform 1 0 42412 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_456
timestamp 1666464484
transform 1 0 43056 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_468
timestamp 1666464484
transform 1 0 44160 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1666464484
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1666464484
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1666464484
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1666464484
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1666464484
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1666464484
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1666464484
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1666464484
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1666464484
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_571
timestamp 1666464484
transform 1 0 53636 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_579
timestamp 1666464484
transform 1 0 54372 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_9
timestamp 1666464484
transform 1 0 1932 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666464484
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666464484
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1666464484
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666464484
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_151
timestamp 1666464484
transform 1 0 14996 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_163
timestamp 1666464484
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1666464484
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666464484
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_229
timestamp 1666464484
transform 1 0 22172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_236
timestamp 1666464484
transform 1 0 22816 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_246
timestamp 1666464484
transform 1 0 23736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_250
timestamp 1666464484
transform 1 0 24104 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_260
timestamp 1666464484
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1666464484
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_292
timestamp 1666464484
transform 1 0 27968 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_298
timestamp 1666464484
transform 1 0 28520 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_304
timestamp 1666464484
transform 1 0 29072 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_310
timestamp 1666464484
transform 1 0 29624 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_317
timestamp 1666464484
transform 1 0 30268 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_321
timestamp 1666464484
transform 1 0 30636 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_328
timestamp 1666464484
transform 1 0 31280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1666464484
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_348
timestamp 1666464484
transform 1 0 33120 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_363
timestamp 1666464484
transform 1 0 34500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_371
timestamp 1666464484
transform 1 0 35236 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_377
timestamp 1666464484
transform 1 0 35788 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1666464484
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1666464484
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_400
timestamp 1666464484
transform 1 0 37904 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_420
timestamp 1666464484
transform 1 0 39744 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_426
timestamp 1666464484
transform 1 0 40296 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_446
timestamp 1666464484
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1666464484
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1666464484
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1666464484
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1666464484
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1666464484
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1666464484
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1666464484
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1666464484
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1666464484
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1666464484
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1666464484
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1666464484
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_561
timestamp 1666464484
transform 1 0 52716 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_571
timestamp 1666464484
transform 1 0 53636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_579
timestamp 1666464484
transform 1 0 54372 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_9
timestamp 1666464484
transform 1 0 1932 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666464484
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666464484
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_149
timestamp 1666464484
transform 1 0 14812 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_155
timestamp 1666464484
transform 1 0 15364 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_167
timestamp 1666464484
transform 1 0 16468 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_179
timestamp 1666464484
transform 1 0 17572 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1666464484
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666464484
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1666464484
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_233
timestamp 1666464484
transform 1 0 22540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_237
timestamp 1666464484
transform 1 0 22908 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_240
timestamp 1666464484
transform 1 0 23184 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1666464484
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_276
timestamp 1666464484
transform 1 0 26496 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_296
timestamp 1666464484
transform 1 0 28336 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_313
timestamp 1666464484
transform 1 0 29900 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_316
timestamp 1666464484
transform 1 0 30176 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_325
timestamp 1666464484
transform 1 0 31004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_334
timestamp 1666464484
transform 1 0 31832 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_341
timestamp 1666464484
transform 1 0 32476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_350
timestamp 1666464484
transform 1 0 33304 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1666464484
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1666464484
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_383
timestamp 1666464484
transform 1 0 36340 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1666464484
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_412
timestamp 1666464484
transform 1 0 39008 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1666464484
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1666464484
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_439
timestamp 1666464484
transform 1 0 41492 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_451
timestamp 1666464484
transform 1 0 42596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_463
timestamp 1666464484
transform 1 0 43700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1666464484
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1666464484
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1666464484
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1666464484
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1666464484
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1666464484
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1666464484
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1666464484
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_557
timestamp 1666464484
transform 1 0 52348 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_565
timestamp 1666464484
transform 1 0 53084 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_571
timestamp 1666464484
transform 1 0 53636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_579
timestamp 1666464484
transform 1 0 54372 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_9
timestamp 1666464484
transform 1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666464484
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666464484
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1666464484
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1666464484
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1666464484
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1666464484
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666464484
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_237
timestamp 1666464484
transform 1 0 22908 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_245
timestamp 1666464484
transform 1 0 23644 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_249
timestamp 1666464484
transform 1 0 24012 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_256
timestamp 1666464484
transform 1 0 24656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_277
timestamp 1666464484
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_299
timestamp 1666464484
transform 1 0 28612 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_307
timestamp 1666464484
transform 1 0 29348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_319
timestamp 1666464484
transform 1 0 30452 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_325
timestamp 1666464484
transform 1 0 31004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1666464484
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666464484
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_343
timestamp 1666464484
transform 1 0 32660 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_349
timestamp 1666464484
transform 1 0 33212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_369
timestamp 1666464484
transform 1 0 35052 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1666464484
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_393
timestamp 1666464484
transform 1 0 37260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_397
timestamp 1666464484
transform 1 0 37628 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_401
timestamp 1666464484
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_421
timestamp 1666464484
transform 1 0 39836 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_430
timestamp 1666464484
transform 1 0 40664 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_442
timestamp 1666464484
transform 1 0 41768 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1666464484
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1666464484
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1666464484
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1666464484
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1666464484
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1666464484
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1666464484
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1666464484
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1666464484
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1666464484
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1666464484
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1666464484
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_561
timestamp 1666464484
transform 1 0 52716 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_571
timestamp 1666464484
transform 1 0 53636 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_579
timestamp 1666464484
transform 1 0 54372 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_8
timestamp 1666464484
transform 1 0 1840 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_14
timestamp 1666464484
transform 1 0 2392 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1666464484
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666464484
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666464484
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666464484
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666464484
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1666464484
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1666464484
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666464484
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666464484
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1666464484
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1666464484
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1666464484
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666464484
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_257
timestamp 1666464484
transform 1 0 24748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_261
timestamp 1666464484
transform 1 0 25116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_272
timestamp 1666464484
transform 1 0 26128 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_295
timestamp 1666464484
transform 1 0 28244 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1666464484
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_321
timestamp 1666464484
transform 1 0 30636 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_327
timestamp 1666464484
transform 1 0 31188 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_330
timestamp 1666464484
transform 1 0 31464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_336
timestamp 1666464484
transform 1 0 32016 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_342
timestamp 1666464484
transform 1 0 32568 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_351
timestamp 1666464484
transform 1 0 33396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1666464484
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_365
timestamp 1666464484
transform 1 0 34684 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_372
timestamp 1666464484
transform 1 0 35328 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_379
timestamp 1666464484
transform 1 0 35972 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_386
timestamp 1666464484
transform 1 0 36616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_392
timestamp 1666464484
transform 1 0 37168 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_398
timestamp 1666464484
transform 1 0 37720 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_404
timestamp 1666464484
transform 1 0 38272 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_408
timestamp 1666464484
transform 1 0 38640 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_415
timestamp 1666464484
transform 1 0 39284 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1666464484
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_421
timestamp 1666464484
transform 1 0 39836 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_425
timestamp 1666464484
transform 1 0 40204 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_437
timestamp 1666464484
transform 1 0 41308 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_449
timestamp 1666464484
transform 1 0 42412 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_461
timestamp 1666464484
transform 1 0 43516 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_473
timestamp 1666464484
transform 1 0 44620 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1666464484
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1666464484
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1666464484
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1666464484
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1666464484
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1666464484
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1666464484
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1666464484
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_557
timestamp 1666464484
transform 1 0 52348 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_563
timestamp 1666464484
transform 1 0 52900 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_571
timestamp 1666464484
transform 1 0 53636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_579
timestamp 1666464484
transform 1 0 54372 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_8
timestamp 1666464484
transform 1 0 1840 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_14
timestamp 1666464484
transform 1 0 2392 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_26
timestamp 1666464484
transform 1 0 3496 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_38
timestamp 1666464484
transform 1 0 4600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1666464484
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666464484
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666464484
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666464484
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666464484
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1666464484
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1666464484
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666464484
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666464484
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_261
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_265
timestamp 1666464484
transform 1 0 25484 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1666464484
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_289
timestamp 1666464484
transform 1 0 27692 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_301
timestamp 1666464484
transform 1 0 28796 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_313
timestamp 1666464484
transform 1 0 29900 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_325
timestamp 1666464484
transform 1 0 31004 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1666464484
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_343
timestamp 1666464484
transform 1 0 32660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_349
timestamp 1666464484
transform 1 0 33212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_355
timestamp 1666464484
transform 1 0 33764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_366
timestamp 1666464484
transform 1 0 34776 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_373
timestamp 1666464484
transform 1 0 35420 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_379
timestamp 1666464484
transform 1 0 35972 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1666464484
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666464484
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 1666464484
transform 1 0 37260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_397
timestamp 1666464484
transform 1 0 37628 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_405
timestamp 1666464484
transform 1 0 38364 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_411
timestamp 1666464484
transform 1 0 38916 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_423
timestamp 1666464484
transform 1 0 40020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_435
timestamp 1666464484
transform 1 0 41124 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1666464484
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1666464484
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1666464484
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1666464484
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1666464484
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1666464484
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1666464484
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1666464484
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1666464484
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1666464484
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1666464484
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_553
timestamp 1666464484
transform 1 0 51980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_558
timestamp 1666464484
transform 1 0 52440 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_561
timestamp 1666464484
transform 1 0 52716 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_565
timestamp 1666464484
transform 1 0 53084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_579
timestamp 1666464484
transform 1 0 54372 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666464484
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666464484
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666464484
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666464484
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1666464484
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1666464484
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666464484
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666464484
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1666464484
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1666464484
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1666464484
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666464484
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_267
timestamp 1666464484
transform 1 0 25668 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_281
timestamp 1666464484
transform 1 0 26956 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_289
timestamp 1666464484
transform 1 0 27692 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_295
timestamp 1666464484
transform 1 0 28244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1666464484
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1666464484
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1666464484
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_345
timestamp 1666464484
transform 1 0 32844 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_349
timestamp 1666464484
transform 1 0 33212 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_352
timestamp 1666464484
transform 1 0 33488 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1666464484
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1666464484
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_369
timestamp 1666464484
transform 1 0 35052 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_375
timestamp 1666464484
transform 1 0 35604 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_381
timestamp 1666464484
transform 1 0 36156 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_387
timestamp 1666464484
transform 1 0 36708 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_393
timestamp 1666464484
transform 1 0 37260 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_405
timestamp 1666464484
transform 1 0 38364 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_417
timestamp 1666464484
transform 1 0 39468 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1666464484
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1666464484
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1666464484
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1666464484
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1666464484
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1666464484
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1666464484
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1666464484
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1666464484
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1666464484
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1666464484
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1666464484
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1666464484
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1666464484
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_557
timestamp 1666464484
transform 1 0 52348 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_563
timestamp 1666464484
transform 1 0 52900 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_571
timestamp 1666464484
transform 1 0 53636 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_579
timestamp 1666464484
transform 1 0 54372 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_21
timestamp 1666464484
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_33
timestamp 1666464484
transform 1 0 4140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1666464484
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1666464484
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666464484
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666464484
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666464484
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666464484
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666464484
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666464484
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666464484
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1666464484
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1666464484
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666464484
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_249
timestamp 1666464484
transform 1 0 24012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_255
timestamp 1666464484
transform 1 0 24564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_261
timestamp 1666464484
transform 1 0 25116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_267
timestamp 1666464484
transform 1 0 25668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1666464484
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_289
timestamp 1666464484
transform 1 0 27692 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_297
timestamp 1666464484
transform 1 0 28428 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_303
timestamp 1666464484
transform 1 0 28980 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_315
timestamp 1666464484
transform 1 0 30084 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_327
timestamp 1666464484
transform 1 0 31188 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1666464484
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1666464484
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_361
timestamp 1666464484
transform 1 0 34316 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_365
timestamp 1666464484
transform 1 0 34684 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_371
timestamp 1666464484
transform 1 0 35236 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_379
timestamp 1666464484
transform 1 0 35972 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1666464484
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1666464484
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1666464484
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1666464484
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1666464484
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1666464484
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1666464484
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1666464484
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1666464484
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1666464484
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1666464484
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1666464484
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666464484
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1666464484
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1666464484
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1666464484
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_541
timestamp 1666464484
transform 1 0 50876 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_549
timestamp 1666464484
transform 1 0 51612 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_552
timestamp 1666464484
transform 1 0 51888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_558
timestamp 1666464484
transform 1 0 52440 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_561
timestamp 1666464484
transform 1 0 52716 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_571
timestamp 1666464484
transform 1 0 53636 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_579
timestamp 1666464484
transform 1 0 54372 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_8
timestamp 1666464484
transform 1 0 1840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_14
timestamp 1666464484
transform 1 0 2392 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1666464484
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666464484
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666464484
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666464484
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666464484
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666464484
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1666464484
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1666464484
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1666464484
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666464484
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1666464484
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666464484
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_245
timestamp 1666464484
transform 1 0 23644 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1666464484
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_259
timestamp 1666464484
transform 1 0 24932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_265
timestamp 1666464484
transform 1 0 25484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_276
timestamp 1666464484
transform 1 0 26496 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_282
timestamp 1666464484
transform 1 0 27048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_291
timestamp 1666464484
transform 1 0 27876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_305
timestamp 1666464484
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_315
timestamp 1666464484
transform 1 0 30084 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_327
timestamp 1666464484
transform 1 0 31188 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_339
timestamp 1666464484
transform 1 0 32292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_351
timestamp 1666464484
transform 1 0 33396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1666464484
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1666464484
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1666464484
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1666464484
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1666464484
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1666464484
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1666464484
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1666464484
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1666464484
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1666464484
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1666464484
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1666464484
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1666464484
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1666464484
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1666464484
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1666464484
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1666464484
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1666464484
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1666464484
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1666464484
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1666464484
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_559
timestamp 1666464484
transform 1 0 52532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_565
timestamp 1666464484
transform 1 0 53084 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_579
timestamp 1666464484
transform 1 0 54372 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666464484
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666464484
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666464484
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666464484
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666464484
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666464484
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666464484
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666464484
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666464484
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666464484
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1666464484
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1666464484
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666464484
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1666464484
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1666464484
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1666464484
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1666464484
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666464484
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_249
timestamp 1666464484
transform 1 0 24012 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_255
timestamp 1666464484
transform 1 0 24564 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_258
timestamp 1666464484
transform 1 0 24840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_264
timestamp 1666464484
transform 1 0 25392 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1666464484
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_291
timestamp 1666464484
transform 1 0 27876 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_300
timestamp 1666464484
transform 1 0 28704 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_306
timestamp 1666464484
transform 1 0 29256 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_318
timestamp 1666464484
transform 1 0 30360 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1666464484
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666464484
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1666464484
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1666464484
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1666464484
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1666464484
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1666464484
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1666464484
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1666464484
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1666464484
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1666464484
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1666464484
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1666464484
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1666464484
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1666464484
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1666464484
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1666464484
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1666464484
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1666464484
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1666464484
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1666464484
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1666464484
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_553
timestamp 1666464484
transform 1 0 51980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_558
timestamp 1666464484
transform 1 0 52440 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_561
timestamp 1666464484
transform 1 0 52716 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_571
timestamp 1666464484
transform 1 0 53636 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_579
timestamp 1666464484
transform 1 0 54372 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_15
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1666464484
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666464484
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666464484
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666464484
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666464484
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_147
timestamp 1666464484
transform 1 0 14628 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_159
timestamp 1666464484
transform 1 0 15732 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_171
timestamp 1666464484
transform 1 0 16836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_183
timestamp 1666464484
transform 1 0 17940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666464484
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666464484
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666464484
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666464484
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666464484
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666464484
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_259
timestamp 1666464484
transform 1 0 24932 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_262
timestamp 1666464484
transform 1 0 25208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_268
timestamp 1666464484
transform 1 0 25760 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_278
timestamp 1666464484
transform 1 0 26680 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_286
timestamp 1666464484
transform 1 0 27416 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_297
timestamp 1666464484
transform 1 0 28428 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_303
timestamp 1666464484
transform 1 0 28980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666464484
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_316
timestamp 1666464484
transform 1 0 30176 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_328
timestamp 1666464484
transform 1 0 31280 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_340
timestamp 1666464484
transform 1 0 32384 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_352
timestamp 1666464484
transform 1 0 33488 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1666464484
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1666464484
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1666464484
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1666464484
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1666464484
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1666464484
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666464484
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666464484
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1666464484
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1666464484
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1666464484
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1666464484
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1666464484
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1666464484
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1666464484
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1666464484
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1666464484
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1666464484
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1666464484
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1666464484
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_557
timestamp 1666464484
transform 1 0 52348 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_563
timestamp 1666464484
transform 1 0 52900 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_571
timestamp 1666464484
transform 1 0 53636 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_579
timestamp 1666464484
transform 1 0 54372 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_21
timestamp 1666464484
transform 1 0 3036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_33
timestamp 1666464484
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1666464484
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1666464484
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666464484
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666464484
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666464484
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666464484
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_137
timestamp 1666464484
transform 1 0 13708 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_145
timestamp 1666464484
transform 1 0 14444 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_151
timestamp 1666464484
transform 1 0 14996 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_163
timestamp 1666464484
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1666464484
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1666464484
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1666464484
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1666464484
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1666464484
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1666464484
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1666464484
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_261
timestamp 1666464484
transform 1 0 25116 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_269
timestamp 1666464484
transform 1 0 25852 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_272
timestamp 1666464484
transform 1 0 26128 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1666464484
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_290
timestamp 1666464484
transform 1 0 27784 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_296
timestamp 1666464484
transform 1 0 28336 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_308
timestamp 1666464484
transform 1 0 29440 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_320
timestamp 1666464484
transform 1 0 30544 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1666464484
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666464484
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666464484
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1666464484
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1666464484
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1666464484
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666464484
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1666464484
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1666464484
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1666464484
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1666464484
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666464484
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1666464484
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1666464484
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1666464484
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1666464484
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1666464484
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1666464484
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1666464484
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1666464484
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1666464484
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1666464484
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1666464484
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1666464484
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_561
timestamp 1666464484
transform 1 0 52716 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_565
timestamp 1666464484
transform 1 0 53084 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_571
timestamp 1666464484
transform 1 0 53636 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_579
timestamp 1666464484
transform 1 0 54372 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_8
timestamp 1666464484
transform 1 0 1840 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_14
timestamp 1666464484
transform 1 0 2392 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_20
timestamp 1666464484
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666464484
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666464484
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666464484
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666464484
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666464484
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666464484
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666464484
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666464484
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666464484
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666464484
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1666464484
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1666464484
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1666464484
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1666464484
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666464484
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1666464484
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_277
timestamp 1666464484
transform 1 0 26588 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_281
timestamp 1666464484
transform 1 0 26956 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_289
timestamp 1666464484
transform 1 0 27692 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_292
timestamp 1666464484
transform 1 0 27968 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1666464484
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1666464484
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1666464484
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1666464484
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1666464484
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666464484
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1666464484
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1666464484
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1666464484
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1666464484
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1666464484
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1666464484
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666464484
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666464484
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1666464484
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1666464484
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1666464484
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1666464484
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1666464484
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1666464484
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1666464484
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1666464484
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1666464484
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1666464484
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1666464484
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1666464484
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1666464484
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_571
timestamp 1666464484
transform 1 0 53636 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_579
timestamp 1666464484
transform 1 0 54372 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666464484
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666464484
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666464484
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666464484
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666464484
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1666464484
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1666464484
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666464484
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666464484
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666464484
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1666464484
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1666464484
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_273
timestamp 1666464484
transform 1 0 26220 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1666464484
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1666464484
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1666464484
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1666464484
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1666464484
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666464484
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1666464484
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1666464484
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1666464484
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1666464484
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1666464484
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1666464484
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1666464484
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1666464484
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1666464484
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1666464484
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1666464484
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1666464484
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1666464484
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1666464484
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1666464484
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1666464484
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1666464484
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1666464484
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1666464484
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1666464484
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1666464484
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1666464484
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1666464484
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_561
timestamp 1666464484
transform 1 0 52716 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_571
timestamp 1666464484
transform 1 0 53636 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_579
timestamp 1666464484
transform 1 0 54372 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1666464484
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666464484
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666464484
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666464484
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666464484
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666464484
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666464484
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666464484
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1666464484
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666464484
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666464484
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1666464484
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1666464484
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1666464484
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1666464484
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666464484
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_265
timestamp 1666464484
transform 1 0 25484 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_271
timestamp 1666464484
transform 1 0 26036 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_274
timestamp 1666464484
transform 1 0 26312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_285
timestamp 1666464484
transform 1 0 27324 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_291
timestamp 1666464484
transform 1 0 27876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1666464484
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666464484
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1666464484
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1666464484
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1666464484
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1666464484
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1666464484
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1666464484
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1666464484
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1666464484
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1666464484
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1666464484
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1666464484
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666464484
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666464484
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1666464484
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1666464484
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1666464484
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1666464484
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1666464484
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1666464484
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1666464484
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1666464484
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1666464484
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1666464484
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1666464484
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1666464484
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1666464484
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1666464484
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_21
timestamp 1666464484
transform 1 0 3036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1666464484
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1666464484
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1666464484
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666464484
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666464484
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666464484
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666464484
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666464484
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1666464484
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1666464484
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666464484
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1666464484
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1666464484
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1666464484
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1666464484
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666464484
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1666464484
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1666464484
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_261
timestamp 1666464484
transform 1 0 25116 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_267
timestamp 1666464484
transform 1 0 25668 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1666464484
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_297
timestamp 1666464484
transform 1 0 28428 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_309
timestamp 1666464484
transform 1 0 29532 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_321
timestamp 1666464484
transform 1 0 30636 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_333
timestamp 1666464484
transform 1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1666464484
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1666464484
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1666464484
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1666464484
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1666464484
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666464484
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1666464484
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1666464484
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1666464484
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1666464484
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1666464484
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1666464484
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1666464484
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1666464484
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1666464484
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1666464484
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1666464484
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1666464484
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1666464484
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1666464484
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1666464484
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1666464484
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1666464484
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1666464484
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_573
timestamp 1666464484
transform 1 0 53820 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_579
timestamp 1666464484
transform 1 0 54372 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_15
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1666464484
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666464484
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666464484
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666464484
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666464484
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666464484
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1666464484
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1666464484
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1666464484
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1666464484
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666464484
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1666464484
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1666464484
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1666464484
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1666464484
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666464484
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_261
timestamp 1666464484
transform 1 0 25116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_267
timestamp 1666464484
transform 1 0 25668 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_273
timestamp 1666464484
transform 1 0 26220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_285
timestamp 1666464484
transform 1 0 27324 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_294
timestamp 1666464484
transform 1 0 28152 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1666464484
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666464484
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666464484
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1666464484
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1666464484
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666464484
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1666464484
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1666464484
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1666464484
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1666464484
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1666464484
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1666464484
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666464484
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1666464484
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1666464484
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1666464484
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1666464484
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1666464484
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1666464484
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1666464484
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1666464484
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1666464484
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1666464484
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1666464484
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1666464484
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1666464484
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1666464484
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_569
timestamp 1666464484
transform 1 0 53452 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_575
timestamp 1666464484
transform 1 0 54004 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_579
timestamp 1666464484
transform 1 0 54372 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666464484
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666464484
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1666464484
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1666464484
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1666464484
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1666464484
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1666464484
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1666464484
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_249
timestamp 1666464484
transform 1 0 24012 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_253
timestamp 1666464484
transform 1 0 24380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_260
timestamp 1666464484
transform 1 0 25024 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_264
timestamp 1666464484
transform 1 0 25392 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1666464484
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_286
timestamp 1666464484
transform 1 0 27416 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_292
timestamp 1666464484
transform 1 0 27968 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_298
timestamp 1666464484
transform 1 0 28520 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_310
timestamp 1666464484
transform 1 0 29624 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_322
timestamp 1666464484
transform 1 0 30728 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1666464484
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1666464484
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1666464484
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1666464484
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1666464484
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1666464484
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1666464484
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1666464484
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1666464484
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1666464484
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1666464484
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1666464484
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1666464484
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1666464484
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1666464484
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1666464484
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1666464484
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1666464484
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1666464484
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1666464484
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1666464484
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1666464484
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1666464484
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1666464484
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1666464484
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_573
timestamp 1666464484
transform 1 0 53820 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_8
timestamp 1666464484
transform 1 0 1840 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_14
timestamp 1666464484
transform 1 0 2392 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_20
timestamp 1666464484
transform 1 0 2944 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666464484
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666464484
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666464484
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666464484
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666464484
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666464484
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666464484
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1666464484
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1666464484
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1666464484
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666464484
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1666464484
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1666464484
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_233
timestamp 1666464484
transform 1 0 22540 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_56_243
timestamp 1666464484
transform 1 0 23460 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666464484
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_257
timestamp 1666464484
transform 1 0 24748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_267
timestamp 1666464484
transform 1 0 25668 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_281
timestamp 1666464484
transform 1 0 26956 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_287
timestamp 1666464484
transform 1 0 27508 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_298
timestamp 1666464484
transform 1 0 28520 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1666464484
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_313
timestamp 1666464484
transform 1 0 29900 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_325
timestamp 1666464484
transform 1 0 31004 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_337
timestamp 1666464484
transform 1 0 32108 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_349
timestamp 1666464484
transform 1 0 33212 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_361
timestamp 1666464484
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1666464484
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1666464484
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1666464484
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1666464484
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1666464484
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1666464484
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1666464484
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1666464484
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1666464484
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1666464484
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1666464484
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1666464484
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1666464484
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1666464484
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1666464484
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1666464484
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1666464484
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1666464484
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1666464484
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1666464484
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1666464484
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_569
timestamp 1666464484
transform 1 0 53452 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_575
timestamp 1666464484
transform 1 0 54004 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_579
timestamp 1666464484
transform 1 0 54372 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1666464484
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1666464484
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1666464484
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1666464484
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666464484
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666464484
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666464484
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666464484
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666464484
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666464484
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666464484
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1666464484
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1666464484
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1666464484
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1666464484
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1666464484
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1666464484
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_237
timestamp 1666464484
transform 1 0 22908 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_241
timestamp 1666464484
transform 1 0 23276 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_252
timestamp 1666464484
transform 1 0 24288 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_260
timestamp 1666464484
transform 1 0 25024 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_264
timestamp 1666464484
transform 1 0 25392 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1666464484
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_293
timestamp 1666464484
transform 1 0 28060 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_299
timestamp 1666464484
transform 1 0 28612 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_316
timestamp 1666464484
transform 1 0 30176 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_322
timestamp 1666464484
transform 1 0 30728 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_328
timestamp 1666464484
transform 1 0 31280 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1666464484
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1666464484
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1666464484
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1666464484
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1666464484
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1666464484
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1666464484
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1666464484
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1666464484
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1666464484
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1666464484
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1666464484
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1666464484
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1666464484
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1666464484
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1666464484
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666464484
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1666464484
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1666464484
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1666464484
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1666464484
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1666464484
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1666464484
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_561
timestamp 1666464484
transform 1 0 52716 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_567
timestamp 1666464484
transform 1 0 53268 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_575
timestamp 1666464484
transform 1 0 54004 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_579
timestamp 1666464484
transform 1 0 54372 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_15
timestamp 1666464484
transform 1 0 2484 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_21
timestamp 1666464484
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666464484
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666464484
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666464484
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666464484
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666464484
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666464484
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666464484
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666464484
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666464484
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666464484
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666464484
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666464484
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666464484
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_141
timestamp 1666464484
transform 1 0 14076 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_149
timestamp 1666464484
transform 1 0 14812 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_161
timestamp 1666464484
transform 1 0 15916 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_173
timestamp 1666464484
transform 1 0 17020 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_185
timestamp 1666464484
transform 1 0 18124 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 1666464484
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1666464484
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1666464484
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_221
timestamp 1666464484
transform 1 0 21436 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_229
timestamp 1666464484
transform 1 0 22172 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_232
timestamp 1666464484
transform 1 0 22448 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_238
timestamp 1666464484
transform 1 0 23000 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_244
timestamp 1666464484
transform 1 0 23552 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1666464484
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1666464484
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_259
timestamp 1666464484
transform 1 0 24932 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_269
timestamp 1666464484
transform 1 0 25852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_281
timestamp 1666464484
transform 1 0 26956 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_288
timestamp 1666464484
transform 1 0 27600 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_298
timestamp 1666464484
transform 1 0 28520 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1666464484
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1666464484
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_319
timestamp 1666464484
transform 1 0 30452 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_325
timestamp 1666464484
transform 1 0 31004 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_331
timestamp 1666464484
transform 1 0 31556 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_337
timestamp 1666464484
transform 1 0 32108 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_349
timestamp 1666464484
transform 1 0 33212 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_361
timestamp 1666464484
transform 1 0 34316 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1666464484
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1666464484
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1666464484
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1666464484
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1666464484
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1666464484
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1666464484
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1666464484
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1666464484
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1666464484
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1666464484
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1666464484
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1666464484
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1666464484
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1666464484
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1666464484
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1666464484
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1666464484
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1666464484
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1666464484
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_557
timestamp 1666464484
transform 1 0 52348 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_563
timestamp 1666464484
transform 1 0 52900 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_575
timestamp 1666464484
transform 1 0 54004 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666464484
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666464484
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666464484
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1666464484
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666464484
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666464484
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666464484
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666464484
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666464484
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666464484
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666464484
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666464484
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_125
timestamp 1666464484
transform 1 0 12604 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_133
timestamp 1666464484
transform 1 0 13340 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_136
timestamp 1666464484
transform 1 0 13616 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_147
timestamp 1666464484
transform 1 0 14628 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_153
timestamp 1666464484
transform 1 0 15180 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_159
timestamp 1666464484
transform 1 0 15732 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666464484
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1666464484
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1666464484
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1666464484
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1666464484
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_217
timestamp 1666464484
transform 1 0 21068 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1666464484
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_225
timestamp 1666464484
transform 1 0 21804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_233
timestamp 1666464484
transform 1 0 22540 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_239
timestamp 1666464484
transform 1 0 23092 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_245
timestamp 1666464484
transform 1 0 23644 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_256
timestamp 1666464484
transform 1 0 24656 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_268
timestamp 1666464484
transform 1 0 25760 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1666464484
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1666464484
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_289
timestamp 1666464484
transform 1 0 27692 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_302
timestamp 1666464484
transform 1 0 28888 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_314
timestamp 1666464484
transform 1 0 29992 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_326
timestamp 1666464484
transform 1 0 31096 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1666464484
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1666464484
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_341
timestamp 1666464484
transform 1 0 32476 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_347
timestamp 1666464484
transform 1 0 33028 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_359
timestamp 1666464484
transform 1 0 34132 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_371
timestamp 1666464484
transform 1 0 35236 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_383
timestamp 1666464484
transform 1 0 36340 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1666464484
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1666464484
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1666464484
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1666464484
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1666464484
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1666464484
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1666464484
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1666464484
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1666464484
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1666464484
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1666464484
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1666464484
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1666464484
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1666464484
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1666464484
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1666464484
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_541
timestamp 1666464484
transform 1 0 50876 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_551
timestamp 1666464484
transform 1 0 51796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_558
timestamp 1666464484
transform 1 0 52440 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_561
timestamp 1666464484
transform 1 0 52716 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_565
timestamp 1666464484
transform 1 0 53084 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_579
timestamp 1666464484
transform 1 0 54372 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_8
timestamp 1666464484
transform 1 0 1840 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_14
timestamp 1666464484
transform 1 0 2392 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_20
timestamp 1666464484
transform 1 0 2944 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666464484
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666464484
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666464484
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666464484
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666464484
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666464484
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666464484
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666464484
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666464484
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666464484
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666464484
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666464484
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1666464484
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_145
timestamp 1666464484
transform 1 0 14444 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_157
timestamp 1666464484
transform 1 0 15548 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_163
timestamp 1666464484
transform 1 0 16100 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_169
timestamp 1666464484
transform 1 0 16652 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_181
timestamp 1666464484
transform 1 0 17756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_193
timestamp 1666464484
transform 1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1666464484
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_209
timestamp 1666464484
transform 1 0 20332 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_219
timestamp 1666464484
transform 1 0 21252 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_225
timestamp 1666464484
transform 1 0 21804 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_231
timestamp 1666464484
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_237
timestamp 1666464484
transform 1 0 22908 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1666464484
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_253
timestamp 1666464484
transform 1 0 24380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_263
timestamp 1666464484
transform 1 0 25300 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_272
timestamp 1666464484
transform 1 0 26128 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_284
timestamp 1666464484
transform 1 0 27232 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_288
timestamp 1666464484
transform 1 0 27600 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_295
timestamp 1666464484
transform 1 0 28244 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1666464484
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_309
timestamp 1666464484
transform 1 0 29532 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_323
timestamp 1666464484
transform 1 0 30820 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_329
timestamp 1666464484
transform 1 0 31372 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_334
timestamp 1666464484
transform 1 0 31832 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_340
timestamp 1666464484
transform 1 0 32384 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_346
timestamp 1666464484
transform 1 0 32936 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_352
timestamp 1666464484
transform 1 0 33488 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1666464484
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1666464484
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1666464484
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1666464484
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1666464484
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1666464484
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1666464484
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1666464484
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1666464484
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1666464484
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1666464484
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1666464484
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1666464484
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1666464484
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1666464484
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1666464484
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1666464484
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1666464484
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1666464484
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1666464484
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_557
timestamp 1666464484
transform 1 0 52348 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_561
timestamp 1666464484
transform 1 0 52716 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_565
timestamp 1666464484
transform 1 0 53084 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_579
timestamp 1666464484
transform 1 0 54372 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_15
timestamp 1666464484
transform 1 0 2484 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_21
timestamp 1666464484
transform 1 0 3036 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_33
timestamp 1666464484
transform 1 0 4140 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_45
timestamp 1666464484
transform 1 0 5244 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1666464484
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666464484
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666464484
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666464484
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666464484
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666464484
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666464484
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666464484
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666464484
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1666464484
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1666464484
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1666464484
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666464484
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1666464484
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1666464484
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1666464484
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_205
timestamp 1666464484
transform 1 0 19964 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_210
timestamp 1666464484
transform 1 0 20424 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_216
timestamp 1666464484
transform 1 0 20976 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1666464484
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1666464484
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_231
timestamp 1666464484
transform 1 0 22356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_234
timestamp 1666464484
transform 1 0 22632 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_240
timestamp 1666464484
transform 1 0 23184 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_252
timestamp 1666464484
transform 1 0 24288 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_264
timestamp 1666464484
transform 1 0 25392 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_270
timestamp 1666464484
transform 1 0 25944 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1666464484
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1666464484
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_291
timestamp 1666464484
transform 1 0 27876 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_301
timestamp 1666464484
transform 1 0 28796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_309
timestamp 1666464484
transform 1 0 29532 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_321
timestamp 1666464484
transform 1 0 30636 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_327
timestamp 1666464484
transform 1 0 31188 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp 1666464484
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1666464484
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_341
timestamp 1666464484
transform 1 0 32476 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_347
timestamp 1666464484
transform 1 0 33028 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_359
timestamp 1666464484
transform 1 0 34132 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_371
timestamp 1666464484
transform 1 0 35236 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_383
timestamp 1666464484
transform 1 0 36340 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1666464484
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1666464484
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1666464484
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1666464484
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1666464484
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1666464484
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1666464484
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1666464484
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1666464484
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1666464484
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1666464484
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1666464484
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1666464484
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1666464484
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1666464484
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1666464484
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1666464484
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_553
timestamp 1666464484
transform 1 0 51980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_558
timestamp 1666464484
transform 1 0 52440 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_561
timestamp 1666464484
transform 1 0 52716 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_565
timestamp 1666464484
transform 1 0 53084 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_579
timestamp 1666464484
transform 1 0 54372 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_15
timestamp 1666464484
transform 1 0 2484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1666464484
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666464484
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666464484
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666464484
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1666464484
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666464484
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1666464484
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666464484
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666464484
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666464484
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666464484
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666464484
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666464484
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666464484
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666464484
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666464484
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1666464484
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1666464484
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1666464484
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1666464484
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1666464484
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_209
timestamp 1666464484
transform 1 0 20332 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_217
timestamp 1666464484
transform 1 0 21068 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_220
timestamp 1666464484
transform 1 0 21344 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_226
timestamp 1666464484
transform 1 0 21896 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_232
timestamp 1666464484
transform 1 0 22448 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_238
timestamp 1666464484
transform 1 0 23000 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_244
timestamp 1666464484
transform 1 0 23552 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1666464484
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_253
timestamp 1666464484
transform 1 0 24380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_258
timestamp 1666464484
transform 1 0 24840 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_270
timestamp 1666464484
transform 1 0 25944 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_279
timestamp 1666464484
transform 1 0 26772 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_290
timestamp 1666464484
transform 1 0 27784 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1666464484
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1666464484
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1666464484
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_313
timestamp 1666464484
transform 1 0 29900 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_319
timestamp 1666464484
transform 1 0 30452 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_325
timestamp 1666464484
transform 1 0 31004 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_331
timestamp 1666464484
transform 1 0 31556 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_337
timestamp 1666464484
transform 1 0 32108 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_343
timestamp 1666464484
transform 1 0 32660 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_355
timestamp 1666464484
transform 1 0 33764 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1666464484
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1666464484
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1666464484
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1666464484
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1666464484
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1666464484
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1666464484
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1666464484
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1666464484
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1666464484
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1666464484
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1666464484
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1666464484
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1666464484
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1666464484
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1666464484
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1666464484
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1666464484
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1666464484
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1666464484
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_545
timestamp 1666464484
transform 1 0 51244 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_549
timestamp 1666464484
transform 1 0 51612 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_552
timestamp 1666464484
transform 1 0 51888 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_558
timestamp 1666464484
transform 1 0 52440 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_565
timestamp 1666464484
transform 1 0 53084 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_579
timestamp 1666464484
transform 1 0 54372 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_15
timestamp 1666464484
transform 1 0 2484 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_21
timestamp 1666464484
transform 1 0 3036 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_33
timestamp 1666464484
transform 1 0 4140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_45
timestamp 1666464484
transform 1 0 5244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 1666464484
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1666464484
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666464484
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666464484
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666464484
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666464484
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666464484
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1666464484
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1666464484
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1666464484
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1666464484
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1666464484
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1666464484
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1666464484
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1666464484
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1666464484
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1666464484
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1666464484
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1666464484
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1666464484
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_229
timestamp 1666464484
transform 1 0 22172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_235
timestamp 1666464484
transform 1 0 22724 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_241
timestamp 1666464484
transform 1 0 23276 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_247
timestamp 1666464484
transform 1 0 23828 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_253
timestamp 1666464484
transform 1 0 24380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_259
timestamp 1666464484
transform 1 0 24932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_265
timestamp 1666464484
transform 1 0 25484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1666464484
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1666464484
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_290
timestamp 1666464484
transform 1 0 27784 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_301
timestamp 1666464484
transform 1 0 28796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_309
timestamp 1666464484
transform 1 0 29532 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_315
timestamp 1666464484
transform 1 0 30084 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_322
timestamp 1666464484
transform 1 0 30728 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_328
timestamp 1666464484
transform 1 0 31280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1666464484
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1666464484
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_341
timestamp 1666464484
transform 1 0 32476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_347
timestamp 1666464484
transform 1 0 33028 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_353
timestamp 1666464484
transform 1 0 33580 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_365
timestamp 1666464484
transform 1 0 34684 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_377
timestamp 1666464484
transform 1 0 35788 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_389
timestamp 1666464484
transform 1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1666464484
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1666464484
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1666464484
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1666464484
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1666464484
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1666464484
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1666464484
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1666464484
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1666464484
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1666464484
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1666464484
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1666464484
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1666464484
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1666464484
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1666464484
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1666464484
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_553
timestamp 1666464484
transform 1 0 51980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_558
timestamp 1666464484
transform 1 0 52440 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_561
timestamp 1666464484
transform 1 0 52716 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_565
timestamp 1666464484
transform 1 0 53084 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_579
timestamp 1666464484
transform 1 0 54372 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1666464484
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666464484
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1666464484
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1666464484
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1666464484
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1666464484
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1666464484
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1666464484
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1666464484
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1666464484
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1666464484
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1666464484
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1666464484
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1666464484
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1666464484
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1666464484
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1666464484
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1666464484
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1666464484
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1666464484
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1666464484
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1666464484
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_221
timestamp 1666464484
transform 1 0 21436 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_229
timestamp 1666464484
transform 1 0 22172 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_232
timestamp 1666464484
transform 1 0 22448 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_238
timestamp 1666464484
transform 1 0 23000 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_244
timestamp 1666464484
transform 1 0 23552 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1666464484
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_253
timestamp 1666464484
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_258
timestamp 1666464484
transform 1 0 24840 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_264
timestamp 1666464484
transform 1 0 25392 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_272
timestamp 1666464484
transform 1 0 26128 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_284
timestamp 1666464484
transform 1 0 27232 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_296
timestamp 1666464484
transform 1 0 28336 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1666464484
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1666464484
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_319
timestamp 1666464484
transform 1 0 30452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_327
timestamp 1666464484
transform 1 0 31188 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_333
timestamp 1666464484
transform 1 0 31740 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_339
timestamp 1666464484
transform 1 0 32292 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_351
timestamp 1666464484
transform 1 0 33396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1666464484
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1666464484
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1666464484
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1666464484
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1666464484
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1666464484
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1666464484
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1666464484
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1666464484
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1666464484
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1666464484
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1666464484
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1666464484
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1666464484
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1666464484
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1666464484
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1666464484
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1666464484
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1666464484
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1666464484
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1666464484
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_545
timestamp 1666464484
transform 1 0 51244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_551
timestamp 1666464484
transform 1 0 51796 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_565
timestamp 1666464484
transform 1 0 53084 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_579
timestamp 1666464484
transform 1 0 54372 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1666464484
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_8
timestamp 1666464484
transform 1 0 1840 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_14
timestamp 1666464484
transform 1 0 2392 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_20
timestamp 1666464484
transform 1 0 2944 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_32
timestamp 1666464484
transform 1 0 4048 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_44
timestamp 1666464484
transform 1 0 5152 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1666464484
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1666464484
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1666464484
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1666464484
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1666464484
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1666464484
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1666464484
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1666464484
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1666464484
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1666464484
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1666464484
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1666464484
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1666464484
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1666464484
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1666464484
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1666464484
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1666464484
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1666464484
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_225
timestamp 1666464484
transform 1 0 21804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_231
timestamp 1666464484
transform 1 0 22356 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_234
timestamp 1666464484
transform 1 0 22632 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_240
timestamp 1666464484
transform 1 0 23184 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_246
timestamp 1666464484
transform 1 0 23736 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_252
timestamp 1666464484
transform 1 0 24288 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_258
timestamp 1666464484
transform 1 0 24840 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_267
timestamp 1666464484
transform 1 0 25668 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_278
timestamp 1666464484
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_281
timestamp 1666464484
transform 1 0 26956 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_292
timestamp 1666464484
transform 1 0 27968 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_298
timestamp 1666464484
transform 1 0 28520 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_302
timestamp 1666464484
transform 1 0 28888 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_311
timestamp 1666464484
transform 1 0 29716 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_323
timestamp 1666464484
transform 1 0 30820 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1666464484
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1666464484
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_337
timestamp 1666464484
transform 1 0 32108 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_345
timestamp 1666464484
transform 1 0 32844 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_351
timestamp 1666464484
transform 1 0 33396 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_357
timestamp 1666464484
transform 1 0 33948 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_363
timestamp 1666464484
transform 1 0 34500 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_369
timestamp 1666464484
transform 1 0 35052 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_381
timestamp 1666464484
transform 1 0 36156 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_389
timestamp 1666464484
transform 1 0 36892 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1666464484
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1666464484
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1666464484
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1666464484
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1666464484
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1666464484
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1666464484
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1666464484
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1666464484
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1666464484
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1666464484
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1666464484
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1666464484
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1666464484
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1666464484
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_541
timestamp 1666464484
transform 1 0 50876 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_544
timestamp 1666464484
transform 1 0 51152 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_558
timestamp 1666464484
transform 1 0 52440 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_561
timestamp 1666464484
transform 1 0 52716 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_565
timestamp 1666464484
transform 1 0 53084 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_579
timestamp 1666464484
transform 1 0 54372 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1666464484
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_9
timestamp 1666464484
transform 1 0 1932 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1666464484
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1666464484
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1666464484
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1666464484
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1666464484
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1666464484
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1666464484
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1666464484
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1666464484
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1666464484
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1666464484
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1666464484
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1666464484
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1666464484
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1666464484
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1666464484
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1666464484
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_177
timestamp 1666464484
transform 1 0 17388 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_180
timestamp 1666464484
transform 1 0 17664 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_192
timestamp 1666464484
transform 1 0 18768 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1666464484
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1666464484
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1666464484
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_233
timestamp 1666464484
transform 1 0 22540 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_238
timestamp 1666464484
transform 1 0 23000 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_244
timestamp 1666464484
transform 1 0 23552 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1666464484
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_253
timestamp 1666464484
transform 1 0 24380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_259
timestamp 1666464484
transform 1 0 24932 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_265
timestamp 1666464484
transform 1 0 25484 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_271
timestamp 1666464484
transform 1 0 26036 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_282
timestamp 1666464484
transform 1 0 27048 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_292
timestamp 1666464484
transform 1 0 27968 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_300
timestamp 1666464484
transform 1 0 28704 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_306
timestamp 1666464484
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_309
timestamp 1666464484
transform 1 0 29532 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_317
timestamp 1666464484
transform 1 0 30268 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_325
timestamp 1666464484
transform 1 0 31004 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_333
timestamp 1666464484
transform 1 0 31740 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_341
timestamp 1666464484
transform 1 0 32476 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_346
timestamp 1666464484
transform 1 0 32936 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_354
timestamp 1666464484
transform 1 0 33672 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_360
timestamp 1666464484
transform 1 0 34224 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1666464484
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1666464484
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1666464484
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1666464484
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1666464484
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1666464484
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1666464484
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1666464484
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1666464484
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1666464484
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1666464484
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1666464484
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1666464484
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1666464484
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1666464484
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1666464484
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1666464484
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1666464484
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_533
timestamp 1666464484
transform 1 0 50140 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_541
timestamp 1666464484
transform 1 0 50876 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_545
timestamp 1666464484
transform 1 0 51244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_551
timestamp 1666464484
transform 1 0 51796 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_565
timestamp 1666464484
transform 1 0 53084 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_579
timestamp 1666464484
transform 1 0 54372 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1666464484
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_15
timestamp 1666464484
transform 1 0 2484 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_21
timestamp 1666464484
transform 1 0 3036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_33
timestamp 1666464484
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1666464484
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1666464484
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1666464484
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1666464484
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1666464484
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1666464484
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1666464484
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666464484
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1666464484
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1666464484
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1666464484
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1666464484
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_161
timestamp 1666464484
transform 1 0 15916 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_166
timestamp 1666464484
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1666464484
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_178
timestamp 1666464484
transform 1 0 17480 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_184
timestamp 1666464484
transform 1 0 18032 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_196
timestamp 1666464484
transform 1 0 19136 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_208
timestamp 1666464484
transform 1 0 20240 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_220
timestamp 1666464484
transform 1 0 21344 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1666464484
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_239
timestamp 1666464484
transform 1 0 23092 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_245
timestamp 1666464484
transform 1 0 23644 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_251
timestamp 1666464484
transform 1 0 24196 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_257
timestamp 1666464484
transform 1 0 24748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_263
timestamp 1666464484
transform 1 0 25300 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_269
timestamp 1666464484
transform 1 0 25852 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_278
timestamp 1666464484
transform 1 0 26680 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 1666464484
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_292
timestamp 1666464484
transform 1 0 27968 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_300
timestamp 1666464484
transform 1 0 28704 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_309
timestamp 1666464484
transform 1 0 29532 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_315
timestamp 1666464484
transform 1 0 30084 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_321
timestamp 1666464484
transform 1 0 30636 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_329
timestamp 1666464484
transform 1 0 31372 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_334
timestamp 1666464484
transform 1 0 31832 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_337
timestamp 1666464484
transform 1 0 32108 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_341
timestamp 1666464484
transform 1 0 32476 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_350
timestamp 1666464484
transform 1 0 33304 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_358
timestamp 1666464484
transform 1 0 34040 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_366
timestamp 1666464484
transform 1 0 34776 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_378
timestamp 1666464484
transform 1 0 35880 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_390
timestamp 1666464484
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1666464484
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1666464484
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1666464484
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1666464484
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1666464484
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1666464484
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1666464484
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1666464484
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1666464484
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1666464484
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1666464484
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1666464484
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1666464484
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1666464484
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1666464484
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_541
timestamp 1666464484
transform 1 0 50876 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_547
timestamp 1666464484
transform 1 0 51428 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_558
timestamp 1666464484
transform 1 0 52440 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_561
timestamp 1666464484
transform 1 0 52716 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_565
timestamp 1666464484
transform 1 0 53084 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_579
timestamp 1666464484
transform 1 0 54372 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1666464484
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_15
timestamp 1666464484
transform 1 0 2484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_21
timestamp 1666464484
transform 1 0 3036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1666464484
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1666464484
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1666464484
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1666464484
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1666464484
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1666464484
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1666464484
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1666464484
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1666464484
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1666464484
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1666464484
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1666464484
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1666464484
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1666464484
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1666464484
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1666464484
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1666464484
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1666464484
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1666464484
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1666464484
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1666464484
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_221
timestamp 1666464484
transform 1 0 21436 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_229
timestamp 1666464484
transform 1 0 22172 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_232
timestamp 1666464484
transform 1 0 22448 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_238
timestamp 1666464484
transform 1 0 23000 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_244
timestamp 1666464484
transform 1 0 23552 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1666464484
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_253
timestamp 1666464484
transform 1 0 24380 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_259
timestamp 1666464484
transform 1 0 24932 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_268
timestamp 1666464484
transform 1 0 25760 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_281
timestamp 1666464484
transform 1 0 26956 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_292
timestamp 1666464484
transform 1 0 27968 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1666464484
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1666464484
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_309
timestamp 1666464484
transform 1 0 29532 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_313
timestamp 1666464484
transform 1 0 29900 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_323
timestamp 1666464484
transform 1 0 30820 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_332
timestamp 1666464484
transform 1 0 31648 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_340
timestamp 1666464484
transform 1 0 32384 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_346
timestamp 1666464484
transform 1 0 32936 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_355
timestamp 1666464484
transform 1 0 33764 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_68_361
timestamp 1666464484
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_365
timestamp 1666464484
transform 1 0 34684 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_371
timestamp 1666464484
transform 1 0 35236 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1666464484
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1666464484
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1666464484
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1666464484
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1666464484
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1666464484
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1666464484
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1666464484
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1666464484
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1666464484
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1666464484
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1666464484
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1666464484
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1666464484
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1666464484
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1666464484
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1666464484
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1666464484
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_545
timestamp 1666464484
transform 1 0 51244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_549
timestamp 1666464484
transform 1 0 51612 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_552
timestamp 1666464484
transform 1 0 51888 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_558
timestamp 1666464484
transform 1 0 52440 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_565
timestamp 1666464484
transform 1 0 53084 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_579
timestamp 1666464484
transform 1 0 54372 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_3
timestamp 1666464484
transform 1 0 1380 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_15
timestamp 1666464484
transform 1 0 2484 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_21
timestamp 1666464484
transform 1 0 3036 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_33
timestamp 1666464484
transform 1 0 4140 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_45
timestamp 1666464484
transform 1 0 5244 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_53
timestamp 1666464484
transform 1 0 5980 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1666464484
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1666464484
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1666464484
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1666464484
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1666464484
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1666464484
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1666464484
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1666464484
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1666464484
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1666464484
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1666464484
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1666464484
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1666464484
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1666464484
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1666464484
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1666464484
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1666464484
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1666464484
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_225
timestamp 1666464484
transform 1 0 21804 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_233
timestamp 1666464484
transform 1 0 22540 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_237
timestamp 1666464484
transform 1 0 22908 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_243
timestamp 1666464484
transform 1 0 23460 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_249
timestamp 1666464484
transform 1 0 24012 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_255
timestamp 1666464484
transform 1 0 24564 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_261
timestamp 1666464484
transform 1 0 25116 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_269
timestamp 1666464484
transform 1 0 25852 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_278
timestamp 1666464484
transform 1 0 26680 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_281
timestamp 1666464484
transform 1 0 26956 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_291
timestamp 1666464484
transform 1 0 27876 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_305
timestamp 1666464484
transform 1 0 29164 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_311
timestamp 1666464484
transform 1 0 29716 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_320
timestamp 1666464484
transform 1 0 30544 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_333
timestamp 1666464484
transform 1 0 31740 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_337
timestamp 1666464484
transform 1 0 32108 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_347
timestamp 1666464484
transform 1 0 33028 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_356
timestamp 1666464484
transform 1 0 33856 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_365
timestamp 1666464484
transform 1 0 34684 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_373
timestamp 1666464484
transform 1 0 35420 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_379
timestamp 1666464484
transform 1 0 35972 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1666464484
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1666464484
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1666464484
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1666464484
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1666464484
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1666464484
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1666464484
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1666464484
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1666464484
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1666464484
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1666464484
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1666464484
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1666464484
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1666464484
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1666464484
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1666464484
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_541
timestamp 1666464484
transform 1 0 50876 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_549
timestamp 1666464484
transform 1 0 51612 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_552
timestamp 1666464484
transform 1 0 51888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_558
timestamp 1666464484
transform 1 0 52440 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_561
timestamp 1666464484
transform 1 0 52716 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_565
timestamp 1666464484
transform 1 0 53084 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_579
timestamp 1666464484
transform 1 0 54372 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1666464484
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_15
timestamp 1666464484
transform 1 0 2484 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_21
timestamp 1666464484
transform 1 0 3036 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1666464484
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1666464484
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1666464484
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1666464484
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1666464484
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1666464484
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1666464484
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1666464484
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1666464484
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1666464484
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1666464484
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1666464484
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1666464484
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1666464484
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1666464484
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1666464484
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1666464484
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1666464484
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1666464484
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1666464484
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1666464484
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1666464484
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_233
timestamp 1666464484
transform 1 0 22540 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_241
timestamp 1666464484
transform 1 0 23276 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_244
timestamp 1666464484
transform 1 0 23552 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 1666464484
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_253
timestamp 1666464484
transform 1 0 24380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_257
timestamp 1666464484
transform 1 0 24748 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_260
timestamp 1666464484
transform 1 0 25024 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_266
timestamp 1666464484
transform 1 0 25576 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_277
timestamp 1666464484
transform 1 0 26588 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_283
timestamp 1666464484
transform 1 0 27140 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_292
timestamp 1666464484
transform 1 0 27968 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_304
timestamp 1666464484
transform 1 0 29072 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_309
timestamp 1666464484
transform 1 0 29532 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_313
timestamp 1666464484
transform 1 0 29900 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_319
timestamp 1666464484
transform 1 0 30452 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_325
timestamp 1666464484
transform 1 0 31004 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_331
timestamp 1666464484
transform 1 0 31556 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_336
timestamp 1666464484
transform 1 0 32016 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_348
timestamp 1666464484
transform 1 0 33120 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1666464484
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1666464484
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_365
timestamp 1666464484
transform 1 0 34684 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_371
timestamp 1666464484
transform 1 0 35236 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_377
timestamp 1666464484
transform 1 0 35788 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_383
timestamp 1666464484
transform 1 0 36340 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_395
timestamp 1666464484
transform 1 0 37444 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_407
timestamp 1666464484
transform 1 0 38548 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1666464484
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1666464484
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1666464484
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1666464484
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1666464484
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1666464484
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1666464484
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1666464484
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1666464484
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1666464484
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1666464484
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1666464484
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1666464484
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1666464484
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_545
timestamp 1666464484
transform 1 0 51244 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_551
timestamp 1666464484
transform 1 0 51796 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_558
timestamp 1666464484
transform 1 0 52440 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_565
timestamp 1666464484
transform 1 0 53084 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_572
timestamp 1666464484
transform 1 0 53728 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_579
timestamp 1666464484
transform 1 0 54372 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1666464484
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_15
timestamp 1666464484
transform 1 0 2484 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_21
timestamp 1666464484
transform 1 0 3036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_33
timestamp 1666464484
transform 1 0 4140 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_45
timestamp 1666464484
transform 1 0 5244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1666464484
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1666464484
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1666464484
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1666464484
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1666464484
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1666464484
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1666464484
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1666464484
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1666464484
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1666464484
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1666464484
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1666464484
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1666464484
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1666464484
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1666464484
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1666464484
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1666464484
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1666464484
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1666464484
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1666464484
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_237
timestamp 1666464484
transform 1 0 22908 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_245
timestamp 1666464484
transform 1 0 23644 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_250
timestamp 1666464484
transform 1 0 24104 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_256
timestamp 1666464484
transform 1 0 24656 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_262
timestamp 1666464484
transform 1 0 25208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_268
timestamp 1666464484
transform 1 0 25760 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_278
timestamp 1666464484
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_281
timestamp 1666464484
transform 1 0 26956 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_290
timestamp 1666464484
transform 1 0 27784 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_294
timestamp 1666464484
transform 1 0 28152 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_302
timestamp 1666464484
transform 1 0 28888 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_314
timestamp 1666464484
transform 1 0 29992 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_320
timestamp 1666464484
transform 1 0 30544 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_326
timestamp 1666464484
transform 1 0 31096 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_332
timestamp 1666464484
transform 1 0 31648 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_337
timestamp 1666464484
transform 1 0 32108 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_343
timestamp 1666464484
transform 1 0 32660 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_352
timestamp 1666464484
transform 1 0 33488 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_361
timestamp 1666464484
transform 1 0 34316 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_367
timestamp 1666464484
transform 1 0 34868 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_373
timestamp 1666464484
transform 1 0 35420 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_379
timestamp 1666464484
transform 1 0 35972 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1666464484
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1666464484
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1666464484
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1666464484
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1666464484
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1666464484
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1666464484
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1666464484
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1666464484
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1666464484
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1666464484
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1666464484
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1666464484
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1666464484
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1666464484
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1666464484
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_541
timestamp 1666464484
transform 1 0 50876 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_549
timestamp 1666464484
transform 1 0 51612 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_552
timestamp 1666464484
transform 1 0 51888 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_558
timestamp 1666464484
transform 1 0 52440 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_561
timestamp 1666464484
transform 1 0 52716 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_565
timestamp 1666464484
transform 1 0 53084 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_579
timestamp 1666464484
transform 1 0 54372 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1666464484
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_15
timestamp 1666464484
transform 1 0 2484 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_21
timestamp 1666464484
transform 1 0 3036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1666464484
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1666464484
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1666464484
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1666464484
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1666464484
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1666464484
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1666464484
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1666464484
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1666464484
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1666464484
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1666464484
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1666464484
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1666464484
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1666464484
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1666464484
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1666464484
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1666464484
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1666464484
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1666464484
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1666464484
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1666464484
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1666464484
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_233
timestamp 1666464484
transform 1 0 22540 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_241
timestamp 1666464484
transform 1 0 23276 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_244
timestamp 1666464484
transform 1 0 23552 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_250
timestamp 1666464484
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 1666464484
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_261
timestamp 1666464484
transform 1 0 25116 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_271
timestamp 1666464484
transform 1 0 26036 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_277
timestamp 1666464484
transform 1 0 26588 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_285
timestamp 1666464484
transform 1 0 27324 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_297
timestamp 1666464484
transform 1 0 28428 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_303
timestamp 1666464484
transform 1 0 28980 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1666464484
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_309
timestamp 1666464484
transform 1 0 29532 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_319
timestamp 1666464484
transform 1 0 30452 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_331
timestamp 1666464484
transform 1 0 31556 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_339
timestamp 1666464484
transform 1 0 32292 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_348
timestamp 1666464484
transform 1 0 33120 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_359
timestamp 1666464484
transform 1 0 34132 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1666464484
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_365
timestamp 1666464484
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_372
timestamp 1666464484
transform 1 0 35328 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_378
timestamp 1666464484
transform 1 0 35880 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_384
timestamp 1666464484
transform 1 0 36432 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_390
timestamp 1666464484
transform 1 0 36984 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_402
timestamp 1666464484
transform 1 0 38088 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_414
timestamp 1666464484
transform 1 0 39192 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1666464484
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1666464484
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1666464484
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1666464484
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1666464484
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1666464484
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1666464484
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1666464484
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1666464484
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1666464484
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1666464484
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1666464484
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1666464484
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_545
timestamp 1666464484
transform 1 0 51244 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_551
timestamp 1666464484
transform 1 0 51796 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_558
timestamp 1666464484
transform 1 0 52440 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_565
timestamp 1666464484
transform 1 0 53084 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_572
timestamp 1666464484
transform 1 0 53728 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_579
timestamp 1666464484
transform 1 0 54372 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_3
timestamp 1666464484
transform 1 0 1380 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_15
timestamp 1666464484
transform 1 0 2484 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_21
timestamp 1666464484
transform 1 0 3036 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_33
timestamp 1666464484
transform 1 0 4140 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_45
timestamp 1666464484
transform 1 0 5244 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_53
timestamp 1666464484
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1666464484
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1666464484
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1666464484
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1666464484
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1666464484
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1666464484
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1666464484
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1666464484
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1666464484
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1666464484
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1666464484
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1666464484
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1666464484
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1666464484
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1666464484
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1666464484
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1666464484
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1666464484
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1666464484
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_237
timestamp 1666464484
transform 1 0 22908 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_245
timestamp 1666464484
transform 1 0 23644 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_248
timestamp 1666464484
transform 1 0 23920 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_254
timestamp 1666464484
transform 1 0 24472 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_265
timestamp 1666464484
transform 1 0 25484 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_278
timestamp 1666464484
transform 1 0 26680 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_281
timestamp 1666464484
transform 1 0 26956 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_287
timestamp 1666464484
transform 1 0 27508 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_290
timestamp 1666464484
transform 1 0 27784 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_302
timestamp 1666464484
transform 1 0 28888 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_308
timestamp 1666464484
transform 1 0 29440 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_314
timestamp 1666464484
transform 1 0 29992 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_323
timestamp 1666464484
transform 1 0 30820 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1666464484
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1666464484
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_337
timestamp 1666464484
transform 1 0 32108 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_349
timestamp 1666464484
transform 1 0 33212 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_360
timestamp 1666464484
transform 1 0 34224 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_366
timestamp 1666464484
transform 1 0 34776 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_372
timestamp 1666464484
transform 1 0 35328 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_378
timestamp 1666464484
transform 1 0 35880 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_384
timestamp 1666464484
transform 1 0 36432 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1666464484
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1666464484
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1666464484
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1666464484
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1666464484
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1666464484
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1666464484
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1666464484
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1666464484
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1666464484
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1666464484
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1666464484
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1666464484
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1666464484
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1666464484
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_541
timestamp 1666464484
transform 1 0 50876 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_549
timestamp 1666464484
transform 1 0 51612 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_552
timestamp 1666464484
transform 1 0 51888 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_558
timestamp 1666464484
transform 1 0 52440 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_561
timestamp 1666464484
transform 1 0 52716 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_565
timestamp 1666464484
transform 1 0 53084 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_579
timestamp 1666464484
transform 1 0 54372 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1666464484
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_15
timestamp 1666464484
transform 1 0 2484 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_21
timestamp 1666464484
transform 1 0 3036 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1666464484
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1666464484
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1666464484
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1666464484
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1666464484
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1666464484
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1666464484
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1666464484
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1666464484
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1666464484
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1666464484
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1666464484
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1666464484
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1666464484
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1666464484
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1666464484
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1666464484
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1666464484
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1666464484
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1666464484
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1666464484
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1666464484
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1666464484
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1666464484
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1666464484
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_253
timestamp 1666464484
transform 1 0 24380 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_261
timestamp 1666464484
transform 1 0 25116 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_267
timestamp 1666464484
transform 1 0 25668 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_273
timestamp 1666464484
transform 1 0 26220 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_279
timestamp 1666464484
transform 1 0 26772 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_285
timestamp 1666464484
transform 1 0 27324 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_291
timestamp 1666464484
transform 1 0 27876 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_297
timestamp 1666464484
transform 1 0 28428 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_303
timestamp 1666464484
transform 1 0 28980 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_306
timestamp 1666464484
transform 1 0 29256 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_309
timestamp 1666464484
transform 1 0 29532 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_318
timestamp 1666464484
transform 1 0 30360 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_324
timestamp 1666464484
transform 1 0 30912 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_330
timestamp 1666464484
transform 1 0 31464 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_336
timestamp 1666464484
transform 1 0 32016 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_340
timestamp 1666464484
transform 1 0 32384 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_349
timestamp 1666464484
transform 1 0 33212 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_358
timestamp 1666464484
transform 1 0 34040 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_365
timestamp 1666464484
transform 1 0 34684 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_369
timestamp 1666464484
transform 1 0 35052 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_375
timestamp 1666464484
transform 1 0 35604 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_387
timestamp 1666464484
transform 1 0 36708 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_399
timestamp 1666464484
transform 1 0 37812 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_411
timestamp 1666464484
transform 1 0 38916 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1666464484
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1666464484
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1666464484
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1666464484
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1666464484
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1666464484
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1666464484
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1666464484
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1666464484
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1666464484
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1666464484
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1666464484
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1666464484
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1666464484
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_545
timestamp 1666464484
transform 1 0 51244 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_549
timestamp 1666464484
transform 1 0 51612 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_552
timestamp 1666464484
transform 1 0 51888 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_558
timestamp 1666464484
transform 1 0 52440 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_565
timestamp 1666464484
transform 1 0 53084 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_579
timestamp 1666464484
transform 1 0 54372 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1666464484
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_15
timestamp 1666464484
transform 1 0 2484 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_21
timestamp 1666464484
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_33
timestamp 1666464484
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1666464484
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1666464484
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1666464484
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1666464484
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1666464484
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1666464484
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1666464484
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1666464484
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1666464484
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1666464484
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1666464484
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1666464484
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1666464484
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1666464484
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1666464484
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1666464484
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1666464484
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1666464484
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1666464484
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1666464484
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1666464484
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1666464484
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1666464484
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_261
timestamp 1666464484
transform 1 0 25116 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_266
timestamp 1666464484
transform 1 0 25576 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_272
timestamp 1666464484
transform 1 0 26128 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_278
timestamp 1666464484
transform 1 0 26680 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_281
timestamp 1666464484
transform 1 0 26956 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_289
timestamp 1666464484
transform 1 0 27692 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_293
timestamp 1666464484
transform 1 0 28060 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_296
timestamp 1666464484
transform 1 0 28336 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_306
timestamp 1666464484
transform 1 0 29256 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_312
timestamp 1666464484
transform 1 0 29808 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_318
timestamp 1666464484
transform 1 0 30360 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_324
timestamp 1666464484
transform 1 0 30912 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_330
timestamp 1666464484
transform 1 0 31464 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1666464484
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_341
timestamp 1666464484
transform 1 0 32476 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_347
timestamp 1666464484
transform 1 0 33028 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_353
timestamp 1666464484
transform 1 0 33580 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_359
timestamp 1666464484
transform 1 0 34132 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_365
timestamp 1666464484
transform 1 0 34684 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_371
timestamp 1666464484
transform 1 0 35236 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_383
timestamp 1666464484
transform 1 0 36340 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1666464484
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1666464484
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1666464484
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1666464484
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1666464484
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1666464484
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1666464484
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1666464484
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1666464484
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1666464484
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1666464484
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1666464484
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1666464484
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1666464484
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1666464484
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1666464484
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1666464484
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_553
timestamp 1666464484
transform 1 0 51980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_558
timestamp 1666464484
transform 1 0 52440 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_561
timestamp 1666464484
transform 1 0 52716 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_565
timestamp 1666464484
transform 1 0 53084 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_579
timestamp 1666464484
transform 1 0 54372 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1666464484
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_15
timestamp 1666464484
transform 1 0 2484 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_21
timestamp 1666464484
transform 1 0 3036 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1666464484
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1666464484
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1666464484
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1666464484
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1666464484
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1666464484
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1666464484
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1666464484
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1666464484
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1666464484
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1666464484
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1666464484
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1666464484
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1666464484
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1666464484
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1666464484
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1666464484
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1666464484
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1666464484
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1666464484
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1666464484
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1666464484
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1666464484
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1666464484
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1666464484
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1666464484
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_265
timestamp 1666464484
transform 1 0 25484 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_269
timestamp 1666464484
transform 1 0 25852 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_272
timestamp 1666464484
transform 1 0 26128 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_278
timestamp 1666464484
transform 1 0 26680 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_290
timestamp 1666464484
transform 1 0 27784 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_296
timestamp 1666464484
transform 1 0 28336 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_299
timestamp 1666464484
transform 1 0 28612 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_305
timestamp 1666464484
transform 1 0 29164 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_309
timestamp 1666464484
transform 1 0 29532 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_313
timestamp 1666464484
transform 1 0 29900 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_319
timestamp 1666464484
transform 1 0 30452 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_325
timestamp 1666464484
transform 1 0 31004 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_331
timestamp 1666464484
transform 1 0 31556 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_337
timestamp 1666464484
transform 1 0 32108 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_343
timestamp 1666464484
transform 1 0 32660 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_349
timestamp 1666464484
transform 1 0 33212 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_355
timestamp 1666464484
transform 1 0 33764 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_361
timestamp 1666464484
transform 1 0 34316 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1666464484
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1666464484
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1666464484
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1666464484
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1666464484
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1666464484
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1666464484
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1666464484
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1666464484
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1666464484
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1666464484
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1666464484
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1666464484
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1666464484
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1666464484
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1666464484
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1666464484
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1666464484
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1666464484
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_545
timestamp 1666464484
transform 1 0 51244 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_551
timestamp 1666464484
transform 1 0 51796 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_557
timestamp 1666464484
transform 1 0 52348 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_565
timestamp 1666464484
transform 1 0 53084 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_579
timestamp 1666464484
transform 1 0 54372 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1666464484
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_15
timestamp 1666464484
transform 1 0 2484 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_21
timestamp 1666464484
transform 1 0 3036 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_33
timestamp 1666464484
transform 1 0 4140 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_45
timestamp 1666464484
transform 1 0 5244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1666464484
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1666464484
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1666464484
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1666464484
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1666464484
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1666464484
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1666464484
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1666464484
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1666464484
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1666464484
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1666464484
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1666464484
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1666464484
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1666464484
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1666464484
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1666464484
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1666464484
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1666464484
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1666464484
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1666464484
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1666464484
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1666464484
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_261
timestamp 1666464484
transform 1 0 25116 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_266
timestamp 1666464484
transform 1 0 25576 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_77_277
timestamp 1666464484
transform 1 0 26588 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_281
timestamp 1666464484
transform 1 0 26956 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_285
timestamp 1666464484
transform 1 0 27324 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_291
timestamp 1666464484
transform 1 0 27876 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_294
timestamp 1666464484
transform 1 0 28152 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_300
timestamp 1666464484
transform 1 0 28704 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_312
timestamp 1666464484
transform 1 0 29808 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_320
timestamp 1666464484
transform 1 0 30544 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_326
timestamp 1666464484
transform 1 0 31096 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_334
timestamp 1666464484
transform 1 0 31832 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_337
timestamp 1666464484
transform 1 0 32108 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_341
timestamp 1666464484
transform 1 0 32476 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_347
timestamp 1666464484
transform 1 0 33028 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_359
timestamp 1666464484
transform 1 0 34132 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_371
timestamp 1666464484
transform 1 0 35236 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_383
timestamp 1666464484
transform 1 0 36340 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1666464484
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1666464484
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1666464484
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1666464484
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1666464484
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1666464484
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1666464484
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1666464484
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1666464484
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1666464484
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1666464484
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1666464484
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1666464484
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1666464484
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1666464484
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1666464484
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_541
timestamp 1666464484
transform 1 0 50876 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_544
timestamp 1666464484
transform 1 0 51152 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_558
timestamp 1666464484
transform 1 0 52440 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_561
timestamp 1666464484
transform 1 0 52716 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_565
timestamp 1666464484
transform 1 0 53084 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_579
timestamp 1666464484
transform 1 0 54372 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1666464484
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_15
timestamp 1666464484
transform 1 0 2484 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_21
timestamp 1666464484
transform 1 0 3036 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1666464484
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1666464484
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1666464484
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1666464484
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1666464484
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1666464484
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1666464484
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1666464484
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1666464484
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1666464484
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1666464484
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1666464484
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1666464484
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1666464484
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1666464484
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1666464484
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1666464484
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1666464484
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1666464484
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1666464484
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1666464484
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1666464484
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1666464484
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1666464484
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1666464484
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1666464484
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1666464484
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_277
timestamp 1666464484
transform 1 0 26588 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_281
timestamp 1666464484
transform 1 0 26956 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_287
timestamp 1666464484
transform 1 0 27508 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_291
timestamp 1666464484
transform 1 0 27876 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_294
timestamp 1666464484
transform 1 0 28152 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_306
timestamp 1666464484
transform 1 0 29256 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1666464484
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1666464484
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1666464484
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1666464484
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1666464484
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1666464484
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1666464484
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1666464484
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1666464484
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1666464484
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1666464484
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1666464484
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1666464484
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1666464484
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1666464484
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1666464484
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1666464484
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1666464484
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1666464484
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1666464484
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1666464484
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1666464484
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1666464484
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1666464484
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_533
timestamp 1666464484
transform 1 0 50140 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_541
timestamp 1666464484
transform 1 0 50876 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_545
timestamp 1666464484
transform 1 0 51244 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_551
timestamp 1666464484
transform 1 0 51796 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_565
timestamp 1666464484
transform 1 0 53084 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_579
timestamp 1666464484
transform 1 0 54372 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1666464484
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_15
timestamp 1666464484
transform 1 0 2484 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_21
timestamp 1666464484
transform 1 0 3036 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_33
timestamp 1666464484
transform 1 0 4140 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_45
timestamp 1666464484
transform 1 0 5244 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_53
timestamp 1666464484
transform 1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1666464484
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1666464484
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1666464484
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1666464484
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1666464484
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1666464484
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1666464484
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1666464484
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1666464484
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1666464484
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1666464484
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1666464484
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1666464484
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1666464484
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1666464484
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1666464484
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1666464484
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1666464484
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1666464484
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1666464484
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1666464484
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1666464484
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1666464484
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1666464484
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1666464484
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1666464484
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1666464484
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1666464484
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1666464484
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1666464484
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_337
timestamp 1666464484
transform 1 0 32108 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_341
timestamp 1666464484
transform 1 0 32476 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_347
timestamp 1666464484
transform 1 0 33028 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_353
timestamp 1666464484
transform 1 0 33580 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_365
timestamp 1666464484
transform 1 0 34684 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_377
timestamp 1666464484
transform 1 0 35788 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_389
timestamp 1666464484
transform 1 0 36892 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1666464484
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1666464484
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1666464484
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1666464484
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1666464484
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1666464484
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1666464484
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1666464484
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1666464484
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1666464484
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1666464484
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1666464484
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1666464484
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1666464484
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1666464484
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_541
timestamp 1666464484
transform 1 0 50876 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_544
timestamp 1666464484
transform 1 0 51152 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_558
timestamp 1666464484
transform 1 0 52440 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_561
timestamp 1666464484
transform 1 0 52716 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_565
timestamp 1666464484
transform 1 0 53084 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_579
timestamp 1666464484
transform 1 0 54372 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1666464484
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_15
timestamp 1666464484
transform 1 0 2484 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1666464484
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1666464484
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1666464484
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1666464484
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1666464484
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1666464484
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1666464484
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1666464484
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1666464484
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1666464484
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1666464484
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1666464484
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1666464484
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1666464484
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1666464484
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1666464484
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1666464484
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1666464484
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1666464484
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1666464484
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1666464484
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1666464484
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1666464484
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1666464484
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1666464484
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1666464484
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1666464484
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1666464484
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1666464484
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1666464484
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1666464484
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1666464484
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1666464484
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_321
timestamp 1666464484
transform 1 0 30636 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_327
timestamp 1666464484
transform 1 0 31188 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_330
timestamp 1666464484
transform 1 0 31464 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_336
timestamp 1666464484
transform 1 0 32016 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_347
timestamp 1666464484
transform 1 0 33028 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_353
timestamp 1666464484
transform 1 0 33580 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_359
timestamp 1666464484
transform 1 0 34132 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1666464484
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_365
timestamp 1666464484
transform 1 0 34684 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_369
timestamp 1666464484
transform 1 0 35052 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_381
timestamp 1666464484
transform 1 0 36156 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_393
timestamp 1666464484
transform 1 0 37260 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_405
timestamp 1666464484
transform 1 0 38364 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_417
timestamp 1666464484
transform 1 0 39468 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1666464484
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1666464484
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1666464484
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1666464484
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1666464484
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1666464484
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1666464484
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1666464484
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1666464484
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1666464484
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1666464484
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1666464484
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_533
timestamp 1666464484
transform 1 0 50140 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_541
timestamp 1666464484
transform 1 0 50876 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_545
timestamp 1666464484
transform 1 0 51244 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_551
timestamp 1666464484
transform 1 0 51796 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_565
timestamp 1666464484
transform 1 0 53084 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_579
timestamp 1666464484
transform 1 0 54372 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_3
timestamp 1666464484
transform 1 0 1380 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_15
timestamp 1666464484
transform 1 0 2484 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_21
timestamp 1666464484
transform 1 0 3036 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_33
timestamp 1666464484
transform 1 0 4140 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_45
timestamp 1666464484
transform 1 0 5244 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_53
timestamp 1666464484
transform 1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1666464484
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1666464484
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1666464484
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1666464484
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1666464484
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1666464484
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1666464484
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1666464484
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1666464484
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1666464484
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1666464484
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1666464484
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1666464484
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1666464484
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1666464484
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1666464484
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1666464484
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1666464484
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1666464484
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1666464484
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1666464484
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1666464484
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1666464484
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1666464484
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1666464484
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1666464484
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_305
timestamp 1666464484
transform 1 0 29164 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_310
timestamp 1666464484
transform 1 0 29624 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_318
timestamp 1666464484
transform 1 0 30360 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_321
timestamp 1666464484
transform 1 0 30636 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_325
timestamp 1666464484
transform 1 0 31004 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_328
timestamp 1666464484
transform 1 0 31280 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_334
timestamp 1666464484
transform 1 0 31832 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_337
timestamp 1666464484
transform 1 0 32108 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_346
timestamp 1666464484
transform 1 0 32936 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_354
timestamp 1666464484
transform 1 0 33672 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_362
timestamp 1666464484
transform 1 0 34408 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_368
timestamp 1666464484
transform 1 0 34960 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_374
timestamp 1666464484
transform 1 0 35512 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_386
timestamp 1666464484
transform 1 0 36616 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1666464484
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1666464484
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1666464484
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1666464484
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1666464484
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1666464484
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1666464484
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1666464484
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1666464484
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1666464484
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1666464484
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1666464484
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1666464484
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1666464484
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_529
timestamp 1666464484
transform 1 0 49772 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_535
timestamp 1666464484
transform 1 0 50324 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_538
timestamp 1666464484
transform 1 0 50600 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_544
timestamp 1666464484
transform 1 0 51152 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_558
timestamp 1666464484
transform 1 0 52440 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_561
timestamp 1666464484
transform 1 0 52716 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_565
timestamp 1666464484
transform 1 0 53084 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_579
timestamp 1666464484
transform 1 0 54372 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1666464484
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_15
timestamp 1666464484
transform 1 0 2484 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1666464484
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1666464484
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1666464484
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1666464484
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1666464484
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1666464484
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1666464484
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1666464484
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1666464484
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1666464484
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1666464484
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1666464484
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1666464484
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1666464484
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1666464484
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1666464484
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1666464484
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1666464484
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1666464484
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1666464484
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1666464484
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1666464484
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1666464484
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1666464484
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1666464484
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1666464484
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1666464484
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1666464484
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1666464484
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1666464484
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_301
timestamp 1666464484
transform 1 0 28796 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_306
timestamp 1666464484
transform 1 0 29256 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_309
timestamp 1666464484
transform 1 0 29532 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_319
timestamp 1666464484
transform 1 0 30452 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_331
timestamp 1666464484
transform 1 0 31556 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_343
timestamp 1666464484
transform 1 0 32660 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_347
timestamp 1666464484
transform 1 0 33028 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_356
timestamp 1666464484
transform 1 0 33856 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_362
timestamp 1666464484
transform 1 0 34408 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_365
timestamp 1666464484
transform 1 0 34684 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_369
timestamp 1666464484
transform 1 0 35052 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_375
timestamp 1666464484
transform 1 0 35604 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_387
timestamp 1666464484
transform 1 0 36708 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_399
timestamp 1666464484
transform 1 0 37812 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_411
timestamp 1666464484
transform 1 0 38916 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1666464484
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1666464484
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1666464484
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1666464484
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1666464484
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1666464484
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1666464484
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1666464484
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1666464484
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1666464484
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1666464484
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_525
timestamp 1666464484
transform 1 0 49404 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_530
timestamp 1666464484
transform 1 0 49864 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_533
timestamp 1666464484
transform 1 0 50140 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_537
timestamp 1666464484
transform 1 0 50508 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_543
timestamp 1666464484
transform 1 0 51060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_554
timestamp 1666464484
transform 1 0 52072 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_565
timestamp 1666464484
transform 1 0 53084 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_579
timestamp 1666464484
transform 1 0 54372 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_3
timestamp 1666464484
transform 1 0 1380 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_15
timestamp 1666464484
transform 1 0 2484 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_21
timestamp 1666464484
transform 1 0 3036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_33
timestamp 1666464484
transform 1 0 4140 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_45
timestamp 1666464484
transform 1 0 5244 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_53
timestamp 1666464484
transform 1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1666464484
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1666464484
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1666464484
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1666464484
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1666464484
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1666464484
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1666464484
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1666464484
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1666464484
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1666464484
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1666464484
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1666464484
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1666464484
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1666464484
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1666464484
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1666464484
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1666464484
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1666464484
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1666464484
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1666464484
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1666464484
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1666464484
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1666464484
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1666464484
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1666464484
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1666464484
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_305
timestamp 1666464484
transform 1 0 29164 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_309
timestamp 1666464484
transform 1 0 29532 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_312
timestamp 1666464484
transform 1 0 29808 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_320
timestamp 1666464484
transform 1 0 30544 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_323
timestamp 1666464484
transform 1 0 30820 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_333
timestamp 1666464484
transform 1 0 31740 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_83_337
timestamp 1666464484
transform 1 0 32108 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_83_341
timestamp 1666464484
transform 1 0 32476 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_355
timestamp 1666464484
transform 1 0 33764 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_366
timestamp 1666464484
transform 1 0 34776 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_372
timestamp 1666464484
transform 1 0 35328 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_378
timestamp 1666464484
transform 1 0 35880 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_384
timestamp 1666464484
transform 1 0 36432 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1666464484
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1666464484
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1666464484
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1666464484
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1666464484
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1666464484
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1666464484
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1666464484
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1666464484
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1666464484
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1666464484
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1666464484
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1666464484
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1666464484
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_529
timestamp 1666464484
transform 1 0 49772 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_534
timestamp 1666464484
transform 1 0 50232 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_540
timestamp 1666464484
transform 1 0 50784 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_547
timestamp 1666464484
transform 1 0 51428 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_558
timestamp 1666464484
transform 1 0 52440 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_561
timestamp 1666464484
transform 1 0 52716 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_565
timestamp 1666464484
transform 1 0 53084 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_579
timestamp 1666464484
transform 1 0 54372 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1666464484
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_15
timestamp 1666464484
transform 1 0 2484 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_21
timestamp 1666464484
transform 1 0 3036 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1666464484
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1666464484
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1666464484
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1666464484
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1666464484
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1666464484
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1666464484
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1666464484
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1666464484
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1666464484
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1666464484
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1666464484
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1666464484
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1666464484
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1666464484
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1666464484
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1666464484
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1666464484
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1666464484
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1666464484
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1666464484
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1666464484
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1666464484
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1666464484
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1666464484
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1666464484
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1666464484
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1666464484
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1666464484
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1666464484
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1666464484
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1666464484
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1666464484
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_335
timestamp 1666464484
transform 1 0 31924 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_341
timestamp 1666464484
transform 1 0 32476 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_355
timestamp 1666464484
transform 1 0 33764 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_84_361
timestamp 1666464484
transform 1 0 34316 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_84_365
timestamp 1666464484
transform 1 0 34684 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_369
timestamp 1666464484
transform 1 0 35052 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_375
timestamp 1666464484
transform 1 0 35604 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_387
timestamp 1666464484
transform 1 0 36708 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_399
timestamp 1666464484
transform 1 0 37812 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_411
timestamp 1666464484
transform 1 0 38916 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1666464484
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1666464484
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1666464484
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1666464484
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1666464484
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1666464484
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1666464484
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1666464484
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1666464484
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1666464484
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1666464484
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1666464484
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1666464484
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_533
timestamp 1666464484
transform 1 0 50140 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_543
timestamp 1666464484
transform 1 0 51060 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_549
timestamp 1666464484
transform 1 0 51612 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_556
timestamp 1666464484
transform 1 0 52256 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_563
timestamp 1666464484
transform 1 0 52900 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_574
timestamp 1666464484
transform 1 0 53912 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_580
timestamp 1666464484
transform 1 0 54464 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_3
timestamp 1666464484
transform 1 0 1380 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_15
timestamp 1666464484
transform 1 0 2484 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_21
timestamp 1666464484
transform 1 0 3036 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_33
timestamp 1666464484
transform 1 0 4140 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_45
timestamp 1666464484
transform 1 0 5244 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_53
timestamp 1666464484
transform 1 0 5980 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1666464484
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1666464484
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1666464484
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1666464484
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1666464484
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1666464484
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1666464484
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1666464484
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1666464484
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1666464484
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1666464484
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1666464484
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1666464484
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1666464484
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1666464484
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1666464484
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1666464484
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1666464484
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1666464484
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1666464484
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1666464484
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1666464484
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1666464484
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1666464484
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1666464484
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1666464484
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1666464484
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1666464484
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1666464484
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1666464484
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_337
timestamp 1666464484
transform 1 0 32108 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_345
timestamp 1666464484
transform 1 0 32844 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_351
timestamp 1666464484
transform 1 0 33396 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_357
timestamp 1666464484
transform 1 0 33948 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_363
timestamp 1666464484
transform 1 0 34500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_375
timestamp 1666464484
transform 1 0 35604 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_387
timestamp 1666464484
transform 1 0 36708 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1666464484
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1666464484
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1666464484
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1666464484
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1666464484
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1666464484
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1666464484
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1666464484
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1666464484
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1666464484
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1666464484
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1666464484
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1666464484
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1666464484
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1666464484
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1666464484
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_541
timestamp 1666464484
transform 1 0 50876 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_545
timestamp 1666464484
transform 1 0 51244 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_551
timestamp 1666464484
transform 1 0 51796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_558
timestamp 1666464484
transform 1 0 52440 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_561
timestamp 1666464484
transform 1 0 52716 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_565
timestamp 1666464484
transform 1 0 53084 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_579
timestamp 1666464484
transform 1 0 54372 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1666464484
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_15
timestamp 1666464484
transform 1 0 2484 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1666464484
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1666464484
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1666464484
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1666464484
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1666464484
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1666464484
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1666464484
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1666464484
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1666464484
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1666464484
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1666464484
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1666464484
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1666464484
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1666464484
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1666464484
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1666464484
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1666464484
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1666464484
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1666464484
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1666464484
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1666464484
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1666464484
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1666464484
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1666464484
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1666464484
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1666464484
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1666464484
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1666464484
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1666464484
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1666464484
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1666464484
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1666464484
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1666464484
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1666464484
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_333
timestamp 1666464484
transform 1 0 31740 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_341
timestamp 1666464484
transform 1 0 32476 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_345
timestamp 1666464484
transform 1 0 32844 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_351
timestamp 1666464484
transform 1 0 33396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1666464484
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1666464484
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1666464484
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1666464484
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1666464484
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1666464484
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1666464484
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1666464484
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1666464484
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1666464484
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1666464484
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1666464484
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1666464484
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1666464484
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1666464484
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1666464484
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1666464484
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1666464484
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1666464484
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1666464484
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_545
timestamp 1666464484
transform 1 0 51244 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_549
timestamp 1666464484
transform 1 0 51612 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_552
timestamp 1666464484
transform 1 0 51888 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_558
timestamp 1666464484
transform 1 0 52440 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_565
timestamp 1666464484
transform 1 0 53084 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_579
timestamp 1666464484
transform 1 0 54372 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_3
timestamp 1666464484
transform 1 0 1380 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_9
timestamp 1666464484
transform 1 0 1932 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1666464484
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1666464484
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1666464484
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1666464484
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1666464484
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1666464484
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1666464484
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1666464484
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1666464484
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1666464484
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1666464484
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1666464484
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1666464484
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1666464484
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1666464484
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1666464484
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1666464484
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1666464484
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1666464484
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1666464484
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1666464484
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1666464484
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1666464484
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1666464484
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1666464484
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1666464484
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1666464484
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1666464484
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1666464484
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1666464484
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1666464484
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1666464484
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1666464484
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1666464484
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1666464484
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1666464484
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1666464484
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1666464484
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1666464484
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1666464484
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1666464484
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1666464484
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1666464484
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1666464484
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1666464484
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1666464484
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1666464484
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1666464484
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1666464484
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1666464484
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1666464484
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1666464484
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1666464484
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1666464484
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1666464484
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1666464484
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1666464484
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_553
timestamp 1666464484
transform 1 0 51980 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_87_558
timestamp 1666464484
transform 1 0 52440 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_561
timestamp 1666464484
transform 1 0 52716 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_565
timestamp 1666464484
transform 1 0 53084 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_572
timestamp 1666464484
transform 1 0 53728 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_579
timestamp 1666464484
transform 1 0 54372 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_3
timestamp 1666464484
transform 1 0 1380 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_15
timestamp 1666464484
transform 1 0 2484 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_88_21
timestamp 1666464484
transform 1 0 3036 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1666464484
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1666464484
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1666464484
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1666464484
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1666464484
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1666464484
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1666464484
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1666464484
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1666464484
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1666464484
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1666464484
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1666464484
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1666464484
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1666464484
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1666464484
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1666464484
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1666464484
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1666464484
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1666464484
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1666464484
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1666464484
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1666464484
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1666464484
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1666464484
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1666464484
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1666464484
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1666464484
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1666464484
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1666464484
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1666464484
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1666464484
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1666464484
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1666464484
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1666464484
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1666464484
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1666464484
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1666464484
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1666464484
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1666464484
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1666464484
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1666464484
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1666464484
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1666464484
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1666464484
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1666464484
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1666464484
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1666464484
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1666464484
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1666464484
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1666464484
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1666464484
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1666464484
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1666464484
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1666464484
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1666464484
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1666464484
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1666464484
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_557
timestamp 1666464484
transform 1 0 52348 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_561
timestamp 1666464484
transform 1 0 52716 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_567
timestamp 1666464484
transform 1 0 53268 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_575
timestamp 1666464484
transform 1 0 54004 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_579
timestamp 1666464484
transform 1 0 54372 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1666464484
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_15
timestamp 1666464484
transform 1 0 2484 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_21
timestamp 1666464484
transform 1 0 3036 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_33
timestamp 1666464484
transform 1 0 4140 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_45
timestamp 1666464484
transform 1 0 5244 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_53
timestamp 1666464484
transform 1 0 5980 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1666464484
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1666464484
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1666464484
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1666464484
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1666464484
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1666464484
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1666464484
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1666464484
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1666464484
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1666464484
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1666464484
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1666464484
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1666464484
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1666464484
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1666464484
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1666464484
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1666464484
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1666464484
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1666464484
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1666464484
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1666464484
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1666464484
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1666464484
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1666464484
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1666464484
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1666464484
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1666464484
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1666464484
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1666464484
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1666464484
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1666464484
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1666464484
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1666464484
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1666464484
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1666464484
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1666464484
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1666464484
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1666464484
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1666464484
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1666464484
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1666464484
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1666464484
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1666464484
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1666464484
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1666464484
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1666464484
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1666464484
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1666464484
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1666464484
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1666464484
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1666464484
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1666464484
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1666464484
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1666464484
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_561
timestamp 1666464484
transform 1 0 52716 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_569
timestamp 1666464484
transform 1 0 53452 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_572
timestamp 1666464484
transform 1 0 53728 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_579
timestamp 1666464484
transform 1 0 54372 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_3
timestamp 1666464484
transform 1 0 1380 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_9
timestamp 1666464484
transform 1 0 1932 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_15
timestamp 1666464484
transform 1 0 2484 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_21
timestamp 1666464484
transform 1 0 3036 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1666464484
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1666464484
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1666464484
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1666464484
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1666464484
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1666464484
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1666464484
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1666464484
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1666464484
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1666464484
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1666464484
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1666464484
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1666464484
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1666464484
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1666464484
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1666464484
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1666464484
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1666464484
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1666464484
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1666464484
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1666464484
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1666464484
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1666464484
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1666464484
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1666464484
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1666464484
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_265
timestamp 1666464484
transform 1 0 25484 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_269
timestamp 1666464484
transform 1 0 25852 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_272
timestamp 1666464484
transform 1 0 26128 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_284
timestamp 1666464484
transform 1 0 27232 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_287
timestamp 1666464484
transform 1 0 27508 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_299
timestamp 1666464484
transform 1 0 28612 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1666464484
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1666464484
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1666464484
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1666464484
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1666464484
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1666464484
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1666464484
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1666464484
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1666464484
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1666464484
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1666464484
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1666464484
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1666464484
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1666464484
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1666464484
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1666464484
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1666464484
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1666464484
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1666464484
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1666464484
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1666464484
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1666464484
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1666464484
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1666464484
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1666464484
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1666464484
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1666464484
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1666464484
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_569
timestamp 1666464484
transform 1 0 53452 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_573
timestamp 1666464484
transform 1 0 53820 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_579
timestamp 1666464484
transform 1 0 54372 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1666464484
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_9
timestamp 1666464484
transform 1 0 1932 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_15
timestamp 1666464484
transform 1 0 2484 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_21
timestamp 1666464484
transform 1 0 3036 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1666464484
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1666464484
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1666464484
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1666464484
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1666464484
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1666464484
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1666464484
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1666464484
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1666464484
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1666464484
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1666464484
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1666464484
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1666464484
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1666464484
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1666464484
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1666464484
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1666464484
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1666464484
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1666464484
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1666464484
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1666464484
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1666464484
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1666464484
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1666464484
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_249
timestamp 1666464484
transform 1 0 24012 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_91_257
timestamp 1666464484
transform 1 0 24748 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_268
timestamp 1666464484
transform 1 0 25760 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_278
timestamp 1666464484
transform 1 0 26680 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_91_281
timestamp 1666464484
transform 1 0 26956 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_294
timestamp 1666464484
transform 1 0 28152 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_306
timestamp 1666464484
transform 1 0 29256 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_318
timestamp 1666464484
transform 1 0 30360 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_330
timestamp 1666464484
transform 1 0 31464 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1666464484
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1666464484
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1666464484
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1666464484
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1666464484
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1666464484
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1666464484
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1666464484
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1666464484
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1666464484
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1666464484
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1666464484
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1666464484
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1666464484
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1666464484
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_485
timestamp 1666464484
transform 1 0 45724 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_488
timestamp 1666464484
transform 1 0 46000 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_500
timestamp 1666464484
transform 1 0 47104 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1666464484
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1666464484
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1666464484
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_541
timestamp 1666464484
transform 1 0 50876 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_91_549
timestamp 1666464484
transform 1 0 51612 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_557
timestamp 1666464484
transform 1 0 52348 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1666464484
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_573
timestamp 1666464484
transform 1 0 53820 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_579
timestamp 1666464484
transform 1 0 54372 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1666464484
transform 1 0 1380 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_9
timestamp 1666464484
transform 1 0 1932 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_17
timestamp 1666464484
transform 1 0 2668 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_23
timestamp 1666464484
transform 1 0 3220 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1666464484
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_29
timestamp 1666464484
transform 1 0 3772 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_33
timestamp 1666464484
transform 1 0 4140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_45
timestamp 1666464484
transform 1 0 5244 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_59
timestamp 1666464484
transform 1 0 6532 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_67
timestamp 1666464484
transform 1 0 7268 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_72
timestamp 1666464484
transform 1 0 7728 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_85
timestamp 1666464484
transform 1 0 8924 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_93
timestamp 1666464484
transform 1 0 9660 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_92_98
timestamp 1666464484
transform 1 0 10120 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_104
timestamp 1666464484
transform 1 0 10672 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_107
timestamp 1666464484
transform 1 0 10948 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1666464484
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_133
timestamp 1666464484
transform 1 0 13340 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_92_138
timestamp 1666464484
transform 1 0 13800 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_141
timestamp 1666464484
transform 1 0 14076 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_92_146
timestamp 1666464484
transform 1 0 14536 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_154
timestamp 1666464484
transform 1 0 15272 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_166
timestamp 1666464484
transform 1 0 16376 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_172
timestamp 1666464484
transform 1 0 16928 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_92_186
timestamp 1666464484
transform 1 0 18216 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_92_194
timestamp 1666464484
transform 1 0 18952 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_92_197
timestamp 1666464484
transform 1 0 19228 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_202
timestamp 1666464484
transform 1 0 19688 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_214
timestamp 1666464484
transform 1 0 20792 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_228
timestamp 1666464484
transform 1 0 22080 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_240
timestamp 1666464484
transform 1 0 23184 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1666464484
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_265
timestamp 1666464484
transform 1 0 25484 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_270
timestamp 1666464484
transform 1 0 25944 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_92_276
timestamp 1666464484
transform 1 0 26496 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_282
timestamp 1666464484
transform 1 0 27048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_285
timestamp 1666464484
transform 1 0 27324 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_293
timestamp 1666464484
transform 1 0 28060 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_305
timestamp 1666464484
transform 1 0 29164 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1666464484
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1666464484
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_333
timestamp 1666464484
transform 1 0 31740 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_341
timestamp 1666464484
transform 1 0 32476 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_92_346
timestamp 1666464484
transform 1 0 32936 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_354
timestamp 1666464484
transform 1 0 33672 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_92_358
timestamp 1666464484
transform 1 0 34040 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1666464484
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_377
timestamp 1666464484
transform 1 0 35788 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_381
timestamp 1666464484
transform 1 0 36156 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_384
timestamp 1666464484
transform 1 0 36432 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_396
timestamp 1666464484
transform 1 0 37536 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_410
timestamp 1666464484
transform 1 0 38824 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_418
timestamp 1666464484
transform 1 0 39560 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1666464484
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1666464484
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_445
timestamp 1666464484
transform 1 0 42044 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_451
timestamp 1666464484
transform 1 0 42596 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_459
timestamp 1666464484
transform 1 0 43332 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_462
timestamp 1666464484
transform 1 0 43608 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_474
timestamp 1666464484
transform 1 0 44712 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_477
timestamp 1666464484
transform 1 0 44988 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_92_481
timestamp 1666464484
transform 1 0 45356 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_487
timestamp 1666464484
transform 1 0 45908 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_498
timestamp 1666464484
transform 1 0 46920 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_506
timestamp 1666464484
transform 1 0 47656 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_510
timestamp 1666464484
transform 1 0 48024 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_524
timestamp 1666464484
transform 1 0 49312 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1666464484
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_545
timestamp 1666464484
transform 1 0 51244 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_549
timestamp 1666464484
transform 1 0 51612 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_92_557
timestamp 1666464484
transform 1 0 52348 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_563
timestamp 1666464484
transform 1 0 52900 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_566
timestamp 1666464484
transform 1 0 53176 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_574
timestamp 1666464484
transform 1 0 53912 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_579
timestamp 1666464484
transform 1 0 54372 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_3
timestamp 1666464484
transform 1 0 1380 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_17
timestamp 1666464484
transform 1 0 2668 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_93_25
timestamp 1666464484
transform 1 0 3404 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_29
timestamp 1666464484
transform 1 0 3772 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_36
timestamp 1666464484
transform 1 0 4416 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_42
timestamp 1666464484
transform 1 0 4968 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_93_50
timestamp 1666464484
transform 1 0 5704 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_93_57
timestamp 1666464484
transform 1 0 6348 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_63
timestamp 1666464484
transform 1 0 6900 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_71
timestamp 1666464484
transform 1 0 7636 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_75
timestamp 1666464484
transform 1 0 8004 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_79
timestamp 1666464484
transform 1 0 8372 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_82
timestamp 1666464484
transform 1 0 8648 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_85
timestamp 1666464484
transform 1 0 8924 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_90
timestamp 1666464484
transform 1 0 9384 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_108
timestamp 1666464484
transform 1 0 11040 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_113
timestamp 1666464484
transform 1 0 11500 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_117
timestamp 1666464484
transform 1 0 11868 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_120
timestamp 1666464484
transform 1 0 12144 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_93_134
timestamp 1666464484
transform 1 0 13432 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_93_141
timestamp 1666464484
transform 1 0 14076 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_152
timestamp 1666464484
transform 1 0 15088 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_166
timestamp 1666464484
transform 1 0 16376 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_169
timestamp 1666464484
transform 1 0 16652 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_173
timestamp 1666464484
transform 1 0 17020 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_181
timestamp 1666464484
transform 1 0 17756 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_194
timestamp 1666464484
transform 1 0 18952 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_197
timestamp 1666464484
transform 1 0 19228 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_201
timestamp 1666464484
transform 1 0 19596 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_205
timestamp 1666464484
transform 1 0 19964 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_211
timestamp 1666464484
transform 1 0 20516 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_93_218
timestamp 1666464484
transform 1 0 21160 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_93_225
timestamp 1666464484
transform 1 0 21804 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_231
timestamp 1666464484
transform 1 0 22356 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_237
timestamp 1666464484
transform 1 0 22908 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_244
timestamp 1666464484
transform 1 0 23552 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_250
timestamp 1666464484
transform 1 0 24104 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_253
timestamp 1666464484
transform 1 0 24380 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_258
timestamp 1666464484
transform 1 0 24840 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_266
timestamp 1666464484
transform 1 0 25576 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_93_270
timestamp 1666464484
transform 1 0 25944 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_93_278
timestamp 1666464484
transform 1 0 26680 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_281
timestamp 1666464484
transform 1 0 26956 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_286
timestamp 1666464484
transform 1 0 27416 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_292
timestamp 1666464484
transform 1 0 27968 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_296
timestamp 1666464484
transform 1 0 28336 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_306
timestamp 1666464484
transform 1 0 29256 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_309
timestamp 1666464484
transform 1 0 29532 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_314
timestamp 1666464484
transform 1 0 29992 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_318
timestamp 1666464484
transform 1 0 30360 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_322
timestamp 1666464484
transform 1 0 30728 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_328
timestamp 1666464484
transform 1 0 31280 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_334
timestamp 1666464484
transform 1 0 31832 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_337
timestamp 1666464484
transform 1 0 32108 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_342
timestamp 1666464484
transform 1 0 32568 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_349
timestamp 1666464484
transform 1 0 33212 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_357
timestamp 1666464484
transform 1 0 33948 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_93_361
timestamp 1666464484
transform 1 0 34316 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_93_365
timestamp 1666464484
transform 1 0 34684 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_374
timestamp 1666464484
transform 1 0 35512 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_380
timestamp 1666464484
transform 1 0 36064 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_387
timestamp 1666464484
transform 1 0 36708 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1666464484
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_393
timestamp 1666464484
transform 1 0 37260 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_400
timestamp 1666464484
transform 1 0 37904 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_406
timestamp 1666464484
transform 1 0 38456 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_93_413
timestamp 1666464484
transform 1 0 39100 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_419
timestamp 1666464484
transform 1 0 39652 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_421
timestamp 1666464484
transform 1 0 39836 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_426
timestamp 1666464484
transform 1 0 40296 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_432
timestamp 1666464484
transform 1 0 40848 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_439
timestamp 1666464484
transform 1 0 41492 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_93_445
timestamp 1666464484
transform 1 0 42044 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_449
timestamp 1666464484
transform 1 0 42412 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_454
timestamp 1666464484
transform 1 0 42872 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_472
timestamp 1666464484
transform 1 0 44528 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_477
timestamp 1666464484
transform 1 0 44988 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_489
timestamp 1666464484
transform 1 0 46092 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_497
timestamp 1666464484
transform 1 0 46828 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_502
timestamp 1666464484
transform 1 0 47288 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_505
timestamp 1666464484
transform 1 0 47564 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_517
timestamp 1666464484
transform 1 0 48668 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_525
timestamp 1666464484
transform 1 0 49404 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_530
timestamp 1666464484
transform 1 0 49864 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_533
timestamp 1666464484
transform 1 0 50140 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_545
timestamp 1666464484
transform 1 0 51244 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1666464484
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1666464484
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_561
timestamp 1666464484
transform 1 0 52716 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_565
timestamp 1666464484
transform 1 0 53084 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_576
timestamp 1666464484
transform 1 0 54096 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_580
timestamp 1666464484
transform 1 0 54464 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 54832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 54832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 54832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 54832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 54832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 54832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 54832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 54832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 54832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 54832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 54832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 54832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 54832 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 54832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 54832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 54832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 54832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 54832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 54832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 54832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 54832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 54832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 54832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 54832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 54832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 54832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 54832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 54832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 54832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 54832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 54832 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 54832 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 54832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 54832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 54832 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 54832 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 54832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 54832 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 54832 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 54832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 54832 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 54832 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 54832 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 54832 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 54832 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 54832 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 54832 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 54832 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 54832 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 54832 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 54832 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 54832 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 54832 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 54832 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 54832 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 54832 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 54832 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 54832 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 54832 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 54832 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 54832 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 54832 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 54832 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 54832 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 54832 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666464484
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666464484
transform -1 0 54832 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666464484
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666464484
transform -1 0 54832 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666464484
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666464484
transform -1 0 54832 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666464484
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666464484
transform -1 0 54832 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666464484
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666464484
transform -1 0 54832 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666464484
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666464484
transform -1 0 54832 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666464484
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666464484
transform -1 0 54832 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666464484
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666464484
transform -1 0 54832 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666464484
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666464484
transform -1 0 54832 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666464484
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666464484
transform -1 0 54832 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666464484
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666464484
transform -1 0 54832 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666464484
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666464484
transform -1 0 54832 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666464484
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666464484
transform -1 0 54832 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666464484
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666464484
transform -1 0 54832 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666464484
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666464484
transform -1 0 54832 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666464484
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666464484
transform -1 0 54832 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666464484
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666464484
transform -1 0 54832 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666464484
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666464484
transform -1 0 54832 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1666464484
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1666464484
transform -1 0 54832 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1666464484
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1666464484
transform -1 0 54832 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1666464484
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1666464484
transform -1 0 54832 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1666464484
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1666464484
transform -1 0 54832 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1666464484
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1666464484
transform -1 0 54832 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1666464484
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1666464484
transform -1 0 54832 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1666464484
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1666464484
transform -1 0 54832 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1666464484
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1666464484
transform -1 0 54832 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1666464484
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1666464484
transform -1 0 54832 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1666464484
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1666464484
transform -1 0 54832 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1666464484
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1666464484
transform -1 0 54832 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666464484
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666464484
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666464484
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666464484
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666464484
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666464484
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666464484
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666464484
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666464484
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666464484
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666464484
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666464484
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666464484
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666464484
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666464484
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666464484
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666464484
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666464484
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666464484
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666464484
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666464484
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666464484
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666464484
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666464484
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666464484
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666464484
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666464484
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666464484
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666464484
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666464484
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666464484
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666464484
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666464484
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666464484
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666464484
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666464484
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666464484
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666464484
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666464484
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666464484
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666464484
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666464484
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666464484
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666464484
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666464484
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666464484
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666464484
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666464484
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666464484
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666464484
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666464484
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666464484
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666464484
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666464484
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666464484
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666464484
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666464484
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666464484
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666464484
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666464484
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666464484
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666464484
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666464484
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666464484
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666464484
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666464484
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666464484
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666464484
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666464484
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666464484
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666464484
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666464484
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666464484
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666464484
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666464484
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666464484
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666464484
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666464484
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666464484
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666464484
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666464484
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666464484
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666464484
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666464484
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666464484
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666464484
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666464484
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666464484
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666464484
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666464484
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666464484
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666464484
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666464484
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666464484
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666464484
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666464484
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666464484
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666464484
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666464484
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666464484
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666464484
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666464484
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666464484
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666464484
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666464484
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666464484
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666464484
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666464484
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666464484
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666464484
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666464484
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666464484
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666464484
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666464484
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666464484
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666464484
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666464484
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666464484
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666464484
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666464484
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666464484
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666464484
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666464484
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666464484
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666464484
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666464484
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666464484
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666464484
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666464484
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666464484
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666464484
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666464484
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666464484
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666464484
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666464484
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666464484
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666464484
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666464484
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666464484
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666464484
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666464484
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666464484
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666464484
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666464484
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666464484
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666464484
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666464484
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666464484
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666464484
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666464484
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666464484
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666464484
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666464484
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666464484
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666464484
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666464484
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666464484
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666464484
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666464484
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666464484
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666464484
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666464484
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666464484
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666464484
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666464484
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666464484
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666464484
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666464484
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666464484
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666464484
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666464484
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666464484
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666464484
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666464484
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666464484
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666464484
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666464484
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666464484
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666464484
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666464484
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666464484
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666464484
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666464484
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666464484
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666464484
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666464484
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666464484
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666464484
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666464484
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666464484
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666464484
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666464484
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666464484
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666464484
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666464484
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666464484
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666464484
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666464484
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666464484
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666464484
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666464484
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666464484
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666464484
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666464484
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666464484
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666464484
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666464484
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666464484
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666464484
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666464484
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666464484
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666464484
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666464484
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666464484
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666464484
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666464484
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666464484
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666464484
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666464484
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666464484
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666464484
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666464484
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666464484
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666464484
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666464484
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1666464484
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1666464484
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1666464484
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1666464484
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1666464484
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1666464484
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1666464484
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1666464484
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1666464484
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1666464484
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1666464484
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1666464484
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1666464484
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1666464484
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1666464484
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1666464484
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1666464484
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1666464484
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1666464484
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1666464484
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1666464484
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1666464484
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1666464484
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1666464484
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1666464484
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1666464484
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1666464484
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1666464484
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1666464484
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1666464484
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1666464484
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1666464484
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1666464484
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1666464484
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1666464484
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1666464484
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1666464484
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1666464484
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1666464484
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1666464484
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1666464484
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1666464484
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1666464484
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1666464484
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1666464484
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1666464484
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1666464484
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1666464484
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1666464484
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1666464484
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1666464484
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1666464484
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1666464484
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1666464484
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1666464484
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1666464484
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1666464484
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1666464484
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1666464484
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1666464484
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1666464484
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1666464484
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1666464484
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1666464484
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1666464484
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1666464484
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1666464484
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1666464484
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1666464484
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1666464484
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1666464484
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1666464484
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1666464484
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1666464484
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1666464484
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1666464484
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1666464484
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1666464484
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1666464484
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1666464484
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1666464484
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1666464484
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1666464484
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1666464484
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1666464484
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1666464484
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1666464484
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1666464484
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1666464484
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1666464484
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1666464484
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1666464484
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1666464484
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1666464484
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1666464484
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1666464484
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1666464484
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1666464484
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1666464484
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1666464484
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1666464484
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1666464484
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1666464484
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1666464484
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1666464484
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1666464484
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1666464484
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1666464484
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1666464484
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1666464484
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1666464484
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1666464484
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1666464484
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1666464484
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1666464484
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1666464484
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1666464484
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1666464484
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1666464484
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1666464484
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1666464484
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1666464484
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1666464484
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1666464484
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1666464484
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1666464484
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1666464484
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1666464484
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1666464484
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1666464484
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1666464484
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1666464484
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1666464484
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1666464484
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1666464484
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1666464484
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1666464484
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1666464484
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1666464484
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1666464484
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1666464484
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1666464484
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1666464484
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1666464484
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1666464484
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1666464484
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1666464484
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1666464484
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1666464484
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1666464484
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1666464484
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1666464484
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1666464484
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1666464484
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1666464484
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1666464484
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1666464484
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1666464484
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1666464484
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1666464484
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1666464484
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1666464484
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1666464484
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1666464484
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1666464484
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1666464484
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1666464484
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1666464484
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1666464484
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1666464484
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1666464484
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1666464484
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1666464484
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1666464484
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1666464484
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1666464484
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1666464484
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1666464484
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1666464484
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1666464484
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1666464484
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1666464484
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1666464484
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1666464484
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1666464484
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1666464484
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1666464484
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1666464484
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1666464484
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1666464484
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1666464484
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1666464484
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1666464484
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1666464484
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1666464484
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1666464484
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1666464484
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1666464484
transform 1 0 3680 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1666464484
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1666464484
transform 1 0 8832 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1666464484
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1666464484
transform 1 0 13984 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1666464484
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1666464484
transform 1 0 19136 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1666464484
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1666464484
transform 1 0 24288 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1666464484
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1666464484
transform 1 0 29440 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1666464484
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1666464484
transform 1 0 34592 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1666464484
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1666464484
transform 1 0 39744 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1666464484
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1666464484
transform 1 0 44896 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1666464484
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1666464484
transform 1 0 50048 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1666464484
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _0574_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 25208 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _0575_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27692 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _0576_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27048 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0577_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28612 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0578_
timestamp 1666464484
transform -1 0 27692 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _0579_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26680 0 -1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _0580_
timestamp 1666464484
transform 1 0 32844 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0581_
timestamp 1666464484
transform 1 0 32292 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0582_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14536 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0583_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0584_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26220 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _0585_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 25668 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0586_
timestamp 1666464484
transform 1 0 27140 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0587_
timestamp 1666464484
transform -1 0 22540 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0588_
timestamp 1666464484
transform 1 0 21252 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0589_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0590_
timestamp 1666464484
transform -1 0 27692 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _0591_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25760 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _0592_
timestamp 1666464484
transform -1 0 26680 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0593_
timestamp 1666464484
transform -1 0 14812 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0594_
timestamp 1666464484
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0595_
timestamp 1666464484
transform 1 0 26036 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 24104 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1666464484
transform 1 0 23000 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_2  _0598_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25760 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _0599_
timestamp 1666464484
transform 1 0 25208 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0600_
timestamp 1666464484
transform -1 0 23184 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0601_
timestamp 1666464484
transform 1 0 21988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _0602_
timestamp 1666464484
transform -1 0 26956 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _0603_
timestamp 1666464484
transform 1 0 26128 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0604_
timestamp 1666464484
transform -1 0 15456 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0605_
timestamp 1666464484
transform 1 0 2300 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0606_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26956 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0607_
timestamp 1666464484
transform 1 0 28244 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0608_
timestamp 1666464484
transform 1 0 30176 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0609_
timestamp 1666464484
transform 1 0 24564 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0610_
timestamp 1666464484
transform -1 0 22908 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0611_
timestamp 1666464484
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0612_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26128 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 24104 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23460 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0615_
timestamp 1666464484
transform -1 0 25024 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0616_
timestamp 1666464484
transform 1 0 23552 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _0617_
timestamp 1666464484
transform -1 0 26956 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _0618_
timestamp 1666464484
transform -1 0 23736 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0619_
timestamp 1666464484
transform 1 0 22540 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_4  _0620_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26496 0 1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__and4bb_2  _0621_
timestamp 1666464484
transform -1 0 28060 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _0622_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 54004 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0623_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28888 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27600 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0625_
timestamp 1666464484
transform 1 0 27876 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0626_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27968 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0627_
timestamp 1666464484
transform -1 0 27416 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_4  _0628_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28704 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__clkinv_2  _0629_
timestamp 1666464484
transform -1 0 30360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0630_
timestamp 1666464484
transform 1 0 22080 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0631_
timestamp 1666464484
transform 1 0 22908 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _0632_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24656 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0633_
timestamp 1666464484
transform 1 0 24472 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0634_
timestamp 1666464484
transform 1 0 14904 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0635_
timestamp 1666464484
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13984 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0637_
timestamp 1666464484
transform 1 0 14260 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _0638_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26588 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _0639_
timestamp 1666464484
transform -1 0 28244 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0640_
timestamp 1666464484
transform 1 0 31372 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0641_
timestamp 1666464484
transform 1 0 26128 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0642_
timestamp 1666464484
transform -1 0 28428 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0644_
timestamp 1666464484
transform 1 0 32292 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0645_
timestamp 1666464484
transform -1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0646_
timestamp 1666464484
transform 1 0 25024 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0647_
timestamp 1666464484
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0648_
timestamp 1666464484
transform 1 0 14904 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0649_
timestamp 1666464484
transform 1 0 15272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _0650_
timestamp 1666464484
transform 1 0 25484 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _0651_
timestamp 1666464484
transform -1 0 18308 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0652_
timestamp 1666464484
transform -1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26772 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0654_
timestamp 1666464484
transform 1 0 25484 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0655_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30820 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0656_
timestamp 1666464484
transform -1 0 27324 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0657_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28612 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0658_
timestamp 1666464484
transform 1 0 29256 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0659_
timestamp 1666464484
transform 1 0 29808 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0660_
timestamp 1666464484
transform 1 0 30820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0661_
timestamp 1666464484
transform -1 0 30360 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0662_
timestamp 1666464484
transform 1 0 31464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0663_
timestamp 1666464484
transform 1 0 28796 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0664_
timestamp 1666464484
transform 1 0 29256 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0665_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29716 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0666_
timestamp 1666464484
transform -1 0 25852 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0667_
timestamp 1666464484
transform 1 0 26496 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0668_
timestamp 1666464484
transform 1 0 29808 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0669_
timestamp 1666464484
transform 1 0 13984 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0670_
timestamp 1666464484
transform 1 0 30084 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0671_
timestamp 1666464484
transform -1 0 31096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0672_
timestamp 1666464484
transform -1 0 30820 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0673_
timestamp 1666464484
transform -1 0 23920 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0674_
timestamp 1666464484
transform 1 0 14812 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0675_
timestamp 1666464484
transform -1 0 30636 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0676_
timestamp 1666464484
transform -1 0 28796 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0677_
timestamp 1666464484
transform 1 0 27140 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0678_
timestamp 1666464484
transform 1 0 28336 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0679_
timestamp 1666464484
transform -1 0 30452 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0680_
timestamp 1666464484
transform 1 0 29716 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0681_
timestamp 1666464484
transform -1 0 30084 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0682_
timestamp 1666464484
transform 1 0 27140 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0683_
timestamp 1666464484
transform -1 0 27876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0684_
timestamp 1666464484
transform 1 0 27140 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0685_
timestamp 1666464484
transform 1 0 27232 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0686_
timestamp 1666464484
transform 1 0 28244 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0687_
timestamp 1666464484
transform 1 0 28244 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0688_
timestamp 1666464484
transform 1 0 13800 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0689_
timestamp 1666464484
transform -1 0 29716 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0690_
timestamp 1666464484
transform 1 0 27324 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0691_
timestamp 1666464484
transform 1 0 27140 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0692_
timestamp 1666464484
transform -1 0 28796 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0693_
timestamp 1666464484
transform 1 0 28704 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0694_
timestamp 1666464484
transform -1 0 29532 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0695_
timestamp 1666464484
transform 1 0 26036 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0696_
timestamp 1666464484
transform -1 0 27232 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0697_
timestamp 1666464484
transform 1 0 25852 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0698_
timestamp 1666464484
transform -1 0 27784 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0699_
timestamp 1666464484
transform 1 0 25944 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0700_
timestamp 1666464484
transform -1 0 25668 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0701_
timestamp 1666464484
transform 1 0 25760 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0702_
timestamp 1666464484
transform 1 0 24012 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0703_
timestamp 1666464484
transform 1 0 23552 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0704_
timestamp 1666464484
transform -1 0 31556 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0705_
timestamp 1666464484
transform -1 0 25484 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0706_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25852 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0707_
timestamp 1666464484
transform -1 0 26588 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0708_
timestamp 1666464484
transform 1 0 24656 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0709_
timestamp 1666464484
transform 1 0 25208 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0710_
timestamp 1666464484
transform -1 0 27876 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0711_
timestamp 1666464484
transform -1 0 26128 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0712_
timestamp 1666464484
transform -1 0 25300 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0713_
timestamp 1666464484
transform 1 0 26680 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0714_
timestamp 1666464484
transform 1 0 28336 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0715_
timestamp 1666464484
transform 1 0 25116 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0716_
timestamp 1666464484
transform 1 0 25852 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0717_
timestamp 1666464484
transform -1 0 28336 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0718_
timestamp 1666464484
transform 1 0 27416 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0719_
timestamp 1666464484
transform -1 0 29532 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0720_
timestamp 1666464484
transform 1 0 26036 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0721_
timestamp 1666464484
transform 1 0 26588 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0722_
timestamp 1666464484
transform 1 0 25024 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0723_
timestamp 1666464484
transform 1 0 27140 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0724_
timestamp 1666464484
transform 1 0 27692 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0725_
timestamp 1666464484
transform -1 0 28428 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0726_
timestamp 1666464484
transform 1 0 23644 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0727_
timestamp 1666464484
transform -1 0 26680 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0728_
timestamp 1666464484
transform 1 0 26404 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0729_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _0730_
timestamp 1666464484
transform 1 0 26128 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0731_
timestamp 1666464484
transform 1 0 16836 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0732_
timestamp 1666464484
transform -1 0 27968 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0733_
timestamp 1666464484
transform -1 0 27784 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0734_
timestamp 1666464484
transform -1 0 26680 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0735_
timestamp 1666464484
transform 1 0 28336 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0736_
timestamp 1666464484
transform 1 0 27508 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0737_
timestamp 1666464484
transform -1 0 30452 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0738_
timestamp 1666464484
transform 1 0 28428 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0739_
timestamp 1666464484
transform -1 0 28888 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0740_
timestamp 1666464484
transform 1 0 27692 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0741_
timestamp 1666464484
transform 1 0 28152 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0742_
timestamp 1666464484
transform 1 0 29808 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0743_
timestamp 1666464484
transform -1 0 33028 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0744_
timestamp 1666464484
transform -1 0 31648 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0745_
timestamp 1666464484
transform -1 0 31004 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0746_
timestamp 1666464484
transform -1 0 53084 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0747_
timestamp 1666464484
transform 1 0 30820 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0748_
timestamp 1666464484
transform 1 0 31280 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0749_
timestamp 1666464484
transform -1 0 31832 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0750_
timestamp 1666464484
transform -1 0 32936 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0751_
timestamp 1666464484
transform -1 0 33120 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0752_
timestamp 1666464484
transform 1 0 32476 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0753_
timestamp 1666464484
transform -1 0 32936 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0754_
timestamp 1666464484
transform 1 0 53268 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0755_
timestamp 1666464484
transform 1 0 31924 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0756_
timestamp 1666464484
transform 1 0 33396 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0757_
timestamp 1666464484
transform -1 0 30820 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0758_
timestamp 1666464484
transform -1 0 34408 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0759_
timestamp 1666464484
transform -1 0 33488 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0760_
timestamp 1666464484
transform 1 0 32844 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0761_
timestamp 1666464484
transform 1 0 34408 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0762_
timestamp 1666464484
transform -1 0 52072 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0763_
timestamp 1666464484
transform 1 0 33028 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0764_
timestamp 1666464484
transform 1 0 33856 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0765_
timestamp 1666464484
transform 1 0 34868 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0766_
timestamp 1666464484
transform 1 0 32384 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0767_
timestamp 1666464484
transform 1 0 33120 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0768_
timestamp 1666464484
transform -1 0 33764 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0769_
timestamp 1666464484
transform -1 0 33672 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0770_
timestamp 1666464484
transform -1 0 52440 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0771_
timestamp 1666464484
transform 1 0 33028 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1666464484
transform 1 0 34224 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0773_
timestamp 1666464484
transform 1 0 35052 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0774_
timestamp 1666464484
transform -1 0 34776 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0775_
timestamp 1666464484
transform -1 0 33120 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0776_
timestamp 1666464484
transform 1 0 33488 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0777_
timestamp 1666464484
transform -1 0 34040 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0778_
timestamp 1666464484
transform -1 0 34224 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0779_
timestamp 1666464484
transform 1 0 32476 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0780_
timestamp 1666464484
transform 1 0 33580 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0781_
timestamp 1666464484
transform 1 0 31648 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0782_
timestamp 1666464484
transform -1 0 34132 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0783_
timestamp 1666464484
transform 1 0 32476 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0784_
timestamp 1666464484
transform 1 0 34868 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0785_
timestamp 1666464484
transform -1 0 35236 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0786_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22264 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0787_
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0788_
timestamp 1666464484
transform -1 0 22908 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0789_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23276 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0790_
timestamp 1666464484
transform 1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0791_
timestamp 1666464484
transform 1 0 14536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0792_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14352 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0793_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14444 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0794_
timestamp 1666464484
transform -1 0 14720 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0795_
timestamp 1666464484
transform 1 0 9476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0796_
timestamp 1666464484
transform 1 0 10396 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0797_
timestamp 1666464484
transform 1 0 10212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0798_
timestamp 1666464484
transform 1 0 10488 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0799_
timestamp 1666464484
transform 1 0 9568 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0800_
timestamp 1666464484
transform 1 0 10488 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0801_
timestamp 1666464484
transform -1 0 13524 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0802_
timestamp 1666464484
transform 1 0 12420 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0803_
timestamp 1666464484
transform 1 0 11960 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0804_
timestamp 1666464484
transform 1 0 13064 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0805_
timestamp 1666464484
transform 1 0 12052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0806_
timestamp 1666464484
transform 1 0 12972 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0807_
timestamp 1666464484
transform 1 0 11224 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0808_
timestamp 1666464484
transform 1 0 13064 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0809_
timestamp 1666464484
transform 1 0 12144 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0810_
timestamp 1666464484
transform 1 0 12420 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0811_
timestamp 1666464484
transform 1 0 12052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0812_
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0813_
timestamp 1666464484
transform -1 0 17112 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0814_
timestamp 1666464484
transform 1 0 13432 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0815_
timestamp 1666464484
transform 1 0 14260 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0816_
timestamp 1666464484
transform -1 0 17204 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0817_
timestamp 1666464484
transform 1 0 13248 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0818_
timestamp 1666464484
transform 1 0 13984 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0819_
timestamp 1666464484
transform 1 0 13064 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0820_
timestamp 1666464484
transform -1 0 15640 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0821_
timestamp 1666464484
transform 1 0 14352 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0822_
timestamp 1666464484
transform 1 0 14996 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0823_
timestamp 1666464484
transform 1 0 13248 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0824_
timestamp 1666464484
transform 1 0 14904 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0825_
timestamp 1666464484
transform 1 0 13984 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0826_
timestamp 1666464484
transform 1 0 14720 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0827_
timestamp 1666464484
transform 1 0 14720 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0828_
timestamp 1666464484
transform 1 0 15732 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0829_
timestamp 1666464484
transform -1 0 17388 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0830_
timestamp 1666464484
transform 1 0 15824 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0831_
timestamp 1666464484
transform 1 0 15640 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0832_
timestamp 1666464484
transform 1 0 15732 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0833_
timestamp 1666464484
transform 1 0 15916 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0834_
timestamp 1666464484
transform 1 0 16008 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0835_
timestamp 1666464484
transform -1 0 17388 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0836_
timestamp 1666464484
transform 1 0 15732 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0837_
timestamp 1666464484
transform 1 0 16836 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0838_
timestamp 1666464484
transform 1 0 16836 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0839_
timestamp 1666464484
transform -1 0 17112 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0840_
timestamp 1666464484
transform 1 0 15548 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0841_
timestamp 1666464484
transform 1 0 16836 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0842_
timestamp 1666464484
transform 1 0 16836 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0843_
timestamp 1666464484
transform -1 0 17572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0844_
timestamp 1666464484
transform 1 0 16560 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0845_
timestamp 1666464484
transform -1 0 17756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0846_
timestamp 1666464484
transform 1 0 16744 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0847_
timestamp 1666464484
transform -1 0 17756 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0848_
timestamp 1666464484
transform 1 0 16836 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0849_
timestamp 1666464484
transform -1 0 41492 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 1666464484
transform 1 0 42504 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 52716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0852_
timestamp 1666464484
transform 1 0 40020 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0853_
timestamp 1666464484
transform 1 0 40020 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0854_
timestamp 1666464484
transform 1 0 39284 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0855_
timestamp 1666464484
transform -1 0 39192 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0856_
timestamp 1666464484
transform -1 0 38640 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1666464484
transform 1 0 39192 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0858_
timestamp 1666464484
transform -1 0 37812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0859_
timestamp 1666464484
transform 1 0 33948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1666464484
transform -1 0 29256 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0861_
timestamp 1666464484
transform 1 0 28888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0862_
timestamp 1666464484
transform 1 0 32568 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0863_
timestamp 1666464484
transform 1 0 32292 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0864_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31372 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _0865_
timestamp 1666464484
transform -1 0 40388 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0866_
timestamp 1666464484
transform 1 0 40020 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0867_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 38180 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30176 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0869_
timestamp 1666464484
transform -1 0 37812 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0870_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 36156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0871_
timestamp 1666464484
transform -1 0 40480 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0872_
timestamp 1666464484
transform 1 0 32660 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0873_
timestamp 1666464484
transform -1 0 30268 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0874_
timestamp 1666464484
transform -1 0 32384 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0875_
timestamp 1666464484
transform 1 0 38364 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0876_
timestamp 1666464484
transform -1 0 40756 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0877_
timestamp 1666464484
transform -1 0 31280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0878_
timestamp 1666464484
transform 1 0 30728 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0879_
timestamp 1666464484
transform -1 0 31280 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0880_
timestamp 1666464484
transform 1 0 40020 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0881_
timestamp 1666464484
transform -1 0 36708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0882_
timestamp 1666464484
transform -1 0 36984 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0883_
timestamp 1666464484
transform -1 0 34408 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0884_
timestamp 1666464484
transform 1 0 36340 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0885_
timestamp 1666464484
transform 1 0 37260 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _0886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35972 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0887_
timestamp 1666464484
transform -1 0 39468 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0888_
timestamp 1666464484
transform -1 0 29256 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0889_
timestamp 1666464484
transform 1 0 29624 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0890_
timestamp 1666464484
transform -1 0 31556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0891_
timestamp 1666464484
transform 1 0 38272 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0892_
timestamp 1666464484
transform -1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1666464484
transform 1 0 28244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0894_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0895_
timestamp 1666464484
transform -1 0 37812 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0896_
timestamp 1666464484
transform 1 0 40112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0897_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 38456 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0898_
timestamp 1666464484
transform 1 0 41216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0899_
timestamp 1666464484
transform 1 0 27508 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0900_
timestamp 1666464484
transform -1 0 39928 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0901_
timestamp 1666464484
transform 1 0 39100 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0902_
timestamp 1666464484
transform 1 0 40756 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0903_
timestamp 1666464484
transform -1 0 24840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0904_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28152 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0905_
timestamp 1666464484
transform -1 0 37628 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0906_
timestamp 1666464484
transform 1 0 41860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0907_
timestamp 1666464484
transform 1 0 40756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0908_
timestamp 1666464484
transform 1 0 27140 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0909_
timestamp 1666464484
transform 1 0 38916 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0910_
timestamp 1666464484
transform 1 0 40296 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 1666464484
transform 1 0 43148 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0912_
timestamp 1666464484
transform 1 0 23644 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0913_
timestamp 1666464484
transform -1 0 27968 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0914_
timestamp 1666464484
transform 1 0 38824 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0915_
timestamp 1666464484
transform 1 0 40664 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0916_
timestamp 1666464484
transform 1 0 41860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1666464484
transform -1 0 30176 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0918_
timestamp 1666464484
transform 1 0 28152 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0919_
timestamp 1666464484
transform 1 0 38640 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0920_
timestamp 1666464484
transform 1 0 37996 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0921_
timestamp 1666464484
transform 1 0 41492 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0922_
timestamp 1666464484
transform -1 0 28612 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0923_
timestamp 1666464484
transform 1 0 32936 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0924_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 36156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0925_
timestamp 1666464484
transform 1 0 37260 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0926_
timestamp 1666464484
transform 1 0 41308 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0927_
timestamp 1666464484
transform -1 0 38456 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0928_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29256 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0929_
timestamp 1666464484
transform 1 0 38732 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0930_
timestamp 1666464484
transform 1 0 40480 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1666464484
transform 1 0 41492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0932_
timestamp 1666464484
transform -1 0 31280 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0933_
timestamp 1666464484
transform -1 0 29164 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0934_
timestamp 1666464484
transform -1 0 41124 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0935_
timestamp 1666464484
transform 1 0 39652 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0936_
timestamp 1666464484
transform 1 0 41492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0937_
timestamp 1666464484
transform -1 0 29164 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0938_
timestamp 1666464484
transform 1 0 38916 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0939_
timestamp 1666464484
transform 1 0 42044 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0940_
timestamp 1666464484
transform 1 0 43240 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0941_
timestamp 1666464484
transform -1 0 30544 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0942_
timestamp 1666464484
transform -1 0 41860 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0943_
timestamp 1666464484
transform 1 0 38180 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0944_
timestamp 1666464484
transform 1 0 42596 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0945_
timestamp 1666464484
transform -1 0 33120 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0946_
timestamp 1666464484
transform 1 0 39468 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0947_
timestamp 1666464484
transform 1 0 41860 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0948_
timestamp 1666464484
transform 1 0 42596 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0949_
timestamp 1666464484
transform -1 0 34316 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0950_
timestamp 1666464484
transform 1 0 40020 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0951_
timestamp 1666464484
transform 1 0 41032 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0952_
timestamp 1666464484
transform 1 0 42780 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0953_
timestamp 1666464484
transform -1 0 33120 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0954_
timestamp 1666464484
transform 1 0 38732 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0955_
timestamp 1666464484
transform 1 0 40020 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0956_
timestamp 1666464484
transform -1 0 40664 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0957_
timestamp 1666464484
transform -1 0 35604 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0958_
timestamp 1666464484
transform 1 0 38548 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0959_
timestamp 1666464484
transform -1 0 40204 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0960_
timestamp 1666464484
transform -1 0 39284 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0961_
timestamp 1666464484
transform -1 0 35696 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0962_
timestamp 1666464484
transform 1 0 37536 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0963_
timestamp 1666464484
transform 1 0 37444 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0964_
timestamp 1666464484
transform -1 0 38640 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0965_
timestamp 1666464484
transform -1 0 35972 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0966_
timestamp 1666464484
transform 1 0 37444 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0967_
timestamp 1666464484
transform -1 0 39008 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0968_
timestamp 1666464484
transform -1 0 37996 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0969_
timestamp 1666464484
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0970_
timestamp 1666464484
transform 1 0 35972 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0971_
timestamp 1666464484
transform -1 0 36800 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0972_
timestamp 1666464484
transform 1 0 35328 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0973_
timestamp 1666464484
transform -1 0 36616 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0974_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 37904 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0975_
timestamp 1666464484
transform -1 0 34316 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0976_
timestamp 1666464484
transform 1 0 32752 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1666464484
transform -1 0 33396 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0978_
timestamp 1666464484
transform 1 0 33764 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0979_
timestamp 1666464484
transform 1 0 34868 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1666464484
transform 1 0 35144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0981_
timestamp 1666464484
transform 1 0 33856 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0982_
timestamp 1666464484
transform 1 0 34316 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1666464484
transform 1 0 35696 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0984_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 35880 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0985_
timestamp 1666464484
transform -1 0 35972 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0986_
timestamp 1666464484
transform -1 0 36616 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0987_
timestamp 1666464484
transform 1 0 33580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0988_
timestamp 1666464484
transform 1 0 34868 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0989_
timestamp 1666464484
transform -1 0 35420 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1666464484
transform -1 0 35052 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0991_
timestamp 1666464484
transform -1 0 34408 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0992_
timestamp 1666464484
transform -1 0 31004 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0993_
timestamp 1666464484
transform 1 0 29900 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1666464484
transform 1 0 37444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0995_
timestamp 1666464484
transform 1 0 32660 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0996_
timestamp 1666464484
transform -1 0 31648 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0997_
timestamp 1666464484
transform 1 0 33396 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0998_
timestamp 1666464484
transform 1 0 31648 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0999_
timestamp 1666464484
transform -1 0 30636 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1666464484
transform -1 0 29256 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1001_
timestamp 1666464484
transform -1 0 29072 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1002_
timestamp 1666464484
transform 1 0 26404 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1003_
timestamp 1666464484
transform -1 0 26588 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1004_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1005_
timestamp 1666464484
transform -1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23460 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1007_
timestamp 1666464484
transform -1 0 25024 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1008_
timestamp 1666464484
transform 1 0 22816 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1009_
timestamp 1666464484
transform 1 0 27140 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1010_
timestamp 1666464484
transform -1 0 29624 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1666464484
transform -1 0 22356 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1012_
timestamp 1666464484
transform 1 0 26864 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1013_
timestamp 1666464484
transform -1 0 22448 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1014_
timestamp 1666464484
transform -1 0 24840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1015_
timestamp 1666464484
transform 1 0 23460 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1016_
timestamp 1666464484
transform 1 0 29072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1017_
timestamp 1666464484
transform 1 0 29716 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1018_
timestamp 1666464484
transform -1 0 28520 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1019_
timestamp 1666464484
transform 1 0 28336 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1020_
timestamp 1666464484
transform -1 0 28704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1666464484
transform -1 0 27784 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1022_
timestamp 1666464484
transform -1 0 27416 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1666464484
transform -1 0 26864 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1024_
timestamp 1666464484
transform -1 0 26036 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1666464484
transform -1 0 24932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1026_
timestamp 1666464484
transform -1 0 27048 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1027_
timestamp 1666464484
transform -1 0 27968 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1028_
timestamp 1666464484
transform 1 0 29716 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1029_
timestamp 1666464484
transform 1 0 27600 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1666464484
transform 1 0 29348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1031_
timestamp 1666464484
transform -1 0 31832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1032_
timestamp 1666464484
transform 1 0 30728 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1033_
timestamp 1666464484
transform -1 0 33856 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1666464484
transform -1 0 29992 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1035_
timestamp 1666464484
transform 1 0 29808 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1036_
timestamp 1666464484
transform -1 0 32936 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1037_
timestamp 1666464484
transform 1 0 33212 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1038_
timestamp 1666464484
transform 1 0 29992 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1666464484
transform 1 0 36708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1040_
timestamp 1666464484
transform -1 0 34040 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1041_
timestamp 1666464484
transform -1 0 40020 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1042_
timestamp 1666464484
transform 1 0 33396 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1043_
timestamp 1666464484
transform -1 0 36984 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1044_
timestamp 1666464484
transform 1 0 35972 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1045_
timestamp 1666464484
transform -1 0 39376 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1046_
timestamp 1666464484
transform 1 0 39284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1047_
timestamp 1666464484
transform -1 0 34408 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _1048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 53360 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1049_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29716 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 1666464484
transform 1 0 27968 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1051_
timestamp 1666464484
transform -1 0 28428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1052_
timestamp 1666464484
transform -1 0 25392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1053_
timestamp 1666464484
transform 1 0 28152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1054_
timestamp 1666464484
transform 1 0 22816 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1055_
timestamp 1666464484
transform -1 0 20240 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1056_
timestamp 1666464484
transform 1 0 26864 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1057_
timestamp 1666464484
transform 1 0 26036 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1058_
timestamp 1666464484
transform -1 0 27416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1059_
timestamp 1666464484
transform -1 0 30176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1060_
timestamp 1666464484
transform -1 0 31648 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1061_
timestamp 1666464484
transform 1 0 30360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1062_
timestamp 1666464484
transform 1 0 29164 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1063_
timestamp 1666464484
transform -1 0 29256 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1064_
timestamp 1666464484
transform -1 0 28152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1065_
timestamp 1666464484
transform 1 0 27232 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1066_
timestamp 1666464484
transform 1 0 27140 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1067_
timestamp 1666464484
transform 1 0 31188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1666464484
transform 1 0 28520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1069_
timestamp 1666464484
transform -1 0 30912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1070_
timestamp 1666464484
transform -1 0 28980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1071_
timestamp 1666464484
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 1666464484
transform -1 0 21528 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1073_
timestamp 1666464484
transform -1 0 49036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1074_
timestamp 1666464484
transform -1 0 41584 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1075_
timestamp 1666464484
transform -1 0 41124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1076_
timestamp 1666464484
transform -1 0 34408 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1077_
timestamp 1666464484
transform 1 0 34868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1078_
timestamp 1666464484
transform -1 0 33764 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1079_
timestamp 1666464484
transform -1 0 33120 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1080_
timestamp 1666464484
transform -1 0 34408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1081_
timestamp 1666464484
transform -1 0 34408 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1082_
timestamp 1666464484
transform 1 0 34868 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1083_
timestamp 1666464484
transform 1 0 35236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1084_
timestamp 1666464484
transform 1 0 33580 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1085_
timestamp 1666464484
transform 1 0 31832 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1666464484
transform 1 0 36064 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1087_
timestamp 1666464484
transform 1 0 31648 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1088_
timestamp 1666464484
transform 1 0 31372 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1089_
timestamp 1666464484
transform -1 0 32568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1090_
timestamp 1666464484
transform -1 0 33764 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1091_
timestamp 1666464484
transform 1 0 37444 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1666464484
transform 1 0 39100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1093_
timestamp 1666464484
transform 1 0 29624 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1094_
timestamp 1666464484
transform 1 0 28796 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1095_
timestamp 1666464484
transform -1 0 29256 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1096_
timestamp 1666464484
transform 1 0 25760 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1097_
timestamp 1666464484
transform -1 0 24380 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1098_
timestamp 1666464484
transform -1 0 22448 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1099_
timestamp 1666464484
transform 1 0 24564 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1100_
timestamp 1666464484
transform 1 0 22540 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1101_
timestamp 1666464484
transform -1 0 24104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1102_
timestamp 1666464484
transform 1 0 23368 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1103_
timestamp 1666464484
transform -1 0 22908 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1104_
timestamp 1666464484
transform -1 0 19688 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1105_
timestamp 1666464484
transform 1 0 23276 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1106_
timestamp 1666464484
transform -1 0 23000 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1107_
timestamp 1666464484
transform -1 0 18952 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1108_
timestamp 1666464484
transform -1 0 33580 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1109_
timestamp 1666464484
transform 1 0 24564 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1110_
timestamp 1666464484
transform -1 0 23552 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1111_
timestamp 1666464484
transform -1 0 22724 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1112_
timestamp 1666464484
transform -1 0 37812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1113_
timestamp 1666464484
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1114_
timestamp 1666464484
transform -1 0 24380 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1115_
timestamp 1666464484
transform -1 0 22724 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1116_
timestamp 1666464484
transform 1 0 31832 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1117_
timestamp 1666464484
transform 1 0 31004 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1118_
timestamp 1666464484
transform 1 0 38088 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1119_
timestamp 1666464484
transform -1 0 30544 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1120_
timestamp 1666464484
transform -1 0 31372 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1121_
timestamp 1666464484
transform -1 0 27508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1122_
timestamp 1666464484
transform 1 0 24012 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1123_
timestamp 1666464484
transform 1 0 23184 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1124_
timestamp 1666464484
transform -1 0 24104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1125_
timestamp 1666464484
transform 1 0 24564 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1126_
timestamp 1666464484
transform -1 0 25024 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1127_
timestamp 1666464484
transform -1 0 23552 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1128_
timestamp 1666464484
transform 1 0 27140 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1129_
timestamp 1666464484
transform 1 0 27324 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1130_
timestamp 1666464484
transform 1 0 28152 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1131_
timestamp 1666464484
transform 1 0 30912 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1132_
timestamp 1666464484
transform 1 0 29532 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1133_
timestamp 1666464484
transform -1 0 30268 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1134_
timestamp 1666464484
transform 1 0 32292 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1135_
timestamp 1666464484
transform 1 0 30544 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1136_
timestamp 1666464484
transform -1 0 31004 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1137_
timestamp 1666464484
transform 1 0 32108 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1138_
timestamp 1666464484
transform 1 0 31372 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1139_
timestamp 1666464484
transform 1 0 32200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1140_
timestamp 1666464484
transform 1 0 34868 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1141_
timestamp 1666464484
transform 1 0 32844 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1142_
timestamp 1666464484
transform 1 0 36708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1143_
timestamp 1666464484
transform 1 0 34868 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1144_
timestamp 1666464484
transform 1 0 34868 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1145_
timestamp 1666464484
transform 1 0 39008 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1146_
timestamp 1666464484
transform 1 0 37628 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1147_
timestamp 1666464484
transform 1 0 36524 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1148_
timestamp 1666464484
transform 1 0 41860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1149_
timestamp 1666464484
transform -1 0 38272 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1150_
timestamp 1666464484
transform 1 0 38640 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1151_
timestamp 1666464484
transform 1 0 40020 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1152_
timestamp 1666464484
transform 1 0 50600 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1153_
timestamp 1666464484
transform -1 0 51888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30084 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1155_
timestamp 1666464484
transform -1 0 23000 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1156_
timestamp 1666464484
transform -1 0 21804 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1157_
timestamp 1666464484
transform 1 0 21988 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1158_
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1159_
timestamp 1666464484
transform 1 0 25116 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1160_
timestamp 1666464484
transform -1 0 22632 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1161_
timestamp 1666464484
transform 1 0 20976 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1162_
timestamp 1666464484
transform -1 0 18952 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1163_
timestamp 1666464484
transform 1 0 21988 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1164_
timestamp 1666464484
transform -1 0 18952 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1165_
timestamp 1666464484
transform 1 0 24564 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1166_
timestamp 1666464484
transform -1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1167_
timestamp 1666464484
transform -1 0 18952 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1168_
timestamp 1666464484
transform -1 0 19596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1169_
timestamp 1666464484
transform 1 0 24564 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1170_
timestamp 1666464484
transform -1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1171_
timestamp 1666464484
transform -1 0 25392 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1172_
timestamp 1666464484
transform 1 0 25760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1173_
timestamp 1666464484
transform 1 0 19228 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1174_
timestamp 1666464484
transform 1 0 18676 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1175_
timestamp 1666464484
transform 1 0 19412 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1176_
timestamp 1666464484
transform -1 0 15548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1177_
timestamp 1666464484
transform -1 0 22540 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1178_
timestamp 1666464484
transform 1 0 19412 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1179_
timestamp 1666464484
transform -1 0 18308 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1180_
timestamp 1666464484
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1666464484
transform -1 0 17756 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1182_
timestamp 1666464484
transform 1 0 20608 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1183_
timestamp 1666464484
transform -1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1184_
timestamp 1666464484
transform 1 0 20516 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1185_
timestamp 1666464484
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1186_
timestamp 1666464484
transform 1 0 18124 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1187_
timestamp 1666464484
transform -1 0 16376 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1188_
timestamp 1666464484
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1189_
timestamp 1666464484
transform -1 0 16376 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1190_
timestamp 1666464484
transform 1 0 20424 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1191_
timestamp 1666464484
transform -1 0 16376 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1192_
timestamp 1666464484
transform 1 0 21252 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1193_
timestamp 1666464484
transform 1 0 20608 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1194_
timestamp 1666464484
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1195_
timestamp 1666464484
transform -1 0 17112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1196_
timestamp 1666464484
transform 1 0 18124 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1197_
timestamp 1666464484
transform -1 0 14904 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1198_
timestamp 1666464484
transform 1 0 21988 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1199_
timestamp 1666464484
transform -1 0 21620 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1200_
timestamp 1666464484
transform -1 0 21528 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1201_
timestamp 1666464484
transform 1 0 21620 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1202_
timestamp 1666464484
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1203_
timestamp 1666464484
transform -1 0 20700 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1204_
timestamp 1666464484
transform 1 0 19596 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1205_
timestamp 1666464484
transform 1 0 19228 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1206_
timestamp 1666464484
transform 1 0 20608 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1207_
timestamp 1666464484
transform -1 0 19688 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1208_
timestamp 1666464484
transform 1 0 21252 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1666464484
transform -1 0 18952 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1210_
timestamp 1666464484
transform 1 0 20516 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1211_
timestamp 1666464484
transform -1 0 17480 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1212_
timestamp 1666464484
transform 1 0 25668 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1213_
timestamp 1666464484
transform -1 0 25024 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1666464484
transform 1 0 25208 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1215_
timestamp 1666464484
transform 1 0 25760 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1216_
timestamp 1666464484
transform 1 0 25300 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1217_
timestamp 1666464484
transform -1 0 25116 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1218_
timestamp 1666464484
transform -1 0 26680 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1219_
timestamp 1666464484
transform 1 0 25852 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1220_
timestamp 1666464484
transform -1 0 24656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1221_
timestamp 1666464484
transform 1 0 27140 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1222_
timestamp 1666464484
transform 1 0 27140 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1223_
timestamp 1666464484
transform 1 0 27048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 37996 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1225_
timestamp 1666464484
transform 1 0 36524 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1226_
timestamp 1666464484
transform 1 0 38180 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1227_
timestamp 1666464484
transform 1 0 38456 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1228_
timestamp 1666464484
transform 1 0 35420 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1229_
timestamp 1666464484
transform 1 0 38272 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1230_
timestamp 1666464484
transform -1 0 38916 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1231_
timestamp 1666464484
transform -1 0 41492 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1232_
timestamp 1666464484
transform -1 0 38916 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1233_
timestamp 1666464484
transform -1 0 41492 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1234_
timestamp 1666464484
transform -1 0 41492 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1235_
timestamp 1666464484
transform -1 0 40296 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1236_
timestamp 1666464484
transform -1 0 38088 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1237_
timestamp 1666464484
transform -1 0 41492 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1238_
timestamp 1666464484
transform -1 0 41676 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1239_
timestamp 1666464484
transform 1 0 40756 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1240_
timestamp 1666464484
transform 1 0 40664 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1241_
timestamp 1666464484
transform 1 0 40664 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1242_
timestamp 1666464484
transform 1 0 40940 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1243_
timestamp 1666464484
transform 1 0 40664 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1244_
timestamp 1666464484
transform 1 0 40020 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1245_
timestamp 1666464484
transform 1 0 38364 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1246_
timestamp 1666464484
transform 1 0 38272 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp 1666464484
transform 1 0 36708 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp 1666464484
transform 1 0 33580 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1249_
timestamp 1666464484
transform 1 0 34868 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1250_
timestamp 1666464484
transform 1 0 35420 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp 1666464484
transform 1 0 34132 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp 1666464484
transform -1 0 36340 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1253_
timestamp 1666464484
transform -1 0 36340 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1254_
timestamp 1666464484
transform -1 0 32844 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1255_
timestamp 1666464484
transform -1 0 33764 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1256_
timestamp 1666464484
transform 1 0 29808 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1257_
timestamp 1666464484
transform -1 0 28612 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1258_
timestamp 1666464484
transform 1 0 25208 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1259_
timestamp 1666464484
transform -1 0 26680 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1260_
timestamp 1666464484
transform 1 0 24564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1261_
timestamp 1666464484
transform -1 0 26680 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1262_
timestamp 1666464484
transform 1 0 24932 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1263_
timestamp 1666464484
transform 1 0 30176 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1264_
timestamp 1666464484
transform 1 0 28336 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1265_
timestamp 1666464484
transform 1 0 25208 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1266_
timestamp 1666464484
transform 1 0 25760 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1267_
timestamp 1666464484
transform -1 0 29256 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1268_
timestamp 1666464484
transform 1 0 30820 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1269_
timestamp 1666464484
transform 1 0 31372 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1270_
timestamp 1666464484
transform -1 0 34132 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1271_
timestamp 1666464484
transform 1 0 34316 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1272_
timestamp 1666464484
transform 1 0 34408 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1273_
timestamp 1666464484
transform -1 0 36340 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1274_
timestamp 1666464484
transform 1 0 34684 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1275_
timestamp 1666464484
transform 1 0 27140 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1276_
timestamp 1666464484
transform 1 0 22172 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27600 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1278_
timestamp 1666464484
transform 1 0 29716 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1279_
timestamp 1666464484
transform 1 0 29348 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1280_
timestamp 1666464484
transform -1 0 28612 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1281_
timestamp 1666464484
transform 1 0 29716 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1282_
timestamp 1666464484
transform 1 0 22264 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1283_
timestamp 1666464484
transform 1 0 48760 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1284_
timestamp 1666464484
transform 1 0 33396 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1285_
timestamp 1666464484
transform 1 0 34592 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1286_
timestamp 1666464484
transform -1 0 35420 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1287_
timestamp 1666464484
transform -1 0 33764 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1288_
timestamp 1666464484
transform -1 0 34316 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1289_
timestamp 1666464484
transform 1 0 29716 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1290_
timestamp 1666464484
transform 1 0 24748 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1291_
timestamp 1666464484
transform 1 0 24564 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1292_
timestamp 1666464484
transform 1 0 22540 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1293_
timestamp 1666464484
transform 1 0 22264 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1294_
timestamp 1666464484
transform 1 0 22724 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1295_
timestamp 1666464484
transform 1 0 23092 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1296_
timestamp 1666464484
transform -1 0 33764 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1297_
timestamp 1666464484
transform -1 0 30360 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1298_
timestamp 1666464484
transform 1 0 24564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1299_
timestamp 1666464484
transform 1 0 23920 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1300_
timestamp 1666464484
transform 1 0 27416 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1301_
timestamp 1666464484
transform 1 0 29808 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1302_
timestamp 1666464484
transform 1 0 31648 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1303_
timestamp 1666464484
transform 1 0 30360 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1304_
timestamp 1666464484
transform -1 0 36340 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1305_
timestamp 1666464484
transform -1 0 35880 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1306_
timestamp 1666464484
transform -1 0 38916 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1307_
timestamp 1666464484
transform -1 0 38916 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1308_
timestamp 1666464484
transform 1 0 52900 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1309_
timestamp 1666464484
transform -1 0 21528 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1310_
timestamp 1666464484
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1311_
timestamp 1666464484
transform 1 0 20056 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1312_
timestamp 1666464484
transform 1 0 19872 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1313_
timestamp 1666464484
transform -1 0 24104 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1314_
timestamp 1666464484
transform -1 0 20884 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1315_
timestamp 1666464484
transform 1 0 23276 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1666464484
transform -1 0 25116 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1317_
timestamp 1666464484
transform 1 0 18216 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp 1666464484
transform 1 0 18216 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1319_
timestamp 1666464484
transform 1 0 18124 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp 1666464484
transform 1 0 17480 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1321_
timestamp 1666464484
transform -1 0 21436 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1322_
timestamp 1666464484
transform 1 0 19872 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp 1666464484
transform 1 0 17848 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp 1666464484
transform 1 0 20056 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1325_
timestamp 1666464484
transform 1 0 19412 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1326_
timestamp 1666464484
transform -1 0 19688 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1666464484
transform -1 0 18952 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1666464484
transform -1 0 19780 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1666464484
transform -1 0 23460 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1330_
timestamp 1666464484
transform -1 0 21344 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1331_
timestamp 1666464484
transform -1 0 22540 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1332_
timestamp 1666464484
transform 1 0 18676 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1333_
timestamp 1666464484
transform 1 0 19412 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1334_
timestamp 1666464484
transform 1 0 19412 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1335_
timestamp 1666464484
transform 1 0 18768 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1336_
timestamp 1666464484
transform 1 0 24932 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1337_
timestamp 1666464484
transform 1 0 25024 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1338_
timestamp 1666464484
transform 1 0 27140 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1339_
timestamp 1666464484
transform 1 0 26864 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _1367_
timestamp 1666464484
transform -1 0 37536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1368_
timestamp 1666464484
transform -1 0 38180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1369_
timestamp 1666464484
transform -1 0 39192 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1370_
timestamp 1666464484
transform -1 0 40296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1371_
timestamp 1666464484
transform -1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1372_
timestamp 1666464484
transform -1 0 42136 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 1666464484
transform -1 0 42964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1374_
timestamp 1666464484
transform -1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1375_
timestamp 1666464484
transform -1 0 44528 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1376_
timestamp 1666464484
transform -1 0 44160 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1377_
timestamp 1666464484
transform -1 0 44804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1378_
timestamp 1666464484
transform -1 0 45448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1379_
timestamp 1666464484
transform -1 0 45448 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1380_
timestamp 1666464484
transform -1 0 46092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1381_
timestamp 1666464484
transform -1 0 45816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1382_
timestamp 1666464484
transform -1 0 46736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net235 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20148 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1666464484
transform -1 0 36984 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net235
timestamp 1666464484
transform 1 0 18216 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net235
timestamp 1666464484
transform 1 0 18216 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1666464484
transform 1 0 23368 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1666464484
transform 1 0 26036 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1666464484
transform 1 0 20792 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1666464484
transform -1 0 25208 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1666464484
transform 1 0 36432 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1666464484
transform 1 0 39008 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1666464484
transform -1 0 38272 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1666464484
transform -1 0 40848 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  fanout355
timestamp 1666464484
transform -1 0 43240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout356
timestamp 1666464484
transform 1 0 15824 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 37168 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1666464484
transform 1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1666464484
transform -1 0 34040 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1666464484
transform -1 0 33028 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1666464484
transform -1 0 32568 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1666464484
transform 1 0 30360 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1666464484
transform 1 0 36248 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1666464484
transform -1 0 35604 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1666464484
transform 1 0 25760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1666464484
transform -1 0 27876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1666464484
transform 1 0 25760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1666464484
transform -1 0 34776 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1666464484
transform 1 0 33580 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1666464484
transform 1 0 25760 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1666464484
transform -1 0 26680 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1666464484
transform -1 0 25484 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1666464484
transform -1 0 26036 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1666464484
transform -1 0 24104 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1666464484
transform 1 0 25392 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1666464484
transform -1 0 33672 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1666464484
transform -1 0 34868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1666464484
transform -1 0 25760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1666464484
transform -1 0 24196 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1666464484
transform -1 0 26496 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1666464484
transform -1 0 36892 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1666464484
transform -1 0 36708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1666464484
transform 1 0 34868 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1666464484
transform 1 0 33672 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1666464484
transform 1 0 27232 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1666464484
transform 1 0 27876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1666464484
transform 1 0 27324 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1666464484
transform -1 0 31556 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1666464484
transform 1 0 30912 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1666464484
transform -1 0 31556 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1666464484
transform -1 0 37720 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1666464484
transform 1 0 36156 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1666464484
transform 1 0 37444 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1666464484
transform -1 0 30452 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1666464484
transform -1 0 28888 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1666464484
transform 1 0 29532 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1666464484
transform -1 0 30452 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1666464484
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1666464484
transform 1 0 32292 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1666464484
transform -1 0 31924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1666464484
transform 1 0 32292 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1666464484
transform -1 0 27324 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1666464484
transform 1 0 32108 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1666464484
transform -1 0 33028 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1666464484
transform 1 0 33212 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1666464484
transform 1 0 24656 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1666464484
transform 1 0 26404 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1666464484
transform -1 0 26312 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1666464484
transform 1 0 31648 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1666464484
transform -1 0 31740 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1666464484
transform -1 0 35420 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1666464484
transform 1 0 53452 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1666464484
transform 1 0 53452 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1666464484
transform -1 0 52440 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1666464484
transform 1 0 53452 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1666464484
transform 1 0 52164 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1666464484
transform 1 0 53452 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1666464484
transform -1 0 52440 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1666464484
transform 1 0 52808 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1666464484
transform 1 0 54096 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666464484
transform 1 0 53452 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1666464484
transform -1 0 53084 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1666464484
transform 1 0 53452 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1666464484
transform 1 0 54096 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1666464484
transform 1 0 52164 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1666464484
transform 1 0 53452 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1666464484
transform 1 0 53452 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1666464484
transform 1 0 52808 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1666464484
transform 1 0 52164 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1666464484
transform 1 0 52808 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1666464484
transform 1 0 52808 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1666464484
transform 1 0 53452 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1666464484
transform 1 0 53452 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1666464484
transform 1 0 53452 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1666464484
transform 1 0 53452 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1666464484
transform 1 0 53452 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1666464484
transform 1 0 53452 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1666464484
transform -1 0 53084 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1666464484
transform 1 0 1564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1666464484
transform 1 0 1564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1666464484
transform -1 0 1840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1666464484
transform -1 0 1840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1666464484
transform -1 0 2484 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1666464484
transform -1 0 2484 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1666464484
transform -1 0 1840 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1666464484
transform -1 0 2484 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1666464484
transform 1 0 53452 0 -1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1666464484
transform 1 0 52164 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1666464484
transform 1 0 53452 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1666464484
transform -1 0 52440 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1666464484
transform 1 0 53452 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1666464484
transform 1 0 52164 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1666464484
transform 1 0 53452 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1666464484
transform -1 0 52440 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1666464484
transform -1 0 52900 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1666464484
transform 1 0 51980 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1666464484
transform -1 0 51428 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1666464484
transform 1 0 53452 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1666464484
transform 1 0 54096 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1666464484
transform 1 0 52808 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1666464484
transform 1 0 52164 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1666464484
transform 1 0 54096 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1666464484
transform 1 0 53452 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1666464484
transform 1 0 53452 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1666464484
transform 1 0 53452 0 -1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1666464484
transform 1 0 53452 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1666464484
transform 1 0 53452 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1666464484
transform 1 0 53452 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1666464484
transform -1 0 53084 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1666464484
transform 1 0 53452 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1666464484
transform 1 0 53452 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1666464484
transform -1 0 52440 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1666464484
transform 1 0 53452 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1666464484
transform -1 0 2484 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1666464484
transform -1 0 2484 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1666464484
transform -1 0 2484 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1666464484
transform -1 0 2484 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1666464484
transform -1 0 2484 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1666464484
transform -1 0 2484 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1666464484
transform -1 0 2484 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1666464484
transform -1 0 2484 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1666464484
transform -1 0 2484 0 1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 1666464484
transform -1 0 2484 0 -1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1666464484
transform -1 0 2484 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1666464484
transform -1 0 2484 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1666464484
transform 1 0 1564 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1666464484
transform -1 0 2484 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1666464484
transform -1 0 2484 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1666464484
transform 1 0 1564 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1666464484
transform 1 0 1564 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1666464484
transform 1 0 1564 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1666464484
transform 1 0 2300 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input82
timestamp 1666464484
transform -1 0 2484 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input83
timestamp 1666464484
transform -1 0 2484 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input84
timestamp 1666464484
transform -1 0 2484 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1666464484
transform -1 0 2484 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1666464484
transform -1 0 2484 0 -1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input87
timestamp 1666464484
transform -1 0 2484 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1666464484
transform -1 0 2484 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input89
timestamp 1666464484
transform -1 0 2484 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input90
timestamp 1666464484
transform 1 0 11316 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1666464484
transform -1 0 23552 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1666464484
transform -1 0 24840 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1666464484
transform -1 0 25944 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1666464484
transform -1 0 27416 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1666464484
transform 1 0 28060 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1666464484
transform 1 0 29716 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1666464484
transform 1 0 30452 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1666464484
transform 1 0 32292 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1666464484
transform 1 0 32936 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1666464484
transform 1 0 34040 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input101
timestamp 1666464484
transform 1 0 12512 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1666464484
transform 1 0 35236 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1666464484
transform 1 0 36432 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1666464484
transform 1 0 37628 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1666464484
transform 1 0 38824 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1666464484
transform 1 0 40020 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1666464484
transform 1 0 41216 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1666464484
transform 1 0 42596 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1666464484
transform 1 0 14260 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1666464484
transform -1 0 15088 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input111
timestamp 1666464484
transform -1 0 16376 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input112
timestamp 1666464484
transform 1 0 17296 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input113
timestamp 1666464484
transform -1 0 18952 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1666464484
transform -1 0 19964 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1666464484
transform -1 0 21160 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1666464484
transform -1 0 22356 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input117
timestamp 1666464484
transform -1 0 48116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 1666464484
transform -1 0 51796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1666464484
transform -1 0 51428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1666464484
transform -1 0 48852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1666464484
transform -1 0 48852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input122
timestamp 1666464484
transform 1 0 49220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input123
timestamp 1666464484
transform -1 0 49588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input124
timestamp 1666464484
transform -1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input125
timestamp 1666464484
transform -1 0 50324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input126
timestamp 1666464484
transform -1 0 51428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input127
timestamp 1666464484
transform -1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input128
timestamp 1666464484
transform -1 0 52164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input129
timestamp 1666464484
transform 1 0 45172 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input130
timestamp 1666464484
transform 1 0 46000 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input131
timestamp 1666464484
transform 1 0 47748 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input132
timestamp 1666464484
transform 1 0 48392 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input133
timestamp 1666464484
transform 1 0 50324 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input134
timestamp 1666464484
transform -1 0 51980 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input135
timestamp 1666464484
transform -1 0 52348 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input136
timestamp 1666464484
transform 1 0 53176 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input137
timestamp 1666464484
transform -1 0 2484 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input138
timestamp 1666464484
transform -1 0 2484 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1666464484
transform -1 0 1840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input140
timestamp 1666464484
transform -1 0 2484 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input141
timestamp 1666464484
transform -1 0 2484 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input142
timestamp 1666464484
transform -1 0 2484 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input143
timestamp 1666464484
transform -1 0 2484 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input144
timestamp 1666464484
transform -1 0 2484 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input145
timestamp 1666464484
transform -1 0 1840 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input146
timestamp 1666464484
transform -1 0 2668 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input147
timestamp 1666464484
transform 1 0 3036 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input148
timestamp 1666464484
transform -1 0 4416 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input149
timestamp 1666464484
transform 1 0 5336 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input150
timestamp 1666464484
transform 1 0 6532 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input151
timestamp 1666464484
transform -1 0 8004 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input152
timestamp 1666464484
transform -1 0 9384 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input153
timestamp 1666464484
transform 1 0 10120 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input154
timestamp 1666464484
transform -1 0 2484 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input155
timestamp 1666464484
transform -1 0 2484 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input156
timestamp 1666464484
transform -1 0 1840 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input157
timestamp 1666464484
transform -1 0 2484 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input158
timestamp 1666464484
transform -1 0 2484 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input159
timestamp 1666464484
transform -1 0 2484 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input160
timestamp 1666464484
transform -1 0 2484 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input161
timestamp 1666464484
transform -1 0 1840 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input162
timestamp 1666464484
transform -1 0 54372 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input163
timestamp 1666464484
transform -1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input164
timestamp 1666464484
transform -1 0 8648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input165
timestamp 1666464484
transform -1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input166
timestamp 1666464484
transform -1 0 9200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input167
timestamp 1666464484
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input168
timestamp 1666464484
transform -1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input169
timestamp 1666464484
transform -1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input170
timestamp 1666464484
transform -1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input171
timestamp 1666464484
transform -1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input172
timestamp 1666464484
transform -1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input173
timestamp 1666464484
transform 1 0 12420 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input174
timestamp 1666464484
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input175
timestamp 1666464484
transform -1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input176
timestamp 1666464484
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input177
timestamp 1666464484
transform -1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input178
timestamp 1666464484
transform -1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input179
timestamp 1666464484
transform -1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input180
timestamp 1666464484
transform -1 0 13800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input181
timestamp 1666464484
transform -1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input182
timestamp 1666464484
transform -1 0 15088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input183
timestamp 1666464484
transform -1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input184
timestamp 1666464484
transform -1 0 16376 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input185
timestamp 1666464484
transform -1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input186
timestamp 1666464484
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input187
timestamp 1666464484
transform 1 0 17572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input188
timestamp 1666464484
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input189
timestamp 1666464484
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input190
timestamp 1666464484
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input191
timestamp 1666464484
transform -1 0 7176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input192
timestamp 1666464484
transform -1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input193
timestamp 1666464484
transform 1 0 7636 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input194
timestamp 1666464484
transform -1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input195
timestamp 1666464484
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input196
timestamp 1666464484
transform -1 0 52440 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input197
timestamp 1666464484
transform 1 0 54096 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input198
timestamp 1666464484
transform 1 0 1564 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input199
timestamp 1666464484
transform 1 0 43608 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input200
timestamp 1666464484
transform -1 0 2484 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input201
timestamp 1666464484
transform -1 0 54372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input202
timestamp 1666464484
transform 1 0 53452 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input203
timestamp 1666464484
transform -1 0 53636 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input204
timestamp 1666464484
transform 1 0 53452 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input205
timestamp 1666464484
transform -1 0 52532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input206
timestamp 1666464484
transform -1 0 53636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input207
timestamp 1666464484
transform -1 0 53636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input208
timestamp 1666464484
transform -1 0 54372 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input209
timestamp 1666464484
transform -1 0 53636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input210
timestamp 1666464484
transform -1 0 54372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input211
timestamp 1666464484
transform -1 0 53636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input212
timestamp 1666464484
transform -1 0 54372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input213
timestamp 1666464484
transform -1 0 53636 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input214
timestamp 1666464484
transform -1 0 54372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input215
timestamp 1666464484
transform -1 0 53636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input216
timestamp 1666464484
transform -1 0 54372 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input217
timestamp 1666464484
transform -1 0 53636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input218
timestamp 1666464484
transform -1 0 54372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input219
timestamp 1666464484
transform -1 0 54372 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input220
timestamp 1666464484
transform -1 0 53636 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input221
timestamp 1666464484
transform -1 0 54372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input222
timestamp 1666464484
transform -1 0 53636 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input223
timestamp 1666464484
transform -1 0 54372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input224
timestamp 1666464484
transform -1 0 54372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input225
timestamp 1666464484
transform -1 0 53636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input226
timestamp 1666464484
transform -1 0 54372 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input227
timestamp 1666464484
transform -1 0 53636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input228
timestamp 1666464484
transform -1 0 54372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input229
timestamp 1666464484
transform -1 0 53636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input230
timestamp 1666464484
transform -1 0 54372 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input231
timestamp 1666464484
transform -1 0 53636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input232
timestamp 1666464484
transform -1 0 54372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input233
timestamp 1666464484
transform 1 0 53176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input234
timestamp 1666464484
transform -1 0 52440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_357 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 19320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_358
timestamp 1666464484
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_359
timestamp 1666464484
transform -1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_360
timestamp 1666464484
transform 1 0 19872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_361
timestamp 1666464484
transform -1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_362
timestamp 1666464484
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_363
timestamp 1666464484
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_364
timestamp 1666464484
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_365
timestamp 1666464484
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_366
timestamp 1666464484
transform 1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_367
timestamp 1666464484
transform -1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_368
timestamp 1666464484
transform 1 0 54096 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_369
timestamp 1666464484
transform 1 0 54096 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_370
timestamp 1666464484
transform 1 0 54096 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_371
timestamp 1666464484
transform 1 0 54096 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_372
timestamp 1666464484
transform 1 0 52808 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_373
timestamp 1666464484
transform 1 0 33764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_374
timestamp 1666464484
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_375
timestamp 1666464484
transform 1 0 34408 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_376
timestamp 1666464484
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_377
timestamp 1666464484
transform 1 0 35052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_378
timestamp 1666464484
transform 1 0 36156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_379
timestamp 1666464484
transform 1 0 35696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_380
timestamp 1666464484
transform 1 0 36340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_381
timestamp 1666464484
transform 1 0 35972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_382
timestamp 1666464484
transform 1 0 36616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_383
timestamp 1666464484
transform 1 0 36708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output235
timestamp 1666464484
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1666464484
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1666464484
transform -1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1666464484
transform -1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1666464484
transform -1 0 1932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1666464484
transform -1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1666464484
transform -1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1666464484
transform -1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1666464484
transform -1 0 1932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1666464484
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1666464484
transform -1 0 1932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1666464484
transform -1 0 1932 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1666464484
transform -1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1666464484
transform -1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1666464484
transform -1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1666464484
transform -1 0 1932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1666464484
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1666464484
transform -1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1666464484
transform -1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1666464484
transform -1 0 1932 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1666464484
transform -1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1666464484
transform -1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1666464484
transform -1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1666464484
transform -1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1666464484
transform -1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1666464484
transform -1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1666464484
transform -1 0 1932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1666464484
transform -1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1666464484
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1666464484
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1666464484
transform -1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1666464484
transform 1 0 38916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1666464484
transform 1 0 38548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1666464484
transform 1 0 39284 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1666464484
transform 1 0 40020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1666464484
transform -1 0 40388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1666464484
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1666464484
transform -1 0 41124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1666464484
transform 1 0 41492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1666464484
transform -1 0 41860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1666464484
transform -1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1666464484
transform 1 0 42596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1666464484
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1666464484
transform -1 0 43700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1666464484
transform 1 0 44068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output280
timestamp 1666464484
transform 1 0 44068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output281
timestamp 1666464484
transform 1 0 45172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output282
timestamp 1666464484
transform 1 0 44804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output283
timestamp 1666464484
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output284
timestamp 1666464484
transform 1 0 45540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output285
timestamp 1666464484
transform 1 0 46644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output286
timestamp 1666464484
transform 1 0 46276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output287
timestamp 1666464484
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output288
timestamp 1666464484
transform 1 0 47748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output289
timestamp 1666464484
transform -1 0 47012 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output290
timestamp 1666464484
transform -1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output291
timestamp 1666464484
transform -1 0 23736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output292
timestamp 1666464484
transform -1 0 23368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output293
timestamp 1666464484
transform -1 0 24472 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output294
timestamp 1666464484
transform 1 0 23736 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output295
timestamp 1666464484
transform -1 0 25300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output296
timestamp 1666464484
transform 1 0 24840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output297
timestamp 1666464484
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output298
timestamp 1666464484
transform 1 0 25576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output299
timestamp 1666464484
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output300
timestamp 1666464484
transform 1 0 26312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output301
timestamp 1666464484
transform 1 0 26312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output302
timestamp 1666464484
transform -1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output303
timestamp 1666464484
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output304
timestamp 1666464484
transform -1 0 28612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output305
timestamp 1666464484
transform 1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output306
timestamp 1666464484
transform -1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output307
timestamp 1666464484
transform -1 0 29256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output308
timestamp 1666464484
transform -1 0 30820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output309
timestamp 1666464484
transform -1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output310
timestamp 1666464484
transform -1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output311
timestamp 1666464484
transform -1 0 31188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output312
timestamp 1666464484
transform -1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output313
timestamp 1666464484
transform -1 0 32660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output314
timestamp 1666464484
transform -1 0 33396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output315
timestamp 1666464484
transform -1 0 33396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output316
timestamp 1666464484
transform -1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output317
timestamp 1666464484
transform -1 0 1932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output318
timestamp 1666464484
transform -1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output319
timestamp 1666464484
transform -1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output320
timestamp 1666464484
transform -1 0 1932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output321
timestamp 1666464484
transform -1 0 1932 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output322
timestamp 1666464484
transform -1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output323
timestamp 1666464484
transform -1 0 1932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output324
timestamp 1666464484
transform -1 0 1932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output325
timestamp 1666464484
transform -1 0 1932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output326
timestamp 1666464484
transform -1 0 1932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output327
timestamp 1666464484
transform -1 0 54372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output328
timestamp 1666464484
transform 1 0 54004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output329
timestamp 1666464484
transform 1 0 54004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output330
timestamp 1666464484
transform 1 0 54004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output331
timestamp 1666464484
transform 1 0 54004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output332
timestamp 1666464484
transform 1 0 54004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output333
timestamp 1666464484
transform 1 0 54004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output334
timestamp 1666464484
transform 1 0 54004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output335
timestamp 1666464484
transform 1 0 54004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output336
timestamp 1666464484
transform 1 0 54004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output337
timestamp 1666464484
transform 1 0 54004 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output338
timestamp 1666464484
transform 1 0 53268 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output339
timestamp 1666464484
transform 1 0 54004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output340
timestamp 1666464484
transform 1 0 53268 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output341
timestamp 1666464484
transform 1 0 54004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output342
timestamp 1666464484
transform 1 0 54004 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output343
timestamp 1666464484
transform 1 0 53268 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output344
timestamp 1666464484
transform 1 0 54004 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output345
timestamp 1666464484
transform 1 0 54004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output346
timestamp 1666464484
transform 1 0 54004 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output347
timestamp 1666464484
transform 1 0 54004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output348
timestamp 1666464484
transform 1 0 54004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output349
timestamp 1666464484
transform 1 0 54004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output350
timestamp 1666464484
transform 1 0 54004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output351
timestamp 1666464484
transform 1 0 54004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output352
timestamp 1666464484
transform 1 0 54004 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output353
timestamp 1666464484
transform 1 0 54004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output354
timestamp 1666464484
transform 1 0 54004 0 -1 16320
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 design_clk_o
port 0 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 dsi_all[0]
port 1 nsew signal tristate
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 dsi_all[10]
port 2 nsew signal tristate
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 dsi_all[11]
port 3 nsew signal tristate
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 dsi_all[12]
port 4 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 dsi_all[13]
port 5 nsew signal tristate
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 dsi_all[14]
port 6 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 dsi_all[15]
port 7 nsew signal tristate
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 dsi_all[16]
port 8 nsew signal tristate
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 dsi_all[17]
port 9 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 dsi_all[18]
port 10 nsew signal tristate
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 dsi_all[19]
port 11 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 dsi_all[1]
port 12 nsew signal tristate
flabel metal3 s 0 14016 800 14136 0 FreeSans 480 0 0 0 dsi_all[20]
port 13 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 dsi_all[21]
port 14 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 dsi_all[22]
port 15 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 dsi_all[23]
port 16 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 dsi_all[24]
port 17 nsew signal tristate
flabel metal3 s 0 16736 800 16856 0 FreeSans 480 0 0 0 dsi_all[25]
port 18 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 dsi_all[26]
port 19 nsew signal tristate
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 dsi_all[2]
port 20 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 dsi_all[3]
port 21 nsew signal tristate
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 dsi_all[4]
port 22 nsew signal tristate
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 dsi_all[5]
port 23 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 dsi_all[6]
port 24 nsew signal tristate
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 dsi_all[7]
port 25 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 dsi_all[8]
port 26 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 dsi_all[9]
port 27 nsew signal tristate
flabel metal3 s 55200 34552 56000 34672 0 FreeSans 480 0 0 0 dso_6502[0]
port 28 nsew signal input
flabel metal3 s 55200 37272 56000 37392 0 FreeSans 480 0 0 0 dso_6502[10]
port 29 nsew signal input
flabel metal3 s 55200 37544 56000 37664 0 FreeSans 480 0 0 0 dso_6502[11]
port 30 nsew signal input
flabel metal3 s 55200 37816 56000 37936 0 FreeSans 480 0 0 0 dso_6502[12]
port 31 nsew signal input
flabel metal3 s 55200 38088 56000 38208 0 FreeSans 480 0 0 0 dso_6502[13]
port 32 nsew signal input
flabel metal3 s 55200 38360 56000 38480 0 FreeSans 480 0 0 0 dso_6502[14]
port 33 nsew signal input
flabel metal3 s 55200 38632 56000 38752 0 FreeSans 480 0 0 0 dso_6502[15]
port 34 nsew signal input
flabel metal3 s 55200 38904 56000 39024 0 FreeSans 480 0 0 0 dso_6502[16]
port 35 nsew signal input
flabel metal3 s 55200 39176 56000 39296 0 FreeSans 480 0 0 0 dso_6502[17]
port 36 nsew signal input
flabel metal3 s 55200 39448 56000 39568 0 FreeSans 480 0 0 0 dso_6502[18]
port 37 nsew signal input
flabel metal3 s 55200 39720 56000 39840 0 FreeSans 480 0 0 0 dso_6502[19]
port 38 nsew signal input
flabel metal3 s 55200 34824 56000 34944 0 FreeSans 480 0 0 0 dso_6502[1]
port 39 nsew signal input
flabel metal3 s 55200 39992 56000 40112 0 FreeSans 480 0 0 0 dso_6502[20]
port 40 nsew signal input
flabel metal3 s 55200 40264 56000 40384 0 FreeSans 480 0 0 0 dso_6502[21]
port 41 nsew signal input
flabel metal3 s 55200 40536 56000 40656 0 FreeSans 480 0 0 0 dso_6502[22]
port 42 nsew signal input
flabel metal3 s 55200 40808 56000 40928 0 FreeSans 480 0 0 0 dso_6502[23]
port 43 nsew signal input
flabel metal3 s 55200 41080 56000 41200 0 FreeSans 480 0 0 0 dso_6502[24]
port 44 nsew signal input
flabel metal3 s 55200 41352 56000 41472 0 FreeSans 480 0 0 0 dso_6502[25]
port 45 nsew signal input
flabel metal3 s 55200 41624 56000 41744 0 FreeSans 480 0 0 0 dso_6502[26]
port 46 nsew signal input
flabel metal3 s 55200 35096 56000 35216 0 FreeSans 480 0 0 0 dso_6502[2]
port 47 nsew signal input
flabel metal3 s 55200 35368 56000 35488 0 FreeSans 480 0 0 0 dso_6502[3]
port 48 nsew signal input
flabel metal3 s 55200 35640 56000 35760 0 FreeSans 480 0 0 0 dso_6502[4]
port 49 nsew signal input
flabel metal3 s 55200 35912 56000 36032 0 FreeSans 480 0 0 0 dso_6502[5]
port 50 nsew signal input
flabel metal3 s 55200 36184 56000 36304 0 FreeSans 480 0 0 0 dso_6502[6]
port 51 nsew signal input
flabel metal3 s 55200 36456 56000 36576 0 FreeSans 480 0 0 0 dso_6502[7]
port 52 nsew signal input
flabel metal3 s 55200 36728 56000 36848 0 FreeSans 480 0 0 0 dso_6502[8]
port 53 nsew signal input
flabel metal3 s 55200 37000 56000 37120 0 FreeSans 480 0 0 0 dso_6502[9]
port 54 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 dso_LCD[0]
port 55 nsew signal input
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 dso_LCD[1]
port 56 nsew signal input
flabel metal3 s 0 24896 800 25016 0 FreeSans 480 0 0 0 dso_LCD[2]
port 57 nsew signal input
flabel metal3 s 0 25440 800 25560 0 FreeSans 480 0 0 0 dso_LCD[3]
port 58 nsew signal input
flabel metal3 s 0 25984 800 26104 0 FreeSans 480 0 0 0 dso_LCD[4]
port 59 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 dso_LCD[5]
port 60 nsew signal input
flabel metal3 s 0 27072 800 27192 0 FreeSans 480 0 0 0 dso_LCD[6]
port 61 nsew signal input
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 dso_LCD[7]
port 62 nsew signal input
flabel metal3 s 55200 41896 56000 42016 0 FreeSans 480 0 0 0 dso_as1802[0]
port 63 nsew signal input
flabel metal3 s 55200 44616 56000 44736 0 FreeSans 480 0 0 0 dso_as1802[10]
port 64 nsew signal input
flabel metal3 s 55200 44888 56000 45008 0 FreeSans 480 0 0 0 dso_as1802[11]
port 65 nsew signal input
flabel metal3 s 55200 45160 56000 45280 0 FreeSans 480 0 0 0 dso_as1802[12]
port 66 nsew signal input
flabel metal3 s 55200 45432 56000 45552 0 FreeSans 480 0 0 0 dso_as1802[13]
port 67 nsew signal input
flabel metal3 s 55200 45704 56000 45824 0 FreeSans 480 0 0 0 dso_as1802[14]
port 68 nsew signal input
flabel metal3 s 55200 45976 56000 46096 0 FreeSans 480 0 0 0 dso_as1802[15]
port 69 nsew signal input
flabel metal3 s 55200 46248 56000 46368 0 FreeSans 480 0 0 0 dso_as1802[16]
port 70 nsew signal input
flabel metal3 s 55200 46520 56000 46640 0 FreeSans 480 0 0 0 dso_as1802[17]
port 71 nsew signal input
flabel metal3 s 55200 46792 56000 46912 0 FreeSans 480 0 0 0 dso_as1802[18]
port 72 nsew signal input
flabel metal3 s 55200 47064 56000 47184 0 FreeSans 480 0 0 0 dso_as1802[19]
port 73 nsew signal input
flabel metal3 s 55200 42168 56000 42288 0 FreeSans 480 0 0 0 dso_as1802[1]
port 74 nsew signal input
flabel metal3 s 55200 47336 56000 47456 0 FreeSans 480 0 0 0 dso_as1802[20]
port 75 nsew signal input
flabel metal3 s 55200 47608 56000 47728 0 FreeSans 480 0 0 0 dso_as1802[21]
port 76 nsew signal input
flabel metal3 s 55200 47880 56000 48000 0 FreeSans 480 0 0 0 dso_as1802[22]
port 77 nsew signal input
flabel metal3 s 55200 48152 56000 48272 0 FreeSans 480 0 0 0 dso_as1802[23]
port 78 nsew signal input
flabel metal3 s 55200 48424 56000 48544 0 FreeSans 480 0 0 0 dso_as1802[24]
port 79 nsew signal input
flabel metal3 s 55200 48696 56000 48816 0 FreeSans 480 0 0 0 dso_as1802[25]
port 80 nsew signal input
flabel metal3 s 55200 48968 56000 49088 0 FreeSans 480 0 0 0 dso_as1802[26]
port 81 nsew signal input
flabel metal3 s 55200 42440 56000 42560 0 FreeSans 480 0 0 0 dso_as1802[2]
port 82 nsew signal input
flabel metal3 s 55200 42712 56000 42832 0 FreeSans 480 0 0 0 dso_as1802[3]
port 83 nsew signal input
flabel metal3 s 55200 42984 56000 43104 0 FreeSans 480 0 0 0 dso_as1802[4]
port 84 nsew signal input
flabel metal3 s 55200 43256 56000 43376 0 FreeSans 480 0 0 0 dso_as1802[5]
port 85 nsew signal input
flabel metal3 s 55200 43528 56000 43648 0 FreeSans 480 0 0 0 dso_as1802[6]
port 86 nsew signal input
flabel metal3 s 55200 43800 56000 43920 0 FreeSans 480 0 0 0 dso_as1802[7]
port 87 nsew signal input
flabel metal3 s 55200 44072 56000 44192 0 FreeSans 480 0 0 0 dso_as1802[8]
port 88 nsew signal input
flabel metal3 s 55200 44344 56000 44464 0 FreeSans 480 0 0 0 dso_as1802[9]
port 89 nsew signal input
flabel metal3 s 0 38496 800 38616 0 FreeSans 480 0 0 0 dso_as2650[0]
port 90 nsew signal input
flabel metal3 s 0 43936 800 44056 0 FreeSans 480 0 0 0 dso_as2650[10]
port 91 nsew signal input
flabel metal3 s 0 44480 800 44600 0 FreeSans 480 0 0 0 dso_as2650[11]
port 92 nsew signal input
flabel metal3 s 0 45024 800 45144 0 FreeSans 480 0 0 0 dso_as2650[12]
port 93 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 dso_as2650[13]
port 94 nsew signal input
flabel metal3 s 0 46112 800 46232 0 FreeSans 480 0 0 0 dso_as2650[14]
port 95 nsew signal input
flabel metal3 s 0 46656 800 46776 0 FreeSans 480 0 0 0 dso_as2650[15]
port 96 nsew signal input
flabel metal3 s 0 47200 800 47320 0 FreeSans 480 0 0 0 dso_as2650[16]
port 97 nsew signal input
flabel metal3 s 0 47744 800 47864 0 FreeSans 480 0 0 0 dso_as2650[17]
port 98 nsew signal input
flabel metal3 s 0 48288 800 48408 0 FreeSans 480 0 0 0 dso_as2650[18]
port 99 nsew signal input
flabel metal3 s 0 48832 800 48952 0 FreeSans 480 0 0 0 dso_as2650[19]
port 100 nsew signal input
flabel metal3 s 0 39040 800 39160 0 FreeSans 480 0 0 0 dso_as2650[1]
port 101 nsew signal input
flabel metal3 s 0 49376 800 49496 0 FreeSans 480 0 0 0 dso_as2650[20]
port 102 nsew signal input
flabel metal3 s 0 49920 800 50040 0 FreeSans 480 0 0 0 dso_as2650[21]
port 103 nsew signal input
flabel metal3 s 0 50464 800 50584 0 FreeSans 480 0 0 0 dso_as2650[22]
port 104 nsew signal input
flabel metal3 s 0 51008 800 51128 0 FreeSans 480 0 0 0 dso_as2650[23]
port 105 nsew signal input
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 dso_as2650[24]
port 106 nsew signal input
flabel metal3 s 0 52096 800 52216 0 FreeSans 480 0 0 0 dso_as2650[25]
port 107 nsew signal input
flabel metal3 s 0 52640 800 52760 0 FreeSans 480 0 0 0 dso_as2650[26]
port 108 nsew signal input
flabel metal3 s 0 39584 800 39704 0 FreeSans 480 0 0 0 dso_as2650[2]
port 109 nsew signal input
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 dso_as2650[3]
port 110 nsew signal input
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 dso_as2650[4]
port 111 nsew signal input
flabel metal3 s 0 41216 800 41336 0 FreeSans 480 0 0 0 dso_as2650[5]
port 112 nsew signal input
flabel metal3 s 0 41760 800 41880 0 FreeSans 480 0 0 0 dso_as2650[6]
port 113 nsew signal input
flabel metal3 s 0 42304 800 42424 0 FreeSans 480 0 0 0 dso_as2650[7]
port 114 nsew signal input
flabel metal3 s 0 42848 800 42968 0 FreeSans 480 0 0 0 dso_as2650[8]
port 115 nsew signal input
flabel metal3 s 0 43392 800 43512 0 FreeSans 480 0 0 0 dso_as2650[9]
port 116 nsew signal input
flabel metal2 s 11242 55200 11298 56000 0 FreeSans 224 90 0 0 dso_as5401[0]
port 117 nsew signal input
flabel metal2 s 23202 55200 23258 56000 0 FreeSans 224 90 0 0 dso_as5401[10]
port 118 nsew signal input
flabel metal2 s 24398 55200 24454 56000 0 FreeSans 224 90 0 0 dso_as5401[11]
port 119 nsew signal input
flabel metal2 s 25594 55200 25650 56000 0 FreeSans 224 90 0 0 dso_as5401[12]
port 120 nsew signal input
flabel metal2 s 26790 55200 26846 56000 0 FreeSans 224 90 0 0 dso_as5401[13]
port 121 nsew signal input
flabel metal2 s 27986 55200 28042 56000 0 FreeSans 224 90 0 0 dso_as5401[14]
port 122 nsew signal input
flabel metal2 s 29182 55200 29238 56000 0 FreeSans 224 90 0 0 dso_as5401[15]
port 123 nsew signal input
flabel metal2 s 30378 55200 30434 56000 0 FreeSans 224 90 0 0 dso_as5401[16]
port 124 nsew signal input
flabel metal2 s 31574 55200 31630 56000 0 FreeSans 224 90 0 0 dso_as5401[17]
port 125 nsew signal input
flabel metal2 s 32770 55200 32826 56000 0 FreeSans 224 90 0 0 dso_as5401[18]
port 126 nsew signal input
flabel metal2 s 33966 55200 34022 56000 0 FreeSans 224 90 0 0 dso_as5401[19]
port 127 nsew signal input
flabel metal2 s 12438 55200 12494 56000 0 FreeSans 224 90 0 0 dso_as5401[1]
port 128 nsew signal input
flabel metal2 s 35162 55200 35218 56000 0 FreeSans 224 90 0 0 dso_as5401[20]
port 129 nsew signal input
flabel metal2 s 36358 55200 36414 56000 0 FreeSans 224 90 0 0 dso_as5401[21]
port 130 nsew signal input
flabel metal2 s 37554 55200 37610 56000 0 FreeSans 224 90 0 0 dso_as5401[22]
port 131 nsew signal input
flabel metal2 s 38750 55200 38806 56000 0 FreeSans 224 90 0 0 dso_as5401[23]
port 132 nsew signal input
flabel metal2 s 39946 55200 40002 56000 0 FreeSans 224 90 0 0 dso_as5401[24]
port 133 nsew signal input
flabel metal2 s 41142 55200 41198 56000 0 FreeSans 224 90 0 0 dso_as5401[25]
port 134 nsew signal input
flabel metal2 s 42338 55200 42394 56000 0 FreeSans 224 90 0 0 dso_as5401[26]
port 135 nsew signal input
flabel metal2 s 13634 55200 13690 56000 0 FreeSans 224 90 0 0 dso_as5401[2]
port 136 nsew signal input
flabel metal2 s 14830 55200 14886 56000 0 FreeSans 224 90 0 0 dso_as5401[3]
port 137 nsew signal input
flabel metal2 s 16026 55200 16082 56000 0 FreeSans 224 90 0 0 dso_as5401[4]
port 138 nsew signal input
flabel metal2 s 17222 55200 17278 56000 0 FreeSans 224 90 0 0 dso_as5401[5]
port 139 nsew signal input
flabel metal2 s 18418 55200 18474 56000 0 FreeSans 224 90 0 0 dso_as5401[6]
port 140 nsew signal input
flabel metal2 s 19614 55200 19670 56000 0 FreeSans 224 90 0 0 dso_as5401[7]
port 141 nsew signal input
flabel metal2 s 20810 55200 20866 56000 0 FreeSans 224 90 0 0 dso_as5401[8]
port 142 nsew signal input
flabel metal2 s 22006 55200 22062 56000 0 FreeSans 224 90 0 0 dso_as5401[9]
port 143 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 dso_counter[0]
port 144 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 dso_counter[10]
port 145 nsew signal input
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 dso_counter[11]
port 146 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 dso_counter[1]
port 147 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 dso_counter[2]
port 148 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 dso_counter[3]
port 149 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 dso_counter[4]
port 150 nsew signal input
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 dso_counter[5]
port 151 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 dso_counter[6]
port 152 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 dso_counter[7]
port 153 nsew signal input
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 dso_counter[8]
port 154 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 dso_counter[9]
port 155 nsew signal input
flabel metal2 s 44730 55200 44786 56000 0 FreeSans 224 90 0 0 dso_diceroll[0]
port 156 nsew signal input
flabel metal2 s 45926 55200 45982 56000 0 FreeSans 224 90 0 0 dso_diceroll[1]
port 157 nsew signal input
flabel metal2 s 47122 55200 47178 56000 0 FreeSans 224 90 0 0 dso_diceroll[2]
port 158 nsew signal input
flabel metal2 s 48318 55200 48374 56000 0 FreeSans 224 90 0 0 dso_diceroll[3]
port 159 nsew signal input
flabel metal2 s 49514 55200 49570 56000 0 FreeSans 224 90 0 0 dso_diceroll[4]
port 160 nsew signal input
flabel metal2 s 50710 55200 50766 56000 0 FreeSans 224 90 0 0 dso_diceroll[5]
port 161 nsew signal input
flabel metal2 s 51906 55200 51962 56000 0 FreeSans 224 90 0 0 dso_diceroll[6]
port 162 nsew signal input
flabel metal2 s 53102 55200 53158 56000 0 FreeSans 224 90 0 0 dso_diceroll[7]
port 163 nsew signal input
flabel metal3 s 0 28160 800 28280 0 FreeSans 480 0 0 0 dso_mc14500[0]
port 164 nsew signal input
flabel metal3 s 0 28704 800 28824 0 FreeSans 480 0 0 0 dso_mc14500[1]
port 165 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 dso_mc14500[2]
port 166 nsew signal input
flabel metal3 s 0 29792 800 29912 0 FreeSans 480 0 0 0 dso_mc14500[3]
port 167 nsew signal input
flabel metal3 s 0 30336 800 30456 0 FreeSans 480 0 0 0 dso_mc14500[4]
port 168 nsew signal input
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 dso_mc14500[5]
port 169 nsew signal input
flabel metal3 s 0 31424 800 31544 0 FreeSans 480 0 0 0 dso_mc14500[6]
port 170 nsew signal input
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 dso_mc14500[7]
port 171 nsew signal input
flabel metal3 s 0 32512 800 32632 0 FreeSans 480 0 0 0 dso_mc14500[8]
port 172 nsew signal input
flabel metal2 s 1674 55200 1730 56000 0 FreeSans 224 90 0 0 dso_multiplier[0]
port 173 nsew signal input
flabel metal2 s 2870 55200 2926 56000 0 FreeSans 224 90 0 0 dso_multiplier[1]
port 174 nsew signal input
flabel metal2 s 4066 55200 4122 56000 0 FreeSans 224 90 0 0 dso_multiplier[2]
port 175 nsew signal input
flabel metal2 s 5262 55200 5318 56000 0 FreeSans 224 90 0 0 dso_multiplier[3]
port 176 nsew signal input
flabel metal2 s 6458 55200 6514 56000 0 FreeSans 224 90 0 0 dso_multiplier[4]
port 177 nsew signal input
flabel metal2 s 7654 55200 7710 56000 0 FreeSans 224 90 0 0 dso_multiplier[5]
port 178 nsew signal input
flabel metal2 s 8850 55200 8906 56000 0 FreeSans 224 90 0 0 dso_multiplier[6]
port 179 nsew signal input
flabel metal2 s 10046 55200 10102 56000 0 FreeSans 224 90 0 0 dso_multiplier[7]
port 180 nsew signal input
flabel metal3 s 0 33600 800 33720 0 FreeSans 480 0 0 0 dso_tbb1143[0]
port 181 nsew signal input
flabel metal3 s 0 34144 800 34264 0 FreeSans 480 0 0 0 dso_tbb1143[1]
port 182 nsew signal input
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 dso_tbb1143[2]
port 183 nsew signal input
flabel metal3 s 0 35232 800 35352 0 FreeSans 480 0 0 0 dso_tbb1143[3]
port 184 nsew signal input
flabel metal3 s 0 35776 800 35896 0 FreeSans 480 0 0 0 dso_tbb1143[4]
port 185 nsew signal input
flabel metal3 s 0 36320 800 36440 0 FreeSans 480 0 0 0 dso_tbb1143[5]
port 186 nsew signal input
flabel metal3 s 0 36864 800 36984 0 FreeSans 480 0 0 0 dso_tbb1143[6]
port 187 nsew signal input
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 dso_tbb1143[7]
port 188 nsew signal input
flabel metal2 s 54298 55200 54354 56000 0 FreeSans 224 90 0 0 dso_tune
port 189 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 io_in[0]
port 190 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 io_in[10]
port 191 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 io_in[11]
port 192 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 io_in[12]
port 193 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 io_in[13]
port 194 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 io_in[14]
port 195 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 io_in[15]
port 196 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 io_in[16]
port 197 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 io_in[17]
port 198 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 io_in[18]
port 199 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 io_in[19]
port 200 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 io_in[1]
port 201 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 io_in[20]
port 202 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 io_in[21]
port 203 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 io_in[22]
port 204 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 io_in[23]
port 205 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 io_in[24]
port 206 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 io_in[25]
port 207 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 io_in[26]
port 208 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 io_in[27]
port 209 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 io_in[28]
port 210 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 io_in[29]
port 211 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 io_in[2]
port 212 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 io_in[30]
port 213 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 io_in[31]
port 214 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 io_in[32]
port 215 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 io_in[33]
port 216 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 io_in[34]
port 217 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 io_in[35]
port 218 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 io_in[36]
port 219 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 io_in[37]
port 220 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 io_in[3]
port 221 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 io_in[4]
port 222 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 io_in[5]
port 223 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 io_in[6]
port 224 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 io_in[7]
port 225 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 io_in[8]
port 226 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 io_in[9]
port 227 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 228 nsew signal tristate
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 229 nsew signal tristate
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 230 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 231 nsew signal tristate
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 232 nsew signal tristate
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 233 nsew signal tristate
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 234 nsew signal tristate
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 235 nsew signal tristate
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 236 nsew signal tristate
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 237 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 238 nsew signal tristate
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 239 nsew signal tristate
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 240 nsew signal tristate
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 241 nsew signal tristate
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 242 nsew signal tristate
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 243 nsew signal tristate
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 244 nsew signal tristate
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 245 nsew signal tristate
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 246 nsew signal tristate
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 247 nsew signal tristate
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 248 nsew signal tristate
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 249 nsew signal tristate
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 250 nsew signal tristate
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 251 nsew signal tristate
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 252 nsew signal tristate
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 253 nsew signal tristate
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 254 nsew signal tristate
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 255 nsew signal tristate
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 256 nsew signal tristate
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 257 nsew signal tristate
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 258 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 259 nsew signal tristate
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 260 nsew signal tristate
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 261 nsew signal tristate
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 262 nsew signal tristate
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 263 nsew signal tristate
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 264 nsew signal tristate
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 265 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 io_out[0]
port 266 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 io_out[10]
port 267 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 io_out[11]
port 268 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 io_out[12]
port 269 nsew signal tristate
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 io_out[13]
port 270 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 io_out[14]
port 271 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 io_out[15]
port 272 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 io_out[16]
port 273 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 io_out[17]
port 274 nsew signal tristate
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 io_out[18]
port 275 nsew signal tristate
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 io_out[19]
port 276 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 io_out[1]
port 277 nsew signal tristate
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 io_out[20]
port 278 nsew signal tristate
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 io_out[21]
port 279 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 io_out[22]
port 280 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 io_out[23]
port 281 nsew signal tristate
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 io_out[24]
port 282 nsew signal tristate
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 io_out[25]
port 283 nsew signal tristate
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 io_out[26]
port 284 nsew signal tristate
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 io_out[27]
port 285 nsew signal tristate
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 io_out[28]
port 286 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 io_out[29]
port 287 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 io_out[2]
port 288 nsew signal tristate
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 io_out[30]
port 289 nsew signal tristate
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 io_out[31]
port 290 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 io_out[32]
port 291 nsew signal tristate
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 io_out[33]
port 292 nsew signal tristate
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 io_out[34]
port 293 nsew signal tristate
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 io_out[35]
port 294 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 io_out[36]
port 295 nsew signal tristate
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 io_out[37]
port 296 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 io_out[3]
port 297 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 io_out[4]
port 298 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 io_out[5]
port 299 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 io_out[6]
port 300 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 io_out[7]
port 301 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 io_out[8]
port 302 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 io_out[9]
port 303 nsew signal tristate
flabel metal3 s 55200 34280 56000 34400 0 FreeSans 480 0 0 0 oeb_6502
port 304 nsew signal input
flabel metal3 s 55200 49240 56000 49360 0 FreeSans 480 0 0 0 oeb_as1802
port 305 nsew signal input
flabel metal3 s 0 37952 800 38072 0 FreeSans 480 0 0 0 oeb_as2650
port 306 nsew signal input
flabel metal2 s 43534 55200 43590 56000 0 FreeSans 224 90 0 0 oeb_as5401
port 307 nsew signal input
flabel metal3 s 0 33056 800 33176 0 FreeSans 480 0 0 0 oeb_mc14500
port 308 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 rst_6502
port 309 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 rst_LCD
port 310 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 rst_as1802
port 311 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 rst_as2650
port 312 nsew signal tristate
flabel metal3 s 0 20544 800 20664 0 FreeSans 480 0 0 0 rst_as5401
port 313 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 rst_counter
port 314 nsew signal tristate
flabel metal3 s 0 21632 800 21752 0 FreeSans 480 0 0 0 rst_diceroll
port 315 nsew signal tristate
flabel metal3 s 0 22176 800 22296 0 FreeSans 480 0 0 0 rst_mc14500
port 316 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 rst_tbb1143
port 317 nsew signal tristate
flabel metal3 s 0 23264 800 23384 0 FreeSans 480 0 0 0 rst_tune
port 318 nsew signal tristate
flabel metal4 s 4208 2128 4528 53360 0 FreeSans 1920 90 0 0 vccd1
port 319 nsew power bidirectional
flabel metal4 s 34928 2128 35248 53360 0 FreeSans 1920 90 0 0 vccd1
port 319 nsew power bidirectional
flabel metal4 s 19568 2128 19888 53360 0 FreeSans 1920 90 0 0 vssd1
port 320 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 53360 0 FreeSans 1920 90 0 0 vssd1
port 320 nsew ground bidirectional
flabel metal3 s 55200 6536 56000 6656 0 FreeSans 480 0 0 0 wb_clk_i
port 321 nsew signal input
flabel metal3 s 55200 6808 56000 6928 0 FreeSans 480 0 0 0 wb_rst_i
port 322 nsew signal input
flabel metal3 s 55200 7080 56000 7200 0 FreeSans 480 0 0 0 wbs_ack_o
port 323 nsew signal tristate
flabel metal3 s 55200 8168 56000 8288 0 FreeSans 480 0 0 0 wbs_adr_i[0]
port 324 nsew signal input
flabel metal3 s 55200 16328 56000 16448 0 FreeSans 480 0 0 0 wbs_adr_i[10]
port 325 nsew signal input
flabel metal3 s 55200 17144 56000 17264 0 FreeSans 480 0 0 0 wbs_adr_i[11]
port 326 nsew signal input
flabel metal3 s 55200 17960 56000 18080 0 FreeSans 480 0 0 0 wbs_adr_i[12]
port 327 nsew signal input
flabel metal3 s 55200 18776 56000 18896 0 FreeSans 480 0 0 0 wbs_adr_i[13]
port 328 nsew signal input
flabel metal3 s 55200 19592 56000 19712 0 FreeSans 480 0 0 0 wbs_adr_i[14]
port 329 nsew signal input
flabel metal3 s 55200 20408 56000 20528 0 FreeSans 480 0 0 0 wbs_adr_i[15]
port 330 nsew signal input
flabel metal3 s 55200 21224 56000 21344 0 FreeSans 480 0 0 0 wbs_adr_i[16]
port 331 nsew signal input
flabel metal3 s 55200 22040 56000 22160 0 FreeSans 480 0 0 0 wbs_adr_i[17]
port 332 nsew signal input
flabel metal3 s 55200 22856 56000 22976 0 FreeSans 480 0 0 0 wbs_adr_i[18]
port 333 nsew signal input
flabel metal3 s 55200 23672 56000 23792 0 FreeSans 480 0 0 0 wbs_adr_i[19]
port 334 nsew signal input
flabel metal3 s 55200 8984 56000 9104 0 FreeSans 480 0 0 0 wbs_adr_i[1]
port 335 nsew signal input
flabel metal3 s 55200 24488 56000 24608 0 FreeSans 480 0 0 0 wbs_adr_i[20]
port 336 nsew signal input
flabel metal3 s 55200 25304 56000 25424 0 FreeSans 480 0 0 0 wbs_adr_i[21]
port 337 nsew signal input
flabel metal3 s 55200 26120 56000 26240 0 FreeSans 480 0 0 0 wbs_adr_i[22]
port 338 nsew signal input
flabel metal3 s 55200 26936 56000 27056 0 FreeSans 480 0 0 0 wbs_adr_i[23]
port 339 nsew signal input
flabel metal3 s 55200 27752 56000 27872 0 FreeSans 480 0 0 0 wbs_adr_i[24]
port 340 nsew signal input
flabel metal3 s 55200 28568 56000 28688 0 FreeSans 480 0 0 0 wbs_adr_i[25]
port 341 nsew signal input
flabel metal3 s 55200 29384 56000 29504 0 FreeSans 480 0 0 0 wbs_adr_i[26]
port 342 nsew signal input
flabel metal3 s 55200 30200 56000 30320 0 FreeSans 480 0 0 0 wbs_adr_i[27]
port 343 nsew signal input
flabel metal3 s 55200 31016 56000 31136 0 FreeSans 480 0 0 0 wbs_adr_i[28]
port 344 nsew signal input
flabel metal3 s 55200 31832 56000 31952 0 FreeSans 480 0 0 0 wbs_adr_i[29]
port 345 nsew signal input
flabel metal3 s 55200 9800 56000 9920 0 FreeSans 480 0 0 0 wbs_adr_i[2]
port 346 nsew signal input
flabel metal3 s 55200 32648 56000 32768 0 FreeSans 480 0 0 0 wbs_adr_i[30]
port 347 nsew signal input
flabel metal3 s 55200 33464 56000 33584 0 FreeSans 480 0 0 0 wbs_adr_i[31]
port 348 nsew signal input
flabel metal3 s 55200 10616 56000 10736 0 FreeSans 480 0 0 0 wbs_adr_i[3]
port 349 nsew signal input
flabel metal3 s 55200 11432 56000 11552 0 FreeSans 480 0 0 0 wbs_adr_i[4]
port 350 nsew signal input
flabel metal3 s 55200 12248 56000 12368 0 FreeSans 480 0 0 0 wbs_adr_i[5]
port 351 nsew signal input
flabel metal3 s 55200 13064 56000 13184 0 FreeSans 480 0 0 0 wbs_adr_i[6]
port 352 nsew signal input
flabel metal3 s 55200 13880 56000 14000 0 FreeSans 480 0 0 0 wbs_adr_i[7]
port 353 nsew signal input
flabel metal3 s 55200 14696 56000 14816 0 FreeSans 480 0 0 0 wbs_adr_i[8]
port 354 nsew signal input
flabel metal3 s 55200 15512 56000 15632 0 FreeSans 480 0 0 0 wbs_adr_i[9]
port 355 nsew signal input
flabel metal3 s 55200 7352 56000 7472 0 FreeSans 480 0 0 0 wbs_cyc_i
port 356 nsew signal input
flabel metal3 s 55200 8440 56000 8560 0 FreeSans 480 0 0 0 wbs_dat_i[0]
port 357 nsew signal input
flabel metal3 s 55200 16600 56000 16720 0 FreeSans 480 0 0 0 wbs_dat_i[10]
port 358 nsew signal input
flabel metal3 s 55200 17416 56000 17536 0 FreeSans 480 0 0 0 wbs_dat_i[11]
port 359 nsew signal input
flabel metal3 s 55200 18232 56000 18352 0 FreeSans 480 0 0 0 wbs_dat_i[12]
port 360 nsew signal input
flabel metal3 s 55200 19048 56000 19168 0 FreeSans 480 0 0 0 wbs_dat_i[13]
port 361 nsew signal input
flabel metal3 s 55200 19864 56000 19984 0 FreeSans 480 0 0 0 wbs_dat_i[14]
port 362 nsew signal input
flabel metal3 s 55200 20680 56000 20800 0 FreeSans 480 0 0 0 wbs_dat_i[15]
port 363 nsew signal input
flabel metal3 s 55200 21496 56000 21616 0 FreeSans 480 0 0 0 wbs_dat_i[16]
port 364 nsew signal input
flabel metal3 s 55200 22312 56000 22432 0 FreeSans 480 0 0 0 wbs_dat_i[17]
port 365 nsew signal input
flabel metal3 s 55200 23128 56000 23248 0 FreeSans 480 0 0 0 wbs_dat_i[18]
port 366 nsew signal input
flabel metal3 s 55200 23944 56000 24064 0 FreeSans 480 0 0 0 wbs_dat_i[19]
port 367 nsew signal input
flabel metal3 s 55200 9256 56000 9376 0 FreeSans 480 0 0 0 wbs_dat_i[1]
port 368 nsew signal input
flabel metal3 s 55200 24760 56000 24880 0 FreeSans 480 0 0 0 wbs_dat_i[20]
port 369 nsew signal input
flabel metal3 s 55200 25576 56000 25696 0 FreeSans 480 0 0 0 wbs_dat_i[21]
port 370 nsew signal input
flabel metal3 s 55200 26392 56000 26512 0 FreeSans 480 0 0 0 wbs_dat_i[22]
port 371 nsew signal input
flabel metal3 s 55200 27208 56000 27328 0 FreeSans 480 0 0 0 wbs_dat_i[23]
port 372 nsew signal input
flabel metal3 s 55200 28024 56000 28144 0 FreeSans 480 0 0 0 wbs_dat_i[24]
port 373 nsew signal input
flabel metal3 s 55200 28840 56000 28960 0 FreeSans 480 0 0 0 wbs_dat_i[25]
port 374 nsew signal input
flabel metal3 s 55200 29656 56000 29776 0 FreeSans 480 0 0 0 wbs_dat_i[26]
port 375 nsew signal input
flabel metal3 s 55200 30472 56000 30592 0 FreeSans 480 0 0 0 wbs_dat_i[27]
port 376 nsew signal input
flabel metal3 s 55200 31288 56000 31408 0 FreeSans 480 0 0 0 wbs_dat_i[28]
port 377 nsew signal input
flabel metal3 s 55200 32104 56000 32224 0 FreeSans 480 0 0 0 wbs_dat_i[29]
port 378 nsew signal input
flabel metal3 s 55200 10072 56000 10192 0 FreeSans 480 0 0 0 wbs_dat_i[2]
port 379 nsew signal input
flabel metal3 s 55200 32920 56000 33040 0 FreeSans 480 0 0 0 wbs_dat_i[30]
port 380 nsew signal input
flabel metal3 s 55200 33736 56000 33856 0 FreeSans 480 0 0 0 wbs_dat_i[31]
port 381 nsew signal input
flabel metal3 s 55200 10888 56000 11008 0 FreeSans 480 0 0 0 wbs_dat_i[3]
port 382 nsew signal input
flabel metal3 s 55200 11704 56000 11824 0 FreeSans 480 0 0 0 wbs_dat_i[4]
port 383 nsew signal input
flabel metal3 s 55200 12520 56000 12640 0 FreeSans 480 0 0 0 wbs_dat_i[5]
port 384 nsew signal input
flabel metal3 s 55200 13336 56000 13456 0 FreeSans 480 0 0 0 wbs_dat_i[6]
port 385 nsew signal input
flabel metal3 s 55200 14152 56000 14272 0 FreeSans 480 0 0 0 wbs_dat_i[7]
port 386 nsew signal input
flabel metal3 s 55200 14968 56000 15088 0 FreeSans 480 0 0 0 wbs_dat_i[8]
port 387 nsew signal input
flabel metal3 s 55200 15784 56000 15904 0 FreeSans 480 0 0 0 wbs_dat_i[9]
port 388 nsew signal input
flabel metal3 s 55200 8712 56000 8832 0 FreeSans 480 0 0 0 wbs_dat_o[0]
port 389 nsew signal tristate
flabel metal3 s 55200 16872 56000 16992 0 FreeSans 480 0 0 0 wbs_dat_o[10]
port 390 nsew signal tristate
flabel metal3 s 55200 17688 56000 17808 0 FreeSans 480 0 0 0 wbs_dat_o[11]
port 391 nsew signal tristate
flabel metal3 s 55200 18504 56000 18624 0 FreeSans 480 0 0 0 wbs_dat_o[12]
port 392 nsew signal tristate
flabel metal3 s 55200 19320 56000 19440 0 FreeSans 480 0 0 0 wbs_dat_o[13]
port 393 nsew signal tristate
flabel metal3 s 55200 20136 56000 20256 0 FreeSans 480 0 0 0 wbs_dat_o[14]
port 394 nsew signal tristate
flabel metal3 s 55200 20952 56000 21072 0 FreeSans 480 0 0 0 wbs_dat_o[15]
port 395 nsew signal tristate
flabel metal3 s 55200 21768 56000 21888 0 FreeSans 480 0 0 0 wbs_dat_o[16]
port 396 nsew signal tristate
flabel metal3 s 55200 22584 56000 22704 0 FreeSans 480 0 0 0 wbs_dat_o[17]
port 397 nsew signal tristate
flabel metal3 s 55200 23400 56000 23520 0 FreeSans 480 0 0 0 wbs_dat_o[18]
port 398 nsew signal tristate
flabel metal3 s 55200 24216 56000 24336 0 FreeSans 480 0 0 0 wbs_dat_o[19]
port 399 nsew signal tristate
flabel metal3 s 55200 9528 56000 9648 0 FreeSans 480 0 0 0 wbs_dat_o[1]
port 400 nsew signal tristate
flabel metal3 s 55200 25032 56000 25152 0 FreeSans 480 0 0 0 wbs_dat_o[20]
port 401 nsew signal tristate
flabel metal3 s 55200 25848 56000 25968 0 FreeSans 480 0 0 0 wbs_dat_o[21]
port 402 nsew signal tristate
flabel metal3 s 55200 26664 56000 26784 0 FreeSans 480 0 0 0 wbs_dat_o[22]
port 403 nsew signal tristate
flabel metal3 s 55200 27480 56000 27600 0 FreeSans 480 0 0 0 wbs_dat_o[23]
port 404 nsew signal tristate
flabel metal3 s 55200 28296 56000 28416 0 FreeSans 480 0 0 0 wbs_dat_o[24]
port 405 nsew signal tristate
flabel metal3 s 55200 29112 56000 29232 0 FreeSans 480 0 0 0 wbs_dat_o[25]
port 406 nsew signal tristate
flabel metal3 s 55200 29928 56000 30048 0 FreeSans 480 0 0 0 wbs_dat_o[26]
port 407 nsew signal tristate
flabel metal3 s 55200 30744 56000 30864 0 FreeSans 480 0 0 0 wbs_dat_o[27]
port 408 nsew signal tristate
flabel metal3 s 55200 31560 56000 31680 0 FreeSans 480 0 0 0 wbs_dat_o[28]
port 409 nsew signal tristate
flabel metal3 s 55200 32376 56000 32496 0 FreeSans 480 0 0 0 wbs_dat_o[29]
port 410 nsew signal tristate
flabel metal3 s 55200 10344 56000 10464 0 FreeSans 480 0 0 0 wbs_dat_o[2]
port 411 nsew signal tristate
flabel metal3 s 55200 33192 56000 33312 0 FreeSans 480 0 0 0 wbs_dat_o[30]
port 412 nsew signal tristate
flabel metal3 s 55200 34008 56000 34128 0 FreeSans 480 0 0 0 wbs_dat_o[31]
port 413 nsew signal tristate
flabel metal3 s 55200 11160 56000 11280 0 FreeSans 480 0 0 0 wbs_dat_o[3]
port 414 nsew signal tristate
flabel metal3 s 55200 11976 56000 12096 0 FreeSans 480 0 0 0 wbs_dat_o[4]
port 415 nsew signal tristate
flabel metal3 s 55200 12792 56000 12912 0 FreeSans 480 0 0 0 wbs_dat_o[5]
port 416 nsew signal tristate
flabel metal3 s 55200 13608 56000 13728 0 FreeSans 480 0 0 0 wbs_dat_o[6]
port 417 nsew signal tristate
flabel metal3 s 55200 14424 56000 14544 0 FreeSans 480 0 0 0 wbs_dat_o[7]
port 418 nsew signal tristate
flabel metal3 s 55200 15240 56000 15360 0 FreeSans 480 0 0 0 wbs_dat_o[8]
port 419 nsew signal tristate
flabel metal3 s 55200 16056 56000 16176 0 FreeSans 480 0 0 0 wbs_dat_o[9]
port 420 nsew signal tristate
flabel metal3 s 55200 7624 56000 7744 0 FreeSans 480 0 0 0 wbs_stb_i
port 421 nsew signal input
flabel metal3 s 55200 7896 56000 8016 0 FreeSans 480 0 0 0 wbs_we_i
port 422 nsew signal input
rlabel metal1 27968 52768 27968 52768 0 vccd1
rlabel metal1 27968 53312 27968 53312 0 vssd1
rlabel metal1 38216 9554 38216 9554 0 _0000_
rlabel metal1 36887 9962 36887 9962 0 _0001_
rlabel metal1 38456 10234 38456 10234 0 _0002_
rlabel metal2 40066 11526 40066 11526 0 _0003_
rlabel metal2 36018 11526 36018 11526 0 _0004_
rlabel metal1 38492 12818 38492 12818 0 _0005_
rlabel metal1 40112 12954 40112 12954 0 _0006_
rlabel metal2 40802 13906 40802 13906 0 _0007_
rlabel metal1 39514 14892 39514 14892 0 _0008_
rlabel metal1 43194 15368 43194 15368 0 _0009_
rlabel metal1 41287 16558 41287 16558 0 _0010_
rlabel metal1 40449 17238 40449 17238 0 _0011_
rlabel metal1 39146 18088 39146 18088 0 _0012_
rlabel metal1 41492 17782 41492 17782 0 _0013_
rlabel metal1 41492 19482 41492 19482 0 _0014_
rlabel metal1 43286 20808 43286 20808 0 _0015_
rlabel metal1 42688 20774 42688 20774 0 _0016_
rlabel metal1 42642 22542 42642 22542 0 _0017_
rlabel metal1 42826 22984 42826 22984 0 _0018_
rlabel metal1 40786 23766 40786 23766 0 _0019_
rlabel metal1 40240 24174 40240 24174 0 _0020_
rlabel via1 38681 24786 38681 24786 0 _0021_
rlabel metal1 38256 23766 38256 23766 0 _0022_
rlabel metal1 36928 24174 36928 24174 0 _0023_
rlabel metal1 33610 24854 33610 24854 0 _0024_
rlabel metal1 35277 24106 35277 24106 0 _0025_
rlabel via1 35737 24854 35737 24854 0 _0026_
rlabel metal2 33810 14620 33810 14620 0 _0027_
rlabel metal1 36294 12954 36294 12954 0 _0028_
rlabel metal1 35976 14314 35976 14314 0 _0029_
rlabel metal1 35021 15402 35021 15402 0 _0030_
rlabel metal1 33948 14586 33948 14586 0 _0031_
rlabel metal1 29654 14314 29654 14314 0 _0032_
rlabel metal1 27462 12716 27462 12716 0 _0033_
rlabel metal1 20056 12070 20056 12070 0 _0034_
rlabel metal1 24058 12240 24058 12240 0 _0035_
rlabel metal1 24456 15402 24456 15402 0 _0036_
rlabel metal2 24702 17476 24702 17476 0 _0037_
rlabel metal1 24978 18802 24978 18802 0 _0038_
rlabel metal2 30314 16422 30314 16422 0 _0039_
rlabel metal1 28556 17170 28556 17170 0 _0040_
rlabel metal1 25116 18938 25116 18938 0 _0041_
rlabel metal2 26542 19108 26542 19108 0 _0042_
rlabel metal1 29256 19482 29256 19482 0 _0043_
rlabel metal1 30268 19414 30268 19414 0 _0044_
rlabel metal1 32522 19278 32522 19278 0 _0045_
rlabel metal1 34561 19754 34561 19754 0 _0046_
rlabel metal1 33534 18190 33534 18190 0 _0047_
rlabel metal1 34270 17782 34270 17782 0 _0048_
rlabel metal1 37306 19958 37306 19958 0 _0049_
rlabel metal2 33810 22066 33810 22066 0 _0050_
rlabel metal1 27360 8466 27360 8466 0 _0051_
rlabel metal2 22494 10268 22494 10268 0 _0052_
rlabel metal1 27324 7514 27324 7514 0 _0053_
rlabel metal2 30406 7650 30406 7650 0 _0054_
rlabel metal1 28796 7242 28796 7242 0 _0055_
rlabel metal1 30958 10166 30958 10166 0 _0056_
rlabel viali 30028 8942 30028 8942 0 _0057_
rlabel metal2 21482 10234 21482 10234 0 _0058_
rlabel metal1 49036 9146 49036 9146 0 _0059_
rlabel metal1 33616 8466 33616 8466 0 _0060_
rlabel metal1 35006 8602 35006 8602 0 _0061_
rlabel metal1 35972 9146 35972 9146 0 _0062_
rlabel metal2 32522 9078 32522 9078 0 _0063_
rlabel metal1 38778 11322 38778 11322 0 _0064_
rlabel metal1 29256 10234 29256 10234 0 _0065_
rlabel metal1 23092 9418 23092 9418 0 _0066_
rlabel metal2 24058 10642 24058 10642 0 _0067_
rlabel metal1 19642 13192 19642 13192 0 _0068_
rlabel metal1 20470 16456 20470 16456 0 _0069_
rlabel metal1 22846 17238 22846 17238 0 _0070_
rlabel metal1 22954 17782 22954 17782 0 _0071_
rlabel metal1 33544 17170 33544 17170 0 _0072_
rlabel metal1 29398 18258 29398 18258 0 _0073_
rlabel metal1 24855 20808 24855 20808 0 _0074_
rlabel metal1 24140 21522 24140 21522 0 _0075_
rlabel metal1 27963 21998 27963 21998 0 _0076_
rlabel metal1 30171 23018 30171 23018 0 _0077_
rlabel metal2 31326 23800 31326 23800 0 _0078_
rlabel metal2 32246 23324 32246 23324 0 _0079_
rlabel metal1 36309 21930 36309 21930 0 _0080_
rlabel metal1 38410 18088 38410 18088 0 _0081_
rlabel metal2 40342 19176 40342 19176 0 _0082_
rlabel metal1 39330 21114 39330 21114 0 _0083_
rlabel metal1 52976 7786 52976 7786 0 _0084_
rlabel metal1 21436 6970 21436 6970 0 _0085_
rlabel metal1 22760 7854 22760 7854 0 _0086_
rlabel metal1 20224 8534 20224 8534 0 _0087_
rlabel metal1 18906 6664 18906 6664 0 _0088_
rlabel metal2 23690 6562 23690 6562 0 _0089_
rlabel metal1 19780 6426 19780 6426 0 _0090_
rlabel metal1 22908 8058 22908 8058 0 _0091_
rlabel metal1 25392 6970 25392 6970 0 _0092_
rlabel metal1 18630 6426 18630 6426 0 _0093_
rlabel metal1 18436 7378 18436 7378 0 _0094_
rlabel metal2 18262 9894 18262 9894 0 _0095_
rlabel metal1 17756 10234 17756 10234 0 _0096_
rlabel metal2 20838 10234 20838 10234 0 _0097_
rlabel metal2 18814 10642 18814 10642 0 _0098_
rlabel metal1 16330 10744 16330 10744 0 _0099_
rlabel via1 20373 12818 20373 12818 0 _0100_
rlabel metal1 19212 14314 19212 14314 0 _0101_
rlabel metal1 19698 12818 19698 12818 0 _0102_
rlabel metal2 17066 13090 17066 13090 0 _0103_
rlabel metal1 14904 13498 14904 13498 0 _0104_
rlabel metal2 21574 19516 21574 19516 0 _0105_
rlabel metal2 21666 16082 21666 16082 0 _0106_
rlabel metal1 20654 18632 20654 18632 0 _0107_
rlabel metal1 19131 19346 19131 19346 0 _0108_
rlabel metal1 19580 17578 19580 17578 0 _0109_
rlabel metal1 19632 15470 19632 15470 0 _0110_
rlabel metal1 17434 16456 17434 16456 0 _0111_
rlabel via1 25249 24106 25249 24106 0 _0112_
rlabel metal1 25192 24854 25192 24854 0 _0113_
rlabel metal1 26026 24786 26026 24786 0 _0114_
rlabel metal1 27140 23290 27140 23290 0 _0115_
rlabel metal1 26266 7412 26266 7412 0 _0116_
rlabel metal1 26818 7378 26818 7378 0 _0117_
rlabel metal1 30774 8466 30774 8466 0 _0118_
rlabel metal1 30912 7378 30912 7378 0 _0119_
rlabel metal1 29118 7514 29118 7514 0 _0120_
rlabel metal1 28152 7378 28152 7378 0 _0121_
rlabel metal2 27370 10812 27370 10812 0 _0122_
rlabel metal1 31418 10064 31418 10064 0 _0123_
rlabel metal1 29670 7446 29670 7446 0 _0124_
rlabel metal1 28842 9452 28842 9452 0 _0125_
rlabel metal2 22126 9724 22126 9724 0 _0126_
rlabel metal2 41078 14348 41078 14348 0 _0127_
rlabel metal2 40894 13821 40894 13821 0 _0128_
rlabel metal1 14490 14042 14490 14042 0 _0129_
rlabel metal1 33534 7888 33534 7888 0 _0130_
rlabel metal2 33350 8500 33350 8500 0 _0131_
rlabel metal2 39238 11951 39238 11951 0 _0132_
rlabel metal1 34454 9146 34454 9146 0 _0133_
rlabel metal2 35466 9180 35466 9180 0 _0134_
rlabel metal1 32062 10064 32062 10064 0 _0135_
rlabel metal1 35006 8942 35006 8942 0 _0136_
rlabel metal2 31694 9350 31694 9350 0 _0137_
rlabel metal1 32062 8466 32062 8466 0 _0138_
rlabel metal1 33810 11254 33810 11254 0 _0139_
rlabel metal1 39284 11118 39284 11118 0 _0140_
rlabel metal2 29670 12036 29670 12036 0 _0141_
rlabel metal2 29026 11186 29026 11186 0 _0142_
rlabel metal2 24932 12580 24932 12580 0 _0143_
rlabel metal2 22218 10540 22218 10540 0 _0144_
rlabel metal1 22908 12682 22908 12682 0 _0145_
rlabel metal2 23874 9690 23874 9690 0 _0146_
rlabel metal2 23414 14518 23414 14518 0 _0147_
rlabel metal2 20930 14280 20930 14280 0 _0148_
rlabel metal1 23046 15130 23046 15130 0 _0149_
rlabel metal1 22356 16218 22356 16218 0 _0150_
rlabel metal1 32752 22066 32752 22066 0 _0151_
rlabel metal2 24610 17170 24610 17170 0 _0152_
rlabel metal1 22816 17850 22816 17850 0 _0153_
rlabel metal1 20654 20502 20654 20502 0 _0154_
rlabel metal1 24380 17850 24380 17850 0 _0155_
rlabel metal1 22540 17646 22540 17646 0 _0156_
rlabel metal2 31878 16796 31878 16796 0 _0157_
rlabel metal1 31740 16014 31740 16014 0 _0158_
rlabel metal1 30820 17646 30820 17646 0 _0159_
rlabel metal2 28014 18054 28014 18054 0 _0160_
rlabel metal1 23736 20434 23736 20434 0 _0161_
rlabel metal1 23736 20570 23736 20570 0 _0162_
rlabel metal1 24702 20026 24702 20026 0 _0163_
rlabel metal1 23506 21522 23506 21522 0 _0164_
rlabel metal1 27370 21658 27370 21658 0 _0165_
rlabel metal1 28060 22610 28060 22610 0 _0166_
rlabel metal2 30958 22440 30958 22440 0 _0167_
rlabel metal1 29992 22746 29992 22746 0 _0168_
rlabel metal2 32338 23426 32338 23426 0 _0169_
rlabel metal2 30958 24582 30958 24582 0 _0170_
rlabel metal1 31878 21862 31878 21862 0 _0171_
rlabel metal1 32108 24174 32108 24174 0 _0172_
rlabel metal1 34776 21114 34776 21114 0 _0173_
rlabel metal2 36938 22049 36938 22049 0 _0174_
rlabel viali 35098 16559 35098 16559 0 _0175_
rlabel metal1 39238 18224 39238 18224 0 _0176_
rlabel metal1 37214 19482 37214 19482 0 _0177_
rlabel metal2 39422 20162 39422 20162 0 _0178_
rlabel via1 38686 21845 38686 21845 0 _0179_
rlabel metal1 40204 20910 40204 20910 0 _0180_
rlabel metal2 51658 9146 51658 9146 0 _0181_
rlabel metal1 23736 13974 23736 13974 0 _0182_
rlabel metal1 21620 16014 21620 16014 0 _0183_
rlabel metal1 19780 9010 19780 9010 0 _0184_
rlabel metal2 21666 6970 21666 6970 0 _0185_
rlabel metal1 25162 8024 25162 8024 0 _0186_
rlabel metal1 19458 8942 19458 8942 0 _0187_
rlabel metal1 18768 6766 18768 6766 0 _0188_
rlabel metal1 24058 6290 24058 6290 0 _0189_
rlabel metal2 19366 7004 19366 7004 0 _0190_
rlabel metal1 23552 6154 23552 6154 0 _0191_
rlabel metal1 25990 6698 25990 6698 0 _0192_
rlabel metal1 18952 6290 18952 6290 0 _0193_
rlabel metal1 19458 8840 19458 8840 0 _0194_
rlabel metal1 21298 13804 21298 13804 0 _0195_
rlabel metal1 18078 8976 18078 8976 0 _0196_
rlabel metal1 17710 10030 17710 10030 0 _0197_
rlabel metal2 20654 9996 20654 9996 0 _0198_
rlabel metal1 18676 9554 18676 9554 0 _0199_
rlabel metal1 17112 10642 17112 10642 0 _0200_
rlabel metal1 20700 13702 20700 13702 0 _0201_
rlabel metal1 19136 14858 19136 14858 0 _0202_
rlabel metal1 21068 10030 21068 10030 0 _0203_
rlabel metal1 16882 12784 16882 12784 0 _0204_
rlabel metal2 14674 13821 14674 13821 0 _0205_
rlabel metal1 21712 19822 21712 19822 0 _0206_
rlabel metal2 21850 16218 21850 16218 0 _0207_
rlabel metal1 20608 18734 20608 18734 0 _0208_
rlabel metal2 19642 20230 19642 20230 0 _0209_
rlabel metal1 20516 18394 20516 18394 0 _0210_
rlabel metal1 20010 17646 20010 17646 0 _0211_
rlabel metal1 18952 16218 18952 16218 0 _0212_
rlabel metal1 25714 17238 25714 17238 0 _0213_
rlabel metal1 25208 23834 25208 23834 0 _0214_
rlabel metal1 25760 8602 25760 8602 0 _0215_
rlabel metal1 25116 22746 25116 22746 0 _0216_
rlabel metal1 26542 10778 26542 10778 0 _0217_
rlabel metal1 25852 23290 25852 23290 0 _0218_
rlabel metal1 27094 9418 27094 9418 0 _0219_
rlabel metal2 27278 23290 27278 23290 0 _0220_
rlabel metal1 14858 22406 14858 22406 0 _0221_
rlabel metal1 26358 33456 26358 33456 0 _0222_
rlabel metal1 26266 28730 26266 28730 0 _0223_
rlabel metal2 29026 25670 29026 25670 0 _0224_
rlabel metal1 26680 32402 26680 32402 0 _0225_
rlabel metal2 25530 51782 25530 51782 0 _0226_
rlabel metal1 33994 48518 33994 48518 0 _0227_
rlabel metal1 14628 22610 14628 22610 0 _0228_
rlabel metal1 14076 22406 14076 22406 0 _0229_
rlabel metal1 27186 32368 27186 32368 0 _0230_
rlabel metal1 26404 40018 26404 40018 0 _0231_
rlabel metal2 22310 21233 22310 21233 0 _0232_
rlabel metal1 21482 21488 21482 21488 0 _0233_
rlabel metal1 26956 32810 26956 32810 0 _0234_
rlabel metal1 26496 34034 26496 34034 0 _0235_
rlabel metal1 26588 28186 26588 28186 0 _0236_
rlabel metal1 15180 24378 15180 24378 0 _0237_
rlabel metal1 14398 24038 14398 24038 0 _0238_
rlabel metal1 27370 32436 27370 32436 0 _0239_
rlabel metal1 23414 23086 23414 23086 0 _0240_
rlabel metal2 25346 35224 25346 35224 0 _0241_
rlabel metal1 27186 20978 27186 20978 0 _0242_
rlabel metal1 22448 20910 22448 20910 0 _0243_
rlabel metal2 26266 35700 26266 35700 0 _0244_
rlabel metal1 16905 22746 16905 22746 0 _0245_
rlabel metal1 4715 22610 4715 22610 0 _0246_
rlabel metal1 26174 34102 26174 34102 0 _0247_
rlabel metal1 32844 49062 32844 49062 0 _0248_
rlabel metal2 31142 47192 31142 47192 0 _0249_
rlabel metal2 31878 41004 31878 41004 0 _0250_
rlabel metal2 22218 21148 22218 21148 0 _0251_
rlabel metal1 25806 23698 25806 23698 0 _0252_
rlabel metal2 23506 22780 23506 22780 0 _0253_
rlabel metal1 24196 22950 24196 22950 0 _0254_
rlabel metal1 27074 35054 27074 35054 0 _0255_
rlabel metal1 23000 23698 23000 23698 0 _0256_
rlabel metal1 52210 33626 52210 33626 0 _0257_
rlabel metal1 53774 33864 53774 33864 0 _0258_
rlabel metal2 53406 33728 53406 33728 0 _0259_
rlabel metal2 29118 33932 29118 33932 0 _0260_
rlabel metal2 28474 33354 28474 33354 0 _0261_
rlabel metal1 27968 33082 27968 33082 0 _0262_
rlabel metal1 28520 32538 28520 32538 0 _0263_
rlabel metal1 30406 33354 30406 33354 0 _0264_
rlabel metal1 22724 3502 22724 3502 0 _0265_
rlabel metal1 24380 33354 24380 33354 0 _0266_
rlabel metal1 14030 29104 14030 29104 0 _0267_
rlabel metal1 17526 12852 17526 12852 0 _0268_
rlabel metal1 14168 12206 14168 12206 0 _0269_
rlabel metal2 48254 46478 48254 46478 0 _0270_
rlabel metal2 26910 37689 26910 37689 0 _0271_
rlabel metal2 26358 41718 26358 41718 0 _0272_
rlabel metal2 29486 18207 29486 18207 0 _0273_
rlabel metal1 28520 15334 28520 15334 0 _0274_
rlabel metal1 28106 26996 28106 26996 0 _0275_
rlabel metal2 15318 13498 15318 13498 0 _0276_
rlabel metal2 26082 51850 26082 51850 0 _0277_
rlabel metal1 17020 16014 17020 16014 0 _0278_
rlabel metal1 25806 36346 25806 36346 0 _0279_
rlabel metal1 25576 39814 25576 39814 0 _0280_
rlabel metal2 30130 38114 30130 38114 0 _0281_
rlabel metal2 27738 40154 27738 40154 0 _0282_
rlabel metal2 29207 38522 29207 38522 0 _0283_
rlabel metal1 29900 38318 29900 38318 0 _0284_
rlabel metal1 30774 37230 30774 37230 0 _0285_
rlabel metal1 29670 42534 29670 42534 0 _0286_
rlabel metal2 28658 41038 28658 41038 0 _0287_
rlabel metal1 29440 38726 29440 38726 0 _0288_
rlabel metal2 30406 34204 30406 34204 0 _0289_
rlabel metal1 26266 34170 26266 34170 0 _0290_
rlabel metal1 26588 40018 26588 40018 0 _0291_
rlabel metal2 30498 37196 30498 37196 0 _0292_
rlabel metal1 14858 34442 14858 34442 0 _0293_
rlabel metal2 30406 34663 30406 34663 0 _0294_
rlabel metal1 30084 41990 30084 41990 0 _0295_
rlabel metal1 15410 34952 15410 34952 0 _0296_
rlabel metal2 26542 35360 26542 35360 0 _0297_
rlabel metal1 27692 27982 27692 27982 0 _0298_
rlabel metal2 27830 28322 27830 28322 0 _0299_
rlabel metal2 30406 37281 30406 37281 0 _0300_
rlabel metal1 29808 37094 29808 37094 0 _0301_
rlabel metal1 30038 27438 30038 27438 0 _0302_
rlabel metal1 27830 36006 27830 36006 0 _0303_
rlabel metal1 27784 27574 27784 27574 0 _0304_
rlabel metal1 28198 27846 28198 27846 0 _0305_
rlabel via3 28267 33116 28267 33116 0 _0306_
rlabel metal1 28474 27506 28474 27506 0 _0307_
rlabel metal1 19251 29070 19251 29070 0 _0308_
rlabel metal2 28842 37383 28842 37383 0 _0309_
rlabel metal1 28474 37434 28474 37434 0 _0310_
rlabel viali 28193 36776 28193 36776 0 _0311_
rlabel metal2 28750 37060 28750 37060 0 _0312_
rlabel metal1 29256 35734 29256 35734 0 _0313_
rlabel metal1 26910 35802 26910 35802 0 _0314_
rlabel metal1 26082 37094 26082 37094 0 _0315_
rlabel metal3 26519 40052 26519 40052 0 _0316_
rlabel metal2 26542 40698 26542 40698 0 _0317_
rlabel metal2 25622 39100 25622 39100 0 _0318_
rlabel metal1 25576 37230 25576 37230 0 _0319_
rlabel metal1 24104 34714 24104 34714 0 _0320_
rlabel metal1 24610 42126 24610 42126 0 _0321_
rlabel metal1 29900 41786 29900 41786 0 _0322_
rlabel metal1 25668 42194 25668 42194 0 _0323_
rlabel metal1 25392 44234 25392 44234 0 _0324_
rlabel metal2 25898 35258 25898 35258 0 _0325_
rlabel metal1 27830 35632 27830 35632 0 _0326_
rlabel metal1 26082 35088 26082 35088 0 _0327_
rlabel metal1 25438 35054 25438 35054 0 _0328_
rlabel metal1 27508 30906 27508 30906 0 _0329_
rlabel metal1 33396 38998 33396 38998 0 _0330_
rlabel metal1 26680 51782 26680 51782 0 _0331_
rlabel metal1 26588 36890 26588 36890 0 _0332_
rlabel metal1 27554 37434 27554 37434 0 _0333_
rlabel metal1 28888 36822 28888 36822 0 _0334_
rlabel metal2 26634 34884 26634 34884 0 _0335_
rlabel metal1 27600 31790 27600 31790 0 _0336_
rlabel metal2 25714 39848 25714 39848 0 _0337_
rlabel metal1 27784 31722 27784 31722 0 _0338_
rlabel metal2 28382 31484 28382 31484 0 _0339_
rlabel metal1 27830 38726 27830 38726 0 _0340_
rlabel metal1 33120 39338 33120 39338 0 _0341_
rlabel metal1 27140 38522 27140 38522 0 _0342_
rlabel metal1 26680 39066 26680 39066 0 _0343_
rlabel metal1 19757 39066 19757 39066 0 _0344_
rlabel metal1 26772 38726 26772 38726 0 _0345_
rlabel metal1 26864 43622 26864 43622 0 _0346_
rlabel metal1 28474 38386 28474 38386 0 _0347_
rlabel metal1 28980 51782 28980 51782 0 _0348_
rlabel metal1 29440 40086 29440 40086 0 _0349_
rlabel metal1 28474 41242 28474 41242 0 _0350_
rlabel metal1 28198 41786 28198 41786 0 _0351_
rlabel metal1 33033 40018 33033 40018 0 _0352_
rlabel metal2 32338 39610 32338 39610 0 _0353_
rlabel metal1 31050 38318 31050 38318 0 _0354_
rlabel metal1 31878 47158 31878 47158 0 _0355_
rlabel metal1 31418 47158 31418 47158 0 _0356_
rlabel metal2 31694 39406 31694 39406 0 _0357_
rlabel metal1 32706 46342 32706 46342 0 _0358_
rlabel metal1 32476 39406 32476 39406 0 _0359_
rlabel metal1 32844 38318 32844 38318 0 _0360_
rlabel metal2 53866 47532 53866 47532 0 _0361_
rlabel metal1 33488 40086 33488 40086 0 _0362_
rlabel metal2 32706 39644 32706 39644 0 _0363_
rlabel metal1 33442 41072 33442 41072 0 _0364_
rlabel metal1 32844 38998 32844 38998 0 _0365_
rlabel metal1 33902 38930 33902 38930 0 _0366_
rlabel metal2 35834 47294 35834 47294 0 _0367_
rlabel metal1 33810 41174 33810 41174 0 _0368_
rlabel metal1 34638 39406 34638 39406 0 _0369_
rlabel metal1 33074 46138 33074 46138 0 _0370_
rlabel metal1 33764 39406 33764 39406 0 _0371_
rlabel metal1 33442 38318 33442 38318 0 _0372_
rlabel metal1 33074 48042 33074 48042 0 _0373_
rlabel metal1 34224 40086 34224 40086 0 _0374_
rlabel metal1 34914 40018 34914 40018 0 _0375_
rlabel metal1 33304 41582 33304 41582 0 _0376_
rlabel metal1 33442 40494 33442 40494 0 _0377_
rlabel metal2 33902 39678 33902 39678 0 _0378_
rlabel metal1 32522 42262 32522 42262 0 _0379_
rlabel metal1 33396 42330 33396 42330 0 _0380_
rlabel metal1 32476 40630 32476 40630 0 _0381_
rlabel metal1 33028 41786 33028 41786 0 _0382_
rlabel metal1 34868 41582 34868 41582 0 _0383_
rlabel metal1 35236 40494 35236 40494 0 _0384_
rlabel metal2 22402 11832 22402 11832 0 _0385_
rlabel metal1 17388 12206 17388 12206 0 _0386_
rlabel metal2 23230 10642 23230 10642 0 _0387_
rlabel metal1 14904 4590 14904 4590 0 _0388_
rlabel metal2 10902 3842 10902 3842 0 _0389_
rlabel metal1 14904 3162 14904 3162 0 _0390_
rlabel metal1 13294 6664 13294 6664 0 _0391_
rlabel via1 10902 3502 10902 3502 0 _0392_
rlabel metal1 10856 3162 10856 3162 0 _0393_
rlabel metal1 10534 4250 10534 4250 0 _0394_
rlabel metal1 12972 4794 12972 4794 0 _0395_
rlabel metal1 13018 4046 13018 4046 0 _0396_
rlabel metal1 12696 4794 12696 4794 0 _0397_
rlabel metal1 13294 5780 13294 5780 0 _0398_
rlabel metal1 12788 5882 12788 5882 0 _0399_
rlabel metal2 12558 6902 12558 6902 0 _0400_
rlabel metal1 16238 12818 16238 12818 0 _0401_
rlabel metal1 14352 5066 14352 5066 0 _0402_
rlabel metal2 17342 10098 17342 10098 0 _0403_
rlabel metal1 14168 9146 14168 9146 0 _0404_
rlabel metal1 14352 9418 14352 9418 0 _0405_
rlabel metal1 15180 8602 15180 8602 0 _0406_
rlabel metal1 14076 10234 14076 10234 0 _0407_
rlabel metal1 14858 10438 14858 10438 0 _0408_
rlabel metal1 15272 11322 15272 11322 0 _0409_
rlabel metal1 16744 10778 16744 10778 0 _0410_
rlabel metal1 16192 11322 16192 11322 0 _0411_
rlabel metal1 16468 9146 16468 9146 0 _0412_
rlabel metal1 16330 13838 16330 13838 0 _0413_
rlabel metal2 17342 13668 17342 13668 0 _0414_
rlabel metal1 16330 10234 16330 10234 0 _0415_
rlabel metal1 17388 13838 17388 13838 0 _0416_
rlabel metal1 17388 14382 17388 14382 0 _0417_
rlabel metal2 17250 11492 17250 11492 0 _0418_
rlabel metal1 17388 8058 17388 8058 0 _0419_
rlabel metal1 40710 10778 40710 10778 0 _0420_
rlabel metal2 40388 14926 40388 14926 0 _0421_
rlabel metal1 40250 10676 40250 10676 0 _0422_
rlabel metal2 40066 13345 40066 13345 0 _0423_
rlabel metal1 41078 17646 41078 17646 0 _0424_
rlabel metal1 39238 13328 39238 13328 0 _0425_
rlabel metal1 38732 9146 38732 9146 0 _0426_
rlabel metal1 38939 12206 38939 12206 0 _0427_
rlabel metal2 37674 12342 37674 12342 0 _0428_
rlabel metal1 37720 12410 37720 12410 0 _0429_
rlabel metal1 29026 7174 29026 7174 0 _0430_
rlabel metal2 29118 13940 29118 13940 0 _0431_
rlabel metal1 35972 9554 35972 9554 0 _0432_
rlabel metal1 32706 10778 32706 10778 0 _0433_
rlabel metal2 32338 11594 32338 11594 0 _0434_
rlabel metal1 31372 10710 31372 10710 0 _0435_
rlabel metal1 34822 15470 34822 15470 0 _0436_
rlabel metal2 39790 11628 39790 11628 0 _0437_
rlabel metal2 30774 10200 30774 10200 0 _0438_
rlabel metal2 36478 10812 36478 10812 0 _0439_
rlabel metal1 39468 10030 39468 10030 0 _0440_
rlabel metal1 31234 10234 31234 10234 0 _0441_
rlabel metal1 30958 10778 30958 10778 0 _0442_
rlabel metal1 38134 10166 38134 10166 0 _0443_
rlabel metal2 40526 11356 40526 11356 0 _0444_
rlabel metal2 31234 12988 31234 12988 0 _0445_
rlabel metal2 30590 12036 30590 12036 0 _0446_
rlabel via2 36478 11237 36478 11237 0 _0447_
rlabel metal1 35507 12206 35507 12206 0 _0448_
rlabel metal2 37122 12784 37122 12784 0 _0449_
rlabel viali 36478 11119 36478 11119 0 _0450_
rlabel metal1 36846 20366 36846 20366 0 _0451_
rlabel metal2 36662 11594 36662 11594 0 _0452_
rlabel metal1 38916 12274 38916 12274 0 _0453_
rlabel via1 29762 12818 29762 12818 0 _0454_
rlabel metal1 30590 11730 30590 11730 0 _0455_
rlabel metal1 36938 12342 36938 12342 0 _0456_
rlabel metal1 26864 14382 26864 14382 0 _0457_
rlabel metal1 28198 13294 28198 13294 0 _0458_
rlabel metal1 33074 13464 33074 13464 0 _0459_
rlabel metal2 40158 13022 40158 13022 0 _0460_
rlabel metal2 36570 16048 36570 16048 0 _0461_
rlabel metal2 39698 15198 39698 15198 0 _0462_
rlabel metal1 39882 15062 39882 15062 0 _0463_
rlabel viali 39340 14382 39340 14382 0 _0464_
rlabel metal1 40848 13294 40848 13294 0 _0465_
rlabel metal1 27968 14994 27968 14994 0 _0466_
rlabel metal1 34822 14552 34822 14552 0 _0467_
rlabel metal2 41538 15028 41538 15028 0 _0468_
rlabel metal1 39882 21590 39882 21590 0 _0469_
rlabel metal2 33166 15708 33166 15708 0 _0470_
rlabel metal2 40526 15198 40526 15198 0 _0471_
rlabel metal2 43378 15232 43378 15232 0 _0472_
rlabel metal1 24104 16762 24104 16762 0 _0473_
rlabel metal1 36202 17272 36202 17272 0 _0474_
rlabel via2 39422 16779 39422 16779 0 _0475_
rlabel metal2 42090 16762 42090 16762 0 _0476_
rlabel metal1 29210 15674 29210 15674 0 _0477_
rlabel metal1 33350 16456 33350 16456 0 _0478_
rlabel metal1 38686 17170 38686 17170 0 _0479_
rlabel metal1 40250 17000 40250 17000 0 _0480_
rlabel metal2 33718 16082 33718 16082 0 _0481_
rlabel metal1 34868 16218 34868 16218 0 _0482_
rlabel metal2 37490 16660 37490 16660 0 _0483_
rlabel metal1 37858 16762 37858 16762 0 _0484_
rlabel metal1 38180 18190 38180 18190 0 _0485_
rlabel metal1 36754 17544 36754 17544 0 _0486_
rlabel metal1 40342 18258 40342 18258 0 _0487_
rlabel metal2 41722 17884 41722 17884 0 _0488_
rlabel metal2 28566 21216 28566 21216 0 _0489_
rlabel metal1 41124 19346 41124 19346 0 _0490_
rlabel metal2 39882 18870 39882 18870 0 _0491_
rlabel metal1 40710 18156 40710 18156 0 _0492_
rlabel metal1 38962 20978 38962 20978 0 _0493_
rlabel metal2 42274 20298 42274 20298 0 _0494_
rlabel metal1 42964 20026 42964 20026 0 _0495_
rlabel metal2 41814 20876 41814 20876 0 _0496_
rlabel metal2 38962 19312 38962 19312 0 _0497_
rlabel metal1 39376 18394 39376 18394 0 _0498_
rlabel metal1 39238 21522 39238 21522 0 _0499_
rlabel metal2 42090 21828 42090 21828 0 _0500_
rlabel metal2 42274 21828 42274 21828 0 _0501_
rlabel metal1 39882 22474 39882 22474 0 _0502_
rlabel metal1 41262 22100 41262 22100 0 _0503_
rlabel metal1 41492 22066 41492 22066 0 _0504_
rlabel metal1 38732 22610 38732 22610 0 _0505_
rlabel metal1 39790 22746 39790 22746 0 _0506_
rlabel metal2 40434 24038 40434 24038 0 _0507_
rlabel via2 35558 22763 35558 22763 0 _0508_
rlabel metal2 39974 22780 39974 22780 0 _0509_
rlabel metal2 39790 23970 39790 23970 0 _0510_
rlabel metal1 37582 23120 37582 23120 0 _0511_
rlabel metal1 37904 23290 37904 23290 0 _0512_
rlabel metal1 38134 23834 38134 23834 0 _0513_
rlabel metal1 36018 21658 36018 21658 0 _0514_
rlabel metal1 38410 22746 38410 22746 0 _0515_
rlabel metal1 38180 24378 38180 24378 0 _0516_
rlabel metal1 38088 13498 38088 13498 0 _0517_
rlabel metal1 36386 22746 36386 22746 0 _0518_
rlabel metal2 35558 23630 35558 23630 0 _0519_
rlabel metal1 35788 23834 35788 23834 0 _0520_
rlabel metal1 36018 12614 36018 12614 0 _0521_
rlabel metal2 33718 24582 33718 24582 0 _0522_
rlabel metal2 33166 25092 33166 25092 0 _0523_
rlabel metal1 35098 25228 35098 25228 0 _0524_
rlabel metal1 35374 25466 35374 25466 0 _0525_
rlabel metal1 34500 23834 34500 23834 0 _0526_
rlabel metal1 35926 25296 35926 25296 0 _0527_
rlabel metal1 36064 10234 36064 10234 0 _0528_
rlabel metal1 31096 13906 31096 13906 0 _0529_
rlabel metal1 34868 15334 34868 15334 0 _0530_
rlabel metal2 34822 11900 34822 11900 0 _0531_
rlabel metal2 32982 12444 32982 12444 0 _0532_
rlabel metal1 30268 13294 30268 13294 0 _0533_
rlabel metal1 30728 13498 30728 13498 0 _0534_
rlabel metal1 32614 13872 32614 13872 0 _0535_
rlabel metal2 15410 14076 15410 14076 0 _0536_
rlabel metal2 31694 14756 31694 14756 0 _0537_
rlabel metal1 29854 10778 29854 10778 0 _0538_
rlabel metal1 26726 16558 26726 16558 0 _0539_
rlabel metal1 19918 12274 19918 12274 0 _0540_
rlabel metal2 24058 13124 24058 13124 0 _0541_
rlabel metal1 25178 16490 25178 16490 0 _0542_
rlabel metal2 29578 15912 29578 15912 0 _0543_
rlabel metal1 26864 15130 26864 15130 0 _0544_
rlabel metal1 29072 15130 29072 15130 0 _0545_
rlabel metal2 29118 16388 29118 16388 0 _0546_
rlabel metal2 22402 16966 22402 16966 0 _0547_
rlabel metal1 29532 16014 29532 16014 0 _0548_
rlabel metal1 27370 20400 27370 20400 0 _0549_
rlabel metal1 28566 18802 28566 18802 0 _0550_
rlabel metal2 28198 17476 28198 17476 0 _0551_
rlabel metal2 27186 21284 27186 21284 0 _0552_
rlabel metal1 25806 21964 25806 21964 0 _0553_
rlabel metal2 24702 20298 24702 20298 0 _0554_
rlabel metal2 27830 19550 27830 19550 0 _0555_
rlabel metal1 30038 20570 30038 20570 0 _0556_
rlabel metal1 28336 19890 28336 19890 0 _0557_
rlabel metal1 30222 19890 30222 19890 0 _0558_
rlabel metal2 33166 18734 33166 18734 0 _0559_
rlabel metal1 32844 19482 32844 19482 0 _0560_
rlabel metal1 38686 18768 38686 18768 0 _0561_
rlabel metal1 32660 18938 32660 18938 0 _0562_
rlabel metal1 32338 20332 32338 20332 0 _0563_
rlabel metal1 34546 17714 34546 17714 0 _0564_
rlabel metal1 36478 21318 36478 21318 0 _0565_
rlabel metal2 36018 19108 36018 19108 0 _0566_
rlabel metal1 38824 19482 38824 19482 0 _0567_
rlabel metal1 53176 9078 53176 9078 0 _0568_
rlabel metal2 29486 10370 29486 10370 0 _0569_
rlabel metal1 28106 9146 28106 9146 0 _0570_
rlabel metal1 25576 8466 25576 8466 0 _0571_
rlabel metal1 26726 8058 26726 8058 0 _0572_
rlabel metal1 20010 10676 20010 10676 0 _0573_
rlabel metal1 18308 16150 18308 16150 0 clknet_0_net235
rlabel metal2 16146 14790 16146 14790 0 clknet_0_wb_clk_i
rlabel metal2 20010 15674 20010 15674 0 clknet_1_0__leaf_net235
rlabel metal1 2070 18258 2070 18258 0 clknet_1_1__leaf_net235
rlabel metal1 19504 12614 19504 12614 0 clknet_3_0__leaf_wb_clk_i
rlabel metal1 33442 8500 33442 8500 0 clknet_3_1__leaf_wb_clk_i
rlabel metal1 20148 12818 20148 12818 0 clknet_3_2__leaf_wb_clk_i
rlabel metal1 18722 19380 18722 19380 0 clknet_3_3__leaf_wb_clk_i
rlabel metal1 39100 9622 39100 9622 0 clknet_3_4__leaf_wb_clk_i
rlabel metal2 52946 7684 52946 7684 0 clknet_3_5__leaf_wb_clk_i
rlabel metal1 36432 20978 36432 20978 0 clknet_3_6__leaf_wb_clk_i
rlabel metal1 40756 20910 40756 20910 0 clknet_3_7__leaf_wb_clk_i
rlabel metal1 26772 33014 26772 33014 0 design_addr\[0\]
rlabel metal1 26266 32776 26266 32776 0 design_addr\[1\]
rlabel metal2 27554 25772 27554 25772 0 design_addr\[2\]
rlabel metal2 28198 24820 28198 24820 0 design_addr\[3\]
rlabel metal3 1142 17884 1142 17884 0 design_clk_o
rlabel metal3 1188 3196 1188 3196 0 dsi_all[0]
rlabel metal3 1188 8636 1188 8636 0 dsi_all[10]
rlabel metal3 1188 9180 1188 9180 0 dsi_all[11]
rlabel metal3 1188 9724 1188 9724 0 dsi_all[12]
rlabel metal3 1188 10268 1188 10268 0 dsi_all[13]
rlabel metal3 1188 10812 1188 10812 0 dsi_all[14]
rlabel metal3 1188 11356 1188 11356 0 dsi_all[15]
rlabel metal3 1188 11900 1188 11900 0 dsi_all[16]
rlabel metal3 1188 12444 1188 12444 0 dsi_all[17]
rlabel metal3 1188 12988 1188 12988 0 dsi_all[18]
rlabel metal3 1188 13532 1188 13532 0 dsi_all[19]
rlabel metal3 1188 3740 1188 3740 0 dsi_all[1]
rlabel metal3 1188 14076 1188 14076 0 dsi_all[20]
rlabel metal3 1188 14620 1188 14620 0 dsi_all[21]
rlabel metal3 1188 15164 1188 15164 0 dsi_all[22]
rlabel metal3 1188 15708 1188 15708 0 dsi_all[23]
rlabel metal2 1702 16337 1702 16337 0 dsi_all[24]
rlabel metal3 1188 16796 1188 16796 0 dsi_all[25]
rlabel metal3 1188 17340 1188 17340 0 dsi_all[26]
rlabel metal3 1188 4284 1188 4284 0 dsi_all[2]
rlabel metal3 1188 4828 1188 4828 0 dsi_all[3]
rlabel metal3 1188 5372 1188 5372 0 dsi_all[4]
rlabel metal3 1188 5916 1188 5916 0 dsi_all[5]
rlabel metal2 1702 6545 1702 6545 0 dsi_all[6]
rlabel metal3 1188 7004 1188 7004 0 dsi_all[7]
rlabel metal3 1188 7548 1188 7548 0 dsi_all[8]
rlabel metal3 1188 8092 1188 8092 0 dsi_all[9]
rlabel metal1 53544 35054 53544 35054 0 dso_6502[0]
rlabel metal1 53452 38862 53452 38862 0 dso_6502[10]
rlabel via2 53038 37621 53038 37621 0 dso_6502[11]
rlabel metal2 53498 38641 53498 38641 0 dso_6502[12]
rlabel metal2 52210 38233 52210 38233 0 dso_6502[13]
rlabel metal1 53544 39950 53544 39950 0 dso_6502[14]
rlabel via2 53038 38709 53038 38709 0 dso_6502[15]
rlabel metal2 53038 39185 53038 39185 0 dso_6502[16]
rlabel metal2 54326 39865 54326 39865 0 dso_6502[17]
rlabel metal2 53682 40001 53682 40001 0 dso_6502[18]
rlabel metal1 52900 40494 52900 40494 0 dso_6502[19]
rlabel metal2 53498 34731 53498 34731 0 dso_6502[1]
rlabel metal3 54840 40052 54840 40052 0 dso_6502[20]
rlabel metal2 52394 40409 52394 40409 0 dso_6502[21]
rlabel metal2 53498 40817 53498 40817 0 dso_6502[22]
rlabel metal3 54472 40868 54472 40868 0 dso_6502[23]
rlabel metal3 54150 41140 54150 41140 0 dso_6502[24]
rlabel metal2 52394 41497 52394 41497 0 dso_6502[25]
rlabel metal2 52394 42109 52394 42109 0 dso_6502[26]
rlabel metal1 52716 36142 52716 36142 0 dso_6502[2]
rlabel metal2 53498 35513 53498 35513 0 dso_6502[3]
rlabel metal1 53682 36142 53682 36142 0 dso_6502[4]
rlabel metal1 53544 36686 53544 36686 0 dso_6502[5]
rlabel metal2 53498 36771 53498 36771 0 dso_6502[6]
rlabel metal1 53590 37774 53590 37774 0 dso_6502[7]
rlabel metal1 53636 38318 53636 38318 0 dso_6502[8]
rlabel metal2 53038 36975 53038 36975 0 dso_6502[9]
rlabel metal2 1702 23987 1702 23987 0 dso_LCD[0]
rlabel metal2 1702 24599 1702 24599 0 dso_LCD[1]
rlabel metal2 1610 25109 1610 25109 0 dso_LCD[2]
rlabel metal2 1610 25687 1610 25687 0 dso_LCD[3]
rlabel metal3 1464 26044 1464 26044 0 dso_LCD[4]
rlabel metal1 2622 26894 2622 26894 0 dso_LCD[5]
rlabel metal2 1610 27285 1610 27285 0 dso_LCD[6]
rlabel via2 2254 27659 2254 27659 0 dso_LCD[7]
rlabel metal2 53498 42041 53498 42041 0 dso_as1802[0]
rlabel metal2 52210 44761 52210 44761 0 dso_as1802[10]
rlabel metal2 53498 45713 53498 45713 0 dso_as1802[11]
rlabel via2 53038 45237 53038 45237 0 dso_as1802[12]
rlabel metal1 53590 47022 53590 47022 0 dso_as1802[13]
rlabel metal2 52210 45849 52210 45849 0 dso_as1802[14]
rlabel metal1 53544 47566 53544 47566 0 dso_as1802[15]
rlabel via2 53038 46325 53038 46325 0 dso_as1802[16]
rlabel metal2 52670 47345 52670 47345 0 dso_as1802[17]
rlabel metal2 52210 47481 52210 47481 0 dso_as1802[18]
rlabel metal1 51336 47634 51336 47634 0 dso_as1802[19]
rlabel metal2 53498 42449 53498 42449 0 dso_as1802[1]
rlabel metal1 54418 49810 54418 49810 0 dso_as1802[20]
rlabel metal1 53084 49198 53084 49198 0 dso_as1802[21]
rlabel metal2 52394 48331 52394 48331 0 dso_as1802[22]
rlabel metal2 54326 49249 54326 49249 0 dso_as1802[23]
rlabel metal2 53682 49147 53682 49147 0 dso_as1802[24]
rlabel metal1 53544 49198 53544 49198 0 dso_as1802[25]
rlabel metal2 53498 48841 53498 48841 0 dso_as1802[26]
rlabel metal1 53590 43214 53590 43214 0 dso_as1802[2]
rlabel metal1 53498 43690 53498 43690 0 dso_as1802[3]
rlabel metal2 53498 43673 53498 43673 0 dso_as1802[4]
rlabel metal2 52946 43503 52946 43503 0 dso_as1802[5]
rlabel metal1 53590 44846 53590 44846 0 dso_as1802[6]
rlabel metal1 53544 45390 53544 45390 0 dso_as1802[7]
rlabel via2 53038 44149 53038 44149 0 dso_as1802[8]
rlabel metal1 53452 45934 53452 45934 0 dso_as1802[9]
rlabel metal1 2622 38862 2622 38862 0 dso_as2650[0]
rlabel metal1 2622 44302 2622 44302 0 dso_as2650[10]
rlabel metal1 2622 44846 2622 44846 0 dso_as2650[11]
rlabel metal1 2622 45390 2622 45390 0 dso_as2650[12]
rlabel metal1 2622 45934 2622 45934 0 dso_as2650[13]
rlabel metal1 2622 46478 2622 46478 0 dso_as2650[14]
rlabel metal1 2622 47022 2622 47022 0 dso_as2650[15]
rlabel metal1 2622 47566 2622 47566 0 dso_as2650[16]
rlabel metal1 2622 48110 2622 48110 0 dso_as2650[17]
rlabel metal1 2622 48654 2622 48654 0 dso_as2650[18]
rlabel metal1 2622 49198 2622 49198 0 dso_as2650[19]
rlabel metal1 2622 39406 2622 39406 0 dso_as2650[1]
rlabel metal2 1702 49623 1702 49623 0 dso_as2650[20]
rlabel metal1 2622 50286 2622 50286 0 dso_as2650[21]
rlabel metal1 2622 50830 2622 50830 0 dso_as2650[22]
rlabel metal2 1702 51187 1702 51187 0 dso_as2650[23]
rlabel metal2 1702 51799 1702 51799 0 dso_as2650[24]
rlabel metal1 1748 52394 1748 52394 0 dso_as2650[25]
rlabel metal1 2622 52394 2622 52394 0 dso_as2650[26]
rlabel metal1 2622 39950 2622 39950 0 dso_as2650[2]
rlabel metal1 2622 40494 2622 40494 0 dso_as2650[3]
rlabel metal1 2622 41038 2622 41038 0 dso_as2650[4]
rlabel metal1 2622 41582 2622 41582 0 dso_as2650[5]
rlabel metal1 2622 42126 2622 42126 0 dso_as2650[6]
rlabel metal1 2622 42670 2622 42670 0 dso_as2650[7]
rlabel metal1 2622 43214 2622 43214 0 dso_as2650[8]
rlabel metal1 2622 43758 2622 43758 0 dso_as2650[9]
rlabel metal2 11362 53907 11362 53907 0 dso_as5401[0]
rlabel metal2 23322 54179 23322 54179 0 dso_as5401[10]
rlabel metal2 24610 54179 24610 54179 0 dso_as5401[11]
rlabel metal2 25714 54179 25714 54179 0 dso_as5401[12]
rlabel metal2 26634 54247 26634 54247 0 dso_as5401[13]
rlabel metal2 28290 54179 28290 54179 0 dso_as5401[14]
rlabel metal2 29210 54240 29210 54240 0 dso_as5401[15]
rlabel metal2 30682 54179 30682 54179 0 dso_as5401[16]
rlabel metal2 31786 53499 31786 53499 0 dso_as5401[17]
rlabel metal1 32982 53074 32982 53074 0 dso_as5401[18]
rlabel metal2 34270 54179 34270 54179 0 dso_as5401[19]
rlabel metal2 12558 54179 12558 54179 0 dso_as5401[1]
rlabel metal2 35466 54179 35466 54179 0 dso_as5401[20]
rlabel metal2 36662 54179 36662 54179 0 dso_as5401[21]
rlabel metal2 37858 54179 37858 54179 0 dso_as5401[22]
rlabel metal2 39054 54179 39054 54179 0 dso_as5401[23]
rlabel metal1 40158 53074 40158 53074 0 dso_as5401[24]
rlabel metal2 41400 53074 41400 53074 0 dso_as5401[25]
rlabel metal1 42596 53074 42596 53074 0 dso_as5401[26]
rlabel metal2 13662 53968 13662 53968 0 dso_as5401[2]
rlabel metal2 14858 54172 14858 54172 0 dso_as5401[3]
rlabel metal2 16330 54179 16330 54179 0 dso_as5401[4]
rlabel metal2 17342 53907 17342 53907 0 dso_as5401[5]
rlabel metal1 18676 53074 18676 53074 0 dso_as5401[6]
rlabel metal1 19596 53074 19596 53074 0 dso_as5401[7]
rlabel metal2 20930 54179 20930 54179 0 dso_as5401[8]
rlabel metal1 22080 53074 22080 53074 0 dso_as5401[9]
rlabel metal1 47610 3026 47610 3026 0 dso_counter[0]
rlabel metal2 51842 3230 51842 3230 0 dso_counter[10]
rlabel metal2 51014 3672 51014 3672 0 dso_counter[11]
rlabel metal1 48024 2346 48024 2346 0 dso_counter[1]
rlabel metal1 48024 3366 48024 3366 0 dso_counter[2]
rlabel metal1 48668 2414 48668 2414 0 dso_counter[3]
rlabel metal1 48944 3026 48944 3026 0 dso_counter[4]
rlabel metal1 49772 2346 49772 2346 0 dso_counter[5]
rlabel metal1 50278 2992 50278 2992 0 dso_counter[6]
rlabel metal1 50508 2414 50508 2414 0 dso_counter[7]
rlabel metal1 51014 2958 51014 2958 0 dso_counter[8]
rlabel metal2 52026 2210 52026 2210 0 dso_counter[9]
rlabel metal1 44988 53074 44988 53074 0 dso_diceroll[0]
rlabel metal2 46046 53907 46046 53907 0 dso_diceroll[1]
rlabel metal2 47150 54240 47150 54240 0 dso_diceroll[2]
rlabel metal2 48438 53907 48438 53907 0 dso_diceroll[3]
rlabel metal2 49726 53431 49726 53431 0 dso_diceroll[4]
rlabel via1 51474 53142 51474 53142 0 dso_diceroll[5]
rlabel metal1 51750 52666 51750 52666 0 dso_diceroll[6]
rlabel metal2 53222 54179 53222 54179 0 dso_diceroll[7]
rlabel metal1 2622 28526 2622 28526 0 dso_mc14500[0]
rlabel metal1 2622 29070 2622 29070 0 dso_mc14500[1]
rlabel metal2 1610 29461 1610 29461 0 dso_mc14500[2]
rlabel via2 2254 29835 2254 29835 0 dso_mc14500[3]
rlabel metal1 2622 30702 2622 30702 0 dso_mc14500[4]
rlabel metal1 2622 31246 2622 31246 0 dso_mc14500[5]
rlabel metal1 2622 31790 2622 31790 0 dso_mc14500[6]
rlabel metal1 2622 32334 2622 32334 0 dso_mc14500[7]
rlabel metal2 1610 32725 1610 32725 0 dso_mc14500[8]
rlabel metal1 2162 53006 2162 53006 0 dso_multiplier[0]
rlabel metal2 3174 54213 3174 54213 0 dso_multiplier[1]
rlabel metal1 4140 53074 4140 53074 0 dso_multiplier[2]
rlabel metal2 5474 54213 5474 54213 0 dso_multiplier[3]
rlabel metal2 6670 54213 6670 54213 0 dso_multiplier[4]
rlabel metal2 7774 54179 7774 54179 0 dso_multiplier[5]
rlabel metal2 8602 54247 8602 54247 0 dso_multiplier[6]
rlabel metal2 10166 54179 10166 54179 0 dso_multiplier[7]
rlabel metal1 2622 33966 2622 33966 0 dso_tbb1143[0]
rlabel metal1 2622 34510 2622 34510 0 dso_tbb1143[1]
rlabel metal2 1610 34901 1610 34901 0 dso_tbb1143[2]
rlabel metal1 2622 35598 2622 35598 0 dso_tbb1143[3]
rlabel metal1 2668 36142 2668 36142 0 dso_tbb1143[4]
rlabel metal1 2622 36686 2622 36686 0 dso_tbb1143[5]
rlabel metal1 2622 37298 2622 37298 0 dso_tbb1143[6]
rlabel metal2 1610 37655 1610 37655 0 dso_tbb1143[7]
rlabel metal1 54280 52394 54280 52394 0 dso_tune
rlabel metal1 7038 2346 7038 2346 0 io_in[10]
rlabel metal2 8418 3298 8418 3298 0 io_in[11]
rlabel metal1 8326 3060 8326 3060 0 io_in[12]
rlabel metal2 9798 1761 9798 1761 0 io_in[13]
rlabel metal1 9752 3026 9752 3026 0 io_in[14]
rlabel metal2 10534 1761 10534 1761 0 io_in[15]
rlabel metal2 5474 2176 5474 2176 0 io_in[16]
rlabel metal1 10626 2414 10626 2414 0 io_in[17]
rlabel metal2 6026 2142 6026 2142 0 io_in[18]
rlabel metal2 12006 1707 12006 1707 0 io_in[19]
rlabel metal2 11638 3978 11638 3978 0 io_in[20]
rlabel metal1 9798 2550 9798 2550 0 io_in[21]
rlabel metal1 12558 2414 12558 2414 0 io_in[22]
rlabel metal2 13754 3706 13754 3706 0 io_in[23]
rlabel metal1 12190 2618 12190 2618 0 io_in[24]
rlabel metal1 13202 2414 13202 2414 0 io_in[25]
rlabel metal1 14168 3026 14168 3026 0 io_in[26]
rlabel viali 13570 2412 13570 2412 0 io_in[27]
rlabel metal2 15318 1761 15318 1761 0 io_in[28]
rlabel metal1 15134 2414 15134 2414 0 io_in[29]
rlabel metal1 15778 2414 15778 2414 0 io_in[30]
rlabel metal1 16284 3026 16284 3026 0 io_in[31]
rlabel metal2 16790 1588 16790 1588 0 io_in[32]
rlabel metal1 17066 2278 17066 2278 0 io_in[33]
rlabel metal2 17802 3196 17802 3196 0 io_in[34]
rlabel metal1 17756 2414 17756 2414 0 io_in[35]
rlabel metal2 18538 3196 18538 3196 0 io_in[36]
rlabel metal1 18446 2414 18446 2414 0 io_in[37]
rlabel metal1 6900 3502 6900 3502 0 io_in[5]
rlabel metal2 7222 1761 7222 1761 0 io_in[6]
rlabel metal1 7636 2414 7636 2414 0 io_in[7]
rlabel metal2 7958 1761 7958 1761 0 io_in[8]
rlabel metal2 7682 3468 7682 3468 0 io_in[9]
rlabel metal2 37030 1520 37030 1520 0 io_oeb[11]
rlabel metal2 37398 1656 37398 1656 0 io_oeb[12]
rlabel metal1 37858 2822 37858 2822 0 io_oeb[13]
rlabel metal2 38134 1520 38134 1520 0 io_oeb[14]
rlabel metal1 38640 2822 38640 2822 0 io_oeb[15]
rlabel metal1 39192 2822 39192 2822 0 io_oeb[16]
rlabel metal2 39238 1520 39238 1520 0 io_oeb[17]
rlabel metal1 39882 2822 39882 2822 0 io_oeb[18]
rlabel metal2 39974 1656 39974 1656 0 io_oeb[19]
rlabel metal1 40618 2822 40618 2822 0 io_oeb[20]
rlabel metal2 40710 1520 40710 1520 0 io_oeb[21]
rlabel metal2 41078 1792 41078 1792 0 io_oeb[22]
rlabel metal2 41446 1656 41446 1656 0 io_oeb[23]
rlabel metal1 42320 2822 42320 2822 0 io_oeb[24]
rlabel metal2 42182 1520 42182 1520 0 io_oeb[25]
rlabel metal1 42780 2890 42780 2890 0 io_oeb[26]
rlabel metal2 42918 1656 42918 1656 0 io_oeb[27]
rlabel metal1 43424 2890 43424 2890 0 io_oeb[28]
rlabel metal2 43654 1520 43654 1520 0 io_oeb[29]
rlabel metal1 44528 2890 44528 2890 0 io_oeb[30]
rlabel metal2 44390 1656 44390 1656 0 io_oeb[31]
rlabel metal1 45264 2822 45264 2822 0 io_oeb[32]
rlabel metal2 45126 1554 45126 1554 0 io_oeb[33]
rlabel metal1 46000 2890 46000 2890 0 io_oeb[34]
rlabel metal1 46000 3366 46000 3366 0 io_oeb[35]
rlabel metal2 46230 1656 46230 1656 0 io_oeb[36]
rlabel metal1 46690 3366 46690 3366 0 io_oeb[37]
rlabel metal2 23046 1520 23046 1520 0 io_out[11]
rlabel metal1 23460 2822 23460 2822 0 io_out[12]
rlabel metal2 23782 1520 23782 1520 0 io_out[13]
rlabel metal1 24196 2822 24196 2822 0 io_out[14]
rlabel metal2 24518 1520 24518 1520 0 io_out[15]
rlabel metal1 24978 3366 24978 3366 0 io_out[16]
rlabel metal1 25162 2822 25162 2822 0 io_out[17]
rlabel metal2 25622 1520 25622 1520 0 io_out[18]
rlabel metal1 25898 2822 25898 2822 0 io_out[19]
rlabel metal2 26358 1520 26358 1520 0 io_out[20]
rlabel metal1 26634 2822 26634 2822 0 io_out[21]
rlabel metal2 27094 1520 27094 1520 0 io_out[22]
rlabel metal1 27554 2822 27554 2822 0 io_out[23]
rlabel metal2 27830 1520 27830 1520 0 io_out[24]
rlabel metal1 28290 2822 28290 2822 0 io_out[25]
rlabel metal2 28566 1520 28566 1520 0 io_out[26]
rlabel metal2 28934 1656 28934 1656 0 io_out[27]
rlabel metal2 29302 1520 29302 1520 0 io_out[28]
rlabel metal2 29670 1520 29670 1520 0 io_out[29]
rlabel metal1 30130 2822 30130 2822 0 io_out[30]
rlabel metal2 30406 1656 30406 1656 0 io_out[31]
rlabel metal1 30866 2822 30866 2822 0 io_out[32]
rlabel metal2 31142 1520 31142 1520 0 io_out[33]
rlabel metal2 31510 1826 31510 1826 0 io_out[34]
rlabel metal2 31878 1656 31878 1656 0 io_out[35]
rlabel metal1 32706 2822 32706 2822 0 io_out[36]
rlabel metal2 32614 1520 32614 1520 0 io_out[37]
rlabel metal1 45540 35190 45540 35190 0 net1
rlabel metal1 53498 40392 53498 40392 0 net10
rlabel metal1 33350 52870 33350 52870 0 net100
rlabel metal2 12834 48450 12834 48450 0 net101
rlabel metal1 34822 52870 34822 52870 0 net102
rlabel metal1 35926 52870 35926 52870 0 net103
rlabel metal1 36202 52938 36202 52938 0 net104
rlabel metal1 36156 48246 36156 48246 0 net105
rlabel metal1 39514 52870 39514 52870 0 net106
rlabel metal2 41262 52734 41262 52734 0 net107
rlabel metal2 42642 52700 42642 52700 0 net108
rlabel metal2 14306 43452 14306 43452 0 net109
rlabel metal1 53130 40698 53130 40698 0 net11
rlabel metal1 15226 35088 15226 35088 0 net110
rlabel metal2 16054 51714 16054 51714 0 net111
rlabel metal1 20240 52462 20240 52462 0 net112
rlabel metal1 20056 53006 20056 53006 0 net113
rlabel metal1 21988 52938 21988 52938 0 net114
rlabel metal1 23368 53210 23368 53210 0 net115
rlabel metal1 24288 44438 24288 44438 0 net116
rlabel metal2 32614 34204 32614 34204 0 net117
rlabel metal2 51566 4658 51566 4658 0 net118
rlabel metal2 51198 17952 51198 17952 0 net119
rlabel metal1 53774 34646 53774 34646 0 net12
rlabel metal2 31786 33592 31786 33592 0 net120
rlabel metal1 41078 28458 41078 28458 0 net121
rlabel metal1 48530 2618 48530 2618 0 net122
rlabel metal2 33810 34238 33810 34238 0 net123
rlabel metal1 50186 2550 50186 2550 0 net124
rlabel metal2 27370 37655 27370 37655 0 net125
rlabel metal2 51106 5134 51106 5134 0 net126
rlabel metal1 23966 34510 23966 34510 0 net127
rlabel via2 51842 2363 51842 2363 0 net128
rlabel metal2 45494 51680 45494 51680 0 net129
rlabel metal1 35328 41990 35328 41990 0 net13
rlabel metal2 46322 45968 46322 45968 0 net130
rlabel metal2 48070 47532 48070 47532 0 net131
rlabel metal2 47058 52870 47058 52870 0 net132
rlabel metal1 50416 53006 50416 53006 0 net133
rlabel metal1 40710 52972 40710 52972 0 net134
rlabel via2 52026 52547 52026 52547 0 net135
rlabel metal2 49542 52360 49542 52360 0 net136
rlabel metal1 2162 28492 2162 28492 0 net137
rlabel metal2 4554 29376 4554 29376 0 net138
rlabel metal1 1794 29512 1794 29512 0 net139
rlabel metal1 52072 40698 52072 40698 0 net14
rlabel via2 26818 37179 26818 37179 0 net140
rlabel metal1 10028 30770 10028 30770 0 net141
rlabel metal1 11500 31314 11500 31314 0 net142
rlabel metal2 2162 31076 2162 31076 0 net143
rlabel metal1 2162 32300 2162 32300 0 net144
rlabel metal1 1794 32776 1794 32776 0 net145
rlabel metal1 3082 53040 3082 53040 0 net146
rlabel metal2 3266 43945 3266 43945 0 net147
rlabel metal1 24564 52122 24564 52122 0 net148
rlabel metal2 5566 45560 5566 45560 0 net149
rlabel metal1 52486 41174 52486 41174 0 net15
rlabel metal2 6762 43180 6762 43180 0 net150
rlabel metal1 9844 52870 9844 52870 0 net151
rlabel metal2 9338 52564 9338 52564 0 net152
rlabel metal2 10442 48654 10442 48654 0 net153
rlabel metal1 22908 36550 22908 36550 0 net154
rlabel metal1 4531 34578 4531 34578 0 net155
rlabel metal2 1794 34816 1794 34816 0 net156
rlabel metal2 15134 35836 15134 35836 0 net157
rlabel metal1 4531 36210 4531 36210 0 net158
rlabel metal2 17250 38284 17250 38284 0 net159
rlabel metal1 53406 41718 53406 41718 0 net16
rlabel metal1 2162 37196 2162 37196 0 net160
rlabel metal2 14858 38284 14858 38284 0 net161
rlabel metal2 54050 44132 54050 44132 0 net162
rlabel metal1 20194 2482 20194 2482 0 net163
rlabel metal1 8602 3434 8602 3434 0 net164
rlabel metal2 8510 3400 8510 3400 0 net165
rlabel metal1 9844 2890 9844 2890 0 net166
rlabel metal2 9798 3570 9798 3570 0 net167
rlabel metal2 13110 4182 13110 4182 0 net168
rlabel metal1 10488 2618 10488 2618 0 net169
rlabel metal1 32981 41616 32981 41616 0 net17
rlabel metal1 10902 2550 10902 2550 0 net170
rlabel metal1 11362 2618 11362 2618 0 net171
rlabel metal2 12926 3536 12926 3536 0 net172
rlabel metal1 12604 3706 12604 3706 0 net173
rlabel metal1 12834 2890 12834 2890 0 net174
rlabel metal1 12880 2278 12880 2278 0 net175
rlabel metal2 13386 6562 13386 6562 0 net176
rlabel metal1 13478 3162 13478 3162 0 net177
rlabel metal2 13110 2689 13110 2689 0 net178
rlabel metal1 14122 3162 14122 3162 0 net179
rlabel metal1 35328 43078 35328 43078 0 net18
rlabel metal1 14030 2618 14030 2618 0 net180
rlabel metal2 15594 6834 15594 6834 0 net181
rlabel metal1 15502 2550 15502 2550 0 net182
rlabel metal1 15962 2618 15962 2618 0 net183
rlabel metal1 16468 3162 16468 3162 0 net184
rlabel metal1 16698 2618 16698 2618 0 net185
rlabel metal1 16836 10166 16836 10166 0 net186
rlabel metal1 17434 8330 17434 8330 0 net187
rlabel metal1 17250 6868 17250 6868 0 net188
rlabel metal1 17710 7242 17710 7242 0 net189
rlabel metal1 45540 41616 45540 41616 0 net19
rlabel metal1 17756 7990 17756 7990 0 net190
rlabel metal2 7130 4420 7130 4420 0 net191
rlabel metal1 9522 3026 9522 3026 0 net192
rlabel metal1 22218 2618 22218 2618 0 net193
rlabel metal2 12466 6222 12466 6222 0 net194
rlabel metal1 15502 2856 15502 2856 0 net195
rlabel metal2 53682 34204 53682 34204 0 net196
rlabel metal1 54050 50694 54050 50694 0 net197
rlabel metal2 4370 37978 4370 37978 0 net198
rlabel metal2 43930 43792 43930 43792 0 net199
rlabel metal1 52210 38896 52210 38896 0 net2
rlabel metal1 52854 36040 52854 36040 0 net20
rlabel metal1 2162 33388 2162 33388 0 net200
rlabel metal1 33396 12818 33396 12818 0 net201
rlabel metal2 53774 20298 53774 20298 0 net202
rlabel metal1 38778 24820 38778 24820 0 net203
rlabel metal1 38502 16014 38502 16014 0 net204
rlabel metal1 52624 8942 52624 8942 0 net205
rlabel metal2 36662 8296 36662 8296 0 net206
rlabel metal2 53314 16847 53314 16847 0 net207
rlabel metal2 54142 17578 54142 17578 0 net208
rlabel metal2 40250 17663 40250 17663 0 net209
rlabel metal1 53774 35564 53774 35564 0 net21
rlabel metal1 32246 16626 32246 16626 0 net210
rlabel via2 53314 20451 53314 20451 0 net211
rlabel metal1 20378 13906 20378 13906 0 net212
rlabel metal2 53314 21743 53314 21743 0 net213
rlabel via2 54050 21947 54050 21947 0 net214
rlabel metal2 18814 22379 18814 22379 0 net215
rlabel metal1 18400 15334 18400 15334 0 net216
rlabel metal2 38686 8738 38686 8738 0 net217
rlabel metal2 54142 23902 54142 23902 0 net218
rlabel metal1 19136 17170 19136 17170 0 net219
rlabel metal2 49634 36414 49634 36414 0 net22
rlabel metal1 20562 19346 20562 19346 0 net220
rlabel metal2 20010 20434 20010 20434 0 net221
rlabel metal1 20654 18326 20654 18326 0 net222
rlabel metal1 18308 18122 18308 18122 0 net223
rlabel via2 20930 16099 20930 16099 0 net224
rlabel metal2 53406 10200 53406 10200 0 net225
rlabel metal2 53360 9660 53360 9660 0 net226
rlabel metal2 52486 9214 52486 9214 0 net227
rlabel metal1 18584 7718 18584 7718 0 net228
rlabel metal2 53314 13634 53314 13634 0 net229
rlabel metal2 53774 36516 53774 36516 0 net23
rlabel metal2 53866 13396 53866 13396 0 net230
rlabel metal2 53314 15776 53314 15776 0 net231
rlabel via2 14766 15011 14766 15011 0 net232
rlabel metal1 53314 8874 53314 8874 0 net233
rlabel metal2 53590 8568 53590 8568 0 net234
rlabel metal1 20746 17238 20746 17238 0 net235
rlabel metal1 1886 3570 1886 3570 0 net236
rlabel metal1 2323 8942 2323 8942 0 net237
rlabel metal1 14030 9520 14030 9520 0 net238
rlabel metal1 15318 9350 15318 9350 0 net239
rlabel metal1 45540 36720 45540 36720 0 net24
rlabel metal2 15042 10438 15042 10438 0 net240
rlabel metal2 11086 10948 11086 10948 0 net241
rlabel metal1 2323 11730 2323 11730 0 net242
rlabel metal2 15778 12070 15778 12070 0 net243
rlabel metal1 4393 12818 4393 12818 0 net244
rlabel metal2 1886 13124 1886 13124 0 net245
rlabel metal2 4370 14110 4370 14110 0 net246
rlabel metal2 10442 3910 10442 3910 0 net247
rlabel metal1 15732 13702 15732 13702 0 net248
rlabel metal2 4646 14722 4646 14722 0 net249
rlabel metal1 49542 37808 49542 37808 0 net25
rlabel metal2 15594 15028 15594 15028 0 net250
rlabel metal1 4393 16082 4393 16082 0 net251
rlabel metal2 16606 15572 16606 15572 0 net252
rlabel metal1 16652 15674 16652 15674 0 net253
rlabel metal1 16146 16218 16146 16218 0 net254
rlabel metal2 10534 4318 10534 4318 0 net255
rlabel metal2 10534 4998 10534 4998 0 net256
rlabel metal2 12466 5508 12466 5508 0 net257
rlabel metal2 13110 6086 13110 6086 0 net258
rlabel metal2 13018 6596 13018 6596 0 net259
rlabel metal2 53774 38964 53774 38964 0 net26
rlabel metal2 11086 7106 11086 7106 0 net260
rlabel metal1 2323 7854 2323 7854 0 net261
rlabel metal2 11086 7990 11086 7990 0 net262
rlabel metal1 37168 2414 37168 2414 0 net263
rlabel metal1 38088 2414 38088 2414 0 net264
rlabel metal2 38134 3196 38134 3196 0 net265
rlabel metal1 38870 2414 38870 2414 0 net266
rlabel metal1 14674 12070 14674 12070 0 net267
rlabel metal2 13754 13124 13754 13124 0 net268
rlabel metal1 39606 3366 39606 3366 0 net269
rlabel metal2 44206 36448 44206 36448 0 net27
rlabel metal1 14858 14450 14858 14450 0 net270
rlabel metal1 40526 3366 40526 3366 0 net271
rlabel metal1 15870 7922 15870 7922 0 net272
rlabel metal1 41216 3638 41216 3638 0 net273
rlabel metal2 14674 8211 14674 8211 0 net274
rlabel metal1 42964 2414 42964 2414 0 net275
rlabel metal1 15226 14246 15226 14246 0 net276
rlabel metal1 43378 2448 43378 2448 0 net277
rlabel metal1 16238 16490 16238 16490 0 net278
rlabel metal1 44022 2414 44022 2414 0 net279
rlabel metal2 1794 23902 1794 23902 0 net28
rlabel metal2 44114 3196 44114 3196 0 net280
rlabel metal1 44850 3366 44850 3366 0 net281
rlabel metal1 44758 3026 44758 3026 0 net282
rlabel metal1 45862 2414 45862 2414 0 net283
rlabel metal2 45586 3196 45586 3196 0 net284
rlabel metal1 46184 2482 46184 2482 0 net285
rlabel metal2 46322 3468 46322 3468 0 net286
rlabel metal2 45954 3978 45954 3978 0 net287
rlabel metal1 47242 3910 47242 3910 0 net288
rlabel metal1 16836 15062 16836 15062 0 net289
rlabel metal2 4094 24208 4094 24208 0 net29
rlabel metal3 32545 13668 32545 13668 0 net290
rlabel via3 30613 15164 30613 15164 0 net291
rlabel metal1 32315 7310 32315 7310 0 net292
rlabel metal2 32246 5508 32246 5508 0 net293
rlabel metal1 23644 2414 23644 2414 0 net294
rlabel metal2 29854 19516 29854 19516 0 net295
rlabel metal1 27629 13294 27629 13294 0 net296
rlabel metal1 24978 2414 24978 2414 0 net297
rlabel metal1 18078 14586 18078 14586 0 net298
rlabel metal1 25760 2414 25760 2414 0 net299
rlabel metal1 52118 37740 52118 37740 0 net3
rlabel metal1 1794 25160 1794 25160 0 net30
rlabel via3 29325 35972 29325 35972 0 net300
rlabel metal1 27002 3434 27002 3434 0 net301
rlabel metal2 28106 15521 28106 15521 0 net302
rlabel metal1 27692 2414 27692 2414 0 net303
rlabel metal2 28796 20876 28796 20876 0 net304
rlabel metal1 28382 2414 28382 2414 0 net305
rlabel metal1 29992 2414 29992 2414 0 net306
rlabel metal1 29440 2414 29440 2414 0 net307
rlabel metal1 30866 2414 30866 2414 0 net308
rlabel metal2 32430 28186 32430 28186 0 net309
rlabel metal1 8188 25738 8188 25738 0 net31
rlabel metal1 31648 2414 31648 2414 0 net310
rlabel metal1 35880 39338 35880 39338 0 net311
rlabel metal1 32752 2414 32752 2414 0 net312
rlabel metal2 36340 17204 36340 17204 0 net313
rlabel metal1 33580 2414 33580 2414 0 net314
rlabel metal1 32062 40358 32062 40358 0 net315
rlabel metal1 34086 2380 34086 2380 0 net316
rlabel metal1 2530 18938 2530 18938 0 net317
rlabel metal2 14306 19516 14306 19516 0 net318
rlabel metal1 2484 20026 2484 20026 0 net319
rlabel metal1 4531 26418 4531 26418 0 net32
rlabel metal1 2162 20434 2162 20434 0 net320
rlabel metal2 13938 21114 13938 21114 0 net321
rlabel metal2 2438 21318 2438 21318 0 net322
rlabel metal2 2438 21828 2438 21828 0 net323
rlabel metal2 1886 22372 1886 22372 0 net324
rlabel metal2 2346 22916 2346 22916 0 net325
rlabel metal1 2162 23698 2162 23698 0 net326
rlabel metal2 54326 7242 54326 7242 0 net327
rlabel metal1 51198 8500 51198 8500 0 net328
rlabel metal1 54050 16490 54050 16490 0 net329
rlabel metal1 2162 26860 2162 26860 0 net33
rlabel metal1 39330 17578 39330 17578 0 net330
rlabel metal2 53498 17408 53498 17408 0 net331
rlabel metal1 54050 19278 54050 19278 0 net332
rlabel metal2 40802 19550 40802 19550 0 net333
rlabel metal1 52555 20910 52555 20910 0 net334
rlabel metal1 52555 21522 52555 21522 0 net335
rlabel metal2 39790 21998 39790 21998 0 net336
rlabel metal1 52555 23086 52555 23086 0 net337
rlabel metal2 40342 23052 40342 23052 0 net338
rlabel metal2 52302 9180 52302 9180 0 net339
rlabel metal1 1794 27336 1794 27336 0 net34
rlabel metal1 40158 22984 40158 22984 0 net340
rlabel metal1 39422 24582 39422 24582 0 net341
rlabel metal1 39330 23494 39330 23494 0 net342
rlabel metal1 37352 26554 37352 26554 0 net343
rlabel metal1 35282 24922 35282 24922 0 net344
rlabel metal1 35742 26486 35742 26486 0 net345
rlabel metal2 37674 27744 37674 27744 0 net346
rlabel metal1 40020 10098 40020 10098 0 net347
rlabel metal2 51106 11458 51106 11458 0 net348
rlabel via2 37766 12291 37766 12291 0 net349
rlabel metal2 2714 27268 2714 27268 0 net35
rlabel metal2 39422 12988 39422 12988 0 net350
rlabel metal2 54050 13498 54050 13498 0 net351
rlabel metal2 54050 14212 54050 14212 0 net352
rlabel metal2 54050 14943 54050 14943 0 net353
rlabel metal2 54050 15878 54050 15878 0 net354
rlabel metal2 42734 3910 42734 3910 0 net355
rlabel metal1 18975 3706 18975 3706 0 net356
rlabel metal1 19044 2822 19044 2822 0 net357
rlabel metal2 19366 1588 19366 1588 0 net358
rlabel metal2 19734 823 19734 823 0 net359
rlabel metal2 52578 42534 52578 42534 0 net36
rlabel metal2 20102 1792 20102 1792 0 net360
rlabel metal1 20516 2822 20516 2822 0 net361
rlabel metal2 20838 1656 20838 1656 0 net362
rlabel metal2 21206 1588 21206 1588 0 net363
rlabel metal1 21528 2822 21528 2822 0 net364
rlabel metal2 21942 1588 21942 1588 0 net365
rlabel metal2 22310 1792 22310 1792 0 net366
rlabel metal1 22724 2822 22724 2822 0 net367
rlabel metal2 54326 30957 54326 30957 0 net368
rlabel metal3 54794 31620 54794 31620 0 net369
rlabel via2 52486 44931 52486 44931 0 net37
rlabel metal2 54326 32657 54326 32657 0 net370
rlabel via2 54326 33269 54326 33269 0 net371
rlabel metal1 53176 35054 53176 35054 0 net372
rlabel metal1 33396 2958 33396 2958 0 net373
rlabel metal2 33350 959 33350 959 0 net374
rlabel metal1 34086 2890 34086 2890 0 net375
rlabel metal2 34086 1588 34086 1588 0 net376
rlabel metal1 34776 3094 34776 3094 0 net377
rlabel metal2 34822 1554 34822 1554 0 net378
rlabel metal2 35190 1163 35190 1163 0 net379
rlabel metal2 47058 45730 47058 45730 0 net38
rlabel metal1 35972 3026 35972 3026 0 net380
rlabel metal1 35972 3366 35972 3366 0 net381
rlabel metal1 36478 3366 36478 3366 0 net382
rlabel metal1 36708 4182 36708 4182 0 net383
rlabel metal1 35328 23086 35328 23086 0 net384
rlabel metal1 34812 20434 34812 20434 0 net385
rlabel metal1 33718 18734 33718 18734 0 net386
rlabel metal2 31694 19040 31694 19040 0 net387
rlabel metal1 29992 16082 29992 16082 0 net388
rlabel metal2 31050 16966 31050 16966 0 net389
rlabel metal1 28704 41786 28704 41786 0 net39
rlabel metal1 35696 18054 35696 18054 0 net390
rlabel metal1 34817 18326 34817 18326 0 net391
rlabel metal1 24334 16694 24334 16694 0 net392
rlabel metal1 24794 17238 24794 17238 0 net393
rlabel metal1 26270 17238 26270 17238 0 net394
rlabel metal2 36294 19040 36294 19040 0 net395
rlabel metal1 34438 19414 34438 19414 0 net396
rlabel metal1 27140 18734 27140 18734 0 net397
rlabel metal1 26036 19482 26036 19482 0 net398
rlabel metal2 23690 18938 23690 18938 0 net399
rlabel metal2 53590 37723 53590 37723 0 net4
rlabel metal2 52946 45968 52946 45968 0 net40
rlabel via1 25249 18258 25249 18258 0 net400
rlabel metal1 24978 13294 24978 13294 0 net401
rlabel metal1 26174 13498 26174 13498 0 net402
rlabel metal2 32890 13940 32890 13940 0 net403
rlabel metal1 33820 14994 33820 14994 0 net404
rlabel metal1 22724 13226 22724 13226 0 net405
rlabel metal1 20930 12614 20930 12614 0 net406
rlabel metal1 25663 13906 25663 13906 0 net407
rlabel metal2 36386 13294 36386 13294 0 net408
rlabel via1 36022 13226 36022 13226 0 net409
rlabel metal1 45540 43656 45540 43656 0 net41
rlabel metal1 35604 10982 35604 10982 0 net410
rlabel via1 34449 13906 34449 13906 0 net411
rlabel metal1 28106 12070 28106 12070 0 net412
rlabel metal2 28842 12988 28842 12988 0 net413
rlabel metal2 28014 13430 28014 13430 0 net414
rlabel metal1 33074 18326 33074 18326 0 net415
rlabel metal1 33442 19278 33442 19278 0 net416
rlabel metal1 29716 16558 29716 16558 0 net417
rlabel metal1 36984 18938 36984 18938 0 net418
rlabel metal1 38226 19210 38226 19210 0 net419
rlabel metal2 52762 45662 52762 45662 0 net42
rlabel metal2 39514 20026 39514 20026 0 net420
rlabel metal1 29026 19278 29026 19278 0 net421
rlabel metal2 28290 17272 28290 17272 0 net422
rlabel metal1 30222 20468 30222 20468 0 net423
rlabel metal1 28888 19958 28888 19958 0 net424
rlabel metal2 29578 19516 29578 19516 0 net425
rlabel metal2 32890 19516 32890 19516 0 net426
rlabel metal1 30268 19210 30268 19210 0 net427
rlabel metal1 36892 19822 36892 19822 0 net428
rlabel metal2 26634 21522 26634 21522 0 net429
rlabel metal1 51612 46478 51612 46478 0 net43
rlabel metal1 33212 12070 33212 12070 0 net430
rlabel metal1 30222 13362 30222 13362 0 net431
rlabel metal1 34316 15674 34316 15674 0 net432
rlabel via2 25346 14909 25346 14909 0 net433
rlabel metal2 29210 15130 29210 15130 0 net434
rlabel metal1 25024 16218 25024 16218 0 net435
rlabel metal2 32154 13940 32154 13940 0 net436
rlabel metal1 30682 14858 30682 14858 0 net437
rlabel metal1 35236 12886 35236 12886 0 net438
rlabel metal2 53038 47498 53038 47498 0 net44
rlabel metal1 33396 46546 33396 46546 0 net45
rlabel metal2 51382 47770 51382 47770 0 net46
rlabel via2 53774 42755 53774 42755 0 net47
rlabel metal2 48162 48110 48162 48110 0 net48
rlabel metal1 52256 47022 52256 47022 0 net49
rlabel metal2 34454 38964 34454 38964 0 net5
rlabel metal1 45540 48552 45540 48552 0 net50
rlabel metal1 52348 47634 52348 47634 0 net51
rlabel metal1 35558 47634 35558 47634 0 net52
rlabel metal1 45540 49232 45540 49232 0 net53
rlabel metal2 38778 45152 38778 45152 0 net54
rlabel metal1 45540 40664 45540 40664 0 net55
rlabel metal1 45540 43248 45540 43248 0 net56
rlabel metal1 45540 41038 45540 41038 0 net57
rlabel metal2 52854 37366 52854 37366 0 net58
rlabel metal1 45540 37910 45540 37910 0 net59
rlabel metal1 46230 39984 46230 39984 0 net6
rlabel via2 53774 45475 53774 45475 0 net60
rlabel metal1 41400 43384 41400 43384 0 net61
rlabel metal2 52670 45220 52670 45220 0 net62
rlabel metal1 4531 38930 4531 38930 0 net63
rlabel metal2 2254 40477 2254 40477 0 net64
rlabel metal1 2162 44812 2162 44812 0 net65
rlabel metal1 2162 45356 2162 45356 0 net66
rlabel metal1 2254 45934 2254 45934 0 net67
rlabel metal1 2392 46546 2392 46546 0 net68
rlabel metal1 2438 47090 2438 47090 0 net69
rlabel via2 52118 38947 52118 38947 0 net7
rlabel metal2 29118 47430 29118 47430 0 net70
rlabel metal1 2162 48076 2162 48076 0 net71
rlabel metal2 2254 47532 2254 47532 0 net72
rlabel metal2 2346 48348 2346 48348 0 net73
rlabel metal1 4531 39474 4531 39474 0 net74
rlabel metal1 1978 49742 1978 49742 0 net75
rlabel metal2 2162 49402 2162 49402 0 net76
rlabel metal2 2438 47685 2438 47685 0 net77
rlabel metal2 2714 49606 2714 49606 0 net78
rlabel metal2 1886 47600 1886 47600 0 net79
rlabel metal1 49496 39610 49496 39610 0 net8
rlabel metal1 1840 52462 1840 52462 0 net80
rlabel metal1 2576 52462 2576 52462 0 net81
rlabel metal1 30020 40018 30020 40018 0 net82
rlabel metal2 2162 39202 2162 39202 0 net83
rlabel metal1 4531 41106 4531 41106 0 net84
rlabel metal2 24518 41446 24518 41446 0 net85
rlabel metal2 2346 39780 2346 39780 0 net86
rlabel metal1 2162 42636 2162 42636 0 net87
rlabel metal1 2346 43282 2346 43282 0 net88
rlabel metal2 2070 38335 2070 38335 0 net89
rlabel metal1 54004 46954 54004 46954 0 net9
rlabel metal2 11638 47821 11638 47821 0 net90
rlabel metal2 25438 52462 25438 52462 0 net91
rlabel metal1 25760 52938 25760 52938 0 net92
rlabel metal1 25944 52870 25944 52870 0 net93
rlabel metal1 27186 52870 27186 52870 0 net94
rlabel metal1 27968 52054 27968 52054 0 net95
rlabel metal1 29256 52870 29256 52870 0 net96
rlabel metal1 30314 52870 30314 52870 0 net97
rlabel metal1 31786 52870 31786 52870 0 net98
rlabel metal1 32568 52938 32568 52938 0 net99
rlabel metal2 53038 34425 53038 34425 0 oeb_6502
rlabel metal1 54096 51306 54096 51306 0 oeb_as1802
rlabel metal2 1702 38131 1702 38131 0 oeb_as2650
rlabel metal2 43654 54179 43654 54179 0 oeb_as5401
rlabel metal1 2622 33422 2622 33422 0 oeb_mc14500
rlabel metal3 1188 18428 1188 18428 0 rst_6502
rlabel metal3 1188 18972 1188 18972 0 rst_LCD
rlabel metal3 1188 19516 1188 19516 0 rst_as1802
rlabel metal3 1188 20060 1188 20060 0 rst_as2650
rlabel metal3 1188 20604 1188 20604 0 rst_as5401
rlabel metal3 1188 21148 1188 21148 0 rst_counter
rlabel metal3 1188 21692 1188 21692 0 rst_diceroll
rlabel metal3 1188 22236 1188 22236 0 rst_mc14500
rlabel metal3 1188 22780 1188 22780 0 rst_tbb1143
rlabel metal3 1188 23324 1188 23324 0 rst_tune
rlabel metal2 51290 6715 51290 6715 0 wb_clk_i
rlabel metal2 23598 11016 23598 11016 0 wb_clk_override
rlabel metal1 35696 14042 35696 14042 0 wb_counter\[0\]
rlabel metal1 25392 16558 25392 16558 0 wb_counter\[10\]
rlabel metal1 27554 18054 27554 18054 0 wb_counter\[11\]
rlabel metal1 32798 16626 32798 16626 0 wb_counter\[12\]
rlabel metal2 28842 17850 28842 17850 0 wb_counter\[13\]
rlabel metal1 25576 20774 25576 20774 0 wb_counter\[14\]
rlabel metal1 25898 21556 25898 21556 0 wb_counter\[15\]
rlabel metal1 27692 21522 27692 21522 0 wb_counter\[16\]
rlabel metal1 32614 21522 32614 21522 0 wb_counter\[17\]
rlabel metal1 33534 21998 33534 21998 0 wb_counter\[18\]
rlabel metal1 32154 21998 32154 21998 0 wb_counter\[19\]
rlabel metal3 36156 13124 36156 13124 0 wb_counter\[1\]
rlabel metal1 35512 20842 35512 20842 0 wb_counter\[20\]
rlabel metal1 36064 18190 36064 18190 0 wb_counter\[21\]
rlabel metal1 37766 18802 37766 18802 0 wb_counter\[22\]
rlabel metal2 37490 20944 37490 20944 0 wb_counter\[23\]
rlabel metal2 35374 13532 35374 13532 0 wb_counter\[2\]
rlabel metal1 32246 9418 32246 9418 0 wb_counter\[3\]
rlabel metal2 33534 14076 33534 14076 0 wb_counter\[4\]
rlabel metal1 31464 13362 31464 13362 0 wb_counter\[5\]
rlabel metal2 20194 13056 20194 13056 0 wb_counter\[6\]
rlabel metal2 26634 14042 26634 14042 0 wb_counter\[7\]
rlabel metal1 26542 14586 26542 14586 0 wb_counter\[8\]
rlabel metal1 26174 15674 26174 15674 0 wb_counter\[9\]
rlabel metal2 31786 9622 31786 9622 0 wb_design_addr_override\[0\]
rlabel metal1 30912 8330 30912 8330 0 wb_design_addr_override\[1\]
rlabel metal1 33994 11288 33994 11288 0 wb_design_addr_override\[2\]
rlabel metal1 31188 9146 31188 9146 0 wb_design_addr_override\[3\]
rlabel metal1 50508 9554 50508 9554 0 wb_feedback_delay
rlabel metal1 19688 7242 19688 7242 0 wb_io_override\[0\]
rlabel metal1 19918 9996 19918 9996 0 wb_io_override\[10\]
rlabel metal1 18768 10982 18768 10982 0 wb_io_override\[11\]
rlabel metal1 20056 10982 20056 10982 0 wb_io_override\[12\]
rlabel metal1 21114 11594 21114 11594 0 wb_io_override\[13\]
rlabel metal1 18400 12206 18400 12206 0 wb_io_override\[14\]
rlabel metal2 21482 12750 21482 12750 0 wb_io_override\[15\]
rlabel metal1 20930 14892 20930 14892 0 wb_io_override\[16\]
rlabel metal2 18262 13464 18262 13464 0 wb_io_override\[17\]
rlabel metal1 17756 13158 17756 13158 0 wb_io_override\[18\]
rlabel metal1 18492 14042 18492 14042 0 wb_io_override\[19\]
rlabel metal2 24978 4250 24978 4250 0 wb_io_override\[1\]
rlabel metal1 21114 19482 21114 19482 0 wb_io_override\[20\]
rlabel metal1 20010 16422 20010 16422 0 wb_io_override\[21\]
rlabel metal2 21206 19074 21206 19074 0 wb_io_override\[22\]
rlabel metal1 18584 19482 18584 19482 0 wb_io_override\[23\]
rlabel metal1 20792 17510 20792 17510 0 wb_io_override\[24\]
rlabel metal1 21298 15606 21298 15606 0 wb_io_override\[25\]
rlabel metal1 20838 16218 20838 16218 0 wb_io_override\[26\]
rlabel metal1 21252 8330 21252 8330 0 wb_io_override\[2\]
rlabel metal2 21298 6188 21298 6188 0 wb_io_override\[3\]
rlabel metal1 22770 6630 22770 6630 0 wb_io_override\[4\]
rlabel metal1 19366 6630 19366 6630 0 wb_io_override\[5\]
rlabel metal1 24610 8330 24610 8330 0 wb_io_override\[6\]
rlabel metal1 20654 6732 20654 6732 0 wb_io_override\[7\]
rlabel metal2 19642 8092 19642 8092 0 wb_io_override\[8\]
rlabel metal1 18492 7174 18492 7174 0 wb_io_override\[9\]
rlabel metal1 23414 9690 23414 9690 0 wb_override
rlabel metal1 54326 7378 54326 7378 0 wb_rst_i
rlabel metal2 32062 8976 32062 8976 0 wb_rst_override
rlabel metal2 23690 10506 23690 10506 0 wb_single_step
rlabel metal2 54142 7055 54142 7055 0 wbs_ack_o
rlabel metal2 53498 25585 53498 25585 0 wbs_adr_i[21]
rlabel metal2 53590 26265 53590 26265 0 wbs_adr_i[22]
rlabel metal2 53498 27217 53498 27217 0 wbs_adr_i[23]
rlabel metal2 52302 7633 52302 7633 0 wbs_cyc_i
rlabel via2 53498 8483 53498 8483 0 wbs_dat_i[0]
rlabel via2 53590 16677 53590 16677 0 wbs_dat_i[10]
rlabel metal2 54234 17357 54234 17357 0 wbs_dat_i[11]
rlabel metal2 53498 18479 53498 18479 0 wbs_dat_i[12]
rlabel metal2 54234 18921 54234 18921 0 wbs_dat_i[13]
rlabel via2 53590 19941 53590 19941 0 wbs_dat_i[14]
rlabel metal2 54234 20621 54234 20621 0 wbs_dat_i[15]
rlabel metal2 53498 21743 53498 21743 0 wbs_dat_i[16]
rlabel metal2 53590 21828 53590 21828 0 wbs_dat_i[17]
rlabel via2 53590 23205 53590 23205 0 wbs_dat_i[18]
rlabel metal2 54234 23885 54234 23885 0 wbs_dat_i[19]
rlabel metal3 54426 9316 54426 9316 0 wbs_dat_i[1]
rlabel metal2 54234 24497 54234 24497 0 wbs_dat_i[20]
rlabel metal1 53912 24786 53912 24786 0 wbs_dat_i[21]
rlabel metal1 53544 26962 53544 26962 0 wbs_dat_i[22]
rlabel metal2 54234 27149 54234 27149 0 wbs_dat_i[23]
rlabel metal2 53498 28271 53498 28271 0 wbs_dat_i[24]
rlabel metal2 54234 28713 54234 28713 0 wbs_dat_i[25]
rlabel metal2 54234 29665 54234 29665 0 wbs_dat_i[26]
rlabel via2 53498 10149 53498 10149 0 wbs_dat_i[2]
rlabel metal2 54234 10829 54234 10829 0 wbs_dat_i[3]
rlabel metal2 53498 11951 53498 11951 0 wbs_dat_i[4]
rlabel metal2 54234 12393 54234 12393 0 wbs_dat_i[5]
rlabel via2 53590 13413 53590 13413 0 wbs_dat_i[6]
rlabel metal2 54234 14093 54234 14093 0 wbs_dat_i[7]
rlabel metal2 53498 15215 53498 15215 0 wbs_dat_i[8]
rlabel metal2 54234 15657 54234 15657 0 wbs_dat_i[9]
rlabel metal2 54234 8687 54234 8687 0 wbs_dat_o[0]
rlabel metal2 54234 16847 54234 16847 0 wbs_dat_o[10]
rlabel via2 54234 17765 54234 17765 0 wbs_dat_o[11]
rlabel metal2 54234 18479 54234 18479 0 wbs_dat_o[12]
rlabel metal2 54234 19431 54234 19431 0 wbs_dat_o[13]
rlabel metal2 54234 20111 54234 20111 0 wbs_dat_o[14]
rlabel via2 54234 21029 54234 21029 0 wbs_dat_o[15]
rlabel metal2 54234 21743 54234 21743 0 wbs_dat_o[16]
rlabel metal2 54234 22695 54234 22695 0 wbs_dat_o[17]
rlabel metal2 54234 23375 54234 23375 0 wbs_dat_o[18]
rlabel metal2 53498 24429 53498 24429 0 wbs_dat_o[19]
rlabel metal2 54234 9503 54234 9503 0 wbs_dat_o[1]
rlabel via2 53498 25109 53498 25109 0 wbs_dat_o[20]
rlabel metal2 54234 25687 54234 25687 0 wbs_dat_o[21]
rlabel metal2 54234 26639 54234 26639 0 wbs_dat_o[22]
rlabel metal2 53498 27693 53498 27693 0 wbs_dat_o[23]
rlabel metal2 54234 28271 54234 28271 0 wbs_dat_o[24]
rlabel metal2 54234 29223 54234 29223 0 wbs_dat_o[25]
rlabel via2 54234 30005 54234 30005 0 wbs_dat_o[26]
rlabel metal2 54234 10319 54234 10319 0 wbs_dat_o[2]
rlabel via2 54234 11237 54234 11237 0 wbs_dat_o[3]
rlabel metal2 54234 11951 54234 11951 0 wbs_dat_o[4]
rlabel metal2 54234 12903 54234 12903 0 wbs_dat_o[5]
rlabel metal2 54234 13583 54234 13583 0 wbs_dat_o[6]
rlabel via2 54234 14501 54234 14501 0 wbs_dat_o[7]
rlabel metal2 54234 15215 54234 15215 0 wbs_dat_o[8]
rlabel metal2 54234 16167 54234 16167 0 wbs_dat_o[9]
rlabel metal2 53406 7531 53406 7531 0 wbs_stb_i
rlabel metal2 52210 8211 52210 8211 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 56000 56000
<< end >>
